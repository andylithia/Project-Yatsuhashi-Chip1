** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA24_2.sch
**.subckt LNA24_2
XM1 n_ds1 vgate1 net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=5 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=12 m=12
Ldeg1 net1 GND 2n m=1
V1 net2 GND 1.8
V2 net3 GND dc 0 ac 0 portnum 1 z0 50
C2 net8 net3 1u m=1
V3 net4 GND dc 0 ac 0 portnum 2 z0 50
C4 net4 net5 0.1p m=1
Ldeg2 net7 net8 7n m=1
R1 vbias1 net7 5k m=1
Lload1 net2 net5 5n m=1
V4 vbias1 GND 1.2
XM2 net5 net2 net6 GND sky130_fd_pr__nfet_01v8 L=0.15 W=15 nf=5 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=12 m=12
Lcpl net6 n_ds1 1n m=1
K1 Ldeg1 Lcpli 0.9
Lcpli vgate1 net7 0 m=1
C1 net1 vgate1 50f m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.param L=0.18
.param Ls=0.5n
.param W=10
.param W2=20
.param NF=1
.param M=1
.op
.plot @m.xm1.msky130_fd_pr__nfet_01v8[vgs]
.plot @m.xm1.msky130_fd_pr__nfet_01v8[vds]
.print @m.xm3.msky130_fd_pr__nfet_01v8[vgs]
.print @m.xm3.msky130_fd_pr__nfet_01v8[vds]
.sp dec 1000 3e9 6e9 0
.control
run
display
plot db(S_1_1) db(S_1_2) db(S_2_2) db(S_2_1)
plot S_1_1 smithgrid
print @m.xm1.msky130_fd_pr__nfet_01v8[id]
print @m.xm1.msky130_fd_pr__nfet_01v8[vgs]
print @m.xm1.msky130_fd_pr__nfet_01v8[vds]
print @m.xm3.msky130_fd_pr__nfet_01v8[vgs]
print @m.xm3.msky130_fd_pr__nfet_01v8[vds]
print @m.xm3.msky130_fd_pr__nfet_01v8[id]
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
