* SPICE3 file created from ./COMMON/mimcap3_W2L5.ext - technology: sky130A

X0 top bot sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=5e+06u
C0 bot top 3.54fF
