magic
tech sky130A
magscale 1 2
timestamp 1658893076
<< metal1 >>
rect 26 1310 1266 1380
rect 26 100 84 1310
rect 140 1240 360 1260
rect 140 1160 160 1240
rect 240 1160 260 1240
rect 340 1160 360 1240
rect 140 1140 360 1160
rect 151 1128 353 1140
rect 420 302 478 1310
rect 530 1240 750 1260
rect 530 1160 550 1240
rect 630 1160 650 1240
rect 730 1160 750 1240
rect 530 1140 750 1160
rect 541 1128 743 1140
rect 814 302 872 1310
rect 930 1240 1150 1260
rect 930 1160 950 1240
rect 1030 1160 1050 1240
rect 1130 1160 1150 1240
rect 930 1140 1150 1160
rect 941 1128 1143 1140
rect 420 110 421 139
rect 814 110 815 139
rect 1208 100 1266 1310
rect 151 60 353 72
rect 541 60 743 72
rect 941 60 1143 72
rect 140 40 360 60
rect 140 -40 160 40
rect 240 -40 260 40
rect 340 -40 360 40
rect 140 -60 360 -40
rect 530 40 750 60
rect 530 -40 550 40
rect 630 -40 650 40
rect 730 -40 750 40
rect 530 -60 750 -40
rect 930 40 1150 60
rect 930 -40 950 40
rect 1030 -40 1050 40
rect 1130 -40 1150 40
rect 930 -60 1150 -40
<< via1 >>
rect 160 1160 240 1240
rect 260 1160 340 1240
rect 550 1160 630 1240
rect 650 1160 730 1240
rect 950 1160 1030 1240
rect 1050 1160 1130 1240
rect 160 -40 240 40
rect 260 -40 340 40
rect 550 -40 630 40
rect 650 -40 730 40
rect 950 -40 1030 40
rect 1050 -40 1130 40
<< metal2 >>
rect 140 1240 360 1260
rect 140 1160 160 1240
rect 240 1160 260 1240
rect 340 1160 360 1240
rect 140 1140 360 1160
rect 530 1240 750 1260
rect 530 1160 550 1240
rect 630 1160 650 1240
rect 730 1160 750 1240
rect 530 1140 750 1160
rect 930 1240 1150 1260
rect 930 1160 950 1240
rect 1030 1160 1050 1240
rect 1130 1160 1150 1240
rect 930 1140 1150 1160
rect 0 622 1292 1094
rect 0 100 1292 572
rect 140 40 360 60
rect 140 -40 160 40
rect 240 -40 260 40
rect 340 -40 360 40
rect 140 -60 360 -40
rect 530 40 750 60
rect 530 -40 550 40
rect 630 -40 650 40
rect 730 -40 750 40
rect 530 -60 750 -40
rect 930 40 1150 60
rect 930 -40 950 40
rect 1030 -40 1050 40
rect 1130 -40 1150 40
rect 930 -60 1150 -40
<< via2 >>
rect 160 1160 230 1240
rect 270 1160 340 1240
rect 550 1160 620 1240
rect 660 1160 730 1240
rect 950 1160 1020 1240
rect 1060 1160 1130 1240
rect 160 -40 230 40
rect 270 -40 340 40
rect 550 -40 620 40
rect 660 -40 730 40
rect 950 -40 1020 40
rect 1060 -40 1130 40
<< metal3 >>
rect 140 1240 1150 1260
rect 140 1160 160 1240
rect 230 1160 270 1240
rect 340 1160 550 1240
rect 620 1160 660 1240
rect 730 1160 950 1240
rect 1020 1160 1060 1240
rect 1130 1160 1150 1240
rect 140 1140 1150 1160
rect 400 60 500 1140
rect 800 60 900 1140
rect 140 40 1150 60
rect 140 -40 160 40
rect 230 -40 270 40
rect 340 -40 550 40
rect 620 -40 660 40
rect 730 -40 950 40
rect 1020 -40 1060 40
rect 1130 -40 1150 40
rect 140 -60 1150 -40
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1658893076
transform 1 0 -10 0 1 -10
box 10 10 514 1204
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1
timestamp 1658893076
transform -1 0 908 0 1 -10
box 10 10 514 1204
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2
timestamp 1658893076
transform 1 0 778 0 1 -10
box 10 10 514 1204
<< labels >>
rlabel metal1 26 1310 1266 1380 1 sub
rlabel metal3 140 1140 1140 1260 1 G
rlabel metal2 0 622 1292 1094 1 D
rlabel metal2 0 100 1292 572 1 S
<< end >>
