magic
tech sky130A
magscale 1 2
timestamp 1663721312
<< viali >>
rect 236 6432 4959 6470
rect 46 236 84 6280
rect 5054 236 5092 6280
rect 236 46 4902 84
<< metal1 >>
rect 30 6470 5110 6480
rect 30 6432 236 6470
rect 4959 6432 5110 6470
rect 30 6422 5110 6432
rect 30 6420 100 6422
rect 5040 6420 5110 6422
rect 232 6290 252 6390
rect 4886 6290 4906 6390
rect 165 6238 231 6258
rect 165 258 231 278
rect 323 6238 389 6258
rect 323 258 389 278
rect 481 6238 547 6258
rect 481 258 547 278
rect 639 6238 705 6258
rect 639 258 705 278
rect 797 6238 863 6258
rect 797 258 863 278
rect 955 6238 1021 6258
rect 955 258 1021 278
rect 1113 6238 1179 6258
rect 1113 258 1179 278
rect 1271 6238 1337 6258
rect 1271 258 1337 278
rect 1429 6238 1495 6258
rect 1429 258 1495 278
rect 1587 6238 1653 6258
rect 1587 258 1653 278
rect 1745 6238 1811 6258
rect 1745 258 1811 278
rect 1903 6238 1969 6258
rect 1903 258 1969 278
rect 2061 6238 2127 6258
rect 2061 258 2127 278
rect 2219 6238 2285 6258
rect 2219 258 2285 278
rect 2377 6238 2443 6258
rect 2377 258 2443 278
rect 2535 6238 2601 6258
rect 2535 258 2601 278
rect 2693 6238 2759 6258
rect 2693 258 2759 278
rect 2851 6238 2917 6258
rect 2851 258 2917 278
rect 3009 6238 3075 6258
rect 3009 258 3075 278
rect 3167 6238 3233 6258
rect 3167 258 3233 278
rect 3325 6238 3391 6258
rect 3325 258 3391 278
rect 3483 6238 3549 6258
rect 3483 258 3549 278
rect 3641 6238 3707 6258
rect 3641 258 3707 278
rect 3799 6238 3865 6258
rect 3799 258 3865 278
rect 3957 6238 4023 6258
rect 3957 258 4023 278
rect 4115 6238 4181 6258
rect 4115 258 4181 278
rect 4273 6238 4339 6258
rect 4273 258 4339 278
rect 4431 6238 4497 6258
rect 4431 258 4497 278
rect 4589 6238 4655 6258
rect 4589 258 4655 278
rect 4747 6238 4813 6258
rect 4747 258 4813 278
rect 4905 6238 4971 6258
rect 4905 258 4971 278
rect 232 126 252 226
rect 4886 126 4906 226
rect 30 94 100 100
rect 5040 94 5110 100
rect 30 84 5110 94
rect 30 46 236 84
rect 4902 46 5110 84
rect 30 30 5110 46
<< via1 >>
rect 30 6280 100 6420
rect 252 6290 4886 6390
rect 30 236 46 6280
rect 46 236 84 6280
rect 84 236 100 6280
rect 5040 6280 5110 6420
rect 165 278 231 6238
rect 323 278 389 6238
rect 481 278 547 6238
rect 639 278 705 6238
rect 797 278 863 6238
rect 955 278 1021 6238
rect 1113 278 1179 6238
rect 1271 278 1337 6238
rect 1429 278 1495 6238
rect 1587 278 1653 6238
rect 1745 278 1811 6238
rect 1903 278 1969 6238
rect 2061 278 2127 6238
rect 2219 278 2285 6238
rect 2377 278 2443 6238
rect 2535 278 2601 6238
rect 2693 278 2759 6238
rect 2851 278 2917 6238
rect 3009 278 3075 6238
rect 3167 278 3233 6238
rect 3325 278 3391 6238
rect 3483 278 3549 6238
rect 3641 278 3707 6238
rect 3799 278 3865 6238
rect 3957 278 4023 6238
rect 4115 278 4181 6238
rect 4273 278 4339 6238
rect 4431 278 4497 6238
rect 4589 278 4655 6238
rect 4747 278 4813 6238
rect 4905 278 4971 6238
rect 30 100 100 236
rect 5040 236 5054 6280
rect 5054 236 5092 6280
rect 5092 236 5110 6280
rect 252 126 4886 226
rect 5040 100 5110 236
<< metal2 >>
rect 30 6420 100 6480
rect 5040 6420 5110 6480
rect 232 6380 252 6390
rect 4886 6380 4906 6390
rect 232 6310 240 6380
rect 4900 6310 4906 6380
rect 232 6290 252 6310
rect 4886 6290 4906 6310
rect 165 6238 231 6258
rect 165 258 231 278
rect 323 6238 389 6258
rect 323 258 389 278
rect 481 6238 547 6258
rect 481 258 547 278
rect 639 6238 705 6258
rect 639 258 705 278
rect 797 6238 863 6258
rect 797 258 863 278
rect 955 6238 1021 6258
rect 955 258 1021 278
rect 1113 6238 1179 6258
rect 1113 258 1179 278
rect 1271 6238 1337 6258
rect 1271 258 1337 278
rect 1429 6238 1495 6258
rect 1429 258 1495 278
rect 1587 6238 1653 6258
rect 1587 258 1653 278
rect 1745 6238 1811 6258
rect 1745 258 1811 278
rect 1903 6238 1969 6258
rect 1903 258 1969 278
rect 2061 6238 2127 6258
rect 2061 258 2127 278
rect 2219 6238 2285 6258
rect 2219 258 2285 278
rect 2377 6238 2443 6258
rect 2377 258 2443 278
rect 2535 6238 2601 6258
rect 2535 258 2601 278
rect 2693 6238 2759 6258
rect 2693 258 2759 278
rect 2851 6238 2917 6258
rect 2851 258 2917 278
rect 3009 6238 3075 6258
rect 3009 258 3075 278
rect 3167 6238 3233 6258
rect 3167 258 3233 278
rect 3325 6238 3391 6258
rect 3325 258 3391 278
rect 3483 6238 3549 6258
rect 3483 258 3549 278
rect 3641 6238 3707 6258
rect 3641 258 3707 278
rect 3799 6238 3865 6258
rect 3799 258 3865 278
rect 3957 6238 4023 6258
rect 3957 258 4023 278
rect 4115 6238 4181 6258
rect 4115 258 4181 278
rect 4273 6238 4339 6258
rect 4273 258 4339 278
rect 4431 6238 4497 6258
rect 4431 258 4497 278
rect 4589 6238 4655 6258
rect 4589 258 4655 278
rect 4747 6238 4813 6258
rect 4747 258 4813 278
rect 4905 6238 4971 6258
rect 4905 258 4971 278
rect 232 210 252 226
rect 4886 210 4906 226
rect 232 140 240 210
rect 4890 140 4906 210
rect 232 126 252 140
rect 4886 126 4906 140
rect 30 30 100 100
rect 5040 30 5110 100
<< via2 >>
rect 240 6310 252 6380
rect 252 6310 4886 6380
rect 4886 6310 4900 6380
rect 165 885 231 2645
rect 323 3885 389 5645
rect 481 885 547 2645
rect 639 3885 705 5645
rect 797 885 863 2645
rect 955 3885 1021 5645
rect 1113 885 1179 2645
rect 1271 3885 1337 5645
rect 1429 885 1495 2645
rect 1587 3885 1653 5645
rect 1745 885 1811 2645
rect 1903 3885 1969 5645
rect 2061 885 2127 2645
rect 2219 3885 2285 5645
rect 2377 885 2443 2645
rect 2535 3885 2601 5645
rect 2693 885 2759 2645
rect 2851 3885 2917 5645
rect 3009 885 3075 2645
rect 3167 3885 3233 5645
rect 3325 885 3391 2645
rect 3483 3885 3549 5645
rect 3641 885 3707 2645
rect 3799 3885 3865 5645
rect 3957 885 4023 2645
rect 4115 3885 4181 5645
rect 4273 885 4339 2645
rect 4431 3885 4497 5645
rect 4589 885 4655 2645
rect 4747 3885 4813 5645
rect 4905 885 4971 2645
rect 240 140 252 210
rect 252 140 4886 210
rect 4886 140 4890 210
<< metal3 >>
rect 100 6380 5100 6500
rect 100 6310 240 6380
rect 4900 6310 5100 6380
rect 100 6300 5100 6310
rect 30 5645 5110 5800
rect 30 3885 323 5645
rect 389 3885 639 5645
rect 705 3885 955 5645
rect 1021 3885 1271 5645
rect 1337 3885 1587 5645
rect 1653 3885 1903 5645
rect 1969 3885 2219 5645
rect 2285 3885 2535 5645
rect 2601 3885 2851 5645
rect 2917 3885 3167 5645
rect 3233 3885 3483 5645
rect 3549 3885 3799 5645
rect 3865 3885 4115 5645
rect 4181 3885 4431 5645
rect 4497 3885 4747 5645
rect 4813 3885 5110 5645
rect 30 3800 5110 3885
rect 30 2645 5110 2800
rect 30 885 165 2645
rect 231 885 481 2645
rect 547 885 797 2645
rect 863 885 1113 2645
rect 1179 885 1429 2645
rect 1495 885 1745 2645
rect 1811 885 2061 2645
rect 2127 885 2377 2645
rect 2443 885 2693 2645
rect 2759 885 3009 2645
rect 3075 885 3325 2645
rect 3391 885 3641 2645
rect 3707 885 3957 2645
rect 4023 885 4273 2645
rect 4339 885 4589 2645
rect 4655 885 4905 2645
rect 4971 885 5110 2645
rect 30 800 5110 885
rect 100 210 5100 230
rect 100 140 240 210
rect 4890 140 5100 210
rect 100 30 5100 140
use sky130_fd_pr__nfet_g5v0d10v5_UDPNFN  sky130_fd_pr__nfet_g5v0d10v5_UDPNFN_0
timestamp 1663719933
transform 1 0 2569 0 1 3258
box -2569 -3258 2569 3258
<< labels >>
rlabel metal2 30 6420 100 6480 1 SUB
rlabel metal3 140 6300 200 6500 1 G
rlabel metal3 220 3810 260 5770 1 SD1
rlabel metal3 190 810 230 2770 1 SD2
<< end >>
