magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< nwell >>
rect -54 -54 312 306
<< scpmos >>
rect 60 0 90 252
rect 168 0 198 252
<< pdiff >>
rect 0 0 60 252
rect 90 0 168 252
rect 198 0 258 252
<< poly >>
rect 60 252 90 278
rect 168 252 198 278
rect 60 -26 90 0
rect 168 -26 198 0
rect 60 -56 198 -26
<< locali >>
rect 8 93 42 159
rect 112 93 146 159
rect 216 93 250 159
use sky130_sram_1r1w_24x128_8_contact_11  sky130_sram_1r1w_24x128_8_contact_11_0
timestamp 1661296025
transform 1 0 208 0 1 93
box -59 -51 109 117
use sky130_sram_1r1w_24x128_8_contact_11  sky130_sram_1r1w_24x128_8_contact_11_1
timestamp 1661296025
transform 1 0 104 0 1 93
box -59 -51 109 117
use sky130_sram_1r1w_24x128_8_contact_11  sky130_sram_1r1w_24x128_8_contact_11_2
timestamp 1661296025
transform 1 0 0 0 1 93
box -59 -51 109 117
<< labels >>
rlabel poly s 129 -41 129 -41 4 G
port 1 nsew
rlabel locali s 233 126 233 126 4 S
port 2 nsew
rlabel locali s 25 126 25 126 4 S
port 2 nsew
rlabel locali s 129 126 129 126 4 D
port 3 nsew
<< properties >>
string FIXED_BBOX -54 -56 312 306
<< end >>
