magic
tech sky130B
magscale 1 2
timestamp 1662238829
<< nwell >>
rect -4811 -1184 4811 1184
<< pmos >>
rect -4615 -964 -4415 1036
rect -4357 -964 -4157 1036
rect -4099 -964 -3899 1036
rect -3841 -964 -3641 1036
rect -3583 -964 -3383 1036
rect -3325 -964 -3125 1036
rect -3067 -964 -2867 1036
rect -2809 -964 -2609 1036
rect -2551 -964 -2351 1036
rect -2293 -964 -2093 1036
rect -2035 -964 -1835 1036
rect -1777 -964 -1577 1036
rect -1519 -964 -1319 1036
rect -1261 -964 -1061 1036
rect -1003 -964 -803 1036
rect -745 -964 -545 1036
rect -487 -964 -287 1036
rect -229 -964 -29 1036
rect 29 -964 229 1036
rect 287 -964 487 1036
rect 545 -964 745 1036
rect 803 -964 1003 1036
rect 1061 -964 1261 1036
rect 1319 -964 1519 1036
rect 1577 -964 1777 1036
rect 1835 -964 2035 1036
rect 2093 -964 2293 1036
rect 2351 -964 2551 1036
rect 2609 -964 2809 1036
rect 2867 -964 3067 1036
rect 3125 -964 3325 1036
rect 3383 -964 3583 1036
rect 3641 -964 3841 1036
rect 3899 -964 4099 1036
rect 4157 -964 4357 1036
rect 4415 -964 4615 1036
<< pdiff >>
rect -4673 1024 -4615 1036
rect -4673 -952 -4661 1024
rect -4627 -952 -4615 1024
rect -4673 -964 -4615 -952
rect -4415 1024 -4357 1036
rect -4415 -952 -4403 1024
rect -4369 -952 -4357 1024
rect -4415 -964 -4357 -952
rect -4157 1024 -4099 1036
rect -4157 -952 -4145 1024
rect -4111 -952 -4099 1024
rect -4157 -964 -4099 -952
rect -3899 1024 -3841 1036
rect -3899 -952 -3887 1024
rect -3853 -952 -3841 1024
rect -3899 -964 -3841 -952
rect -3641 1024 -3583 1036
rect -3641 -952 -3629 1024
rect -3595 -952 -3583 1024
rect -3641 -964 -3583 -952
rect -3383 1024 -3325 1036
rect -3383 -952 -3371 1024
rect -3337 -952 -3325 1024
rect -3383 -964 -3325 -952
rect -3125 1024 -3067 1036
rect -3125 -952 -3113 1024
rect -3079 -952 -3067 1024
rect -3125 -964 -3067 -952
rect -2867 1024 -2809 1036
rect -2867 -952 -2855 1024
rect -2821 -952 -2809 1024
rect -2867 -964 -2809 -952
rect -2609 1024 -2551 1036
rect -2609 -952 -2597 1024
rect -2563 -952 -2551 1024
rect -2609 -964 -2551 -952
rect -2351 1024 -2293 1036
rect -2351 -952 -2339 1024
rect -2305 -952 -2293 1024
rect -2351 -964 -2293 -952
rect -2093 1024 -2035 1036
rect -2093 -952 -2081 1024
rect -2047 -952 -2035 1024
rect -2093 -964 -2035 -952
rect -1835 1024 -1777 1036
rect -1835 -952 -1823 1024
rect -1789 -952 -1777 1024
rect -1835 -964 -1777 -952
rect -1577 1024 -1519 1036
rect -1577 -952 -1565 1024
rect -1531 -952 -1519 1024
rect -1577 -964 -1519 -952
rect -1319 1024 -1261 1036
rect -1319 -952 -1307 1024
rect -1273 -952 -1261 1024
rect -1319 -964 -1261 -952
rect -1061 1024 -1003 1036
rect -1061 -952 -1049 1024
rect -1015 -952 -1003 1024
rect -1061 -964 -1003 -952
rect -803 1024 -745 1036
rect -803 -952 -791 1024
rect -757 -952 -745 1024
rect -803 -964 -745 -952
rect -545 1024 -487 1036
rect -545 -952 -533 1024
rect -499 -952 -487 1024
rect -545 -964 -487 -952
rect -287 1024 -229 1036
rect -287 -952 -275 1024
rect -241 -952 -229 1024
rect -287 -964 -229 -952
rect -29 1024 29 1036
rect -29 -952 -17 1024
rect 17 -952 29 1024
rect -29 -964 29 -952
rect 229 1024 287 1036
rect 229 -952 241 1024
rect 275 -952 287 1024
rect 229 -964 287 -952
rect 487 1024 545 1036
rect 487 -952 499 1024
rect 533 -952 545 1024
rect 487 -964 545 -952
rect 745 1024 803 1036
rect 745 -952 757 1024
rect 791 -952 803 1024
rect 745 -964 803 -952
rect 1003 1024 1061 1036
rect 1003 -952 1015 1024
rect 1049 -952 1061 1024
rect 1003 -964 1061 -952
rect 1261 1024 1319 1036
rect 1261 -952 1273 1024
rect 1307 -952 1319 1024
rect 1261 -964 1319 -952
rect 1519 1024 1577 1036
rect 1519 -952 1531 1024
rect 1565 -952 1577 1024
rect 1519 -964 1577 -952
rect 1777 1024 1835 1036
rect 1777 -952 1789 1024
rect 1823 -952 1835 1024
rect 1777 -964 1835 -952
rect 2035 1024 2093 1036
rect 2035 -952 2047 1024
rect 2081 -952 2093 1024
rect 2035 -964 2093 -952
rect 2293 1024 2351 1036
rect 2293 -952 2305 1024
rect 2339 -952 2351 1024
rect 2293 -964 2351 -952
rect 2551 1024 2609 1036
rect 2551 -952 2563 1024
rect 2597 -952 2609 1024
rect 2551 -964 2609 -952
rect 2809 1024 2867 1036
rect 2809 -952 2821 1024
rect 2855 -952 2867 1024
rect 2809 -964 2867 -952
rect 3067 1024 3125 1036
rect 3067 -952 3079 1024
rect 3113 -952 3125 1024
rect 3067 -964 3125 -952
rect 3325 1024 3383 1036
rect 3325 -952 3337 1024
rect 3371 -952 3383 1024
rect 3325 -964 3383 -952
rect 3583 1024 3641 1036
rect 3583 -952 3595 1024
rect 3629 -952 3641 1024
rect 3583 -964 3641 -952
rect 3841 1024 3899 1036
rect 3841 -952 3853 1024
rect 3887 -952 3899 1024
rect 3841 -964 3899 -952
rect 4099 1024 4157 1036
rect 4099 -952 4111 1024
rect 4145 -952 4157 1024
rect 4099 -964 4157 -952
rect 4357 1024 4415 1036
rect 4357 -952 4369 1024
rect 4403 -952 4415 1024
rect 4357 -964 4415 -952
rect 4615 1024 4673 1036
rect 4615 -952 4627 1024
rect 4661 -952 4673 1024
rect 4615 -964 4673 -952
<< pdiffc >>
rect -4661 -952 -4627 1024
rect -4403 -952 -4369 1024
rect -4145 -952 -4111 1024
rect -3887 -952 -3853 1024
rect -3629 -952 -3595 1024
rect -3371 -952 -3337 1024
rect -3113 -952 -3079 1024
rect -2855 -952 -2821 1024
rect -2597 -952 -2563 1024
rect -2339 -952 -2305 1024
rect -2081 -952 -2047 1024
rect -1823 -952 -1789 1024
rect -1565 -952 -1531 1024
rect -1307 -952 -1273 1024
rect -1049 -952 -1015 1024
rect -791 -952 -757 1024
rect -533 -952 -499 1024
rect -275 -952 -241 1024
rect -17 -952 17 1024
rect 241 -952 275 1024
rect 499 -952 533 1024
rect 757 -952 791 1024
rect 1015 -952 1049 1024
rect 1273 -952 1307 1024
rect 1531 -952 1565 1024
rect 1789 -952 1823 1024
rect 2047 -952 2081 1024
rect 2305 -952 2339 1024
rect 2563 -952 2597 1024
rect 2821 -952 2855 1024
rect 3079 -952 3113 1024
rect 3337 -952 3371 1024
rect 3595 -952 3629 1024
rect 3853 -952 3887 1024
rect 4111 -952 4145 1024
rect 4369 -952 4403 1024
rect 4627 -952 4661 1024
<< nsubdiff >>
rect -4775 1114 -4679 1148
rect 4679 1114 4775 1148
rect -4775 1051 -4741 1114
rect 4741 1051 4775 1114
rect -4775 -1114 -4741 -1051
rect 4741 -1114 4775 -1051
rect -4775 -1148 -4679 -1114
rect 4679 -1148 4775 -1114
<< nsubdiffcont >>
rect -4679 1114 4679 1148
rect -4775 -1051 -4741 1051
rect 4741 -1051 4775 1051
rect -4679 -1148 4679 -1114
<< poly >>
rect -4615 1036 -4415 1062
rect -4357 1036 -4157 1062
rect -4099 1036 -3899 1062
rect -3841 1036 -3641 1062
rect -3583 1036 -3383 1062
rect -3325 1036 -3125 1062
rect -3067 1036 -2867 1062
rect -2809 1036 -2609 1062
rect -2551 1036 -2351 1062
rect -2293 1036 -2093 1062
rect -2035 1036 -1835 1062
rect -1777 1036 -1577 1062
rect -1519 1036 -1319 1062
rect -1261 1036 -1061 1062
rect -1003 1036 -803 1062
rect -745 1036 -545 1062
rect -487 1036 -287 1062
rect -229 1036 -29 1062
rect 29 1036 229 1062
rect 287 1036 487 1062
rect 545 1036 745 1062
rect 803 1036 1003 1062
rect 1061 1036 1261 1062
rect 1319 1036 1519 1062
rect 1577 1036 1777 1062
rect 1835 1036 2035 1062
rect 2093 1036 2293 1062
rect 2351 1036 2551 1062
rect 2609 1036 2809 1062
rect 2867 1036 3067 1062
rect 3125 1036 3325 1062
rect 3383 1036 3583 1062
rect 3641 1036 3841 1062
rect 3899 1036 4099 1062
rect 4157 1036 4357 1062
rect 4415 1036 4615 1062
rect -4615 -1011 -4415 -964
rect -4615 -1045 -4599 -1011
rect -4431 -1045 -4415 -1011
rect -4615 -1061 -4415 -1045
rect -4357 -1011 -4157 -964
rect -4357 -1045 -4341 -1011
rect -4173 -1045 -4157 -1011
rect -4357 -1061 -4157 -1045
rect -4099 -1011 -3899 -964
rect -4099 -1045 -4083 -1011
rect -3915 -1045 -3899 -1011
rect -4099 -1061 -3899 -1045
rect -3841 -1011 -3641 -964
rect -3841 -1045 -3825 -1011
rect -3657 -1045 -3641 -1011
rect -3841 -1061 -3641 -1045
rect -3583 -1011 -3383 -964
rect -3583 -1045 -3567 -1011
rect -3399 -1045 -3383 -1011
rect -3583 -1061 -3383 -1045
rect -3325 -1011 -3125 -964
rect -3325 -1045 -3309 -1011
rect -3141 -1045 -3125 -1011
rect -3325 -1061 -3125 -1045
rect -3067 -1011 -2867 -964
rect -3067 -1045 -3051 -1011
rect -2883 -1045 -2867 -1011
rect -3067 -1061 -2867 -1045
rect -2809 -1011 -2609 -964
rect -2809 -1045 -2793 -1011
rect -2625 -1045 -2609 -1011
rect -2809 -1061 -2609 -1045
rect -2551 -1011 -2351 -964
rect -2551 -1045 -2535 -1011
rect -2367 -1045 -2351 -1011
rect -2551 -1061 -2351 -1045
rect -2293 -1011 -2093 -964
rect -2293 -1045 -2277 -1011
rect -2109 -1045 -2093 -1011
rect -2293 -1061 -2093 -1045
rect -2035 -1011 -1835 -964
rect -2035 -1045 -2019 -1011
rect -1851 -1045 -1835 -1011
rect -2035 -1061 -1835 -1045
rect -1777 -1011 -1577 -964
rect -1777 -1045 -1761 -1011
rect -1593 -1045 -1577 -1011
rect -1777 -1061 -1577 -1045
rect -1519 -1011 -1319 -964
rect -1519 -1045 -1503 -1011
rect -1335 -1045 -1319 -1011
rect -1519 -1061 -1319 -1045
rect -1261 -1011 -1061 -964
rect -1261 -1045 -1245 -1011
rect -1077 -1045 -1061 -1011
rect -1261 -1061 -1061 -1045
rect -1003 -1011 -803 -964
rect -1003 -1045 -987 -1011
rect -819 -1045 -803 -1011
rect -1003 -1061 -803 -1045
rect -745 -1011 -545 -964
rect -745 -1045 -729 -1011
rect -561 -1045 -545 -1011
rect -745 -1061 -545 -1045
rect -487 -1011 -287 -964
rect -487 -1045 -471 -1011
rect -303 -1045 -287 -1011
rect -487 -1061 -287 -1045
rect -229 -1011 -29 -964
rect -229 -1045 -213 -1011
rect -45 -1045 -29 -1011
rect -229 -1061 -29 -1045
rect 29 -1011 229 -964
rect 29 -1045 45 -1011
rect 213 -1045 229 -1011
rect 29 -1061 229 -1045
rect 287 -1011 487 -964
rect 287 -1045 303 -1011
rect 471 -1045 487 -1011
rect 287 -1061 487 -1045
rect 545 -1011 745 -964
rect 545 -1045 561 -1011
rect 729 -1045 745 -1011
rect 545 -1061 745 -1045
rect 803 -1011 1003 -964
rect 803 -1045 819 -1011
rect 987 -1045 1003 -1011
rect 803 -1061 1003 -1045
rect 1061 -1011 1261 -964
rect 1061 -1045 1077 -1011
rect 1245 -1045 1261 -1011
rect 1061 -1061 1261 -1045
rect 1319 -1011 1519 -964
rect 1319 -1045 1335 -1011
rect 1503 -1045 1519 -1011
rect 1319 -1061 1519 -1045
rect 1577 -1011 1777 -964
rect 1577 -1045 1593 -1011
rect 1761 -1045 1777 -1011
rect 1577 -1061 1777 -1045
rect 1835 -1011 2035 -964
rect 1835 -1045 1851 -1011
rect 2019 -1045 2035 -1011
rect 1835 -1061 2035 -1045
rect 2093 -1011 2293 -964
rect 2093 -1045 2109 -1011
rect 2277 -1045 2293 -1011
rect 2093 -1061 2293 -1045
rect 2351 -1011 2551 -964
rect 2351 -1045 2367 -1011
rect 2535 -1045 2551 -1011
rect 2351 -1061 2551 -1045
rect 2609 -1011 2809 -964
rect 2609 -1045 2625 -1011
rect 2793 -1045 2809 -1011
rect 2609 -1061 2809 -1045
rect 2867 -1011 3067 -964
rect 2867 -1045 2883 -1011
rect 3051 -1045 3067 -1011
rect 2867 -1061 3067 -1045
rect 3125 -1011 3325 -964
rect 3125 -1045 3141 -1011
rect 3309 -1045 3325 -1011
rect 3125 -1061 3325 -1045
rect 3383 -1011 3583 -964
rect 3383 -1045 3399 -1011
rect 3567 -1045 3583 -1011
rect 3383 -1061 3583 -1045
rect 3641 -1011 3841 -964
rect 3641 -1045 3657 -1011
rect 3825 -1045 3841 -1011
rect 3641 -1061 3841 -1045
rect 3899 -1011 4099 -964
rect 3899 -1045 3915 -1011
rect 4083 -1045 4099 -1011
rect 3899 -1061 4099 -1045
rect 4157 -1011 4357 -964
rect 4157 -1045 4173 -1011
rect 4341 -1045 4357 -1011
rect 4157 -1061 4357 -1045
rect 4415 -1011 4615 -964
rect 4415 -1045 4431 -1011
rect 4599 -1045 4615 -1011
rect 4415 -1061 4615 -1045
<< polycont >>
rect -4599 -1045 -4431 -1011
rect -4341 -1045 -4173 -1011
rect -4083 -1045 -3915 -1011
rect -3825 -1045 -3657 -1011
rect -3567 -1045 -3399 -1011
rect -3309 -1045 -3141 -1011
rect -3051 -1045 -2883 -1011
rect -2793 -1045 -2625 -1011
rect -2535 -1045 -2367 -1011
rect -2277 -1045 -2109 -1011
rect -2019 -1045 -1851 -1011
rect -1761 -1045 -1593 -1011
rect -1503 -1045 -1335 -1011
rect -1245 -1045 -1077 -1011
rect -987 -1045 -819 -1011
rect -729 -1045 -561 -1011
rect -471 -1045 -303 -1011
rect -213 -1045 -45 -1011
rect 45 -1045 213 -1011
rect 303 -1045 471 -1011
rect 561 -1045 729 -1011
rect 819 -1045 987 -1011
rect 1077 -1045 1245 -1011
rect 1335 -1045 1503 -1011
rect 1593 -1045 1761 -1011
rect 1851 -1045 2019 -1011
rect 2109 -1045 2277 -1011
rect 2367 -1045 2535 -1011
rect 2625 -1045 2793 -1011
rect 2883 -1045 3051 -1011
rect 3141 -1045 3309 -1011
rect 3399 -1045 3567 -1011
rect 3657 -1045 3825 -1011
rect 3915 -1045 4083 -1011
rect 4173 -1045 4341 -1011
rect 4431 -1045 4599 -1011
<< locali >>
rect -4775 1114 -4679 1148
rect 4679 1114 4775 1148
rect -4775 1051 -4741 1114
rect 4741 1051 4775 1114
rect -4661 1024 -4627 1040
rect -4661 -968 -4627 -952
rect -4403 1024 -4369 1040
rect -4403 -968 -4369 -952
rect -4145 1024 -4111 1040
rect -4145 -968 -4111 -952
rect -3887 1024 -3853 1040
rect -3887 -968 -3853 -952
rect -3629 1024 -3595 1040
rect -3629 -968 -3595 -952
rect -3371 1024 -3337 1040
rect -3371 -968 -3337 -952
rect -3113 1024 -3079 1040
rect -3113 -968 -3079 -952
rect -2855 1024 -2821 1040
rect -2855 -968 -2821 -952
rect -2597 1024 -2563 1040
rect -2597 -968 -2563 -952
rect -2339 1024 -2305 1040
rect -2339 -968 -2305 -952
rect -2081 1024 -2047 1040
rect -2081 -968 -2047 -952
rect -1823 1024 -1789 1040
rect -1823 -968 -1789 -952
rect -1565 1024 -1531 1040
rect -1565 -968 -1531 -952
rect -1307 1024 -1273 1040
rect -1307 -968 -1273 -952
rect -1049 1024 -1015 1040
rect -1049 -968 -1015 -952
rect -791 1024 -757 1040
rect -791 -968 -757 -952
rect -533 1024 -499 1040
rect -533 -968 -499 -952
rect -275 1024 -241 1040
rect -275 -968 -241 -952
rect -17 1024 17 1040
rect -17 -968 17 -952
rect 241 1024 275 1040
rect 241 -968 275 -952
rect 499 1024 533 1040
rect 499 -968 533 -952
rect 757 1024 791 1040
rect 757 -968 791 -952
rect 1015 1024 1049 1040
rect 1015 -968 1049 -952
rect 1273 1024 1307 1040
rect 1273 -968 1307 -952
rect 1531 1024 1565 1040
rect 1531 -968 1565 -952
rect 1789 1024 1823 1040
rect 1789 -968 1823 -952
rect 2047 1024 2081 1040
rect 2047 -968 2081 -952
rect 2305 1024 2339 1040
rect 2305 -968 2339 -952
rect 2563 1024 2597 1040
rect 2563 -968 2597 -952
rect 2821 1024 2855 1040
rect 2821 -968 2855 -952
rect 3079 1024 3113 1040
rect 3079 -968 3113 -952
rect 3337 1024 3371 1040
rect 3337 -968 3371 -952
rect 3595 1024 3629 1040
rect 3595 -968 3629 -952
rect 3853 1024 3887 1040
rect 3853 -968 3887 -952
rect 4111 1024 4145 1040
rect 4111 -968 4145 -952
rect 4369 1024 4403 1040
rect 4369 -968 4403 -952
rect 4627 1024 4661 1040
rect 4627 -968 4661 -952
rect -4615 -1045 -4599 -1011
rect -4431 -1045 -4415 -1011
rect -4357 -1045 -4341 -1011
rect -4173 -1045 -4157 -1011
rect -4099 -1045 -4083 -1011
rect -3915 -1045 -3899 -1011
rect -3841 -1045 -3825 -1011
rect -3657 -1045 -3641 -1011
rect -3583 -1045 -3567 -1011
rect -3399 -1045 -3383 -1011
rect -3325 -1045 -3309 -1011
rect -3141 -1045 -3125 -1011
rect -3067 -1045 -3051 -1011
rect -2883 -1045 -2867 -1011
rect -2809 -1045 -2793 -1011
rect -2625 -1045 -2609 -1011
rect -2551 -1045 -2535 -1011
rect -2367 -1045 -2351 -1011
rect -2293 -1045 -2277 -1011
rect -2109 -1045 -2093 -1011
rect -2035 -1045 -2019 -1011
rect -1851 -1045 -1835 -1011
rect -1777 -1045 -1761 -1011
rect -1593 -1045 -1577 -1011
rect -1519 -1045 -1503 -1011
rect -1335 -1045 -1319 -1011
rect -1261 -1045 -1245 -1011
rect -1077 -1045 -1061 -1011
rect -1003 -1045 -987 -1011
rect -819 -1045 -803 -1011
rect -745 -1045 -729 -1011
rect -561 -1045 -545 -1011
rect -487 -1045 -471 -1011
rect -303 -1045 -287 -1011
rect -229 -1045 -213 -1011
rect -45 -1045 -29 -1011
rect 29 -1045 45 -1011
rect 213 -1045 229 -1011
rect 287 -1045 303 -1011
rect 471 -1045 487 -1011
rect 545 -1045 561 -1011
rect 729 -1045 745 -1011
rect 803 -1045 819 -1011
rect 987 -1045 1003 -1011
rect 1061 -1045 1077 -1011
rect 1245 -1045 1261 -1011
rect 1319 -1045 1335 -1011
rect 1503 -1045 1519 -1011
rect 1577 -1045 1593 -1011
rect 1761 -1045 1777 -1011
rect 1835 -1045 1851 -1011
rect 2019 -1045 2035 -1011
rect 2093 -1045 2109 -1011
rect 2277 -1045 2293 -1011
rect 2351 -1045 2367 -1011
rect 2535 -1045 2551 -1011
rect 2609 -1045 2625 -1011
rect 2793 -1045 2809 -1011
rect 2867 -1045 2883 -1011
rect 3051 -1045 3067 -1011
rect 3125 -1045 3141 -1011
rect 3309 -1045 3325 -1011
rect 3383 -1045 3399 -1011
rect 3567 -1045 3583 -1011
rect 3641 -1045 3657 -1011
rect 3825 -1045 3841 -1011
rect 3899 -1045 3915 -1011
rect 4083 -1045 4099 -1011
rect 4157 -1045 4173 -1011
rect 4341 -1045 4357 -1011
rect 4415 -1045 4431 -1011
rect 4599 -1045 4615 -1011
rect -4775 -1114 -4741 -1051
rect 4741 -1114 4775 -1051
rect -4775 -1148 -4679 -1114
rect 4679 -1148 4775 -1114
<< viali >>
rect -4661 -952 -4627 1024
rect -4403 -952 -4369 1024
rect -4145 -952 -4111 1024
rect -3887 -952 -3853 1024
rect -3629 -952 -3595 1024
rect -3371 -952 -3337 1024
rect -3113 -952 -3079 1024
rect -2855 -952 -2821 1024
rect -2597 -952 -2563 1024
rect -2339 -952 -2305 1024
rect -2081 -952 -2047 1024
rect -1823 -952 -1789 1024
rect -1565 -952 -1531 1024
rect -1307 -952 -1273 1024
rect -1049 -952 -1015 1024
rect -791 -952 -757 1024
rect -533 -952 -499 1024
rect -275 -952 -241 1024
rect -17 -952 17 1024
rect 241 -952 275 1024
rect 499 -952 533 1024
rect 757 -952 791 1024
rect 1015 -952 1049 1024
rect 1273 -952 1307 1024
rect 1531 -952 1565 1024
rect 1789 -952 1823 1024
rect 2047 -952 2081 1024
rect 2305 -952 2339 1024
rect 2563 -952 2597 1024
rect 2821 -952 2855 1024
rect 3079 -952 3113 1024
rect 3337 -952 3371 1024
rect 3595 -952 3629 1024
rect 3853 -952 3887 1024
rect 4111 -952 4145 1024
rect 4369 -952 4403 1024
rect 4627 -952 4661 1024
rect -4599 -1045 -4431 -1011
rect -4341 -1045 -4173 -1011
rect -4083 -1045 -3915 -1011
rect -3825 -1045 -3657 -1011
rect -3567 -1045 -3399 -1011
rect -3309 -1045 -3141 -1011
rect -3051 -1045 -2883 -1011
rect -2793 -1045 -2625 -1011
rect -2535 -1045 -2367 -1011
rect -2277 -1045 -2109 -1011
rect -2019 -1045 -1851 -1011
rect -1761 -1045 -1593 -1011
rect -1503 -1045 -1335 -1011
rect -1245 -1045 -1077 -1011
rect -987 -1045 -819 -1011
rect -729 -1045 -561 -1011
rect -471 -1045 -303 -1011
rect -213 -1045 -45 -1011
rect 45 -1045 213 -1011
rect 303 -1045 471 -1011
rect 561 -1045 729 -1011
rect 819 -1045 987 -1011
rect 1077 -1045 1245 -1011
rect 1335 -1045 1503 -1011
rect 1593 -1045 1761 -1011
rect 1851 -1045 2019 -1011
rect 2109 -1045 2277 -1011
rect 2367 -1045 2535 -1011
rect 2625 -1045 2793 -1011
rect 2883 -1045 3051 -1011
rect 3141 -1045 3309 -1011
rect 3399 -1045 3567 -1011
rect 3657 -1045 3825 -1011
rect 3915 -1045 4083 -1011
rect 4173 -1045 4341 -1011
rect 4431 -1045 4599 -1011
<< metal1 >>
rect -4667 1024 -4621 1036
rect -4667 -952 -4661 1024
rect -4627 -952 -4621 1024
rect -4667 -964 -4621 -952
rect -4409 1024 -4363 1036
rect -4409 -952 -4403 1024
rect -4369 -952 -4363 1024
rect -4409 -964 -4363 -952
rect -4151 1024 -4105 1036
rect -4151 -952 -4145 1024
rect -4111 -952 -4105 1024
rect -4151 -964 -4105 -952
rect -3893 1024 -3847 1036
rect -3893 -952 -3887 1024
rect -3853 -952 -3847 1024
rect -3893 -964 -3847 -952
rect -3635 1024 -3589 1036
rect -3635 -952 -3629 1024
rect -3595 -952 -3589 1024
rect -3635 -964 -3589 -952
rect -3377 1024 -3331 1036
rect -3377 -952 -3371 1024
rect -3337 -952 -3331 1024
rect -3377 -964 -3331 -952
rect -3119 1024 -3073 1036
rect -3119 -952 -3113 1024
rect -3079 -952 -3073 1024
rect -3119 -964 -3073 -952
rect -2861 1024 -2815 1036
rect -2861 -952 -2855 1024
rect -2821 -952 -2815 1024
rect -2861 -964 -2815 -952
rect -2603 1024 -2557 1036
rect -2603 -952 -2597 1024
rect -2563 -952 -2557 1024
rect -2603 -964 -2557 -952
rect -2345 1024 -2299 1036
rect -2345 -952 -2339 1024
rect -2305 -952 -2299 1024
rect -2345 -964 -2299 -952
rect -2087 1024 -2041 1036
rect -2087 -952 -2081 1024
rect -2047 -952 -2041 1024
rect -2087 -964 -2041 -952
rect -1829 1024 -1783 1036
rect -1829 -952 -1823 1024
rect -1789 -952 -1783 1024
rect -1829 -964 -1783 -952
rect -1571 1024 -1525 1036
rect -1571 -952 -1565 1024
rect -1531 -952 -1525 1024
rect -1571 -964 -1525 -952
rect -1313 1024 -1267 1036
rect -1313 -952 -1307 1024
rect -1273 -952 -1267 1024
rect -1313 -964 -1267 -952
rect -1055 1024 -1009 1036
rect -1055 -952 -1049 1024
rect -1015 -952 -1009 1024
rect -1055 -964 -1009 -952
rect -797 1024 -751 1036
rect -797 -952 -791 1024
rect -757 -952 -751 1024
rect -797 -964 -751 -952
rect -539 1024 -493 1036
rect -539 -952 -533 1024
rect -499 -952 -493 1024
rect -539 -964 -493 -952
rect -281 1024 -235 1036
rect -281 -952 -275 1024
rect -241 -952 -235 1024
rect -281 -964 -235 -952
rect -23 1024 23 1036
rect -23 -952 -17 1024
rect 17 -952 23 1024
rect -23 -964 23 -952
rect 235 1024 281 1036
rect 235 -952 241 1024
rect 275 -952 281 1024
rect 235 -964 281 -952
rect 493 1024 539 1036
rect 493 -952 499 1024
rect 533 -952 539 1024
rect 493 -964 539 -952
rect 751 1024 797 1036
rect 751 -952 757 1024
rect 791 -952 797 1024
rect 751 -964 797 -952
rect 1009 1024 1055 1036
rect 1009 -952 1015 1024
rect 1049 -952 1055 1024
rect 1009 -964 1055 -952
rect 1267 1024 1313 1036
rect 1267 -952 1273 1024
rect 1307 -952 1313 1024
rect 1267 -964 1313 -952
rect 1525 1024 1571 1036
rect 1525 -952 1531 1024
rect 1565 -952 1571 1024
rect 1525 -964 1571 -952
rect 1783 1024 1829 1036
rect 1783 -952 1789 1024
rect 1823 -952 1829 1024
rect 1783 -964 1829 -952
rect 2041 1024 2087 1036
rect 2041 -952 2047 1024
rect 2081 -952 2087 1024
rect 2041 -964 2087 -952
rect 2299 1024 2345 1036
rect 2299 -952 2305 1024
rect 2339 -952 2345 1024
rect 2299 -964 2345 -952
rect 2557 1024 2603 1036
rect 2557 -952 2563 1024
rect 2597 -952 2603 1024
rect 2557 -964 2603 -952
rect 2815 1024 2861 1036
rect 2815 -952 2821 1024
rect 2855 -952 2861 1024
rect 2815 -964 2861 -952
rect 3073 1024 3119 1036
rect 3073 -952 3079 1024
rect 3113 -952 3119 1024
rect 3073 -964 3119 -952
rect 3331 1024 3377 1036
rect 3331 -952 3337 1024
rect 3371 -952 3377 1024
rect 3331 -964 3377 -952
rect 3589 1024 3635 1036
rect 3589 -952 3595 1024
rect 3629 -952 3635 1024
rect 3589 -964 3635 -952
rect 3847 1024 3893 1036
rect 3847 -952 3853 1024
rect 3887 -952 3893 1024
rect 3847 -964 3893 -952
rect 4105 1024 4151 1036
rect 4105 -952 4111 1024
rect 4145 -952 4151 1024
rect 4105 -964 4151 -952
rect 4363 1024 4409 1036
rect 4363 -952 4369 1024
rect 4403 -952 4409 1024
rect 4363 -964 4409 -952
rect 4621 1024 4667 1036
rect 4621 -952 4627 1024
rect 4661 -952 4667 1024
rect 4621 -964 4667 -952
rect -4611 -1011 -4419 -1005
rect -4611 -1045 -4599 -1011
rect -4431 -1045 -4419 -1011
rect -4611 -1051 -4419 -1045
rect -4353 -1011 -4161 -1005
rect -4353 -1045 -4341 -1011
rect -4173 -1045 -4161 -1011
rect -4353 -1051 -4161 -1045
rect -4095 -1011 -3903 -1005
rect -4095 -1045 -4083 -1011
rect -3915 -1045 -3903 -1011
rect -4095 -1051 -3903 -1045
rect -3837 -1011 -3645 -1005
rect -3837 -1045 -3825 -1011
rect -3657 -1045 -3645 -1011
rect -3837 -1051 -3645 -1045
rect -3579 -1011 -3387 -1005
rect -3579 -1045 -3567 -1011
rect -3399 -1045 -3387 -1011
rect -3579 -1051 -3387 -1045
rect -3321 -1011 -3129 -1005
rect -3321 -1045 -3309 -1011
rect -3141 -1045 -3129 -1011
rect -3321 -1051 -3129 -1045
rect -3063 -1011 -2871 -1005
rect -3063 -1045 -3051 -1011
rect -2883 -1045 -2871 -1011
rect -3063 -1051 -2871 -1045
rect -2805 -1011 -2613 -1005
rect -2805 -1045 -2793 -1011
rect -2625 -1045 -2613 -1011
rect -2805 -1051 -2613 -1045
rect -2547 -1011 -2355 -1005
rect -2547 -1045 -2535 -1011
rect -2367 -1045 -2355 -1011
rect -2547 -1051 -2355 -1045
rect -2289 -1011 -2097 -1005
rect -2289 -1045 -2277 -1011
rect -2109 -1045 -2097 -1011
rect -2289 -1051 -2097 -1045
rect -2031 -1011 -1839 -1005
rect -2031 -1045 -2019 -1011
rect -1851 -1045 -1839 -1011
rect -2031 -1051 -1839 -1045
rect -1773 -1011 -1581 -1005
rect -1773 -1045 -1761 -1011
rect -1593 -1045 -1581 -1011
rect -1773 -1051 -1581 -1045
rect -1515 -1011 -1323 -1005
rect -1515 -1045 -1503 -1011
rect -1335 -1045 -1323 -1011
rect -1515 -1051 -1323 -1045
rect -1257 -1011 -1065 -1005
rect -1257 -1045 -1245 -1011
rect -1077 -1045 -1065 -1011
rect -1257 -1051 -1065 -1045
rect -999 -1011 -807 -1005
rect -999 -1045 -987 -1011
rect -819 -1045 -807 -1011
rect -999 -1051 -807 -1045
rect -741 -1011 -549 -1005
rect -741 -1045 -729 -1011
rect -561 -1045 -549 -1011
rect -741 -1051 -549 -1045
rect -483 -1011 -291 -1005
rect -483 -1045 -471 -1011
rect -303 -1045 -291 -1011
rect -483 -1051 -291 -1045
rect -225 -1011 -33 -1005
rect -225 -1045 -213 -1011
rect -45 -1045 -33 -1011
rect -225 -1051 -33 -1045
rect 33 -1011 225 -1005
rect 33 -1045 45 -1011
rect 213 -1045 225 -1011
rect 33 -1051 225 -1045
rect 291 -1011 483 -1005
rect 291 -1045 303 -1011
rect 471 -1045 483 -1011
rect 291 -1051 483 -1045
rect 549 -1011 741 -1005
rect 549 -1045 561 -1011
rect 729 -1045 741 -1011
rect 549 -1051 741 -1045
rect 807 -1011 999 -1005
rect 807 -1045 819 -1011
rect 987 -1045 999 -1011
rect 807 -1051 999 -1045
rect 1065 -1011 1257 -1005
rect 1065 -1045 1077 -1011
rect 1245 -1045 1257 -1011
rect 1065 -1051 1257 -1045
rect 1323 -1011 1515 -1005
rect 1323 -1045 1335 -1011
rect 1503 -1045 1515 -1011
rect 1323 -1051 1515 -1045
rect 1581 -1011 1773 -1005
rect 1581 -1045 1593 -1011
rect 1761 -1045 1773 -1011
rect 1581 -1051 1773 -1045
rect 1839 -1011 2031 -1005
rect 1839 -1045 1851 -1011
rect 2019 -1045 2031 -1011
rect 1839 -1051 2031 -1045
rect 2097 -1011 2289 -1005
rect 2097 -1045 2109 -1011
rect 2277 -1045 2289 -1011
rect 2097 -1051 2289 -1045
rect 2355 -1011 2547 -1005
rect 2355 -1045 2367 -1011
rect 2535 -1045 2547 -1011
rect 2355 -1051 2547 -1045
rect 2613 -1011 2805 -1005
rect 2613 -1045 2625 -1011
rect 2793 -1045 2805 -1011
rect 2613 -1051 2805 -1045
rect 2871 -1011 3063 -1005
rect 2871 -1045 2883 -1011
rect 3051 -1045 3063 -1011
rect 2871 -1051 3063 -1045
rect 3129 -1011 3321 -1005
rect 3129 -1045 3141 -1011
rect 3309 -1045 3321 -1011
rect 3129 -1051 3321 -1045
rect 3387 -1011 3579 -1005
rect 3387 -1045 3399 -1011
rect 3567 -1045 3579 -1011
rect 3387 -1051 3579 -1045
rect 3645 -1011 3837 -1005
rect 3645 -1045 3657 -1011
rect 3825 -1045 3837 -1011
rect 3645 -1051 3837 -1045
rect 3903 -1011 4095 -1005
rect 3903 -1045 3915 -1011
rect 4083 -1045 4095 -1011
rect 3903 -1051 4095 -1045
rect 4161 -1011 4353 -1005
rect 4161 -1045 4173 -1011
rect 4341 -1045 4353 -1011
rect 4161 -1051 4353 -1045
rect 4419 -1011 4611 -1005
rect 4419 -1045 4431 -1011
rect 4599 -1045 4611 -1011
rect 4419 -1051 4611 -1045
<< properties >>
string FIXED_BBOX -4758 -1131 4758 1131
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 1 m 1 nf 36 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
