magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< nwell >>
rect -36 679 728 1471
<< poly >>
rect 114 703 144 907
rect 81 637 144 703
rect 114 359 144 637
<< locali >>
rect 0 1397 692 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 486 1130 520 1397
rect 590 1297 624 1397
rect 64 637 98 703
rect 274 687 308 1096
rect 274 653 325 687
rect 274 244 308 653
rect 62 17 96 144
rect 274 17 308 144
rect 486 17 520 144
rect 590 17 624 104
rect 0 -17 692 17
use sky130_sram_1r1w_24x128_8_contact_15  sky130_sram_1r1w_24x128_8_contact_15_0
timestamp 1661296025
transform 1 0 48 0 1 637
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_28  sky130_sram_1r1w_24x128_8_contact_28_0
timestamp 1661296025
transform 1 0 582 0 1 1256
box -59 -43 109 125
use sky130_sram_1r1w_24x128_8_contact_29  sky130_sram_1r1w_24x128_8_contact_29_0
timestamp 1661296025
transform 1 0 582 0 1 63
box -26 -26 76 108
use sky130_sram_1r1w_24x128_8_nmos_m4_w1_260_sli_dli_da_p  sky130_sram_1r1w_24x128_8_nmos_m4_w1_260_sli_dli_da_p_0
timestamp 1661296025
transform 1 0 54 0 1 51
box -26 -26 500 308
use sky130_sram_1r1w_24x128_8_pmos_m4_w2_000_sli_dli_da_p  sky130_sram_1r1w_24x128_8_pmos_m4_w2_000_sli_dli_da_p_0
timestamp 1661296025
transform 1 0 54 0 1 963
box -59 -56 533 454
<< labels >>
rlabel locali s 81 670 81 670 4 A
port 1 nsew
rlabel locali s 308 670 308 670 4 Z
port 2 nsew
rlabel locali s 346 0 346 0 4 gnd
port 3 nsew
rlabel locali s 346 1414 346 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 692 1414
<< end >>
