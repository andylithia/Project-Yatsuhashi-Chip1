magic
tech sky130B
magscale 1 2
timestamp 1662238829
<< nwell >>
rect -4811 -1219 4811 1219
<< pmos >>
rect -4615 -1000 -4415 1000
rect -4357 -1000 -4157 1000
rect -4099 -1000 -3899 1000
rect -3841 -1000 -3641 1000
rect -3583 -1000 -3383 1000
rect -3325 -1000 -3125 1000
rect -3067 -1000 -2867 1000
rect -2809 -1000 -2609 1000
rect -2551 -1000 -2351 1000
rect -2293 -1000 -2093 1000
rect -2035 -1000 -1835 1000
rect -1777 -1000 -1577 1000
rect -1519 -1000 -1319 1000
rect -1261 -1000 -1061 1000
rect -1003 -1000 -803 1000
rect -745 -1000 -545 1000
rect -487 -1000 -287 1000
rect -229 -1000 -29 1000
rect 29 -1000 229 1000
rect 287 -1000 487 1000
rect 545 -1000 745 1000
rect 803 -1000 1003 1000
rect 1061 -1000 1261 1000
rect 1319 -1000 1519 1000
rect 1577 -1000 1777 1000
rect 1835 -1000 2035 1000
rect 2093 -1000 2293 1000
rect 2351 -1000 2551 1000
rect 2609 -1000 2809 1000
rect 2867 -1000 3067 1000
rect 3125 -1000 3325 1000
rect 3383 -1000 3583 1000
rect 3641 -1000 3841 1000
rect 3899 -1000 4099 1000
rect 4157 -1000 4357 1000
rect 4415 -1000 4615 1000
<< pdiff >>
rect -4673 988 -4615 1000
rect -4673 -988 -4661 988
rect -4627 -988 -4615 988
rect -4673 -1000 -4615 -988
rect -4415 988 -4357 1000
rect -4415 -988 -4403 988
rect -4369 -988 -4357 988
rect -4415 -1000 -4357 -988
rect -4157 988 -4099 1000
rect -4157 -988 -4145 988
rect -4111 -988 -4099 988
rect -4157 -1000 -4099 -988
rect -3899 988 -3841 1000
rect -3899 -988 -3887 988
rect -3853 -988 -3841 988
rect -3899 -1000 -3841 -988
rect -3641 988 -3583 1000
rect -3641 -988 -3629 988
rect -3595 -988 -3583 988
rect -3641 -1000 -3583 -988
rect -3383 988 -3325 1000
rect -3383 -988 -3371 988
rect -3337 -988 -3325 988
rect -3383 -1000 -3325 -988
rect -3125 988 -3067 1000
rect -3125 -988 -3113 988
rect -3079 -988 -3067 988
rect -3125 -1000 -3067 -988
rect -2867 988 -2809 1000
rect -2867 -988 -2855 988
rect -2821 -988 -2809 988
rect -2867 -1000 -2809 -988
rect -2609 988 -2551 1000
rect -2609 -988 -2597 988
rect -2563 -988 -2551 988
rect -2609 -1000 -2551 -988
rect -2351 988 -2293 1000
rect -2351 -988 -2339 988
rect -2305 -988 -2293 988
rect -2351 -1000 -2293 -988
rect -2093 988 -2035 1000
rect -2093 -988 -2081 988
rect -2047 -988 -2035 988
rect -2093 -1000 -2035 -988
rect -1835 988 -1777 1000
rect -1835 -988 -1823 988
rect -1789 -988 -1777 988
rect -1835 -1000 -1777 -988
rect -1577 988 -1519 1000
rect -1577 -988 -1565 988
rect -1531 -988 -1519 988
rect -1577 -1000 -1519 -988
rect -1319 988 -1261 1000
rect -1319 -988 -1307 988
rect -1273 -988 -1261 988
rect -1319 -1000 -1261 -988
rect -1061 988 -1003 1000
rect -1061 -988 -1049 988
rect -1015 -988 -1003 988
rect -1061 -1000 -1003 -988
rect -803 988 -745 1000
rect -803 -988 -791 988
rect -757 -988 -745 988
rect -803 -1000 -745 -988
rect -545 988 -487 1000
rect -545 -988 -533 988
rect -499 -988 -487 988
rect -545 -1000 -487 -988
rect -287 988 -229 1000
rect -287 -988 -275 988
rect -241 -988 -229 988
rect -287 -1000 -229 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 229 988 287 1000
rect 229 -988 241 988
rect 275 -988 287 988
rect 229 -1000 287 -988
rect 487 988 545 1000
rect 487 -988 499 988
rect 533 -988 545 988
rect 487 -1000 545 -988
rect 745 988 803 1000
rect 745 -988 757 988
rect 791 -988 803 988
rect 745 -1000 803 -988
rect 1003 988 1061 1000
rect 1003 -988 1015 988
rect 1049 -988 1061 988
rect 1003 -1000 1061 -988
rect 1261 988 1319 1000
rect 1261 -988 1273 988
rect 1307 -988 1319 988
rect 1261 -1000 1319 -988
rect 1519 988 1577 1000
rect 1519 -988 1531 988
rect 1565 -988 1577 988
rect 1519 -1000 1577 -988
rect 1777 988 1835 1000
rect 1777 -988 1789 988
rect 1823 -988 1835 988
rect 1777 -1000 1835 -988
rect 2035 988 2093 1000
rect 2035 -988 2047 988
rect 2081 -988 2093 988
rect 2035 -1000 2093 -988
rect 2293 988 2351 1000
rect 2293 -988 2305 988
rect 2339 -988 2351 988
rect 2293 -1000 2351 -988
rect 2551 988 2609 1000
rect 2551 -988 2563 988
rect 2597 -988 2609 988
rect 2551 -1000 2609 -988
rect 2809 988 2867 1000
rect 2809 -988 2821 988
rect 2855 -988 2867 988
rect 2809 -1000 2867 -988
rect 3067 988 3125 1000
rect 3067 -988 3079 988
rect 3113 -988 3125 988
rect 3067 -1000 3125 -988
rect 3325 988 3383 1000
rect 3325 -988 3337 988
rect 3371 -988 3383 988
rect 3325 -1000 3383 -988
rect 3583 988 3641 1000
rect 3583 -988 3595 988
rect 3629 -988 3641 988
rect 3583 -1000 3641 -988
rect 3841 988 3899 1000
rect 3841 -988 3853 988
rect 3887 -988 3899 988
rect 3841 -1000 3899 -988
rect 4099 988 4157 1000
rect 4099 -988 4111 988
rect 4145 -988 4157 988
rect 4099 -1000 4157 -988
rect 4357 988 4415 1000
rect 4357 -988 4369 988
rect 4403 -988 4415 988
rect 4357 -1000 4415 -988
rect 4615 988 4673 1000
rect 4615 -988 4627 988
rect 4661 -988 4673 988
rect 4615 -1000 4673 -988
<< pdiffc >>
rect -4661 -988 -4627 988
rect -4403 -988 -4369 988
rect -4145 -988 -4111 988
rect -3887 -988 -3853 988
rect -3629 -988 -3595 988
rect -3371 -988 -3337 988
rect -3113 -988 -3079 988
rect -2855 -988 -2821 988
rect -2597 -988 -2563 988
rect -2339 -988 -2305 988
rect -2081 -988 -2047 988
rect -1823 -988 -1789 988
rect -1565 -988 -1531 988
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
rect 1531 -988 1565 988
rect 1789 -988 1823 988
rect 2047 -988 2081 988
rect 2305 -988 2339 988
rect 2563 -988 2597 988
rect 2821 -988 2855 988
rect 3079 -988 3113 988
rect 3337 -988 3371 988
rect 3595 -988 3629 988
rect 3853 -988 3887 988
rect 4111 -988 4145 988
rect 4369 -988 4403 988
rect 4627 -988 4661 988
<< nsubdiff >>
rect -4775 1149 -4679 1183
rect 4679 1149 4775 1183
rect -4775 1087 -4741 1149
rect 4741 1087 4775 1149
rect -4775 -1149 -4741 -1087
rect 4741 -1149 4775 -1087
rect -4775 -1183 -4679 -1149
rect 4679 -1183 4775 -1149
<< nsubdiffcont >>
rect -4679 1149 4679 1183
rect -4775 -1087 -4741 1087
rect 4741 -1087 4775 1087
rect -4679 -1183 4679 -1149
<< poly >>
rect -4615 1081 -4415 1097
rect -4615 1047 -4599 1081
rect -4431 1047 -4415 1081
rect -4615 1000 -4415 1047
rect -4357 1081 -4157 1097
rect -4357 1047 -4341 1081
rect -4173 1047 -4157 1081
rect -4357 1000 -4157 1047
rect -4099 1081 -3899 1097
rect -4099 1047 -4083 1081
rect -3915 1047 -3899 1081
rect -4099 1000 -3899 1047
rect -3841 1081 -3641 1097
rect -3841 1047 -3825 1081
rect -3657 1047 -3641 1081
rect -3841 1000 -3641 1047
rect -3583 1081 -3383 1097
rect -3583 1047 -3567 1081
rect -3399 1047 -3383 1081
rect -3583 1000 -3383 1047
rect -3325 1081 -3125 1097
rect -3325 1047 -3309 1081
rect -3141 1047 -3125 1081
rect -3325 1000 -3125 1047
rect -3067 1081 -2867 1097
rect -3067 1047 -3051 1081
rect -2883 1047 -2867 1081
rect -3067 1000 -2867 1047
rect -2809 1081 -2609 1097
rect -2809 1047 -2793 1081
rect -2625 1047 -2609 1081
rect -2809 1000 -2609 1047
rect -2551 1081 -2351 1097
rect -2551 1047 -2535 1081
rect -2367 1047 -2351 1081
rect -2551 1000 -2351 1047
rect -2293 1081 -2093 1097
rect -2293 1047 -2277 1081
rect -2109 1047 -2093 1081
rect -2293 1000 -2093 1047
rect -2035 1081 -1835 1097
rect -2035 1047 -2019 1081
rect -1851 1047 -1835 1081
rect -2035 1000 -1835 1047
rect -1777 1081 -1577 1097
rect -1777 1047 -1761 1081
rect -1593 1047 -1577 1081
rect -1777 1000 -1577 1047
rect -1519 1081 -1319 1097
rect -1519 1047 -1503 1081
rect -1335 1047 -1319 1081
rect -1519 1000 -1319 1047
rect -1261 1081 -1061 1097
rect -1261 1047 -1245 1081
rect -1077 1047 -1061 1081
rect -1261 1000 -1061 1047
rect -1003 1081 -803 1097
rect -1003 1047 -987 1081
rect -819 1047 -803 1081
rect -1003 1000 -803 1047
rect -745 1081 -545 1097
rect -745 1047 -729 1081
rect -561 1047 -545 1081
rect -745 1000 -545 1047
rect -487 1081 -287 1097
rect -487 1047 -471 1081
rect -303 1047 -287 1081
rect -487 1000 -287 1047
rect -229 1081 -29 1097
rect -229 1047 -213 1081
rect -45 1047 -29 1081
rect -229 1000 -29 1047
rect 29 1081 229 1097
rect 29 1047 45 1081
rect 213 1047 229 1081
rect 29 1000 229 1047
rect 287 1081 487 1097
rect 287 1047 303 1081
rect 471 1047 487 1081
rect 287 1000 487 1047
rect 545 1081 745 1097
rect 545 1047 561 1081
rect 729 1047 745 1081
rect 545 1000 745 1047
rect 803 1081 1003 1097
rect 803 1047 819 1081
rect 987 1047 1003 1081
rect 803 1000 1003 1047
rect 1061 1081 1261 1097
rect 1061 1047 1077 1081
rect 1245 1047 1261 1081
rect 1061 1000 1261 1047
rect 1319 1081 1519 1097
rect 1319 1047 1335 1081
rect 1503 1047 1519 1081
rect 1319 1000 1519 1047
rect 1577 1081 1777 1097
rect 1577 1047 1593 1081
rect 1761 1047 1777 1081
rect 1577 1000 1777 1047
rect 1835 1081 2035 1097
rect 1835 1047 1851 1081
rect 2019 1047 2035 1081
rect 1835 1000 2035 1047
rect 2093 1081 2293 1097
rect 2093 1047 2109 1081
rect 2277 1047 2293 1081
rect 2093 1000 2293 1047
rect 2351 1081 2551 1097
rect 2351 1047 2367 1081
rect 2535 1047 2551 1081
rect 2351 1000 2551 1047
rect 2609 1081 2809 1097
rect 2609 1047 2625 1081
rect 2793 1047 2809 1081
rect 2609 1000 2809 1047
rect 2867 1081 3067 1097
rect 2867 1047 2883 1081
rect 3051 1047 3067 1081
rect 2867 1000 3067 1047
rect 3125 1081 3325 1097
rect 3125 1047 3141 1081
rect 3309 1047 3325 1081
rect 3125 1000 3325 1047
rect 3383 1081 3583 1097
rect 3383 1047 3399 1081
rect 3567 1047 3583 1081
rect 3383 1000 3583 1047
rect 3641 1081 3841 1097
rect 3641 1047 3657 1081
rect 3825 1047 3841 1081
rect 3641 1000 3841 1047
rect 3899 1081 4099 1097
rect 3899 1047 3915 1081
rect 4083 1047 4099 1081
rect 3899 1000 4099 1047
rect 4157 1081 4357 1097
rect 4157 1047 4173 1081
rect 4341 1047 4357 1081
rect 4157 1000 4357 1047
rect 4415 1081 4615 1097
rect 4415 1047 4431 1081
rect 4599 1047 4615 1081
rect 4415 1000 4615 1047
rect -4615 -1047 -4415 -1000
rect -4615 -1081 -4599 -1047
rect -4431 -1081 -4415 -1047
rect -4615 -1097 -4415 -1081
rect -4357 -1047 -4157 -1000
rect -4357 -1081 -4341 -1047
rect -4173 -1081 -4157 -1047
rect -4357 -1097 -4157 -1081
rect -4099 -1047 -3899 -1000
rect -4099 -1081 -4083 -1047
rect -3915 -1081 -3899 -1047
rect -4099 -1097 -3899 -1081
rect -3841 -1047 -3641 -1000
rect -3841 -1081 -3825 -1047
rect -3657 -1081 -3641 -1047
rect -3841 -1097 -3641 -1081
rect -3583 -1047 -3383 -1000
rect -3583 -1081 -3567 -1047
rect -3399 -1081 -3383 -1047
rect -3583 -1097 -3383 -1081
rect -3325 -1047 -3125 -1000
rect -3325 -1081 -3309 -1047
rect -3141 -1081 -3125 -1047
rect -3325 -1097 -3125 -1081
rect -3067 -1047 -2867 -1000
rect -3067 -1081 -3051 -1047
rect -2883 -1081 -2867 -1047
rect -3067 -1097 -2867 -1081
rect -2809 -1047 -2609 -1000
rect -2809 -1081 -2793 -1047
rect -2625 -1081 -2609 -1047
rect -2809 -1097 -2609 -1081
rect -2551 -1047 -2351 -1000
rect -2551 -1081 -2535 -1047
rect -2367 -1081 -2351 -1047
rect -2551 -1097 -2351 -1081
rect -2293 -1047 -2093 -1000
rect -2293 -1081 -2277 -1047
rect -2109 -1081 -2093 -1047
rect -2293 -1097 -2093 -1081
rect -2035 -1047 -1835 -1000
rect -2035 -1081 -2019 -1047
rect -1851 -1081 -1835 -1047
rect -2035 -1097 -1835 -1081
rect -1777 -1047 -1577 -1000
rect -1777 -1081 -1761 -1047
rect -1593 -1081 -1577 -1047
rect -1777 -1097 -1577 -1081
rect -1519 -1047 -1319 -1000
rect -1519 -1081 -1503 -1047
rect -1335 -1081 -1319 -1047
rect -1519 -1097 -1319 -1081
rect -1261 -1047 -1061 -1000
rect -1261 -1081 -1245 -1047
rect -1077 -1081 -1061 -1047
rect -1261 -1097 -1061 -1081
rect -1003 -1047 -803 -1000
rect -1003 -1081 -987 -1047
rect -819 -1081 -803 -1047
rect -1003 -1097 -803 -1081
rect -745 -1047 -545 -1000
rect -745 -1081 -729 -1047
rect -561 -1081 -545 -1047
rect -745 -1097 -545 -1081
rect -487 -1047 -287 -1000
rect -487 -1081 -471 -1047
rect -303 -1081 -287 -1047
rect -487 -1097 -287 -1081
rect -229 -1047 -29 -1000
rect -229 -1081 -213 -1047
rect -45 -1081 -29 -1047
rect -229 -1097 -29 -1081
rect 29 -1047 229 -1000
rect 29 -1081 45 -1047
rect 213 -1081 229 -1047
rect 29 -1097 229 -1081
rect 287 -1047 487 -1000
rect 287 -1081 303 -1047
rect 471 -1081 487 -1047
rect 287 -1097 487 -1081
rect 545 -1047 745 -1000
rect 545 -1081 561 -1047
rect 729 -1081 745 -1047
rect 545 -1097 745 -1081
rect 803 -1047 1003 -1000
rect 803 -1081 819 -1047
rect 987 -1081 1003 -1047
rect 803 -1097 1003 -1081
rect 1061 -1047 1261 -1000
rect 1061 -1081 1077 -1047
rect 1245 -1081 1261 -1047
rect 1061 -1097 1261 -1081
rect 1319 -1047 1519 -1000
rect 1319 -1081 1335 -1047
rect 1503 -1081 1519 -1047
rect 1319 -1097 1519 -1081
rect 1577 -1047 1777 -1000
rect 1577 -1081 1593 -1047
rect 1761 -1081 1777 -1047
rect 1577 -1097 1777 -1081
rect 1835 -1047 2035 -1000
rect 1835 -1081 1851 -1047
rect 2019 -1081 2035 -1047
rect 1835 -1097 2035 -1081
rect 2093 -1047 2293 -1000
rect 2093 -1081 2109 -1047
rect 2277 -1081 2293 -1047
rect 2093 -1097 2293 -1081
rect 2351 -1047 2551 -1000
rect 2351 -1081 2367 -1047
rect 2535 -1081 2551 -1047
rect 2351 -1097 2551 -1081
rect 2609 -1047 2809 -1000
rect 2609 -1081 2625 -1047
rect 2793 -1081 2809 -1047
rect 2609 -1097 2809 -1081
rect 2867 -1047 3067 -1000
rect 2867 -1081 2883 -1047
rect 3051 -1081 3067 -1047
rect 2867 -1097 3067 -1081
rect 3125 -1047 3325 -1000
rect 3125 -1081 3141 -1047
rect 3309 -1081 3325 -1047
rect 3125 -1097 3325 -1081
rect 3383 -1047 3583 -1000
rect 3383 -1081 3399 -1047
rect 3567 -1081 3583 -1047
rect 3383 -1097 3583 -1081
rect 3641 -1047 3841 -1000
rect 3641 -1081 3657 -1047
rect 3825 -1081 3841 -1047
rect 3641 -1097 3841 -1081
rect 3899 -1047 4099 -1000
rect 3899 -1081 3915 -1047
rect 4083 -1081 4099 -1047
rect 3899 -1097 4099 -1081
rect 4157 -1047 4357 -1000
rect 4157 -1081 4173 -1047
rect 4341 -1081 4357 -1047
rect 4157 -1097 4357 -1081
rect 4415 -1047 4615 -1000
rect 4415 -1081 4431 -1047
rect 4599 -1081 4615 -1047
rect 4415 -1097 4615 -1081
<< polycont >>
rect -4599 1047 -4431 1081
rect -4341 1047 -4173 1081
rect -4083 1047 -3915 1081
rect -3825 1047 -3657 1081
rect -3567 1047 -3399 1081
rect -3309 1047 -3141 1081
rect -3051 1047 -2883 1081
rect -2793 1047 -2625 1081
rect -2535 1047 -2367 1081
rect -2277 1047 -2109 1081
rect -2019 1047 -1851 1081
rect -1761 1047 -1593 1081
rect -1503 1047 -1335 1081
rect -1245 1047 -1077 1081
rect -987 1047 -819 1081
rect -729 1047 -561 1081
rect -471 1047 -303 1081
rect -213 1047 -45 1081
rect 45 1047 213 1081
rect 303 1047 471 1081
rect 561 1047 729 1081
rect 819 1047 987 1081
rect 1077 1047 1245 1081
rect 1335 1047 1503 1081
rect 1593 1047 1761 1081
rect 1851 1047 2019 1081
rect 2109 1047 2277 1081
rect 2367 1047 2535 1081
rect 2625 1047 2793 1081
rect 2883 1047 3051 1081
rect 3141 1047 3309 1081
rect 3399 1047 3567 1081
rect 3657 1047 3825 1081
rect 3915 1047 4083 1081
rect 4173 1047 4341 1081
rect 4431 1047 4599 1081
rect -4599 -1081 -4431 -1047
rect -4341 -1081 -4173 -1047
rect -4083 -1081 -3915 -1047
rect -3825 -1081 -3657 -1047
rect -3567 -1081 -3399 -1047
rect -3309 -1081 -3141 -1047
rect -3051 -1081 -2883 -1047
rect -2793 -1081 -2625 -1047
rect -2535 -1081 -2367 -1047
rect -2277 -1081 -2109 -1047
rect -2019 -1081 -1851 -1047
rect -1761 -1081 -1593 -1047
rect -1503 -1081 -1335 -1047
rect -1245 -1081 -1077 -1047
rect -987 -1081 -819 -1047
rect -729 -1081 -561 -1047
rect -471 -1081 -303 -1047
rect -213 -1081 -45 -1047
rect 45 -1081 213 -1047
rect 303 -1081 471 -1047
rect 561 -1081 729 -1047
rect 819 -1081 987 -1047
rect 1077 -1081 1245 -1047
rect 1335 -1081 1503 -1047
rect 1593 -1081 1761 -1047
rect 1851 -1081 2019 -1047
rect 2109 -1081 2277 -1047
rect 2367 -1081 2535 -1047
rect 2625 -1081 2793 -1047
rect 2883 -1081 3051 -1047
rect 3141 -1081 3309 -1047
rect 3399 -1081 3567 -1047
rect 3657 -1081 3825 -1047
rect 3915 -1081 4083 -1047
rect 4173 -1081 4341 -1047
rect 4431 -1081 4599 -1047
<< locali >>
rect -4775 1149 -4679 1183
rect 4679 1149 4775 1183
rect -4775 1087 -4741 1149
rect 4741 1087 4775 1149
rect -4615 1047 -4599 1081
rect -4431 1047 -4415 1081
rect -4357 1047 -4341 1081
rect -4173 1047 -4157 1081
rect -4099 1047 -4083 1081
rect -3915 1047 -3899 1081
rect -3841 1047 -3825 1081
rect -3657 1047 -3641 1081
rect -3583 1047 -3567 1081
rect -3399 1047 -3383 1081
rect -3325 1047 -3309 1081
rect -3141 1047 -3125 1081
rect -3067 1047 -3051 1081
rect -2883 1047 -2867 1081
rect -2809 1047 -2793 1081
rect -2625 1047 -2609 1081
rect -2551 1047 -2535 1081
rect -2367 1047 -2351 1081
rect -2293 1047 -2277 1081
rect -2109 1047 -2093 1081
rect -2035 1047 -2019 1081
rect -1851 1047 -1835 1081
rect -1777 1047 -1761 1081
rect -1593 1047 -1577 1081
rect -1519 1047 -1503 1081
rect -1335 1047 -1319 1081
rect -1261 1047 -1245 1081
rect -1077 1047 -1061 1081
rect -1003 1047 -987 1081
rect -819 1047 -803 1081
rect -745 1047 -729 1081
rect -561 1047 -545 1081
rect -487 1047 -471 1081
rect -303 1047 -287 1081
rect -229 1047 -213 1081
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect 213 1047 229 1081
rect 287 1047 303 1081
rect 471 1047 487 1081
rect 545 1047 561 1081
rect 729 1047 745 1081
rect 803 1047 819 1081
rect 987 1047 1003 1081
rect 1061 1047 1077 1081
rect 1245 1047 1261 1081
rect 1319 1047 1335 1081
rect 1503 1047 1519 1081
rect 1577 1047 1593 1081
rect 1761 1047 1777 1081
rect 1835 1047 1851 1081
rect 2019 1047 2035 1081
rect 2093 1047 2109 1081
rect 2277 1047 2293 1081
rect 2351 1047 2367 1081
rect 2535 1047 2551 1081
rect 2609 1047 2625 1081
rect 2793 1047 2809 1081
rect 2867 1047 2883 1081
rect 3051 1047 3067 1081
rect 3125 1047 3141 1081
rect 3309 1047 3325 1081
rect 3383 1047 3399 1081
rect 3567 1047 3583 1081
rect 3641 1047 3657 1081
rect 3825 1047 3841 1081
rect 3899 1047 3915 1081
rect 4083 1047 4099 1081
rect 4157 1047 4173 1081
rect 4341 1047 4357 1081
rect 4415 1047 4431 1081
rect 4599 1047 4615 1081
rect -4661 988 -4627 1004
rect -4661 -1004 -4627 -988
rect -4403 988 -4369 1004
rect -4403 -1004 -4369 -988
rect -4145 988 -4111 1004
rect -4145 -1004 -4111 -988
rect -3887 988 -3853 1004
rect -3887 -1004 -3853 -988
rect -3629 988 -3595 1004
rect -3629 -1004 -3595 -988
rect -3371 988 -3337 1004
rect -3371 -1004 -3337 -988
rect -3113 988 -3079 1004
rect -3113 -1004 -3079 -988
rect -2855 988 -2821 1004
rect -2855 -1004 -2821 -988
rect -2597 988 -2563 1004
rect -2597 -1004 -2563 -988
rect -2339 988 -2305 1004
rect -2339 -1004 -2305 -988
rect -2081 988 -2047 1004
rect -2081 -1004 -2047 -988
rect -1823 988 -1789 1004
rect -1823 -1004 -1789 -988
rect -1565 988 -1531 1004
rect -1565 -1004 -1531 -988
rect -1307 988 -1273 1004
rect -1307 -1004 -1273 -988
rect -1049 988 -1015 1004
rect -1049 -1004 -1015 -988
rect -791 988 -757 1004
rect -791 -1004 -757 -988
rect -533 988 -499 1004
rect -533 -1004 -499 -988
rect -275 988 -241 1004
rect -275 -1004 -241 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 241 988 275 1004
rect 241 -1004 275 -988
rect 499 988 533 1004
rect 499 -1004 533 -988
rect 757 988 791 1004
rect 757 -1004 791 -988
rect 1015 988 1049 1004
rect 1015 -1004 1049 -988
rect 1273 988 1307 1004
rect 1273 -1004 1307 -988
rect 1531 988 1565 1004
rect 1531 -1004 1565 -988
rect 1789 988 1823 1004
rect 1789 -1004 1823 -988
rect 2047 988 2081 1004
rect 2047 -1004 2081 -988
rect 2305 988 2339 1004
rect 2305 -1004 2339 -988
rect 2563 988 2597 1004
rect 2563 -1004 2597 -988
rect 2821 988 2855 1004
rect 2821 -1004 2855 -988
rect 3079 988 3113 1004
rect 3079 -1004 3113 -988
rect 3337 988 3371 1004
rect 3337 -1004 3371 -988
rect 3595 988 3629 1004
rect 3595 -1004 3629 -988
rect 3853 988 3887 1004
rect 3853 -1004 3887 -988
rect 4111 988 4145 1004
rect 4111 -1004 4145 -988
rect 4369 988 4403 1004
rect 4369 -1004 4403 -988
rect 4627 988 4661 1004
rect 4627 -1004 4661 -988
rect -4615 -1081 -4599 -1047
rect -4431 -1081 -4415 -1047
rect -4357 -1081 -4341 -1047
rect -4173 -1081 -4157 -1047
rect -4099 -1081 -4083 -1047
rect -3915 -1081 -3899 -1047
rect -3841 -1081 -3825 -1047
rect -3657 -1081 -3641 -1047
rect -3583 -1081 -3567 -1047
rect -3399 -1081 -3383 -1047
rect -3325 -1081 -3309 -1047
rect -3141 -1081 -3125 -1047
rect -3067 -1081 -3051 -1047
rect -2883 -1081 -2867 -1047
rect -2809 -1081 -2793 -1047
rect -2625 -1081 -2609 -1047
rect -2551 -1081 -2535 -1047
rect -2367 -1081 -2351 -1047
rect -2293 -1081 -2277 -1047
rect -2109 -1081 -2093 -1047
rect -2035 -1081 -2019 -1047
rect -1851 -1081 -1835 -1047
rect -1777 -1081 -1761 -1047
rect -1593 -1081 -1577 -1047
rect -1519 -1081 -1503 -1047
rect -1335 -1081 -1319 -1047
rect -1261 -1081 -1245 -1047
rect -1077 -1081 -1061 -1047
rect -1003 -1081 -987 -1047
rect -819 -1081 -803 -1047
rect -745 -1081 -729 -1047
rect -561 -1081 -545 -1047
rect -487 -1081 -471 -1047
rect -303 -1081 -287 -1047
rect -229 -1081 -213 -1047
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect 213 -1081 229 -1047
rect 287 -1081 303 -1047
rect 471 -1081 487 -1047
rect 545 -1081 561 -1047
rect 729 -1081 745 -1047
rect 803 -1081 819 -1047
rect 987 -1081 1003 -1047
rect 1061 -1081 1077 -1047
rect 1245 -1081 1261 -1047
rect 1319 -1081 1335 -1047
rect 1503 -1081 1519 -1047
rect 1577 -1081 1593 -1047
rect 1761 -1081 1777 -1047
rect 1835 -1081 1851 -1047
rect 2019 -1081 2035 -1047
rect 2093 -1081 2109 -1047
rect 2277 -1081 2293 -1047
rect 2351 -1081 2367 -1047
rect 2535 -1081 2551 -1047
rect 2609 -1081 2625 -1047
rect 2793 -1081 2809 -1047
rect 2867 -1081 2883 -1047
rect 3051 -1081 3067 -1047
rect 3125 -1081 3141 -1047
rect 3309 -1081 3325 -1047
rect 3383 -1081 3399 -1047
rect 3567 -1081 3583 -1047
rect 3641 -1081 3657 -1047
rect 3825 -1081 3841 -1047
rect 3899 -1081 3915 -1047
rect 4083 -1081 4099 -1047
rect 4157 -1081 4173 -1047
rect 4341 -1081 4357 -1047
rect 4415 -1081 4431 -1047
rect 4599 -1081 4615 -1047
rect -4775 -1149 -4741 -1087
rect 4741 -1149 4775 -1087
rect -4775 -1183 -4679 -1149
rect 4679 -1183 4775 -1149
<< viali >>
rect -4599 1047 -4431 1081
rect -4341 1047 -4173 1081
rect -4083 1047 -3915 1081
rect -3825 1047 -3657 1081
rect -3567 1047 -3399 1081
rect -3309 1047 -3141 1081
rect -3051 1047 -2883 1081
rect -2793 1047 -2625 1081
rect -2535 1047 -2367 1081
rect -2277 1047 -2109 1081
rect -2019 1047 -1851 1081
rect -1761 1047 -1593 1081
rect -1503 1047 -1335 1081
rect -1245 1047 -1077 1081
rect -987 1047 -819 1081
rect -729 1047 -561 1081
rect -471 1047 -303 1081
rect -213 1047 -45 1081
rect 45 1047 213 1081
rect 303 1047 471 1081
rect 561 1047 729 1081
rect 819 1047 987 1081
rect 1077 1047 1245 1081
rect 1335 1047 1503 1081
rect 1593 1047 1761 1081
rect 1851 1047 2019 1081
rect 2109 1047 2277 1081
rect 2367 1047 2535 1081
rect 2625 1047 2793 1081
rect 2883 1047 3051 1081
rect 3141 1047 3309 1081
rect 3399 1047 3567 1081
rect 3657 1047 3825 1081
rect 3915 1047 4083 1081
rect 4173 1047 4341 1081
rect 4431 1047 4599 1081
rect -4661 -988 -4627 988
rect -4403 -988 -4369 988
rect -4145 -988 -4111 988
rect -3887 -988 -3853 988
rect -3629 -988 -3595 988
rect -3371 -988 -3337 988
rect -3113 -988 -3079 988
rect -2855 -988 -2821 988
rect -2597 -988 -2563 988
rect -2339 -988 -2305 988
rect -2081 -988 -2047 988
rect -1823 -988 -1789 988
rect -1565 -988 -1531 988
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
rect 1531 -988 1565 988
rect 1789 -988 1823 988
rect 2047 -988 2081 988
rect 2305 -988 2339 988
rect 2563 -988 2597 988
rect 2821 -988 2855 988
rect 3079 -988 3113 988
rect 3337 -988 3371 988
rect 3595 -988 3629 988
rect 3853 -988 3887 988
rect 4111 -988 4145 988
rect 4369 -988 4403 988
rect 4627 -988 4661 988
rect -4599 -1081 -4431 -1047
rect -4341 -1081 -4173 -1047
rect -4083 -1081 -3915 -1047
rect -3825 -1081 -3657 -1047
rect -3567 -1081 -3399 -1047
rect -3309 -1081 -3141 -1047
rect -3051 -1081 -2883 -1047
rect -2793 -1081 -2625 -1047
rect -2535 -1081 -2367 -1047
rect -2277 -1081 -2109 -1047
rect -2019 -1081 -1851 -1047
rect -1761 -1081 -1593 -1047
rect -1503 -1081 -1335 -1047
rect -1245 -1081 -1077 -1047
rect -987 -1081 -819 -1047
rect -729 -1081 -561 -1047
rect -471 -1081 -303 -1047
rect -213 -1081 -45 -1047
rect 45 -1081 213 -1047
rect 303 -1081 471 -1047
rect 561 -1081 729 -1047
rect 819 -1081 987 -1047
rect 1077 -1081 1245 -1047
rect 1335 -1081 1503 -1047
rect 1593 -1081 1761 -1047
rect 1851 -1081 2019 -1047
rect 2109 -1081 2277 -1047
rect 2367 -1081 2535 -1047
rect 2625 -1081 2793 -1047
rect 2883 -1081 3051 -1047
rect 3141 -1081 3309 -1047
rect 3399 -1081 3567 -1047
rect 3657 -1081 3825 -1047
rect 3915 -1081 4083 -1047
rect 4173 -1081 4341 -1047
rect 4431 -1081 4599 -1047
<< metal1 >>
rect -4611 1081 -4419 1087
rect -4611 1047 -4599 1081
rect -4431 1047 -4419 1081
rect -4611 1041 -4419 1047
rect -4353 1081 -4161 1087
rect -4353 1047 -4341 1081
rect -4173 1047 -4161 1081
rect -4353 1041 -4161 1047
rect -4095 1081 -3903 1087
rect -4095 1047 -4083 1081
rect -3915 1047 -3903 1081
rect -4095 1041 -3903 1047
rect -3837 1081 -3645 1087
rect -3837 1047 -3825 1081
rect -3657 1047 -3645 1081
rect -3837 1041 -3645 1047
rect -3579 1081 -3387 1087
rect -3579 1047 -3567 1081
rect -3399 1047 -3387 1081
rect -3579 1041 -3387 1047
rect -3321 1081 -3129 1087
rect -3321 1047 -3309 1081
rect -3141 1047 -3129 1081
rect -3321 1041 -3129 1047
rect -3063 1081 -2871 1087
rect -3063 1047 -3051 1081
rect -2883 1047 -2871 1081
rect -3063 1041 -2871 1047
rect -2805 1081 -2613 1087
rect -2805 1047 -2793 1081
rect -2625 1047 -2613 1081
rect -2805 1041 -2613 1047
rect -2547 1081 -2355 1087
rect -2547 1047 -2535 1081
rect -2367 1047 -2355 1081
rect -2547 1041 -2355 1047
rect -2289 1081 -2097 1087
rect -2289 1047 -2277 1081
rect -2109 1047 -2097 1081
rect -2289 1041 -2097 1047
rect -2031 1081 -1839 1087
rect -2031 1047 -2019 1081
rect -1851 1047 -1839 1081
rect -2031 1041 -1839 1047
rect -1773 1081 -1581 1087
rect -1773 1047 -1761 1081
rect -1593 1047 -1581 1081
rect -1773 1041 -1581 1047
rect -1515 1081 -1323 1087
rect -1515 1047 -1503 1081
rect -1335 1047 -1323 1081
rect -1515 1041 -1323 1047
rect -1257 1081 -1065 1087
rect -1257 1047 -1245 1081
rect -1077 1047 -1065 1081
rect -1257 1041 -1065 1047
rect -999 1081 -807 1087
rect -999 1047 -987 1081
rect -819 1047 -807 1081
rect -999 1041 -807 1047
rect -741 1081 -549 1087
rect -741 1047 -729 1081
rect -561 1047 -549 1081
rect -741 1041 -549 1047
rect -483 1081 -291 1087
rect -483 1047 -471 1081
rect -303 1047 -291 1081
rect -483 1041 -291 1047
rect -225 1081 -33 1087
rect -225 1047 -213 1081
rect -45 1047 -33 1081
rect -225 1041 -33 1047
rect 33 1081 225 1087
rect 33 1047 45 1081
rect 213 1047 225 1081
rect 33 1041 225 1047
rect 291 1081 483 1087
rect 291 1047 303 1081
rect 471 1047 483 1081
rect 291 1041 483 1047
rect 549 1081 741 1087
rect 549 1047 561 1081
rect 729 1047 741 1081
rect 549 1041 741 1047
rect 807 1081 999 1087
rect 807 1047 819 1081
rect 987 1047 999 1081
rect 807 1041 999 1047
rect 1065 1081 1257 1087
rect 1065 1047 1077 1081
rect 1245 1047 1257 1081
rect 1065 1041 1257 1047
rect 1323 1081 1515 1087
rect 1323 1047 1335 1081
rect 1503 1047 1515 1081
rect 1323 1041 1515 1047
rect 1581 1081 1773 1087
rect 1581 1047 1593 1081
rect 1761 1047 1773 1081
rect 1581 1041 1773 1047
rect 1839 1081 2031 1087
rect 1839 1047 1851 1081
rect 2019 1047 2031 1081
rect 1839 1041 2031 1047
rect 2097 1081 2289 1087
rect 2097 1047 2109 1081
rect 2277 1047 2289 1081
rect 2097 1041 2289 1047
rect 2355 1081 2547 1087
rect 2355 1047 2367 1081
rect 2535 1047 2547 1081
rect 2355 1041 2547 1047
rect 2613 1081 2805 1087
rect 2613 1047 2625 1081
rect 2793 1047 2805 1081
rect 2613 1041 2805 1047
rect 2871 1081 3063 1087
rect 2871 1047 2883 1081
rect 3051 1047 3063 1081
rect 2871 1041 3063 1047
rect 3129 1081 3321 1087
rect 3129 1047 3141 1081
rect 3309 1047 3321 1081
rect 3129 1041 3321 1047
rect 3387 1081 3579 1087
rect 3387 1047 3399 1081
rect 3567 1047 3579 1081
rect 3387 1041 3579 1047
rect 3645 1081 3837 1087
rect 3645 1047 3657 1081
rect 3825 1047 3837 1081
rect 3645 1041 3837 1047
rect 3903 1081 4095 1087
rect 3903 1047 3915 1081
rect 4083 1047 4095 1081
rect 3903 1041 4095 1047
rect 4161 1081 4353 1087
rect 4161 1047 4173 1081
rect 4341 1047 4353 1081
rect 4161 1041 4353 1047
rect 4419 1081 4611 1087
rect 4419 1047 4431 1081
rect 4599 1047 4611 1081
rect 4419 1041 4611 1047
rect -4667 988 -4621 1000
rect -4667 -988 -4661 988
rect -4627 -988 -4621 988
rect -4667 -1000 -4621 -988
rect -4409 988 -4363 1000
rect -4409 -988 -4403 988
rect -4369 -988 -4363 988
rect -4409 -1000 -4363 -988
rect -4151 988 -4105 1000
rect -4151 -988 -4145 988
rect -4111 -988 -4105 988
rect -4151 -1000 -4105 -988
rect -3893 988 -3847 1000
rect -3893 -988 -3887 988
rect -3853 -988 -3847 988
rect -3893 -1000 -3847 -988
rect -3635 988 -3589 1000
rect -3635 -988 -3629 988
rect -3595 -988 -3589 988
rect -3635 -1000 -3589 -988
rect -3377 988 -3331 1000
rect -3377 -988 -3371 988
rect -3337 -988 -3331 988
rect -3377 -1000 -3331 -988
rect -3119 988 -3073 1000
rect -3119 -988 -3113 988
rect -3079 -988 -3073 988
rect -3119 -1000 -3073 -988
rect -2861 988 -2815 1000
rect -2861 -988 -2855 988
rect -2821 -988 -2815 988
rect -2861 -1000 -2815 -988
rect -2603 988 -2557 1000
rect -2603 -988 -2597 988
rect -2563 -988 -2557 988
rect -2603 -1000 -2557 -988
rect -2345 988 -2299 1000
rect -2345 -988 -2339 988
rect -2305 -988 -2299 988
rect -2345 -1000 -2299 -988
rect -2087 988 -2041 1000
rect -2087 -988 -2081 988
rect -2047 -988 -2041 988
rect -2087 -1000 -2041 -988
rect -1829 988 -1783 1000
rect -1829 -988 -1823 988
rect -1789 -988 -1783 988
rect -1829 -1000 -1783 -988
rect -1571 988 -1525 1000
rect -1571 -988 -1565 988
rect -1531 -988 -1525 988
rect -1571 -1000 -1525 -988
rect -1313 988 -1267 1000
rect -1313 -988 -1307 988
rect -1273 -988 -1267 988
rect -1313 -1000 -1267 -988
rect -1055 988 -1009 1000
rect -1055 -988 -1049 988
rect -1015 -988 -1009 988
rect -1055 -1000 -1009 -988
rect -797 988 -751 1000
rect -797 -988 -791 988
rect -757 -988 -751 988
rect -797 -1000 -751 -988
rect -539 988 -493 1000
rect -539 -988 -533 988
rect -499 -988 -493 988
rect -539 -1000 -493 -988
rect -281 988 -235 1000
rect -281 -988 -275 988
rect -241 -988 -235 988
rect -281 -1000 -235 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 235 988 281 1000
rect 235 -988 241 988
rect 275 -988 281 988
rect 235 -1000 281 -988
rect 493 988 539 1000
rect 493 -988 499 988
rect 533 -988 539 988
rect 493 -1000 539 -988
rect 751 988 797 1000
rect 751 -988 757 988
rect 791 -988 797 988
rect 751 -1000 797 -988
rect 1009 988 1055 1000
rect 1009 -988 1015 988
rect 1049 -988 1055 988
rect 1009 -1000 1055 -988
rect 1267 988 1313 1000
rect 1267 -988 1273 988
rect 1307 -988 1313 988
rect 1267 -1000 1313 -988
rect 1525 988 1571 1000
rect 1525 -988 1531 988
rect 1565 -988 1571 988
rect 1525 -1000 1571 -988
rect 1783 988 1829 1000
rect 1783 -988 1789 988
rect 1823 -988 1829 988
rect 1783 -1000 1829 -988
rect 2041 988 2087 1000
rect 2041 -988 2047 988
rect 2081 -988 2087 988
rect 2041 -1000 2087 -988
rect 2299 988 2345 1000
rect 2299 -988 2305 988
rect 2339 -988 2345 988
rect 2299 -1000 2345 -988
rect 2557 988 2603 1000
rect 2557 -988 2563 988
rect 2597 -988 2603 988
rect 2557 -1000 2603 -988
rect 2815 988 2861 1000
rect 2815 -988 2821 988
rect 2855 -988 2861 988
rect 2815 -1000 2861 -988
rect 3073 988 3119 1000
rect 3073 -988 3079 988
rect 3113 -988 3119 988
rect 3073 -1000 3119 -988
rect 3331 988 3377 1000
rect 3331 -988 3337 988
rect 3371 -988 3377 988
rect 3331 -1000 3377 -988
rect 3589 988 3635 1000
rect 3589 -988 3595 988
rect 3629 -988 3635 988
rect 3589 -1000 3635 -988
rect 3847 988 3893 1000
rect 3847 -988 3853 988
rect 3887 -988 3893 988
rect 3847 -1000 3893 -988
rect 4105 988 4151 1000
rect 4105 -988 4111 988
rect 4145 -988 4151 988
rect 4105 -1000 4151 -988
rect 4363 988 4409 1000
rect 4363 -988 4369 988
rect 4403 -988 4409 988
rect 4363 -1000 4409 -988
rect 4621 988 4667 1000
rect 4621 -988 4627 988
rect 4661 -988 4667 988
rect 4621 -1000 4667 -988
rect -4611 -1047 -4419 -1041
rect -4611 -1081 -4599 -1047
rect -4431 -1081 -4419 -1047
rect -4611 -1087 -4419 -1081
rect -4353 -1047 -4161 -1041
rect -4353 -1081 -4341 -1047
rect -4173 -1081 -4161 -1047
rect -4353 -1087 -4161 -1081
rect -4095 -1047 -3903 -1041
rect -4095 -1081 -4083 -1047
rect -3915 -1081 -3903 -1047
rect -4095 -1087 -3903 -1081
rect -3837 -1047 -3645 -1041
rect -3837 -1081 -3825 -1047
rect -3657 -1081 -3645 -1047
rect -3837 -1087 -3645 -1081
rect -3579 -1047 -3387 -1041
rect -3579 -1081 -3567 -1047
rect -3399 -1081 -3387 -1047
rect -3579 -1087 -3387 -1081
rect -3321 -1047 -3129 -1041
rect -3321 -1081 -3309 -1047
rect -3141 -1081 -3129 -1047
rect -3321 -1087 -3129 -1081
rect -3063 -1047 -2871 -1041
rect -3063 -1081 -3051 -1047
rect -2883 -1081 -2871 -1047
rect -3063 -1087 -2871 -1081
rect -2805 -1047 -2613 -1041
rect -2805 -1081 -2793 -1047
rect -2625 -1081 -2613 -1047
rect -2805 -1087 -2613 -1081
rect -2547 -1047 -2355 -1041
rect -2547 -1081 -2535 -1047
rect -2367 -1081 -2355 -1047
rect -2547 -1087 -2355 -1081
rect -2289 -1047 -2097 -1041
rect -2289 -1081 -2277 -1047
rect -2109 -1081 -2097 -1047
rect -2289 -1087 -2097 -1081
rect -2031 -1047 -1839 -1041
rect -2031 -1081 -2019 -1047
rect -1851 -1081 -1839 -1047
rect -2031 -1087 -1839 -1081
rect -1773 -1047 -1581 -1041
rect -1773 -1081 -1761 -1047
rect -1593 -1081 -1581 -1047
rect -1773 -1087 -1581 -1081
rect -1515 -1047 -1323 -1041
rect -1515 -1081 -1503 -1047
rect -1335 -1081 -1323 -1047
rect -1515 -1087 -1323 -1081
rect -1257 -1047 -1065 -1041
rect -1257 -1081 -1245 -1047
rect -1077 -1081 -1065 -1047
rect -1257 -1087 -1065 -1081
rect -999 -1047 -807 -1041
rect -999 -1081 -987 -1047
rect -819 -1081 -807 -1047
rect -999 -1087 -807 -1081
rect -741 -1047 -549 -1041
rect -741 -1081 -729 -1047
rect -561 -1081 -549 -1047
rect -741 -1087 -549 -1081
rect -483 -1047 -291 -1041
rect -483 -1081 -471 -1047
rect -303 -1081 -291 -1047
rect -483 -1087 -291 -1081
rect -225 -1047 -33 -1041
rect -225 -1081 -213 -1047
rect -45 -1081 -33 -1047
rect -225 -1087 -33 -1081
rect 33 -1047 225 -1041
rect 33 -1081 45 -1047
rect 213 -1081 225 -1047
rect 33 -1087 225 -1081
rect 291 -1047 483 -1041
rect 291 -1081 303 -1047
rect 471 -1081 483 -1047
rect 291 -1087 483 -1081
rect 549 -1047 741 -1041
rect 549 -1081 561 -1047
rect 729 -1081 741 -1047
rect 549 -1087 741 -1081
rect 807 -1047 999 -1041
rect 807 -1081 819 -1047
rect 987 -1081 999 -1047
rect 807 -1087 999 -1081
rect 1065 -1047 1257 -1041
rect 1065 -1081 1077 -1047
rect 1245 -1081 1257 -1047
rect 1065 -1087 1257 -1081
rect 1323 -1047 1515 -1041
rect 1323 -1081 1335 -1047
rect 1503 -1081 1515 -1047
rect 1323 -1087 1515 -1081
rect 1581 -1047 1773 -1041
rect 1581 -1081 1593 -1047
rect 1761 -1081 1773 -1047
rect 1581 -1087 1773 -1081
rect 1839 -1047 2031 -1041
rect 1839 -1081 1851 -1047
rect 2019 -1081 2031 -1047
rect 1839 -1087 2031 -1081
rect 2097 -1047 2289 -1041
rect 2097 -1081 2109 -1047
rect 2277 -1081 2289 -1047
rect 2097 -1087 2289 -1081
rect 2355 -1047 2547 -1041
rect 2355 -1081 2367 -1047
rect 2535 -1081 2547 -1047
rect 2355 -1087 2547 -1081
rect 2613 -1047 2805 -1041
rect 2613 -1081 2625 -1047
rect 2793 -1081 2805 -1047
rect 2613 -1087 2805 -1081
rect 2871 -1047 3063 -1041
rect 2871 -1081 2883 -1047
rect 3051 -1081 3063 -1047
rect 2871 -1087 3063 -1081
rect 3129 -1047 3321 -1041
rect 3129 -1081 3141 -1047
rect 3309 -1081 3321 -1047
rect 3129 -1087 3321 -1081
rect 3387 -1047 3579 -1041
rect 3387 -1081 3399 -1047
rect 3567 -1081 3579 -1047
rect 3387 -1087 3579 -1081
rect 3645 -1047 3837 -1041
rect 3645 -1081 3657 -1047
rect 3825 -1081 3837 -1047
rect 3645 -1087 3837 -1081
rect 3903 -1047 4095 -1041
rect 3903 -1081 3915 -1047
rect 4083 -1081 4095 -1047
rect 3903 -1087 4095 -1081
rect 4161 -1047 4353 -1041
rect 4161 -1081 4173 -1047
rect 4341 -1081 4353 -1047
rect 4161 -1087 4353 -1081
rect 4419 -1047 4611 -1041
rect 4419 -1081 4431 -1047
rect 4599 -1081 4611 -1047
rect 4419 -1087 4611 -1081
<< properties >>
string FIXED_BBOX -4758 -1166 4758 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 1 m 1 nf 36 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
