magic
tech sky130A
magscale 1 2
timestamp 1664247789
<< pwell >>
rect 1400 0 6538 6516
rect 7700 0 12838 6516
rect 14000 0 19138 6516
rect 20300 0 25438 6516
rect 1400 -7000 6538 -484
rect 7700 -7000 12838 -484
rect 14000 -7000 19138 -484
rect 20300 -7000 25438 -484
<< mvnmos >>
rect 1628 258 1728 6258
rect 1786 258 1886 6258
rect 1944 258 2044 6258
rect 2102 258 2202 6258
rect 2260 258 2360 6258
rect 2418 258 2518 6258
rect 2576 258 2676 6258
rect 2734 258 2834 6258
rect 2892 258 2992 6258
rect 3050 258 3150 6258
rect 3208 258 3308 6258
rect 3366 258 3466 6258
rect 3524 258 3624 6258
rect 3682 258 3782 6258
rect 3840 258 3940 6258
rect 3998 258 4098 6258
rect 4156 258 4256 6258
rect 4314 258 4414 6258
rect 4472 258 4572 6258
rect 4630 258 4730 6258
rect 4788 258 4888 6258
rect 4946 258 5046 6258
rect 5104 258 5204 6258
rect 5262 258 5362 6258
rect 5420 258 5520 6258
rect 5578 258 5678 6258
rect 5736 258 5836 6258
rect 5894 258 5994 6258
rect 6052 258 6152 6258
rect 6210 258 6310 6258
rect 7928 258 8028 6258
rect 8086 258 8186 6258
rect 8244 258 8344 6258
rect 8402 258 8502 6258
rect 8560 258 8660 6258
rect 8718 258 8818 6258
rect 8876 258 8976 6258
rect 9034 258 9134 6258
rect 9192 258 9292 6258
rect 9350 258 9450 6258
rect 9508 258 9608 6258
rect 9666 258 9766 6258
rect 9824 258 9924 6258
rect 9982 258 10082 6258
rect 10140 258 10240 6258
rect 10298 258 10398 6258
rect 10456 258 10556 6258
rect 10614 258 10714 6258
rect 10772 258 10872 6258
rect 10930 258 11030 6258
rect 11088 258 11188 6258
rect 11246 258 11346 6258
rect 11404 258 11504 6258
rect 11562 258 11662 6258
rect 11720 258 11820 6258
rect 11878 258 11978 6258
rect 12036 258 12136 6258
rect 12194 258 12294 6258
rect 12352 258 12452 6258
rect 12510 258 12610 6258
rect 14228 258 14328 6258
rect 14386 258 14486 6258
rect 14544 258 14644 6258
rect 14702 258 14802 6258
rect 14860 258 14960 6258
rect 15018 258 15118 6258
rect 15176 258 15276 6258
rect 15334 258 15434 6258
rect 15492 258 15592 6258
rect 15650 258 15750 6258
rect 15808 258 15908 6258
rect 15966 258 16066 6258
rect 16124 258 16224 6258
rect 16282 258 16382 6258
rect 16440 258 16540 6258
rect 16598 258 16698 6258
rect 16756 258 16856 6258
rect 16914 258 17014 6258
rect 17072 258 17172 6258
rect 17230 258 17330 6258
rect 17388 258 17488 6258
rect 17546 258 17646 6258
rect 17704 258 17804 6258
rect 17862 258 17962 6258
rect 18020 258 18120 6258
rect 18178 258 18278 6258
rect 18336 258 18436 6258
rect 18494 258 18594 6258
rect 18652 258 18752 6258
rect 18810 258 18910 6258
rect 20528 258 20628 6258
rect 20686 258 20786 6258
rect 20844 258 20944 6258
rect 21002 258 21102 6258
rect 21160 258 21260 6258
rect 21318 258 21418 6258
rect 21476 258 21576 6258
rect 21634 258 21734 6258
rect 21792 258 21892 6258
rect 21950 258 22050 6258
rect 22108 258 22208 6258
rect 22266 258 22366 6258
rect 22424 258 22524 6258
rect 22582 258 22682 6258
rect 22740 258 22840 6258
rect 22898 258 22998 6258
rect 23056 258 23156 6258
rect 23214 258 23314 6258
rect 23372 258 23472 6258
rect 23530 258 23630 6258
rect 23688 258 23788 6258
rect 23846 258 23946 6258
rect 24004 258 24104 6258
rect 24162 258 24262 6258
rect 24320 258 24420 6258
rect 24478 258 24578 6258
rect 24636 258 24736 6258
rect 24794 258 24894 6258
rect 24952 258 25052 6258
rect 25110 258 25210 6258
rect 1628 -6742 1728 -742
rect 1786 -6742 1886 -742
rect 1944 -6742 2044 -742
rect 2102 -6742 2202 -742
rect 2260 -6742 2360 -742
rect 2418 -6742 2518 -742
rect 2576 -6742 2676 -742
rect 2734 -6742 2834 -742
rect 2892 -6742 2992 -742
rect 3050 -6742 3150 -742
rect 3208 -6742 3308 -742
rect 3366 -6742 3466 -742
rect 3524 -6742 3624 -742
rect 3682 -6742 3782 -742
rect 3840 -6742 3940 -742
rect 3998 -6742 4098 -742
rect 4156 -6742 4256 -742
rect 4314 -6742 4414 -742
rect 4472 -6742 4572 -742
rect 4630 -6742 4730 -742
rect 4788 -6742 4888 -742
rect 4946 -6742 5046 -742
rect 5104 -6742 5204 -742
rect 5262 -6742 5362 -742
rect 5420 -6742 5520 -742
rect 5578 -6742 5678 -742
rect 5736 -6742 5836 -742
rect 5894 -6742 5994 -742
rect 6052 -6742 6152 -742
rect 6210 -6742 6310 -742
rect 7928 -6742 8028 -742
rect 8086 -6742 8186 -742
rect 8244 -6742 8344 -742
rect 8402 -6742 8502 -742
rect 8560 -6742 8660 -742
rect 8718 -6742 8818 -742
rect 8876 -6742 8976 -742
rect 9034 -6742 9134 -742
rect 9192 -6742 9292 -742
rect 9350 -6742 9450 -742
rect 9508 -6742 9608 -742
rect 9666 -6742 9766 -742
rect 9824 -6742 9924 -742
rect 9982 -6742 10082 -742
rect 10140 -6742 10240 -742
rect 10298 -6742 10398 -742
rect 10456 -6742 10556 -742
rect 10614 -6742 10714 -742
rect 10772 -6742 10872 -742
rect 10930 -6742 11030 -742
rect 11088 -6742 11188 -742
rect 11246 -6742 11346 -742
rect 11404 -6742 11504 -742
rect 11562 -6742 11662 -742
rect 11720 -6742 11820 -742
rect 11878 -6742 11978 -742
rect 12036 -6742 12136 -742
rect 12194 -6742 12294 -742
rect 12352 -6742 12452 -742
rect 12510 -6742 12610 -742
rect 14228 -6742 14328 -742
rect 14386 -6742 14486 -742
rect 14544 -6742 14644 -742
rect 14702 -6742 14802 -742
rect 14860 -6742 14960 -742
rect 15018 -6742 15118 -742
rect 15176 -6742 15276 -742
rect 15334 -6742 15434 -742
rect 15492 -6742 15592 -742
rect 15650 -6742 15750 -742
rect 15808 -6742 15908 -742
rect 15966 -6742 16066 -742
rect 16124 -6742 16224 -742
rect 16282 -6742 16382 -742
rect 16440 -6742 16540 -742
rect 16598 -6742 16698 -742
rect 16756 -6742 16856 -742
rect 16914 -6742 17014 -742
rect 17072 -6742 17172 -742
rect 17230 -6742 17330 -742
rect 17388 -6742 17488 -742
rect 17546 -6742 17646 -742
rect 17704 -6742 17804 -742
rect 17862 -6742 17962 -742
rect 18020 -6742 18120 -742
rect 18178 -6742 18278 -742
rect 18336 -6742 18436 -742
rect 18494 -6742 18594 -742
rect 18652 -6742 18752 -742
rect 18810 -6742 18910 -742
rect 20528 -6742 20628 -742
rect 20686 -6742 20786 -742
rect 20844 -6742 20944 -742
rect 21002 -6742 21102 -742
rect 21160 -6742 21260 -742
rect 21318 -6742 21418 -742
rect 21476 -6742 21576 -742
rect 21634 -6742 21734 -742
rect 21792 -6742 21892 -742
rect 21950 -6742 22050 -742
rect 22108 -6742 22208 -742
rect 22266 -6742 22366 -742
rect 22424 -6742 22524 -742
rect 22582 -6742 22682 -742
rect 22740 -6742 22840 -742
rect 22898 -6742 22998 -742
rect 23056 -6742 23156 -742
rect 23214 -6742 23314 -742
rect 23372 -6742 23472 -742
rect 23530 -6742 23630 -742
rect 23688 -6742 23788 -742
rect 23846 -6742 23946 -742
rect 24004 -6742 24104 -742
rect 24162 -6742 24262 -742
rect 24320 -6742 24420 -742
rect 24478 -6742 24578 -742
rect 24636 -6742 24736 -742
rect 24794 -6742 24894 -742
rect 24952 -6742 25052 -742
rect 25110 -6742 25210 -742
<< mvndiff >>
rect 1570 6246 1628 6258
rect 1570 270 1582 6246
rect 1616 270 1628 6246
rect 1570 258 1628 270
rect 1728 6246 1786 6258
rect 1728 270 1740 6246
rect 1774 270 1786 6246
rect 1728 258 1786 270
rect 1886 6246 1944 6258
rect 1886 270 1898 6246
rect 1932 270 1944 6246
rect 1886 258 1944 270
rect 2044 6246 2102 6258
rect 2044 270 2056 6246
rect 2090 270 2102 6246
rect 2044 258 2102 270
rect 2202 6246 2260 6258
rect 2202 270 2214 6246
rect 2248 270 2260 6246
rect 2202 258 2260 270
rect 2360 6246 2418 6258
rect 2360 270 2372 6246
rect 2406 270 2418 6246
rect 2360 258 2418 270
rect 2518 6246 2576 6258
rect 2518 270 2530 6246
rect 2564 270 2576 6246
rect 2518 258 2576 270
rect 2676 6246 2734 6258
rect 2676 270 2688 6246
rect 2722 270 2734 6246
rect 2676 258 2734 270
rect 2834 6246 2892 6258
rect 2834 270 2846 6246
rect 2880 270 2892 6246
rect 2834 258 2892 270
rect 2992 6246 3050 6258
rect 2992 270 3004 6246
rect 3038 270 3050 6246
rect 2992 258 3050 270
rect 3150 6246 3208 6258
rect 3150 270 3162 6246
rect 3196 270 3208 6246
rect 3150 258 3208 270
rect 3308 6246 3366 6258
rect 3308 270 3320 6246
rect 3354 270 3366 6246
rect 3308 258 3366 270
rect 3466 6246 3524 6258
rect 3466 270 3478 6246
rect 3512 270 3524 6246
rect 3466 258 3524 270
rect 3624 6246 3682 6258
rect 3624 270 3636 6246
rect 3670 270 3682 6246
rect 3624 258 3682 270
rect 3782 6246 3840 6258
rect 3782 270 3794 6246
rect 3828 270 3840 6246
rect 3782 258 3840 270
rect 3940 6246 3998 6258
rect 3940 270 3952 6246
rect 3986 270 3998 6246
rect 3940 258 3998 270
rect 4098 6246 4156 6258
rect 4098 270 4110 6246
rect 4144 270 4156 6246
rect 4098 258 4156 270
rect 4256 6246 4314 6258
rect 4256 270 4268 6246
rect 4302 270 4314 6246
rect 4256 258 4314 270
rect 4414 6246 4472 6258
rect 4414 270 4426 6246
rect 4460 270 4472 6246
rect 4414 258 4472 270
rect 4572 6246 4630 6258
rect 4572 270 4584 6246
rect 4618 270 4630 6246
rect 4572 258 4630 270
rect 4730 6246 4788 6258
rect 4730 270 4742 6246
rect 4776 270 4788 6246
rect 4730 258 4788 270
rect 4888 6246 4946 6258
rect 4888 270 4900 6246
rect 4934 270 4946 6246
rect 4888 258 4946 270
rect 5046 6246 5104 6258
rect 5046 270 5058 6246
rect 5092 270 5104 6246
rect 5046 258 5104 270
rect 5204 6246 5262 6258
rect 5204 270 5216 6246
rect 5250 270 5262 6246
rect 5204 258 5262 270
rect 5362 6246 5420 6258
rect 5362 270 5374 6246
rect 5408 270 5420 6246
rect 5362 258 5420 270
rect 5520 6246 5578 6258
rect 5520 270 5532 6246
rect 5566 270 5578 6246
rect 5520 258 5578 270
rect 5678 6246 5736 6258
rect 5678 270 5690 6246
rect 5724 270 5736 6246
rect 5678 258 5736 270
rect 5836 6246 5894 6258
rect 5836 270 5848 6246
rect 5882 270 5894 6246
rect 5836 258 5894 270
rect 5994 6246 6052 6258
rect 5994 270 6006 6246
rect 6040 270 6052 6246
rect 5994 258 6052 270
rect 6152 6246 6210 6258
rect 6152 270 6164 6246
rect 6198 270 6210 6246
rect 6152 258 6210 270
rect 6310 6246 6368 6258
rect 6310 270 6322 6246
rect 6356 270 6368 6246
rect 6310 258 6368 270
rect 7870 6246 7928 6258
rect 7870 270 7882 6246
rect 7916 270 7928 6246
rect 7870 258 7928 270
rect 8028 6246 8086 6258
rect 8028 270 8040 6246
rect 8074 270 8086 6246
rect 8028 258 8086 270
rect 8186 6246 8244 6258
rect 8186 270 8198 6246
rect 8232 270 8244 6246
rect 8186 258 8244 270
rect 8344 6246 8402 6258
rect 8344 270 8356 6246
rect 8390 270 8402 6246
rect 8344 258 8402 270
rect 8502 6246 8560 6258
rect 8502 270 8514 6246
rect 8548 270 8560 6246
rect 8502 258 8560 270
rect 8660 6246 8718 6258
rect 8660 270 8672 6246
rect 8706 270 8718 6246
rect 8660 258 8718 270
rect 8818 6246 8876 6258
rect 8818 270 8830 6246
rect 8864 270 8876 6246
rect 8818 258 8876 270
rect 8976 6246 9034 6258
rect 8976 270 8988 6246
rect 9022 270 9034 6246
rect 8976 258 9034 270
rect 9134 6246 9192 6258
rect 9134 270 9146 6246
rect 9180 270 9192 6246
rect 9134 258 9192 270
rect 9292 6246 9350 6258
rect 9292 270 9304 6246
rect 9338 270 9350 6246
rect 9292 258 9350 270
rect 9450 6246 9508 6258
rect 9450 270 9462 6246
rect 9496 270 9508 6246
rect 9450 258 9508 270
rect 9608 6246 9666 6258
rect 9608 270 9620 6246
rect 9654 270 9666 6246
rect 9608 258 9666 270
rect 9766 6246 9824 6258
rect 9766 270 9778 6246
rect 9812 270 9824 6246
rect 9766 258 9824 270
rect 9924 6246 9982 6258
rect 9924 270 9936 6246
rect 9970 270 9982 6246
rect 9924 258 9982 270
rect 10082 6246 10140 6258
rect 10082 270 10094 6246
rect 10128 270 10140 6246
rect 10082 258 10140 270
rect 10240 6246 10298 6258
rect 10240 270 10252 6246
rect 10286 270 10298 6246
rect 10240 258 10298 270
rect 10398 6246 10456 6258
rect 10398 270 10410 6246
rect 10444 270 10456 6246
rect 10398 258 10456 270
rect 10556 6246 10614 6258
rect 10556 270 10568 6246
rect 10602 270 10614 6246
rect 10556 258 10614 270
rect 10714 6246 10772 6258
rect 10714 270 10726 6246
rect 10760 270 10772 6246
rect 10714 258 10772 270
rect 10872 6246 10930 6258
rect 10872 270 10884 6246
rect 10918 270 10930 6246
rect 10872 258 10930 270
rect 11030 6246 11088 6258
rect 11030 270 11042 6246
rect 11076 270 11088 6246
rect 11030 258 11088 270
rect 11188 6246 11246 6258
rect 11188 270 11200 6246
rect 11234 270 11246 6246
rect 11188 258 11246 270
rect 11346 6246 11404 6258
rect 11346 270 11358 6246
rect 11392 270 11404 6246
rect 11346 258 11404 270
rect 11504 6246 11562 6258
rect 11504 270 11516 6246
rect 11550 270 11562 6246
rect 11504 258 11562 270
rect 11662 6246 11720 6258
rect 11662 270 11674 6246
rect 11708 270 11720 6246
rect 11662 258 11720 270
rect 11820 6246 11878 6258
rect 11820 270 11832 6246
rect 11866 270 11878 6246
rect 11820 258 11878 270
rect 11978 6246 12036 6258
rect 11978 270 11990 6246
rect 12024 270 12036 6246
rect 11978 258 12036 270
rect 12136 6246 12194 6258
rect 12136 270 12148 6246
rect 12182 270 12194 6246
rect 12136 258 12194 270
rect 12294 6246 12352 6258
rect 12294 270 12306 6246
rect 12340 270 12352 6246
rect 12294 258 12352 270
rect 12452 6246 12510 6258
rect 12452 270 12464 6246
rect 12498 270 12510 6246
rect 12452 258 12510 270
rect 12610 6246 12668 6258
rect 12610 270 12622 6246
rect 12656 270 12668 6246
rect 12610 258 12668 270
rect 14170 6246 14228 6258
rect 14170 270 14182 6246
rect 14216 270 14228 6246
rect 14170 258 14228 270
rect 14328 6246 14386 6258
rect 14328 270 14340 6246
rect 14374 270 14386 6246
rect 14328 258 14386 270
rect 14486 6246 14544 6258
rect 14486 270 14498 6246
rect 14532 270 14544 6246
rect 14486 258 14544 270
rect 14644 6246 14702 6258
rect 14644 270 14656 6246
rect 14690 270 14702 6246
rect 14644 258 14702 270
rect 14802 6246 14860 6258
rect 14802 270 14814 6246
rect 14848 270 14860 6246
rect 14802 258 14860 270
rect 14960 6246 15018 6258
rect 14960 270 14972 6246
rect 15006 270 15018 6246
rect 14960 258 15018 270
rect 15118 6246 15176 6258
rect 15118 270 15130 6246
rect 15164 270 15176 6246
rect 15118 258 15176 270
rect 15276 6246 15334 6258
rect 15276 270 15288 6246
rect 15322 270 15334 6246
rect 15276 258 15334 270
rect 15434 6246 15492 6258
rect 15434 270 15446 6246
rect 15480 270 15492 6246
rect 15434 258 15492 270
rect 15592 6246 15650 6258
rect 15592 270 15604 6246
rect 15638 270 15650 6246
rect 15592 258 15650 270
rect 15750 6246 15808 6258
rect 15750 270 15762 6246
rect 15796 270 15808 6246
rect 15750 258 15808 270
rect 15908 6246 15966 6258
rect 15908 270 15920 6246
rect 15954 270 15966 6246
rect 15908 258 15966 270
rect 16066 6246 16124 6258
rect 16066 270 16078 6246
rect 16112 270 16124 6246
rect 16066 258 16124 270
rect 16224 6246 16282 6258
rect 16224 270 16236 6246
rect 16270 270 16282 6246
rect 16224 258 16282 270
rect 16382 6246 16440 6258
rect 16382 270 16394 6246
rect 16428 270 16440 6246
rect 16382 258 16440 270
rect 16540 6246 16598 6258
rect 16540 270 16552 6246
rect 16586 270 16598 6246
rect 16540 258 16598 270
rect 16698 6246 16756 6258
rect 16698 270 16710 6246
rect 16744 270 16756 6246
rect 16698 258 16756 270
rect 16856 6246 16914 6258
rect 16856 270 16868 6246
rect 16902 270 16914 6246
rect 16856 258 16914 270
rect 17014 6246 17072 6258
rect 17014 270 17026 6246
rect 17060 270 17072 6246
rect 17014 258 17072 270
rect 17172 6246 17230 6258
rect 17172 270 17184 6246
rect 17218 270 17230 6246
rect 17172 258 17230 270
rect 17330 6246 17388 6258
rect 17330 270 17342 6246
rect 17376 270 17388 6246
rect 17330 258 17388 270
rect 17488 6246 17546 6258
rect 17488 270 17500 6246
rect 17534 270 17546 6246
rect 17488 258 17546 270
rect 17646 6246 17704 6258
rect 17646 270 17658 6246
rect 17692 270 17704 6246
rect 17646 258 17704 270
rect 17804 6246 17862 6258
rect 17804 270 17816 6246
rect 17850 270 17862 6246
rect 17804 258 17862 270
rect 17962 6246 18020 6258
rect 17962 270 17974 6246
rect 18008 270 18020 6246
rect 17962 258 18020 270
rect 18120 6246 18178 6258
rect 18120 270 18132 6246
rect 18166 270 18178 6246
rect 18120 258 18178 270
rect 18278 6246 18336 6258
rect 18278 270 18290 6246
rect 18324 270 18336 6246
rect 18278 258 18336 270
rect 18436 6246 18494 6258
rect 18436 270 18448 6246
rect 18482 270 18494 6246
rect 18436 258 18494 270
rect 18594 6246 18652 6258
rect 18594 270 18606 6246
rect 18640 270 18652 6246
rect 18594 258 18652 270
rect 18752 6246 18810 6258
rect 18752 270 18764 6246
rect 18798 270 18810 6246
rect 18752 258 18810 270
rect 18910 6246 18968 6258
rect 18910 270 18922 6246
rect 18956 270 18968 6246
rect 18910 258 18968 270
rect 20470 6246 20528 6258
rect 20470 270 20482 6246
rect 20516 270 20528 6246
rect 20470 258 20528 270
rect 20628 6246 20686 6258
rect 20628 270 20640 6246
rect 20674 270 20686 6246
rect 20628 258 20686 270
rect 20786 6246 20844 6258
rect 20786 270 20798 6246
rect 20832 270 20844 6246
rect 20786 258 20844 270
rect 20944 6246 21002 6258
rect 20944 270 20956 6246
rect 20990 270 21002 6246
rect 20944 258 21002 270
rect 21102 6246 21160 6258
rect 21102 270 21114 6246
rect 21148 270 21160 6246
rect 21102 258 21160 270
rect 21260 6246 21318 6258
rect 21260 270 21272 6246
rect 21306 270 21318 6246
rect 21260 258 21318 270
rect 21418 6246 21476 6258
rect 21418 270 21430 6246
rect 21464 270 21476 6246
rect 21418 258 21476 270
rect 21576 6246 21634 6258
rect 21576 270 21588 6246
rect 21622 270 21634 6246
rect 21576 258 21634 270
rect 21734 6246 21792 6258
rect 21734 270 21746 6246
rect 21780 270 21792 6246
rect 21734 258 21792 270
rect 21892 6246 21950 6258
rect 21892 270 21904 6246
rect 21938 270 21950 6246
rect 21892 258 21950 270
rect 22050 6246 22108 6258
rect 22050 270 22062 6246
rect 22096 270 22108 6246
rect 22050 258 22108 270
rect 22208 6246 22266 6258
rect 22208 270 22220 6246
rect 22254 270 22266 6246
rect 22208 258 22266 270
rect 22366 6246 22424 6258
rect 22366 270 22378 6246
rect 22412 270 22424 6246
rect 22366 258 22424 270
rect 22524 6246 22582 6258
rect 22524 270 22536 6246
rect 22570 270 22582 6246
rect 22524 258 22582 270
rect 22682 6246 22740 6258
rect 22682 270 22694 6246
rect 22728 270 22740 6246
rect 22682 258 22740 270
rect 22840 6246 22898 6258
rect 22840 270 22852 6246
rect 22886 270 22898 6246
rect 22840 258 22898 270
rect 22998 6246 23056 6258
rect 22998 270 23010 6246
rect 23044 270 23056 6246
rect 22998 258 23056 270
rect 23156 6246 23214 6258
rect 23156 270 23168 6246
rect 23202 270 23214 6246
rect 23156 258 23214 270
rect 23314 6246 23372 6258
rect 23314 270 23326 6246
rect 23360 270 23372 6246
rect 23314 258 23372 270
rect 23472 6246 23530 6258
rect 23472 270 23484 6246
rect 23518 270 23530 6246
rect 23472 258 23530 270
rect 23630 6246 23688 6258
rect 23630 270 23642 6246
rect 23676 270 23688 6246
rect 23630 258 23688 270
rect 23788 6246 23846 6258
rect 23788 270 23800 6246
rect 23834 270 23846 6246
rect 23788 258 23846 270
rect 23946 6246 24004 6258
rect 23946 270 23958 6246
rect 23992 270 24004 6246
rect 23946 258 24004 270
rect 24104 6246 24162 6258
rect 24104 270 24116 6246
rect 24150 270 24162 6246
rect 24104 258 24162 270
rect 24262 6246 24320 6258
rect 24262 270 24274 6246
rect 24308 270 24320 6246
rect 24262 258 24320 270
rect 24420 6246 24478 6258
rect 24420 270 24432 6246
rect 24466 270 24478 6246
rect 24420 258 24478 270
rect 24578 6246 24636 6258
rect 24578 270 24590 6246
rect 24624 270 24636 6246
rect 24578 258 24636 270
rect 24736 6246 24794 6258
rect 24736 270 24748 6246
rect 24782 270 24794 6246
rect 24736 258 24794 270
rect 24894 6246 24952 6258
rect 24894 270 24906 6246
rect 24940 270 24952 6246
rect 24894 258 24952 270
rect 25052 6246 25110 6258
rect 25052 270 25064 6246
rect 25098 270 25110 6246
rect 25052 258 25110 270
rect 25210 6246 25268 6258
rect 25210 270 25222 6246
rect 25256 270 25268 6246
rect 25210 258 25268 270
rect 1570 -754 1628 -742
rect 1570 -6730 1582 -754
rect 1616 -6730 1628 -754
rect 1570 -6742 1628 -6730
rect 1728 -754 1786 -742
rect 1728 -6730 1740 -754
rect 1774 -6730 1786 -754
rect 1728 -6742 1786 -6730
rect 1886 -754 1944 -742
rect 1886 -6730 1898 -754
rect 1932 -6730 1944 -754
rect 1886 -6742 1944 -6730
rect 2044 -754 2102 -742
rect 2044 -6730 2056 -754
rect 2090 -6730 2102 -754
rect 2044 -6742 2102 -6730
rect 2202 -754 2260 -742
rect 2202 -6730 2214 -754
rect 2248 -6730 2260 -754
rect 2202 -6742 2260 -6730
rect 2360 -754 2418 -742
rect 2360 -6730 2372 -754
rect 2406 -6730 2418 -754
rect 2360 -6742 2418 -6730
rect 2518 -754 2576 -742
rect 2518 -6730 2530 -754
rect 2564 -6730 2576 -754
rect 2518 -6742 2576 -6730
rect 2676 -754 2734 -742
rect 2676 -6730 2688 -754
rect 2722 -6730 2734 -754
rect 2676 -6742 2734 -6730
rect 2834 -754 2892 -742
rect 2834 -6730 2846 -754
rect 2880 -6730 2892 -754
rect 2834 -6742 2892 -6730
rect 2992 -754 3050 -742
rect 2992 -6730 3004 -754
rect 3038 -6730 3050 -754
rect 2992 -6742 3050 -6730
rect 3150 -754 3208 -742
rect 3150 -6730 3162 -754
rect 3196 -6730 3208 -754
rect 3150 -6742 3208 -6730
rect 3308 -754 3366 -742
rect 3308 -6730 3320 -754
rect 3354 -6730 3366 -754
rect 3308 -6742 3366 -6730
rect 3466 -754 3524 -742
rect 3466 -6730 3478 -754
rect 3512 -6730 3524 -754
rect 3466 -6742 3524 -6730
rect 3624 -754 3682 -742
rect 3624 -6730 3636 -754
rect 3670 -6730 3682 -754
rect 3624 -6742 3682 -6730
rect 3782 -754 3840 -742
rect 3782 -6730 3794 -754
rect 3828 -6730 3840 -754
rect 3782 -6742 3840 -6730
rect 3940 -754 3998 -742
rect 3940 -6730 3952 -754
rect 3986 -6730 3998 -754
rect 3940 -6742 3998 -6730
rect 4098 -754 4156 -742
rect 4098 -6730 4110 -754
rect 4144 -6730 4156 -754
rect 4098 -6742 4156 -6730
rect 4256 -754 4314 -742
rect 4256 -6730 4268 -754
rect 4302 -6730 4314 -754
rect 4256 -6742 4314 -6730
rect 4414 -754 4472 -742
rect 4414 -6730 4426 -754
rect 4460 -6730 4472 -754
rect 4414 -6742 4472 -6730
rect 4572 -754 4630 -742
rect 4572 -6730 4584 -754
rect 4618 -6730 4630 -754
rect 4572 -6742 4630 -6730
rect 4730 -754 4788 -742
rect 4730 -6730 4742 -754
rect 4776 -6730 4788 -754
rect 4730 -6742 4788 -6730
rect 4888 -754 4946 -742
rect 4888 -6730 4900 -754
rect 4934 -6730 4946 -754
rect 4888 -6742 4946 -6730
rect 5046 -754 5104 -742
rect 5046 -6730 5058 -754
rect 5092 -6730 5104 -754
rect 5046 -6742 5104 -6730
rect 5204 -754 5262 -742
rect 5204 -6730 5216 -754
rect 5250 -6730 5262 -754
rect 5204 -6742 5262 -6730
rect 5362 -754 5420 -742
rect 5362 -6730 5374 -754
rect 5408 -6730 5420 -754
rect 5362 -6742 5420 -6730
rect 5520 -754 5578 -742
rect 5520 -6730 5532 -754
rect 5566 -6730 5578 -754
rect 5520 -6742 5578 -6730
rect 5678 -754 5736 -742
rect 5678 -6730 5690 -754
rect 5724 -6730 5736 -754
rect 5678 -6742 5736 -6730
rect 5836 -754 5894 -742
rect 5836 -6730 5848 -754
rect 5882 -6730 5894 -754
rect 5836 -6742 5894 -6730
rect 5994 -754 6052 -742
rect 5994 -6730 6006 -754
rect 6040 -6730 6052 -754
rect 5994 -6742 6052 -6730
rect 6152 -754 6210 -742
rect 6152 -6730 6164 -754
rect 6198 -6730 6210 -754
rect 6152 -6742 6210 -6730
rect 6310 -754 6368 -742
rect 6310 -6730 6322 -754
rect 6356 -6730 6368 -754
rect 6310 -6742 6368 -6730
rect 7870 -754 7928 -742
rect 7870 -6730 7882 -754
rect 7916 -6730 7928 -754
rect 7870 -6742 7928 -6730
rect 8028 -754 8086 -742
rect 8028 -6730 8040 -754
rect 8074 -6730 8086 -754
rect 8028 -6742 8086 -6730
rect 8186 -754 8244 -742
rect 8186 -6730 8198 -754
rect 8232 -6730 8244 -754
rect 8186 -6742 8244 -6730
rect 8344 -754 8402 -742
rect 8344 -6730 8356 -754
rect 8390 -6730 8402 -754
rect 8344 -6742 8402 -6730
rect 8502 -754 8560 -742
rect 8502 -6730 8514 -754
rect 8548 -6730 8560 -754
rect 8502 -6742 8560 -6730
rect 8660 -754 8718 -742
rect 8660 -6730 8672 -754
rect 8706 -6730 8718 -754
rect 8660 -6742 8718 -6730
rect 8818 -754 8876 -742
rect 8818 -6730 8830 -754
rect 8864 -6730 8876 -754
rect 8818 -6742 8876 -6730
rect 8976 -754 9034 -742
rect 8976 -6730 8988 -754
rect 9022 -6730 9034 -754
rect 8976 -6742 9034 -6730
rect 9134 -754 9192 -742
rect 9134 -6730 9146 -754
rect 9180 -6730 9192 -754
rect 9134 -6742 9192 -6730
rect 9292 -754 9350 -742
rect 9292 -6730 9304 -754
rect 9338 -6730 9350 -754
rect 9292 -6742 9350 -6730
rect 9450 -754 9508 -742
rect 9450 -6730 9462 -754
rect 9496 -6730 9508 -754
rect 9450 -6742 9508 -6730
rect 9608 -754 9666 -742
rect 9608 -6730 9620 -754
rect 9654 -6730 9666 -754
rect 9608 -6742 9666 -6730
rect 9766 -754 9824 -742
rect 9766 -6730 9778 -754
rect 9812 -6730 9824 -754
rect 9766 -6742 9824 -6730
rect 9924 -754 9982 -742
rect 9924 -6730 9936 -754
rect 9970 -6730 9982 -754
rect 9924 -6742 9982 -6730
rect 10082 -754 10140 -742
rect 10082 -6730 10094 -754
rect 10128 -6730 10140 -754
rect 10082 -6742 10140 -6730
rect 10240 -754 10298 -742
rect 10240 -6730 10252 -754
rect 10286 -6730 10298 -754
rect 10240 -6742 10298 -6730
rect 10398 -754 10456 -742
rect 10398 -6730 10410 -754
rect 10444 -6730 10456 -754
rect 10398 -6742 10456 -6730
rect 10556 -754 10614 -742
rect 10556 -6730 10568 -754
rect 10602 -6730 10614 -754
rect 10556 -6742 10614 -6730
rect 10714 -754 10772 -742
rect 10714 -6730 10726 -754
rect 10760 -6730 10772 -754
rect 10714 -6742 10772 -6730
rect 10872 -754 10930 -742
rect 10872 -6730 10884 -754
rect 10918 -6730 10930 -754
rect 10872 -6742 10930 -6730
rect 11030 -754 11088 -742
rect 11030 -6730 11042 -754
rect 11076 -6730 11088 -754
rect 11030 -6742 11088 -6730
rect 11188 -754 11246 -742
rect 11188 -6730 11200 -754
rect 11234 -6730 11246 -754
rect 11188 -6742 11246 -6730
rect 11346 -754 11404 -742
rect 11346 -6730 11358 -754
rect 11392 -6730 11404 -754
rect 11346 -6742 11404 -6730
rect 11504 -754 11562 -742
rect 11504 -6730 11516 -754
rect 11550 -6730 11562 -754
rect 11504 -6742 11562 -6730
rect 11662 -754 11720 -742
rect 11662 -6730 11674 -754
rect 11708 -6730 11720 -754
rect 11662 -6742 11720 -6730
rect 11820 -754 11878 -742
rect 11820 -6730 11832 -754
rect 11866 -6730 11878 -754
rect 11820 -6742 11878 -6730
rect 11978 -754 12036 -742
rect 11978 -6730 11990 -754
rect 12024 -6730 12036 -754
rect 11978 -6742 12036 -6730
rect 12136 -754 12194 -742
rect 12136 -6730 12148 -754
rect 12182 -6730 12194 -754
rect 12136 -6742 12194 -6730
rect 12294 -754 12352 -742
rect 12294 -6730 12306 -754
rect 12340 -6730 12352 -754
rect 12294 -6742 12352 -6730
rect 12452 -754 12510 -742
rect 12452 -6730 12464 -754
rect 12498 -6730 12510 -754
rect 12452 -6742 12510 -6730
rect 12610 -754 12668 -742
rect 12610 -6730 12622 -754
rect 12656 -6730 12668 -754
rect 12610 -6742 12668 -6730
rect 14170 -754 14228 -742
rect 14170 -6730 14182 -754
rect 14216 -6730 14228 -754
rect 14170 -6742 14228 -6730
rect 14328 -754 14386 -742
rect 14328 -6730 14340 -754
rect 14374 -6730 14386 -754
rect 14328 -6742 14386 -6730
rect 14486 -754 14544 -742
rect 14486 -6730 14498 -754
rect 14532 -6730 14544 -754
rect 14486 -6742 14544 -6730
rect 14644 -754 14702 -742
rect 14644 -6730 14656 -754
rect 14690 -6730 14702 -754
rect 14644 -6742 14702 -6730
rect 14802 -754 14860 -742
rect 14802 -6730 14814 -754
rect 14848 -6730 14860 -754
rect 14802 -6742 14860 -6730
rect 14960 -754 15018 -742
rect 14960 -6730 14972 -754
rect 15006 -6730 15018 -754
rect 14960 -6742 15018 -6730
rect 15118 -754 15176 -742
rect 15118 -6730 15130 -754
rect 15164 -6730 15176 -754
rect 15118 -6742 15176 -6730
rect 15276 -754 15334 -742
rect 15276 -6730 15288 -754
rect 15322 -6730 15334 -754
rect 15276 -6742 15334 -6730
rect 15434 -754 15492 -742
rect 15434 -6730 15446 -754
rect 15480 -6730 15492 -754
rect 15434 -6742 15492 -6730
rect 15592 -754 15650 -742
rect 15592 -6730 15604 -754
rect 15638 -6730 15650 -754
rect 15592 -6742 15650 -6730
rect 15750 -754 15808 -742
rect 15750 -6730 15762 -754
rect 15796 -6730 15808 -754
rect 15750 -6742 15808 -6730
rect 15908 -754 15966 -742
rect 15908 -6730 15920 -754
rect 15954 -6730 15966 -754
rect 15908 -6742 15966 -6730
rect 16066 -754 16124 -742
rect 16066 -6730 16078 -754
rect 16112 -6730 16124 -754
rect 16066 -6742 16124 -6730
rect 16224 -754 16282 -742
rect 16224 -6730 16236 -754
rect 16270 -6730 16282 -754
rect 16224 -6742 16282 -6730
rect 16382 -754 16440 -742
rect 16382 -6730 16394 -754
rect 16428 -6730 16440 -754
rect 16382 -6742 16440 -6730
rect 16540 -754 16598 -742
rect 16540 -6730 16552 -754
rect 16586 -6730 16598 -754
rect 16540 -6742 16598 -6730
rect 16698 -754 16756 -742
rect 16698 -6730 16710 -754
rect 16744 -6730 16756 -754
rect 16698 -6742 16756 -6730
rect 16856 -754 16914 -742
rect 16856 -6730 16868 -754
rect 16902 -6730 16914 -754
rect 16856 -6742 16914 -6730
rect 17014 -754 17072 -742
rect 17014 -6730 17026 -754
rect 17060 -6730 17072 -754
rect 17014 -6742 17072 -6730
rect 17172 -754 17230 -742
rect 17172 -6730 17184 -754
rect 17218 -6730 17230 -754
rect 17172 -6742 17230 -6730
rect 17330 -754 17388 -742
rect 17330 -6730 17342 -754
rect 17376 -6730 17388 -754
rect 17330 -6742 17388 -6730
rect 17488 -754 17546 -742
rect 17488 -6730 17500 -754
rect 17534 -6730 17546 -754
rect 17488 -6742 17546 -6730
rect 17646 -754 17704 -742
rect 17646 -6730 17658 -754
rect 17692 -6730 17704 -754
rect 17646 -6742 17704 -6730
rect 17804 -754 17862 -742
rect 17804 -6730 17816 -754
rect 17850 -6730 17862 -754
rect 17804 -6742 17862 -6730
rect 17962 -754 18020 -742
rect 17962 -6730 17974 -754
rect 18008 -6730 18020 -754
rect 17962 -6742 18020 -6730
rect 18120 -754 18178 -742
rect 18120 -6730 18132 -754
rect 18166 -6730 18178 -754
rect 18120 -6742 18178 -6730
rect 18278 -754 18336 -742
rect 18278 -6730 18290 -754
rect 18324 -6730 18336 -754
rect 18278 -6742 18336 -6730
rect 18436 -754 18494 -742
rect 18436 -6730 18448 -754
rect 18482 -6730 18494 -754
rect 18436 -6742 18494 -6730
rect 18594 -754 18652 -742
rect 18594 -6730 18606 -754
rect 18640 -6730 18652 -754
rect 18594 -6742 18652 -6730
rect 18752 -754 18810 -742
rect 18752 -6730 18764 -754
rect 18798 -6730 18810 -754
rect 18752 -6742 18810 -6730
rect 18910 -754 18968 -742
rect 18910 -6730 18922 -754
rect 18956 -6730 18968 -754
rect 18910 -6742 18968 -6730
rect 20470 -754 20528 -742
rect 20470 -6730 20482 -754
rect 20516 -6730 20528 -754
rect 20470 -6742 20528 -6730
rect 20628 -754 20686 -742
rect 20628 -6730 20640 -754
rect 20674 -6730 20686 -754
rect 20628 -6742 20686 -6730
rect 20786 -754 20844 -742
rect 20786 -6730 20798 -754
rect 20832 -6730 20844 -754
rect 20786 -6742 20844 -6730
rect 20944 -754 21002 -742
rect 20944 -6730 20956 -754
rect 20990 -6730 21002 -754
rect 20944 -6742 21002 -6730
rect 21102 -754 21160 -742
rect 21102 -6730 21114 -754
rect 21148 -6730 21160 -754
rect 21102 -6742 21160 -6730
rect 21260 -754 21318 -742
rect 21260 -6730 21272 -754
rect 21306 -6730 21318 -754
rect 21260 -6742 21318 -6730
rect 21418 -754 21476 -742
rect 21418 -6730 21430 -754
rect 21464 -6730 21476 -754
rect 21418 -6742 21476 -6730
rect 21576 -754 21634 -742
rect 21576 -6730 21588 -754
rect 21622 -6730 21634 -754
rect 21576 -6742 21634 -6730
rect 21734 -754 21792 -742
rect 21734 -6730 21746 -754
rect 21780 -6730 21792 -754
rect 21734 -6742 21792 -6730
rect 21892 -754 21950 -742
rect 21892 -6730 21904 -754
rect 21938 -6730 21950 -754
rect 21892 -6742 21950 -6730
rect 22050 -754 22108 -742
rect 22050 -6730 22062 -754
rect 22096 -6730 22108 -754
rect 22050 -6742 22108 -6730
rect 22208 -754 22266 -742
rect 22208 -6730 22220 -754
rect 22254 -6730 22266 -754
rect 22208 -6742 22266 -6730
rect 22366 -754 22424 -742
rect 22366 -6730 22378 -754
rect 22412 -6730 22424 -754
rect 22366 -6742 22424 -6730
rect 22524 -754 22582 -742
rect 22524 -6730 22536 -754
rect 22570 -6730 22582 -754
rect 22524 -6742 22582 -6730
rect 22682 -754 22740 -742
rect 22682 -6730 22694 -754
rect 22728 -6730 22740 -754
rect 22682 -6742 22740 -6730
rect 22840 -754 22898 -742
rect 22840 -6730 22852 -754
rect 22886 -6730 22898 -754
rect 22840 -6742 22898 -6730
rect 22998 -754 23056 -742
rect 22998 -6730 23010 -754
rect 23044 -6730 23056 -754
rect 22998 -6742 23056 -6730
rect 23156 -754 23214 -742
rect 23156 -6730 23168 -754
rect 23202 -6730 23214 -754
rect 23156 -6742 23214 -6730
rect 23314 -754 23372 -742
rect 23314 -6730 23326 -754
rect 23360 -6730 23372 -754
rect 23314 -6742 23372 -6730
rect 23472 -754 23530 -742
rect 23472 -6730 23484 -754
rect 23518 -6730 23530 -754
rect 23472 -6742 23530 -6730
rect 23630 -754 23688 -742
rect 23630 -6730 23642 -754
rect 23676 -6730 23688 -754
rect 23630 -6742 23688 -6730
rect 23788 -754 23846 -742
rect 23788 -6730 23800 -754
rect 23834 -6730 23846 -754
rect 23788 -6742 23846 -6730
rect 23946 -754 24004 -742
rect 23946 -6730 23958 -754
rect 23992 -6730 24004 -754
rect 23946 -6742 24004 -6730
rect 24104 -754 24162 -742
rect 24104 -6730 24116 -754
rect 24150 -6730 24162 -754
rect 24104 -6742 24162 -6730
rect 24262 -754 24320 -742
rect 24262 -6730 24274 -754
rect 24308 -6730 24320 -754
rect 24262 -6742 24320 -6730
rect 24420 -754 24478 -742
rect 24420 -6730 24432 -754
rect 24466 -6730 24478 -754
rect 24420 -6742 24478 -6730
rect 24578 -754 24636 -742
rect 24578 -6730 24590 -754
rect 24624 -6730 24636 -754
rect 24578 -6742 24636 -6730
rect 24736 -754 24794 -742
rect 24736 -6730 24748 -754
rect 24782 -6730 24794 -754
rect 24736 -6742 24794 -6730
rect 24894 -754 24952 -742
rect 24894 -6730 24906 -754
rect 24940 -6730 24952 -754
rect 24894 -6742 24952 -6730
rect 25052 -754 25110 -742
rect 25052 -6730 25064 -754
rect 25098 -6730 25110 -754
rect 25052 -6742 25110 -6730
rect 25210 -754 25268 -742
rect 25210 -6730 25222 -754
rect 25256 -6730 25268 -754
rect 25210 -6742 25268 -6730
<< mvndiffc >>
rect 1582 270 1616 6246
rect 1740 270 1774 6246
rect 1898 270 1932 6246
rect 2056 270 2090 6246
rect 2214 270 2248 6246
rect 2372 270 2406 6246
rect 2530 270 2564 6246
rect 2688 270 2722 6246
rect 2846 270 2880 6246
rect 3004 270 3038 6246
rect 3162 270 3196 6246
rect 3320 270 3354 6246
rect 3478 270 3512 6246
rect 3636 270 3670 6246
rect 3794 270 3828 6246
rect 3952 270 3986 6246
rect 4110 270 4144 6246
rect 4268 270 4302 6246
rect 4426 270 4460 6246
rect 4584 270 4618 6246
rect 4742 270 4776 6246
rect 4900 270 4934 6246
rect 5058 270 5092 6246
rect 5216 270 5250 6246
rect 5374 270 5408 6246
rect 5532 270 5566 6246
rect 5690 270 5724 6246
rect 5848 270 5882 6246
rect 6006 270 6040 6246
rect 6164 270 6198 6246
rect 6322 270 6356 6246
rect 7882 270 7916 6246
rect 8040 270 8074 6246
rect 8198 270 8232 6246
rect 8356 270 8390 6246
rect 8514 270 8548 6246
rect 8672 270 8706 6246
rect 8830 270 8864 6246
rect 8988 270 9022 6246
rect 9146 270 9180 6246
rect 9304 270 9338 6246
rect 9462 270 9496 6246
rect 9620 270 9654 6246
rect 9778 270 9812 6246
rect 9936 270 9970 6246
rect 10094 270 10128 6246
rect 10252 270 10286 6246
rect 10410 270 10444 6246
rect 10568 270 10602 6246
rect 10726 270 10760 6246
rect 10884 270 10918 6246
rect 11042 270 11076 6246
rect 11200 270 11234 6246
rect 11358 270 11392 6246
rect 11516 270 11550 6246
rect 11674 270 11708 6246
rect 11832 270 11866 6246
rect 11990 270 12024 6246
rect 12148 270 12182 6246
rect 12306 270 12340 6246
rect 12464 270 12498 6246
rect 12622 270 12656 6246
rect 14182 270 14216 6246
rect 14340 270 14374 6246
rect 14498 270 14532 6246
rect 14656 270 14690 6246
rect 14814 270 14848 6246
rect 14972 270 15006 6246
rect 15130 270 15164 6246
rect 15288 270 15322 6246
rect 15446 270 15480 6246
rect 15604 270 15638 6246
rect 15762 270 15796 6246
rect 15920 270 15954 6246
rect 16078 270 16112 6246
rect 16236 270 16270 6246
rect 16394 270 16428 6246
rect 16552 270 16586 6246
rect 16710 270 16744 6246
rect 16868 270 16902 6246
rect 17026 270 17060 6246
rect 17184 270 17218 6246
rect 17342 270 17376 6246
rect 17500 270 17534 6246
rect 17658 270 17692 6246
rect 17816 270 17850 6246
rect 17974 270 18008 6246
rect 18132 270 18166 6246
rect 18290 270 18324 6246
rect 18448 270 18482 6246
rect 18606 270 18640 6246
rect 18764 270 18798 6246
rect 18922 270 18956 6246
rect 20482 270 20516 6246
rect 20640 270 20674 6246
rect 20798 270 20832 6246
rect 20956 270 20990 6246
rect 21114 270 21148 6246
rect 21272 270 21306 6246
rect 21430 270 21464 6246
rect 21588 270 21622 6246
rect 21746 270 21780 6246
rect 21904 270 21938 6246
rect 22062 270 22096 6246
rect 22220 270 22254 6246
rect 22378 270 22412 6246
rect 22536 270 22570 6246
rect 22694 270 22728 6246
rect 22852 270 22886 6246
rect 23010 270 23044 6246
rect 23168 270 23202 6246
rect 23326 270 23360 6246
rect 23484 270 23518 6246
rect 23642 270 23676 6246
rect 23800 270 23834 6246
rect 23958 270 23992 6246
rect 24116 270 24150 6246
rect 24274 270 24308 6246
rect 24432 270 24466 6246
rect 24590 270 24624 6246
rect 24748 270 24782 6246
rect 24906 270 24940 6246
rect 25064 270 25098 6246
rect 25222 270 25256 6246
rect 1582 -6730 1616 -754
rect 1740 -6730 1774 -754
rect 1898 -6730 1932 -754
rect 2056 -6730 2090 -754
rect 2214 -6730 2248 -754
rect 2372 -6730 2406 -754
rect 2530 -6730 2564 -754
rect 2688 -6730 2722 -754
rect 2846 -6730 2880 -754
rect 3004 -6730 3038 -754
rect 3162 -6730 3196 -754
rect 3320 -6730 3354 -754
rect 3478 -6730 3512 -754
rect 3636 -6730 3670 -754
rect 3794 -6730 3828 -754
rect 3952 -6730 3986 -754
rect 4110 -6730 4144 -754
rect 4268 -6730 4302 -754
rect 4426 -6730 4460 -754
rect 4584 -6730 4618 -754
rect 4742 -6730 4776 -754
rect 4900 -6730 4934 -754
rect 5058 -6730 5092 -754
rect 5216 -6730 5250 -754
rect 5374 -6730 5408 -754
rect 5532 -6730 5566 -754
rect 5690 -6730 5724 -754
rect 5848 -6730 5882 -754
rect 6006 -6730 6040 -754
rect 6164 -6730 6198 -754
rect 6322 -6730 6356 -754
rect 7882 -6730 7916 -754
rect 8040 -6730 8074 -754
rect 8198 -6730 8232 -754
rect 8356 -6730 8390 -754
rect 8514 -6730 8548 -754
rect 8672 -6730 8706 -754
rect 8830 -6730 8864 -754
rect 8988 -6730 9022 -754
rect 9146 -6730 9180 -754
rect 9304 -6730 9338 -754
rect 9462 -6730 9496 -754
rect 9620 -6730 9654 -754
rect 9778 -6730 9812 -754
rect 9936 -6730 9970 -754
rect 10094 -6730 10128 -754
rect 10252 -6730 10286 -754
rect 10410 -6730 10444 -754
rect 10568 -6730 10602 -754
rect 10726 -6730 10760 -754
rect 10884 -6730 10918 -754
rect 11042 -6730 11076 -754
rect 11200 -6730 11234 -754
rect 11358 -6730 11392 -754
rect 11516 -6730 11550 -754
rect 11674 -6730 11708 -754
rect 11832 -6730 11866 -754
rect 11990 -6730 12024 -754
rect 12148 -6730 12182 -754
rect 12306 -6730 12340 -754
rect 12464 -6730 12498 -754
rect 12622 -6730 12656 -754
rect 14182 -6730 14216 -754
rect 14340 -6730 14374 -754
rect 14498 -6730 14532 -754
rect 14656 -6730 14690 -754
rect 14814 -6730 14848 -754
rect 14972 -6730 15006 -754
rect 15130 -6730 15164 -754
rect 15288 -6730 15322 -754
rect 15446 -6730 15480 -754
rect 15604 -6730 15638 -754
rect 15762 -6730 15796 -754
rect 15920 -6730 15954 -754
rect 16078 -6730 16112 -754
rect 16236 -6730 16270 -754
rect 16394 -6730 16428 -754
rect 16552 -6730 16586 -754
rect 16710 -6730 16744 -754
rect 16868 -6730 16902 -754
rect 17026 -6730 17060 -754
rect 17184 -6730 17218 -754
rect 17342 -6730 17376 -754
rect 17500 -6730 17534 -754
rect 17658 -6730 17692 -754
rect 17816 -6730 17850 -754
rect 17974 -6730 18008 -754
rect 18132 -6730 18166 -754
rect 18290 -6730 18324 -754
rect 18448 -6730 18482 -754
rect 18606 -6730 18640 -754
rect 18764 -6730 18798 -754
rect 18922 -6730 18956 -754
rect 20482 -6730 20516 -754
rect 20640 -6730 20674 -754
rect 20798 -6730 20832 -754
rect 20956 -6730 20990 -754
rect 21114 -6730 21148 -754
rect 21272 -6730 21306 -754
rect 21430 -6730 21464 -754
rect 21588 -6730 21622 -754
rect 21746 -6730 21780 -754
rect 21904 -6730 21938 -754
rect 22062 -6730 22096 -754
rect 22220 -6730 22254 -754
rect 22378 -6730 22412 -754
rect 22536 -6730 22570 -754
rect 22694 -6730 22728 -754
rect 22852 -6730 22886 -754
rect 23010 -6730 23044 -754
rect 23168 -6730 23202 -754
rect 23326 -6730 23360 -754
rect 23484 -6730 23518 -754
rect 23642 -6730 23676 -754
rect 23800 -6730 23834 -754
rect 23958 -6730 23992 -754
rect 24116 -6730 24150 -754
rect 24274 -6730 24308 -754
rect 24432 -6730 24466 -754
rect 24590 -6730 24624 -754
rect 24748 -6730 24782 -754
rect 24906 -6730 24940 -754
rect 25064 -6730 25098 -754
rect 25222 -6730 25256 -754
<< mvpsubdiff >>
rect 1436 6468 6502 6480
rect 1436 6434 1544 6468
rect 6394 6434 6502 6468
rect 1436 6422 6502 6434
rect 1436 6372 1494 6422
rect 1436 144 1448 6372
rect 1482 144 1494 6372
rect 6444 6372 6502 6422
rect 1436 94 1494 144
rect 6444 144 6456 6372
rect 6490 144 6502 6372
rect 6444 94 6502 144
rect 1436 82 6502 94
rect 1436 48 1544 82
rect 6394 48 6502 82
rect 1436 36 6502 48
rect 7736 6468 12802 6480
rect 7736 6434 7844 6468
rect 12694 6434 12802 6468
rect 7736 6422 12802 6434
rect 7736 6372 7794 6422
rect 7736 144 7748 6372
rect 7782 144 7794 6372
rect 12744 6372 12802 6422
rect 7736 94 7794 144
rect 12744 144 12756 6372
rect 12790 144 12802 6372
rect 12744 94 12802 144
rect 7736 82 12802 94
rect 7736 48 7844 82
rect 12694 48 12802 82
rect 7736 36 12802 48
rect 14036 6468 19102 6480
rect 14036 6434 14144 6468
rect 18994 6434 19102 6468
rect 14036 6422 19102 6434
rect 14036 6372 14094 6422
rect 14036 144 14048 6372
rect 14082 144 14094 6372
rect 19044 6372 19102 6422
rect 14036 94 14094 144
rect 19044 144 19056 6372
rect 19090 144 19102 6372
rect 19044 94 19102 144
rect 14036 82 19102 94
rect 14036 48 14144 82
rect 18994 48 19102 82
rect 14036 36 19102 48
rect 20336 6468 25402 6480
rect 20336 6434 20444 6468
rect 25294 6434 25402 6468
rect 20336 6422 25402 6434
rect 20336 6372 20394 6422
rect 20336 144 20348 6372
rect 20382 144 20394 6372
rect 25344 6372 25402 6422
rect 20336 94 20394 144
rect 25344 144 25356 6372
rect 25390 144 25402 6372
rect 25344 94 25402 144
rect 20336 82 25402 94
rect 20336 48 20444 82
rect 25294 48 25402 82
rect 20336 36 25402 48
rect 1436 -532 6502 -520
rect 1436 -566 1544 -532
rect 6394 -566 6502 -532
rect 1436 -578 6502 -566
rect 1436 -628 1494 -578
rect 1436 -6856 1448 -628
rect 1482 -6856 1494 -628
rect 6444 -628 6502 -578
rect 1436 -6906 1494 -6856
rect 6444 -6856 6456 -628
rect 6490 -6856 6502 -628
rect 6444 -6906 6502 -6856
rect 1436 -6918 6502 -6906
rect 1436 -6952 1544 -6918
rect 6394 -6952 6502 -6918
rect 1436 -6964 6502 -6952
rect 7736 -532 12802 -520
rect 7736 -566 7844 -532
rect 12694 -566 12802 -532
rect 7736 -578 12802 -566
rect 7736 -628 7794 -578
rect 7736 -6856 7748 -628
rect 7782 -6856 7794 -628
rect 12744 -628 12802 -578
rect 7736 -6906 7794 -6856
rect 12744 -6856 12756 -628
rect 12790 -6856 12802 -628
rect 12744 -6906 12802 -6856
rect 7736 -6918 12802 -6906
rect 7736 -6952 7844 -6918
rect 12694 -6952 12802 -6918
rect 7736 -6964 12802 -6952
rect 14036 -532 19102 -520
rect 14036 -566 14144 -532
rect 18994 -566 19102 -532
rect 14036 -578 19102 -566
rect 14036 -628 14094 -578
rect 14036 -6856 14048 -628
rect 14082 -6856 14094 -628
rect 19044 -628 19102 -578
rect 14036 -6906 14094 -6856
rect 19044 -6856 19056 -628
rect 19090 -6856 19102 -628
rect 19044 -6906 19102 -6856
rect 14036 -6918 19102 -6906
rect 14036 -6952 14144 -6918
rect 18994 -6952 19102 -6918
rect 14036 -6964 19102 -6952
rect 20336 -532 25402 -520
rect 20336 -566 20444 -532
rect 25294 -566 25402 -532
rect 20336 -578 25402 -566
rect 20336 -628 20394 -578
rect 20336 -6856 20348 -628
rect 20382 -6856 20394 -628
rect 25344 -628 25402 -578
rect 20336 -6906 20394 -6856
rect 25344 -6856 25356 -628
rect 25390 -6856 25402 -628
rect 25344 -6906 25402 -6856
rect 20336 -6918 25402 -6906
rect 20336 -6952 20444 -6918
rect 25294 -6952 25402 -6918
rect 20336 -6964 25402 -6952
<< mvpsubdiffcont >>
rect 1544 6434 6394 6468
rect 1448 144 1482 6372
rect 6456 144 6490 6372
rect 1544 48 6394 82
rect 7844 6434 12694 6468
rect 7748 144 7782 6372
rect 12756 144 12790 6372
rect 7844 48 12694 82
rect 14144 6434 18994 6468
rect 14048 144 14082 6372
rect 19056 144 19090 6372
rect 14144 48 18994 82
rect 20444 6434 25294 6468
rect 20348 144 20382 6372
rect 25356 144 25390 6372
rect 20444 48 25294 82
rect 1544 -566 6394 -532
rect 1448 -6856 1482 -628
rect 6456 -6856 6490 -628
rect 1544 -6952 6394 -6918
rect 7844 -566 12694 -532
rect 7748 -6856 7782 -628
rect 12756 -6856 12790 -628
rect 7844 -6952 12694 -6918
rect 14144 -566 18994 -532
rect 14048 -6856 14082 -628
rect 19056 -6856 19090 -628
rect 14144 -6952 18994 -6918
rect 20444 -566 25294 -532
rect 20348 -6856 20382 -628
rect 25356 -6856 25390 -628
rect 20444 -6952 25294 -6918
<< poly >>
rect 1628 6330 1728 6346
rect 1628 6296 1644 6330
rect 1712 6296 1728 6330
rect 1628 6258 1728 6296
rect 1786 6330 1886 6346
rect 1786 6296 1802 6330
rect 1870 6296 1886 6330
rect 1786 6258 1886 6296
rect 1944 6330 2044 6346
rect 1944 6296 1960 6330
rect 2028 6296 2044 6330
rect 1944 6258 2044 6296
rect 2102 6330 2202 6346
rect 2102 6296 2118 6330
rect 2186 6296 2202 6330
rect 2102 6258 2202 6296
rect 2260 6330 2360 6346
rect 2260 6296 2276 6330
rect 2344 6296 2360 6330
rect 2260 6258 2360 6296
rect 2418 6330 2518 6346
rect 2418 6296 2434 6330
rect 2502 6296 2518 6330
rect 2418 6258 2518 6296
rect 2576 6330 2676 6346
rect 2576 6296 2592 6330
rect 2660 6296 2676 6330
rect 2576 6258 2676 6296
rect 2734 6330 2834 6346
rect 2734 6296 2750 6330
rect 2818 6296 2834 6330
rect 2734 6258 2834 6296
rect 2892 6330 2992 6346
rect 2892 6296 2908 6330
rect 2976 6296 2992 6330
rect 2892 6258 2992 6296
rect 3050 6330 3150 6346
rect 3050 6296 3066 6330
rect 3134 6296 3150 6330
rect 3050 6258 3150 6296
rect 3208 6330 3308 6346
rect 3208 6296 3224 6330
rect 3292 6296 3308 6330
rect 3208 6258 3308 6296
rect 3366 6330 3466 6346
rect 3366 6296 3382 6330
rect 3450 6296 3466 6330
rect 3366 6258 3466 6296
rect 3524 6330 3624 6346
rect 3524 6296 3540 6330
rect 3608 6296 3624 6330
rect 3524 6258 3624 6296
rect 3682 6330 3782 6346
rect 3682 6296 3698 6330
rect 3766 6296 3782 6330
rect 3682 6258 3782 6296
rect 3840 6330 3940 6346
rect 3840 6296 3856 6330
rect 3924 6296 3940 6330
rect 3840 6258 3940 6296
rect 3998 6330 4098 6346
rect 3998 6296 4014 6330
rect 4082 6296 4098 6330
rect 3998 6258 4098 6296
rect 4156 6330 4256 6346
rect 4156 6296 4172 6330
rect 4240 6296 4256 6330
rect 4156 6258 4256 6296
rect 4314 6330 4414 6346
rect 4314 6296 4330 6330
rect 4398 6296 4414 6330
rect 4314 6258 4414 6296
rect 4472 6330 4572 6346
rect 4472 6296 4488 6330
rect 4556 6296 4572 6330
rect 4472 6258 4572 6296
rect 4630 6330 4730 6346
rect 4630 6296 4646 6330
rect 4714 6296 4730 6330
rect 4630 6258 4730 6296
rect 4788 6330 4888 6346
rect 4788 6296 4804 6330
rect 4872 6296 4888 6330
rect 4788 6258 4888 6296
rect 4946 6330 5046 6346
rect 4946 6296 4962 6330
rect 5030 6296 5046 6330
rect 4946 6258 5046 6296
rect 5104 6330 5204 6346
rect 5104 6296 5120 6330
rect 5188 6296 5204 6330
rect 5104 6258 5204 6296
rect 5262 6330 5362 6346
rect 5262 6296 5278 6330
rect 5346 6296 5362 6330
rect 5262 6258 5362 6296
rect 5420 6330 5520 6346
rect 5420 6296 5436 6330
rect 5504 6296 5520 6330
rect 5420 6258 5520 6296
rect 5578 6330 5678 6346
rect 5578 6296 5594 6330
rect 5662 6296 5678 6330
rect 5578 6258 5678 6296
rect 5736 6330 5836 6346
rect 5736 6296 5752 6330
rect 5820 6296 5836 6330
rect 5736 6258 5836 6296
rect 5894 6330 5994 6346
rect 5894 6296 5910 6330
rect 5978 6296 5994 6330
rect 5894 6258 5994 6296
rect 6052 6330 6152 6346
rect 6052 6296 6068 6330
rect 6136 6296 6152 6330
rect 6052 6258 6152 6296
rect 6210 6330 6310 6346
rect 6210 6296 6226 6330
rect 6294 6296 6310 6330
rect 6210 6258 6310 6296
rect 1628 220 1728 258
rect 1628 186 1644 220
rect 1712 186 1728 220
rect 1628 170 1728 186
rect 1786 220 1886 258
rect 1786 186 1802 220
rect 1870 186 1886 220
rect 1786 170 1886 186
rect 1944 220 2044 258
rect 1944 186 1960 220
rect 2028 186 2044 220
rect 1944 170 2044 186
rect 2102 220 2202 258
rect 2102 186 2118 220
rect 2186 186 2202 220
rect 2102 170 2202 186
rect 2260 220 2360 258
rect 2260 186 2276 220
rect 2344 186 2360 220
rect 2260 170 2360 186
rect 2418 220 2518 258
rect 2418 186 2434 220
rect 2502 186 2518 220
rect 2418 170 2518 186
rect 2576 220 2676 258
rect 2576 186 2592 220
rect 2660 186 2676 220
rect 2576 170 2676 186
rect 2734 220 2834 258
rect 2734 186 2750 220
rect 2818 186 2834 220
rect 2734 170 2834 186
rect 2892 220 2992 258
rect 2892 186 2908 220
rect 2976 186 2992 220
rect 2892 170 2992 186
rect 3050 220 3150 258
rect 3050 186 3066 220
rect 3134 186 3150 220
rect 3050 170 3150 186
rect 3208 220 3308 258
rect 3208 186 3224 220
rect 3292 186 3308 220
rect 3208 170 3308 186
rect 3366 220 3466 258
rect 3366 186 3382 220
rect 3450 186 3466 220
rect 3366 170 3466 186
rect 3524 220 3624 258
rect 3524 186 3540 220
rect 3608 186 3624 220
rect 3524 170 3624 186
rect 3682 220 3782 258
rect 3682 186 3698 220
rect 3766 186 3782 220
rect 3682 170 3782 186
rect 3840 220 3940 258
rect 3840 186 3856 220
rect 3924 186 3940 220
rect 3840 170 3940 186
rect 3998 220 4098 258
rect 3998 186 4014 220
rect 4082 186 4098 220
rect 3998 170 4098 186
rect 4156 220 4256 258
rect 4156 186 4172 220
rect 4240 186 4256 220
rect 4156 170 4256 186
rect 4314 220 4414 258
rect 4314 186 4330 220
rect 4398 186 4414 220
rect 4314 170 4414 186
rect 4472 220 4572 258
rect 4472 186 4488 220
rect 4556 186 4572 220
rect 4472 170 4572 186
rect 4630 220 4730 258
rect 4630 186 4646 220
rect 4714 186 4730 220
rect 4630 170 4730 186
rect 4788 220 4888 258
rect 4788 186 4804 220
rect 4872 186 4888 220
rect 4788 170 4888 186
rect 4946 220 5046 258
rect 4946 186 4962 220
rect 5030 186 5046 220
rect 4946 170 5046 186
rect 5104 220 5204 258
rect 5104 186 5120 220
rect 5188 186 5204 220
rect 5104 170 5204 186
rect 5262 220 5362 258
rect 5262 186 5278 220
rect 5346 186 5362 220
rect 5262 170 5362 186
rect 5420 220 5520 258
rect 5420 186 5436 220
rect 5504 186 5520 220
rect 5420 170 5520 186
rect 5578 220 5678 258
rect 5578 186 5594 220
rect 5662 186 5678 220
rect 5578 170 5678 186
rect 5736 220 5836 258
rect 5736 186 5752 220
rect 5820 186 5836 220
rect 5736 170 5836 186
rect 5894 220 5994 258
rect 5894 186 5910 220
rect 5978 186 5994 220
rect 5894 170 5994 186
rect 6052 220 6152 258
rect 6052 186 6068 220
rect 6136 186 6152 220
rect 6052 170 6152 186
rect 6210 220 6310 258
rect 6210 186 6226 220
rect 6294 186 6310 220
rect 6210 170 6310 186
rect 7928 6330 8028 6346
rect 7928 6296 7944 6330
rect 8012 6296 8028 6330
rect 7928 6258 8028 6296
rect 8086 6330 8186 6346
rect 8086 6296 8102 6330
rect 8170 6296 8186 6330
rect 8086 6258 8186 6296
rect 8244 6330 8344 6346
rect 8244 6296 8260 6330
rect 8328 6296 8344 6330
rect 8244 6258 8344 6296
rect 8402 6330 8502 6346
rect 8402 6296 8418 6330
rect 8486 6296 8502 6330
rect 8402 6258 8502 6296
rect 8560 6330 8660 6346
rect 8560 6296 8576 6330
rect 8644 6296 8660 6330
rect 8560 6258 8660 6296
rect 8718 6330 8818 6346
rect 8718 6296 8734 6330
rect 8802 6296 8818 6330
rect 8718 6258 8818 6296
rect 8876 6330 8976 6346
rect 8876 6296 8892 6330
rect 8960 6296 8976 6330
rect 8876 6258 8976 6296
rect 9034 6330 9134 6346
rect 9034 6296 9050 6330
rect 9118 6296 9134 6330
rect 9034 6258 9134 6296
rect 9192 6330 9292 6346
rect 9192 6296 9208 6330
rect 9276 6296 9292 6330
rect 9192 6258 9292 6296
rect 9350 6330 9450 6346
rect 9350 6296 9366 6330
rect 9434 6296 9450 6330
rect 9350 6258 9450 6296
rect 9508 6330 9608 6346
rect 9508 6296 9524 6330
rect 9592 6296 9608 6330
rect 9508 6258 9608 6296
rect 9666 6330 9766 6346
rect 9666 6296 9682 6330
rect 9750 6296 9766 6330
rect 9666 6258 9766 6296
rect 9824 6330 9924 6346
rect 9824 6296 9840 6330
rect 9908 6296 9924 6330
rect 9824 6258 9924 6296
rect 9982 6330 10082 6346
rect 9982 6296 9998 6330
rect 10066 6296 10082 6330
rect 9982 6258 10082 6296
rect 10140 6330 10240 6346
rect 10140 6296 10156 6330
rect 10224 6296 10240 6330
rect 10140 6258 10240 6296
rect 10298 6330 10398 6346
rect 10298 6296 10314 6330
rect 10382 6296 10398 6330
rect 10298 6258 10398 6296
rect 10456 6330 10556 6346
rect 10456 6296 10472 6330
rect 10540 6296 10556 6330
rect 10456 6258 10556 6296
rect 10614 6330 10714 6346
rect 10614 6296 10630 6330
rect 10698 6296 10714 6330
rect 10614 6258 10714 6296
rect 10772 6330 10872 6346
rect 10772 6296 10788 6330
rect 10856 6296 10872 6330
rect 10772 6258 10872 6296
rect 10930 6330 11030 6346
rect 10930 6296 10946 6330
rect 11014 6296 11030 6330
rect 10930 6258 11030 6296
rect 11088 6330 11188 6346
rect 11088 6296 11104 6330
rect 11172 6296 11188 6330
rect 11088 6258 11188 6296
rect 11246 6330 11346 6346
rect 11246 6296 11262 6330
rect 11330 6296 11346 6330
rect 11246 6258 11346 6296
rect 11404 6330 11504 6346
rect 11404 6296 11420 6330
rect 11488 6296 11504 6330
rect 11404 6258 11504 6296
rect 11562 6330 11662 6346
rect 11562 6296 11578 6330
rect 11646 6296 11662 6330
rect 11562 6258 11662 6296
rect 11720 6330 11820 6346
rect 11720 6296 11736 6330
rect 11804 6296 11820 6330
rect 11720 6258 11820 6296
rect 11878 6330 11978 6346
rect 11878 6296 11894 6330
rect 11962 6296 11978 6330
rect 11878 6258 11978 6296
rect 12036 6330 12136 6346
rect 12036 6296 12052 6330
rect 12120 6296 12136 6330
rect 12036 6258 12136 6296
rect 12194 6330 12294 6346
rect 12194 6296 12210 6330
rect 12278 6296 12294 6330
rect 12194 6258 12294 6296
rect 12352 6330 12452 6346
rect 12352 6296 12368 6330
rect 12436 6296 12452 6330
rect 12352 6258 12452 6296
rect 12510 6330 12610 6346
rect 12510 6296 12526 6330
rect 12594 6296 12610 6330
rect 12510 6258 12610 6296
rect 7928 220 8028 258
rect 7928 186 7944 220
rect 8012 186 8028 220
rect 7928 170 8028 186
rect 8086 220 8186 258
rect 8086 186 8102 220
rect 8170 186 8186 220
rect 8086 170 8186 186
rect 8244 220 8344 258
rect 8244 186 8260 220
rect 8328 186 8344 220
rect 8244 170 8344 186
rect 8402 220 8502 258
rect 8402 186 8418 220
rect 8486 186 8502 220
rect 8402 170 8502 186
rect 8560 220 8660 258
rect 8560 186 8576 220
rect 8644 186 8660 220
rect 8560 170 8660 186
rect 8718 220 8818 258
rect 8718 186 8734 220
rect 8802 186 8818 220
rect 8718 170 8818 186
rect 8876 220 8976 258
rect 8876 186 8892 220
rect 8960 186 8976 220
rect 8876 170 8976 186
rect 9034 220 9134 258
rect 9034 186 9050 220
rect 9118 186 9134 220
rect 9034 170 9134 186
rect 9192 220 9292 258
rect 9192 186 9208 220
rect 9276 186 9292 220
rect 9192 170 9292 186
rect 9350 220 9450 258
rect 9350 186 9366 220
rect 9434 186 9450 220
rect 9350 170 9450 186
rect 9508 220 9608 258
rect 9508 186 9524 220
rect 9592 186 9608 220
rect 9508 170 9608 186
rect 9666 220 9766 258
rect 9666 186 9682 220
rect 9750 186 9766 220
rect 9666 170 9766 186
rect 9824 220 9924 258
rect 9824 186 9840 220
rect 9908 186 9924 220
rect 9824 170 9924 186
rect 9982 220 10082 258
rect 9982 186 9998 220
rect 10066 186 10082 220
rect 9982 170 10082 186
rect 10140 220 10240 258
rect 10140 186 10156 220
rect 10224 186 10240 220
rect 10140 170 10240 186
rect 10298 220 10398 258
rect 10298 186 10314 220
rect 10382 186 10398 220
rect 10298 170 10398 186
rect 10456 220 10556 258
rect 10456 186 10472 220
rect 10540 186 10556 220
rect 10456 170 10556 186
rect 10614 220 10714 258
rect 10614 186 10630 220
rect 10698 186 10714 220
rect 10614 170 10714 186
rect 10772 220 10872 258
rect 10772 186 10788 220
rect 10856 186 10872 220
rect 10772 170 10872 186
rect 10930 220 11030 258
rect 10930 186 10946 220
rect 11014 186 11030 220
rect 10930 170 11030 186
rect 11088 220 11188 258
rect 11088 186 11104 220
rect 11172 186 11188 220
rect 11088 170 11188 186
rect 11246 220 11346 258
rect 11246 186 11262 220
rect 11330 186 11346 220
rect 11246 170 11346 186
rect 11404 220 11504 258
rect 11404 186 11420 220
rect 11488 186 11504 220
rect 11404 170 11504 186
rect 11562 220 11662 258
rect 11562 186 11578 220
rect 11646 186 11662 220
rect 11562 170 11662 186
rect 11720 220 11820 258
rect 11720 186 11736 220
rect 11804 186 11820 220
rect 11720 170 11820 186
rect 11878 220 11978 258
rect 11878 186 11894 220
rect 11962 186 11978 220
rect 11878 170 11978 186
rect 12036 220 12136 258
rect 12036 186 12052 220
rect 12120 186 12136 220
rect 12036 170 12136 186
rect 12194 220 12294 258
rect 12194 186 12210 220
rect 12278 186 12294 220
rect 12194 170 12294 186
rect 12352 220 12452 258
rect 12352 186 12368 220
rect 12436 186 12452 220
rect 12352 170 12452 186
rect 12510 220 12610 258
rect 12510 186 12526 220
rect 12594 186 12610 220
rect 12510 170 12610 186
rect 14228 6330 14328 6346
rect 14228 6296 14244 6330
rect 14312 6296 14328 6330
rect 14228 6258 14328 6296
rect 14386 6330 14486 6346
rect 14386 6296 14402 6330
rect 14470 6296 14486 6330
rect 14386 6258 14486 6296
rect 14544 6330 14644 6346
rect 14544 6296 14560 6330
rect 14628 6296 14644 6330
rect 14544 6258 14644 6296
rect 14702 6330 14802 6346
rect 14702 6296 14718 6330
rect 14786 6296 14802 6330
rect 14702 6258 14802 6296
rect 14860 6330 14960 6346
rect 14860 6296 14876 6330
rect 14944 6296 14960 6330
rect 14860 6258 14960 6296
rect 15018 6330 15118 6346
rect 15018 6296 15034 6330
rect 15102 6296 15118 6330
rect 15018 6258 15118 6296
rect 15176 6330 15276 6346
rect 15176 6296 15192 6330
rect 15260 6296 15276 6330
rect 15176 6258 15276 6296
rect 15334 6330 15434 6346
rect 15334 6296 15350 6330
rect 15418 6296 15434 6330
rect 15334 6258 15434 6296
rect 15492 6330 15592 6346
rect 15492 6296 15508 6330
rect 15576 6296 15592 6330
rect 15492 6258 15592 6296
rect 15650 6330 15750 6346
rect 15650 6296 15666 6330
rect 15734 6296 15750 6330
rect 15650 6258 15750 6296
rect 15808 6330 15908 6346
rect 15808 6296 15824 6330
rect 15892 6296 15908 6330
rect 15808 6258 15908 6296
rect 15966 6330 16066 6346
rect 15966 6296 15982 6330
rect 16050 6296 16066 6330
rect 15966 6258 16066 6296
rect 16124 6330 16224 6346
rect 16124 6296 16140 6330
rect 16208 6296 16224 6330
rect 16124 6258 16224 6296
rect 16282 6330 16382 6346
rect 16282 6296 16298 6330
rect 16366 6296 16382 6330
rect 16282 6258 16382 6296
rect 16440 6330 16540 6346
rect 16440 6296 16456 6330
rect 16524 6296 16540 6330
rect 16440 6258 16540 6296
rect 16598 6330 16698 6346
rect 16598 6296 16614 6330
rect 16682 6296 16698 6330
rect 16598 6258 16698 6296
rect 16756 6330 16856 6346
rect 16756 6296 16772 6330
rect 16840 6296 16856 6330
rect 16756 6258 16856 6296
rect 16914 6330 17014 6346
rect 16914 6296 16930 6330
rect 16998 6296 17014 6330
rect 16914 6258 17014 6296
rect 17072 6330 17172 6346
rect 17072 6296 17088 6330
rect 17156 6296 17172 6330
rect 17072 6258 17172 6296
rect 17230 6330 17330 6346
rect 17230 6296 17246 6330
rect 17314 6296 17330 6330
rect 17230 6258 17330 6296
rect 17388 6330 17488 6346
rect 17388 6296 17404 6330
rect 17472 6296 17488 6330
rect 17388 6258 17488 6296
rect 17546 6330 17646 6346
rect 17546 6296 17562 6330
rect 17630 6296 17646 6330
rect 17546 6258 17646 6296
rect 17704 6330 17804 6346
rect 17704 6296 17720 6330
rect 17788 6296 17804 6330
rect 17704 6258 17804 6296
rect 17862 6330 17962 6346
rect 17862 6296 17878 6330
rect 17946 6296 17962 6330
rect 17862 6258 17962 6296
rect 18020 6330 18120 6346
rect 18020 6296 18036 6330
rect 18104 6296 18120 6330
rect 18020 6258 18120 6296
rect 18178 6330 18278 6346
rect 18178 6296 18194 6330
rect 18262 6296 18278 6330
rect 18178 6258 18278 6296
rect 18336 6330 18436 6346
rect 18336 6296 18352 6330
rect 18420 6296 18436 6330
rect 18336 6258 18436 6296
rect 18494 6330 18594 6346
rect 18494 6296 18510 6330
rect 18578 6296 18594 6330
rect 18494 6258 18594 6296
rect 18652 6330 18752 6346
rect 18652 6296 18668 6330
rect 18736 6296 18752 6330
rect 18652 6258 18752 6296
rect 18810 6330 18910 6346
rect 18810 6296 18826 6330
rect 18894 6296 18910 6330
rect 18810 6258 18910 6296
rect 14228 220 14328 258
rect 14228 186 14244 220
rect 14312 186 14328 220
rect 14228 170 14328 186
rect 14386 220 14486 258
rect 14386 186 14402 220
rect 14470 186 14486 220
rect 14386 170 14486 186
rect 14544 220 14644 258
rect 14544 186 14560 220
rect 14628 186 14644 220
rect 14544 170 14644 186
rect 14702 220 14802 258
rect 14702 186 14718 220
rect 14786 186 14802 220
rect 14702 170 14802 186
rect 14860 220 14960 258
rect 14860 186 14876 220
rect 14944 186 14960 220
rect 14860 170 14960 186
rect 15018 220 15118 258
rect 15018 186 15034 220
rect 15102 186 15118 220
rect 15018 170 15118 186
rect 15176 220 15276 258
rect 15176 186 15192 220
rect 15260 186 15276 220
rect 15176 170 15276 186
rect 15334 220 15434 258
rect 15334 186 15350 220
rect 15418 186 15434 220
rect 15334 170 15434 186
rect 15492 220 15592 258
rect 15492 186 15508 220
rect 15576 186 15592 220
rect 15492 170 15592 186
rect 15650 220 15750 258
rect 15650 186 15666 220
rect 15734 186 15750 220
rect 15650 170 15750 186
rect 15808 220 15908 258
rect 15808 186 15824 220
rect 15892 186 15908 220
rect 15808 170 15908 186
rect 15966 220 16066 258
rect 15966 186 15982 220
rect 16050 186 16066 220
rect 15966 170 16066 186
rect 16124 220 16224 258
rect 16124 186 16140 220
rect 16208 186 16224 220
rect 16124 170 16224 186
rect 16282 220 16382 258
rect 16282 186 16298 220
rect 16366 186 16382 220
rect 16282 170 16382 186
rect 16440 220 16540 258
rect 16440 186 16456 220
rect 16524 186 16540 220
rect 16440 170 16540 186
rect 16598 220 16698 258
rect 16598 186 16614 220
rect 16682 186 16698 220
rect 16598 170 16698 186
rect 16756 220 16856 258
rect 16756 186 16772 220
rect 16840 186 16856 220
rect 16756 170 16856 186
rect 16914 220 17014 258
rect 16914 186 16930 220
rect 16998 186 17014 220
rect 16914 170 17014 186
rect 17072 220 17172 258
rect 17072 186 17088 220
rect 17156 186 17172 220
rect 17072 170 17172 186
rect 17230 220 17330 258
rect 17230 186 17246 220
rect 17314 186 17330 220
rect 17230 170 17330 186
rect 17388 220 17488 258
rect 17388 186 17404 220
rect 17472 186 17488 220
rect 17388 170 17488 186
rect 17546 220 17646 258
rect 17546 186 17562 220
rect 17630 186 17646 220
rect 17546 170 17646 186
rect 17704 220 17804 258
rect 17704 186 17720 220
rect 17788 186 17804 220
rect 17704 170 17804 186
rect 17862 220 17962 258
rect 17862 186 17878 220
rect 17946 186 17962 220
rect 17862 170 17962 186
rect 18020 220 18120 258
rect 18020 186 18036 220
rect 18104 186 18120 220
rect 18020 170 18120 186
rect 18178 220 18278 258
rect 18178 186 18194 220
rect 18262 186 18278 220
rect 18178 170 18278 186
rect 18336 220 18436 258
rect 18336 186 18352 220
rect 18420 186 18436 220
rect 18336 170 18436 186
rect 18494 220 18594 258
rect 18494 186 18510 220
rect 18578 186 18594 220
rect 18494 170 18594 186
rect 18652 220 18752 258
rect 18652 186 18668 220
rect 18736 186 18752 220
rect 18652 170 18752 186
rect 18810 220 18910 258
rect 18810 186 18826 220
rect 18894 186 18910 220
rect 18810 170 18910 186
rect 20528 6330 20628 6346
rect 20528 6296 20544 6330
rect 20612 6296 20628 6330
rect 20528 6258 20628 6296
rect 20686 6330 20786 6346
rect 20686 6296 20702 6330
rect 20770 6296 20786 6330
rect 20686 6258 20786 6296
rect 20844 6330 20944 6346
rect 20844 6296 20860 6330
rect 20928 6296 20944 6330
rect 20844 6258 20944 6296
rect 21002 6330 21102 6346
rect 21002 6296 21018 6330
rect 21086 6296 21102 6330
rect 21002 6258 21102 6296
rect 21160 6330 21260 6346
rect 21160 6296 21176 6330
rect 21244 6296 21260 6330
rect 21160 6258 21260 6296
rect 21318 6330 21418 6346
rect 21318 6296 21334 6330
rect 21402 6296 21418 6330
rect 21318 6258 21418 6296
rect 21476 6330 21576 6346
rect 21476 6296 21492 6330
rect 21560 6296 21576 6330
rect 21476 6258 21576 6296
rect 21634 6330 21734 6346
rect 21634 6296 21650 6330
rect 21718 6296 21734 6330
rect 21634 6258 21734 6296
rect 21792 6330 21892 6346
rect 21792 6296 21808 6330
rect 21876 6296 21892 6330
rect 21792 6258 21892 6296
rect 21950 6330 22050 6346
rect 21950 6296 21966 6330
rect 22034 6296 22050 6330
rect 21950 6258 22050 6296
rect 22108 6330 22208 6346
rect 22108 6296 22124 6330
rect 22192 6296 22208 6330
rect 22108 6258 22208 6296
rect 22266 6330 22366 6346
rect 22266 6296 22282 6330
rect 22350 6296 22366 6330
rect 22266 6258 22366 6296
rect 22424 6330 22524 6346
rect 22424 6296 22440 6330
rect 22508 6296 22524 6330
rect 22424 6258 22524 6296
rect 22582 6330 22682 6346
rect 22582 6296 22598 6330
rect 22666 6296 22682 6330
rect 22582 6258 22682 6296
rect 22740 6330 22840 6346
rect 22740 6296 22756 6330
rect 22824 6296 22840 6330
rect 22740 6258 22840 6296
rect 22898 6330 22998 6346
rect 22898 6296 22914 6330
rect 22982 6296 22998 6330
rect 22898 6258 22998 6296
rect 23056 6330 23156 6346
rect 23056 6296 23072 6330
rect 23140 6296 23156 6330
rect 23056 6258 23156 6296
rect 23214 6330 23314 6346
rect 23214 6296 23230 6330
rect 23298 6296 23314 6330
rect 23214 6258 23314 6296
rect 23372 6330 23472 6346
rect 23372 6296 23388 6330
rect 23456 6296 23472 6330
rect 23372 6258 23472 6296
rect 23530 6330 23630 6346
rect 23530 6296 23546 6330
rect 23614 6296 23630 6330
rect 23530 6258 23630 6296
rect 23688 6330 23788 6346
rect 23688 6296 23704 6330
rect 23772 6296 23788 6330
rect 23688 6258 23788 6296
rect 23846 6330 23946 6346
rect 23846 6296 23862 6330
rect 23930 6296 23946 6330
rect 23846 6258 23946 6296
rect 24004 6330 24104 6346
rect 24004 6296 24020 6330
rect 24088 6296 24104 6330
rect 24004 6258 24104 6296
rect 24162 6330 24262 6346
rect 24162 6296 24178 6330
rect 24246 6296 24262 6330
rect 24162 6258 24262 6296
rect 24320 6330 24420 6346
rect 24320 6296 24336 6330
rect 24404 6296 24420 6330
rect 24320 6258 24420 6296
rect 24478 6330 24578 6346
rect 24478 6296 24494 6330
rect 24562 6296 24578 6330
rect 24478 6258 24578 6296
rect 24636 6330 24736 6346
rect 24636 6296 24652 6330
rect 24720 6296 24736 6330
rect 24636 6258 24736 6296
rect 24794 6330 24894 6346
rect 24794 6296 24810 6330
rect 24878 6296 24894 6330
rect 24794 6258 24894 6296
rect 24952 6330 25052 6346
rect 24952 6296 24968 6330
rect 25036 6296 25052 6330
rect 24952 6258 25052 6296
rect 25110 6330 25210 6346
rect 25110 6296 25126 6330
rect 25194 6296 25210 6330
rect 25110 6258 25210 6296
rect 20528 220 20628 258
rect 20528 186 20544 220
rect 20612 186 20628 220
rect 20528 170 20628 186
rect 20686 220 20786 258
rect 20686 186 20702 220
rect 20770 186 20786 220
rect 20686 170 20786 186
rect 20844 220 20944 258
rect 20844 186 20860 220
rect 20928 186 20944 220
rect 20844 170 20944 186
rect 21002 220 21102 258
rect 21002 186 21018 220
rect 21086 186 21102 220
rect 21002 170 21102 186
rect 21160 220 21260 258
rect 21160 186 21176 220
rect 21244 186 21260 220
rect 21160 170 21260 186
rect 21318 220 21418 258
rect 21318 186 21334 220
rect 21402 186 21418 220
rect 21318 170 21418 186
rect 21476 220 21576 258
rect 21476 186 21492 220
rect 21560 186 21576 220
rect 21476 170 21576 186
rect 21634 220 21734 258
rect 21634 186 21650 220
rect 21718 186 21734 220
rect 21634 170 21734 186
rect 21792 220 21892 258
rect 21792 186 21808 220
rect 21876 186 21892 220
rect 21792 170 21892 186
rect 21950 220 22050 258
rect 21950 186 21966 220
rect 22034 186 22050 220
rect 21950 170 22050 186
rect 22108 220 22208 258
rect 22108 186 22124 220
rect 22192 186 22208 220
rect 22108 170 22208 186
rect 22266 220 22366 258
rect 22266 186 22282 220
rect 22350 186 22366 220
rect 22266 170 22366 186
rect 22424 220 22524 258
rect 22424 186 22440 220
rect 22508 186 22524 220
rect 22424 170 22524 186
rect 22582 220 22682 258
rect 22582 186 22598 220
rect 22666 186 22682 220
rect 22582 170 22682 186
rect 22740 220 22840 258
rect 22740 186 22756 220
rect 22824 186 22840 220
rect 22740 170 22840 186
rect 22898 220 22998 258
rect 22898 186 22914 220
rect 22982 186 22998 220
rect 22898 170 22998 186
rect 23056 220 23156 258
rect 23056 186 23072 220
rect 23140 186 23156 220
rect 23056 170 23156 186
rect 23214 220 23314 258
rect 23214 186 23230 220
rect 23298 186 23314 220
rect 23214 170 23314 186
rect 23372 220 23472 258
rect 23372 186 23388 220
rect 23456 186 23472 220
rect 23372 170 23472 186
rect 23530 220 23630 258
rect 23530 186 23546 220
rect 23614 186 23630 220
rect 23530 170 23630 186
rect 23688 220 23788 258
rect 23688 186 23704 220
rect 23772 186 23788 220
rect 23688 170 23788 186
rect 23846 220 23946 258
rect 23846 186 23862 220
rect 23930 186 23946 220
rect 23846 170 23946 186
rect 24004 220 24104 258
rect 24004 186 24020 220
rect 24088 186 24104 220
rect 24004 170 24104 186
rect 24162 220 24262 258
rect 24162 186 24178 220
rect 24246 186 24262 220
rect 24162 170 24262 186
rect 24320 220 24420 258
rect 24320 186 24336 220
rect 24404 186 24420 220
rect 24320 170 24420 186
rect 24478 220 24578 258
rect 24478 186 24494 220
rect 24562 186 24578 220
rect 24478 170 24578 186
rect 24636 220 24736 258
rect 24636 186 24652 220
rect 24720 186 24736 220
rect 24636 170 24736 186
rect 24794 220 24894 258
rect 24794 186 24810 220
rect 24878 186 24894 220
rect 24794 170 24894 186
rect 24952 220 25052 258
rect 24952 186 24968 220
rect 25036 186 25052 220
rect 24952 170 25052 186
rect 25110 220 25210 258
rect 25110 186 25126 220
rect 25194 186 25210 220
rect 25110 170 25210 186
rect 1628 -670 1728 -654
rect 1628 -704 1644 -670
rect 1712 -704 1728 -670
rect 1628 -742 1728 -704
rect 1786 -670 1886 -654
rect 1786 -704 1802 -670
rect 1870 -704 1886 -670
rect 1786 -742 1886 -704
rect 1944 -670 2044 -654
rect 1944 -704 1960 -670
rect 2028 -704 2044 -670
rect 1944 -742 2044 -704
rect 2102 -670 2202 -654
rect 2102 -704 2118 -670
rect 2186 -704 2202 -670
rect 2102 -742 2202 -704
rect 2260 -670 2360 -654
rect 2260 -704 2276 -670
rect 2344 -704 2360 -670
rect 2260 -742 2360 -704
rect 2418 -670 2518 -654
rect 2418 -704 2434 -670
rect 2502 -704 2518 -670
rect 2418 -742 2518 -704
rect 2576 -670 2676 -654
rect 2576 -704 2592 -670
rect 2660 -704 2676 -670
rect 2576 -742 2676 -704
rect 2734 -670 2834 -654
rect 2734 -704 2750 -670
rect 2818 -704 2834 -670
rect 2734 -742 2834 -704
rect 2892 -670 2992 -654
rect 2892 -704 2908 -670
rect 2976 -704 2992 -670
rect 2892 -742 2992 -704
rect 3050 -670 3150 -654
rect 3050 -704 3066 -670
rect 3134 -704 3150 -670
rect 3050 -742 3150 -704
rect 3208 -670 3308 -654
rect 3208 -704 3224 -670
rect 3292 -704 3308 -670
rect 3208 -742 3308 -704
rect 3366 -670 3466 -654
rect 3366 -704 3382 -670
rect 3450 -704 3466 -670
rect 3366 -742 3466 -704
rect 3524 -670 3624 -654
rect 3524 -704 3540 -670
rect 3608 -704 3624 -670
rect 3524 -742 3624 -704
rect 3682 -670 3782 -654
rect 3682 -704 3698 -670
rect 3766 -704 3782 -670
rect 3682 -742 3782 -704
rect 3840 -670 3940 -654
rect 3840 -704 3856 -670
rect 3924 -704 3940 -670
rect 3840 -742 3940 -704
rect 3998 -670 4098 -654
rect 3998 -704 4014 -670
rect 4082 -704 4098 -670
rect 3998 -742 4098 -704
rect 4156 -670 4256 -654
rect 4156 -704 4172 -670
rect 4240 -704 4256 -670
rect 4156 -742 4256 -704
rect 4314 -670 4414 -654
rect 4314 -704 4330 -670
rect 4398 -704 4414 -670
rect 4314 -742 4414 -704
rect 4472 -670 4572 -654
rect 4472 -704 4488 -670
rect 4556 -704 4572 -670
rect 4472 -742 4572 -704
rect 4630 -670 4730 -654
rect 4630 -704 4646 -670
rect 4714 -704 4730 -670
rect 4630 -742 4730 -704
rect 4788 -670 4888 -654
rect 4788 -704 4804 -670
rect 4872 -704 4888 -670
rect 4788 -742 4888 -704
rect 4946 -670 5046 -654
rect 4946 -704 4962 -670
rect 5030 -704 5046 -670
rect 4946 -742 5046 -704
rect 5104 -670 5204 -654
rect 5104 -704 5120 -670
rect 5188 -704 5204 -670
rect 5104 -742 5204 -704
rect 5262 -670 5362 -654
rect 5262 -704 5278 -670
rect 5346 -704 5362 -670
rect 5262 -742 5362 -704
rect 5420 -670 5520 -654
rect 5420 -704 5436 -670
rect 5504 -704 5520 -670
rect 5420 -742 5520 -704
rect 5578 -670 5678 -654
rect 5578 -704 5594 -670
rect 5662 -704 5678 -670
rect 5578 -742 5678 -704
rect 5736 -670 5836 -654
rect 5736 -704 5752 -670
rect 5820 -704 5836 -670
rect 5736 -742 5836 -704
rect 5894 -670 5994 -654
rect 5894 -704 5910 -670
rect 5978 -704 5994 -670
rect 5894 -742 5994 -704
rect 6052 -670 6152 -654
rect 6052 -704 6068 -670
rect 6136 -704 6152 -670
rect 6052 -742 6152 -704
rect 6210 -670 6310 -654
rect 6210 -704 6226 -670
rect 6294 -704 6310 -670
rect 6210 -742 6310 -704
rect 1628 -6780 1728 -6742
rect 1628 -6814 1644 -6780
rect 1712 -6814 1728 -6780
rect 1628 -6830 1728 -6814
rect 1786 -6780 1886 -6742
rect 1786 -6814 1802 -6780
rect 1870 -6814 1886 -6780
rect 1786 -6830 1886 -6814
rect 1944 -6780 2044 -6742
rect 1944 -6814 1960 -6780
rect 2028 -6814 2044 -6780
rect 1944 -6830 2044 -6814
rect 2102 -6780 2202 -6742
rect 2102 -6814 2118 -6780
rect 2186 -6814 2202 -6780
rect 2102 -6830 2202 -6814
rect 2260 -6780 2360 -6742
rect 2260 -6814 2276 -6780
rect 2344 -6814 2360 -6780
rect 2260 -6830 2360 -6814
rect 2418 -6780 2518 -6742
rect 2418 -6814 2434 -6780
rect 2502 -6814 2518 -6780
rect 2418 -6830 2518 -6814
rect 2576 -6780 2676 -6742
rect 2576 -6814 2592 -6780
rect 2660 -6814 2676 -6780
rect 2576 -6830 2676 -6814
rect 2734 -6780 2834 -6742
rect 2734 -6814 2750 -6780
rect 2818 -6814 2834 -6780
rect 2734 -6830 2834 -6814
rect 2892 -6780 2992 -6742
rect 2892 -6814 2908 -6780
rect 2976 -6814 2992 -6780
rect 2892 -6830 2992 -6814
rect 3050 -6780 3150 -6742
rect 3050 -6814 3066 -6780
rect 3134 -6814 3150 -6780
rect 3050 -6830 3150 -6814
rect 3208 -6780 3308 -6742
rect 3208 -6814 3224 -6780
rect 3292 -6814 3308 -6780
rect 3208 -6830 3308 -6814
rect 3366 -6780 3466 -6742
rect 3366 -6814 3382 -6780
rect 3450 -6814 3466 -6780
rect 3366 -6830 3466 -6814
rect 3524 -6780 3624 -6742
rect 3524 -6814 3540 -6780
rect 3608 -6814 3624 -6780
rect 3524 -6830 3624 -6814
rect 3682 -6780 3782 -6742
rect 3682 -6814 3698 -6780
rect 3766 -6814 3782 -6780
rect 3682 -6830 3782 -6814
rect 3840 -6780 3940 -6742
rect 3840 -6814 3856 -6780
rect 3924 -6814 3940 -6780
rect 3840 -6830 3940 -6814
rect 3998 -6780 4098 -6742
rect 3998 -6814 4014 -6780
rect 4082 -6814 4098 -6780
rect 3998 -6830 4098 -6814
rect 4156 -6780 4256 -6742
rect 4156 -6814 4172 -6780
rect 4240 -6814 4256 -6780
rect 4156 -6830 4256 -6814
rect 4314 -6780 4414 -6742
rect 4314 -6814 4330 -6780
rect 4398 -6814 4414 -6780
rect 4314 -6830 4414 -6814
rect 4472 -6780 4572 -6742
rect 4472 -6814 4488 -6780
rect 4556 -6814 4572 -6780
rect 4472 -6830 4572 -6814
rect 4630 -6780 4730 -6742
rect 4630 -6814 4646 -6780
rect 4714 -6814 4730 -6780
rect 4630 -6830 4730 -6814
rect 4788 -6780 4888 -6742
rect 4788 -6814 4804 -6780
rect 4872 -6814 4888 -6780
rect 4788 -6830 4888 -6814
rect 4946 -6780 5046 -6742
rect 4946 -6814 4962 -6780
rect 5030 -6814 5046 -6780
rect 4946 -6830 5046 -6814
rect 5104 -6780 5204 -6742
rect 5104 -6814 5120 -6780
rect 5188 -6814 5204 -6780
rect 5104 -6830 5204 -6814
rect 5262 -6780 5362 -6742
rect 5262 -6814 5278 -6780
rect 5346 -6814 5362 -6780
rect 5262 -6830 5362 -6814
rect 5420 -6780 5520 -6742
rect 5420 -6814 5436 -6780
rect 5504 -6814 5520 -6780
rect 5420 -6830 5520 -6814
rect 5578 -6780 5678 -6742
rect 5578 -6814 5594 -6780
rect 5662 -6814 5678 -6780
rect 5578 -6830 5678 -6814
rect 5736 -6780 5836 -6742
rect 5736 -6814 5752 -6780
rect 5820 -6814 5836 -6780
rect 5736 -6830 5836 -6814
rect 5894 -6780 5994 -6742
rect 5894 -6814 5910 -6780
rect 5978 -6814 5994 -6780
rect 5894 -6830 5994 -6814
rect 6052 -6780 6152 -6742
rect 6052 -6814 6068 -6780
rect 6136 -6814 6152 -6780
rect 6052 -6830 6152 -6814
rect 6210 -6780 6310 -6742
rect 6210 -6814 6226 -6780
rect 6294 -6814 6310 -6780
rect 6210 -6830 6310 -6814
rect 7928 -670 8028 -654
rect 7928 -704 7944 -670
rect 8012 -704 8028 -670
rect 7928 -742 8028 -704
rect 8086 -670 8186 -654
rect 8086 -704 8102 -670
rect 8170 -704 8186 -670
rect 8086 -742 8186 -704
rect 8244 -670 8344 -654
rect 8244 -704 8260 -670
rect 8328 -704 8344 -670
rect 8244 -742 8344 -704
rect 8402 -670 8502 -654
rect 8402 -704 8418 -670
rect 8486 -704 8502 -670
rect 8402 -742 8502 -704
rect 8560 -670 8660 -654
rect 8560 -704 8576 -670
rect 8644 -704 8660 -670
rect 8560 -742 8660 -704
rect 8718 -670 8818 -654
rect 8718 -704 8734 -670
rect 8802 -704 8818 -670
rect 8718 -742 8818 -704
rect 8876 -670 8976 -654
rect 8876 -704 8892 -670
rect 8960 -704 8976 -670
rect 8876 -742 8976 -704
rect 9034 -670 9134 -654
rect 9034 -704 9050 -670
rect 9118 -704 9134 -670
rect 9034 -742 9134 -704
rect 9192 -670 9292 -654
rect 9192 -704 9208 -670
rect 9276 -704 9292 -670
rect 9192 -742 9292 -704
rect 9350 -670 9450 -654
rect 9350 -704 9366 -670
rect 9434 -704 9450 -670
rect 9350 -742 9450 -704
rect 9508 -670 9608 -654
rect 9508 -704 9524 -670
rect 9592 -704 9608 -670
rect 9508 -742 9608 -704
rect 9666 -670 9766 -654
rect 9666 -704 9682 -670
rect 9750 -704 9766 -670
rect 9666 -742 9766 -704
rect 9824 -670 9924 -654
rect 9824 -704 9840 -670
rect 9908 -704 9924 -670
rect 9824 -742 9924 -704
rect 9982 -670 10082 -654
rect 9982 -704 9998 -670
rect 10066 -704 10082 -670
rect 9982 -742 10082 -704
rect 10140 -670 10240 -654
rect 10140 -704 10156 -670
rect 10224 -704 10240 -670
rect 10140 -742 10240 -704
rect 10298 -670 10398 -654
rect 10298 -704 10314 -670
rect 10382 -704 10398 -670
rect 10298 -742 10398 -704
rect 10456 -670 10556 -654
rect 10456 -704 10472 -670
rect 10540 -704 10556 -670
rect 10456 -742 10556 -704
rect 10614 -670 10714 -654
rect 10614 -704 10630 -670
rect 10698 -704 10714 -670
rect 10614 -742 10714 -704
rect 10772 -670 10872 -654
rect 10772 -704 10788 -670
rect 10856 -704 10872 -670
rect 10772 -742 10872 -704
rect 10930 -670 11030 -654
rect 10930 -704 10946 -670
rect 11014 -704 11030 -670
rect 10930 -742 11030 -704
rect 11088 -670 11188 -654
rect 11088 -704 11104 -670
rect 11172 -704 11188 -670
rect 11088 -742 11188 -704
rect 11246 -670 11346 -654
rect 11246 -704 11262 -670
rect 11330 -704 11346 -670
rect 11246 -742 11346 -704
rect 11404 -670 11504 -654
rect 11404 -704 11420 -670
rect 11488 -704 11504 -670
rect 11404 -742 11504 -704
rect 11562 -670 11662 -654
rect 11562 -704 11578 -670
rect 11646 -704 11662 -670
rect 11562 -742 11662 -704
rect 11720 -670 11820 -654
rect 11720 -704 11736 -670
rect 11804 -704 11820 -670
rect 11720 -742 11820 -704
rect 11878 -670 11978 -654
rect 11878 -704 11894 -670
rect 11962 -704 11978 -670
rect 11878 -742 11978 -704
rect 12036 -670 12136 -654
rect 12036 -704 12052 -670
rect 12120 -704 12136 -670
rect 12036 -742 12136 -704
rect 12194 -670 12294 -654
rect 12194 -704 12210 -670
rect 12278 -704 12294 -670
rect 12194 -742 12294 -704
rect 12352 -670 12452 -654
rect 12352 -704 12368 -670
rect 12436 -704 12452 -670
rect 12352 -742 12452 -704
rect 12510 -670 12610 -654
rect 12510 -704 12526 -670
rect 12594 -704 12610 -670
rect 12510 -742 12610 -704
rect 7928 -6780 8028 -6742
rect 7928 -6814 7944 -6780
rect 8012 -6814 8028 -6780
rect 7928 -6830 8028 -6814
rect 8086 -6780 8186 -6742
rect 8086 -6814 8102 -6780
rect 8170 -6814 8186 -6780
rect 8086 -6830 8186 -6814
rect 8244 -6780 8344 -6742
rect 8244 -6814 8260 -6780
rect 8328 -6814 8344 -6780
rect 8244 -6830 8344 -6814
rect 8402 -6780 8502 -6742
rect 8402 -6814 8418 -6780
rect 8486 -6814 8502 -6780
rect 8402 -6830 8502 -6814
rect 8560 -6780 8660 -6742
rect 8560 -6814 8576 -6780
rect 8644 -6814 8660 -6780
rect 8560 -6830 8660 -6814
rect 8718 -6780 8818 -6742
rect 8718 -6814 8734 -6780
rect 8802 -6814 8818 -6780
rect 8718 -6830 8818 -6814
rect 8876 -6780 8976 -6742
rect 8876 -6814 8892 -6780
rect 8960 -6814 8976 -6780
rect 8876 -6830 8976 -6814
rect 9034 -6780 9134 -6742
rect 9034 -6814 9050 -6780
rect 9118 -6814 9134 -6780
rect 9034 -6830 9134 -6814
rect 9192 -6780 9292 -6742
rect 9192 -6814 9208 -6780
rect 9276 -6814 9292 -6780
rect 9192 -6830 9292 -6814
rect 9350 -6780 9450 -6742
rect 9350 -6814 9366 -6780
rect 9434 -6814 9450 -6780
rect 9350 -6830 9450 -6814
rect 9508 -6780 9608 -6742
rect 9508 -6814 9524 -6780
rect 9592 -6814 9608 -6780
rect 9508 -6830 9608 -6814
rect 9666 -6780 9766 -6742
rect 9666 -6814 9682 -6780
rect 9750 -6814 9766 -6780
rect 9666 -6830 9766 -6814
rect 9824 -6780 9924 -6742
rect 9824 -6814 9840 -6780
rect 9908 -6814 9924 -6780
rect 9824 -6830 9924 -6814
rect 9982 -6780 10082 -6742
rect 9982 -6814 9998 -6780
rect 10066 -6814 10082 -6780
rect 9982 -6830 10082 -6814
rect 10140 -6780 10240 -6742
rect 10140 -6814 10156 -6780
rect 10224 -6814 10240 -6780
rect 10140 -6830 10240 -6814
rect 10298 -6780 10398 -6742
rect 10298 -6814 10314 -6780
rect 10382 -6814 10398 -6780
rect 10298 -6830 10398 -6814
rect 10456 -6780 10556 -6742
rect 10456 -6814 10472 -6780
rect 10540 -6814 10556 -6780
rect 10456 -6830 10556 -6814
rect 10614 -6780 10714 -6742
rect 10614 -6814 10630 -6780
rect 10698 -6814 10714 -6780
rect 10614 -6830 10714 -6814
rect 10772 -6780 10872 -6742
rect 10772 -6814 10788 -6780
rect 10856 -6814 10872 -6780
rect 10772 -6830 10872 -6814
rect 10930 -6780 11030 -6742
rect 10930 -6814 10946 -6780
rect 11014 -6814 11030 -6780
rect 10930 -6830 11030 -6814
rect 11088 -6780 11188 -6742
rect 11088 -6814 11104 -6780
rect 11172 -6814 11188 -6780
rect 11088 -6830 11188 -6814
rect 11246 -6780 11346 -6742
rect 11246 -6814 11262 -6780
rect 11330 -6814 11346 -6780
rect 11246 -6830 11346 -6814
rect 11404 -6780 11504 -6742
rect 11404 -6814 11420 -6780
rect 11488 -6814 11504 -6780
rect 11404 -6830 11504 -6814
rect 11562 -6780 11662 -6742
rect 11562 -6814 11578 -6780
rect 11646 -6814 11662 -6780
rect 11562 -6830 11662 -6814
rect 11720 -6780 11820 -6742
rect 11720 -6814 11736 -6780
rect 11804 -6814 11820 -6780
rect 11720 -6830 11820 -6814
rect 11878 -6780 11978 -6742
rect 11878 -6814 11894 -6780
rect 11962 -6814 11978 -6780
rect 11878 -6830 11978 -6814
rect 12036 -6780 12136 -6742
rect 12036 -6814 12052 -6780
rect 12120 -6814 12136 -6780
rect 12036 -6830 12136 -6814
rect 12194 -6780 12294 -6742
rect 12194 -6814 12210 -6780
rect 12278 -6814 12294 -6780
rect 12194 -6830 12294 -6814
rect 12352 -6780 12452 -6742
rect 12352 -6814 12368 -6780
rect 12436 -6814 12452 -6780
rect 12352 -6830 12452 -6814
rect 12510 -6780 12610 -6742
rect 12510 -6814 12526 -6780
rect 12594 -6814 12610 -6780
rect 12510 -6830 12610 -6814
rect 14228 -670 14328 -654
rect 14228 -704 14244 -670
rect 14312 -704 14328 -670
rect 14228 -742 14328 -704
rect 14386 -670 14486 -654
rect 14386 -704 14402 -670
rect 14470 -704 14486 -670
rect 14386 -742 14486 -704
rect 14544 -670 14644 -654
rect 14544 -704 14560 -670
rect 14628 -704 14644 -670
rect 14544 -742 14644 -704
rect 14702 -670 14802 -654
rect 14702 -704 14718 -670
rect 14786 -704 14802 -670
rect 14702 -742 14802 -704
rect 14860 -670 14960 -654
rect 14860 -704 14876 -670
rect 14944 -704 14960 -670
rect 14860 -742 14960 -704
rect 15018 -670 15118 -654
rect 15018 -704 15034 -670
rect 15102 -704 15118 -670
rect 15018 -742 15118 -704
rect 15176 -670 15276 -654
rect 15176 -704 15192 -670
rect 15260 -704 15276 -670
rect 15176 -742 15276 -704
rect 15334 -670 15434 -654
rect 15334 -704 15350 -670
rect 15418 -704 15434 -670
rect 15334 -742 15434 -704
rect 15492 -670 15592 -654
rect 15492 -704 15508 -670
rect 15576 -704 15592 -670
rect 15492 -742 15592 -704
rect 15650 -670 15750 -654
rect 15650 -704 15666 -670
rect 15734 -704 15750 -670
rect 15650 -742 15750 -704
rect 15808 -670 15908 -654
rect 15808 -704 15824 -670
rect 15892 -704 15908 -670
rect 15808 -742 15908 -704
rect 15966 -670 16066 -654
rect 15966 -704 15982 -670
rect 16050 -704 16066 -670
rect 15966 -742 16066 -704
rect 16124 -670 16224 -654
rect 16124 -704 16140 -670
rect 16208 -704 16224 -670
rect 16124 -742 16224 -704
rect 16282 -670 16382 -654
rect 16282 -704 16298 -670
rect 16366 -704 16382 -670
rect 16282 -742 16382 -704
rect 16440 -670 16540 -654
rect 16440 -704 16456 -670
rect 16524 -704 16540 -670
rect 16440 -742 16540 -704
rect 16598 -670 16698 -654
rect 16598 -704 16614 -670
rect 16682 -704 16698 -670
rect 16598 -742 16698 -704
rect 16756 -670 16856 -654
rect 16756 -704 16772 -670
rect 16840 -704 16856 -670
rect 16756 -742 16856 -704
rect 16914 -670 17014 -654
rect 16914 -704 16930 -670
rect 16998 -704 17014 -670
rect 16914 -742 17014 -704
rect 17072 -670 17172 -654
rect 17072 -704 17088 -670
rect 17156 -704 17172 -670
rect 17072 -742 17172 -704
rect 17230 -670 17330 -654
rect 17230 -704 17246 -670
rect 17314 -704 17330 -670
rect 17230 -742 17330 -704
rect 17388 -670 17488 -654
rect 17388 -704 17404 -670
rect 17472 -704 17488 -670
rect 17388 -742 17488 -704
rect 17546 -670 17646 -654
rect 17546 -704 17562 -670
rect 17630 -704 17646 -670
rect 17546 -742 17646 -704
rect 17704 -670 17804 -654
rect 17704 -704 17720 -670
rect 17788 -704 17804 -670
rect 17704 -742 17804 -704
rect 17862 -670 17962 -654
rect 17862 -704 17878 -670
rect 17946 -704 17962 -670
rect 17862 -742 17962 -704
rect 18020 -670 18120 -654
rect 18020 -704 18036 -670
rect 18104 -704 18120 -670
rect 18020 -742 18120 -704
rect 18178 -670 18278 -654
rect 18178 -704 18194 -670
rect 18262 -704 18278 -670
rect 18178 -742 18278 -704
rect 18336 -670 18436 -654
rect 18336 -704 18352 -670
rect 18420 -704 18436 -670
rect 18336 -742 18436 -704
rect 18494 -670 18594 -654
rect 18494 -704 18510 -670
rect 18578 -704 18594 -670
rect 18494 -742 18594 -704
rect 18652 -670 18752 -654
rect 18652 -704 18668 -670
rect 18736 -704 18752 -670
rect 18652 -742 18752 -704
rect 18810 -670 18910 -654
rect 18810 -704 18826 -670
rect 18894 -704 18910 -670
rect 18810 -742 18910 -704
rect 14228 -6780 14328 -6742
rect 14228 -6814 14244 -6780
rect 14312 -6814 14328 -6780
rect 14228 -6830 14328 -6814
rect 14386 -6780 14486 -6742
rect 14386 -6814 14402 -6780
rect 14470 -6814 14486 -6780
rect 14386 -6830 14486 -6814
rect 14544 -6780 14644 -6742
rect 14544 -6814 14560 -6780
rect 14628 -6814 14644 -6780
rect 14544 -6830 14644 -6814
rect 14702 -6780 14802 -6742
rect 14702 -6814 14718 -6780
rect 14786 -6814 14802 -6780
rect 14702 -6830 14802 -6814
rect 14860 -6780 14960 -6742
rect 14860 -6814 14876 -6780
rect 14944 -6814 14960 -6780
rect 14860 -6830 14960 -6814
rect 15018 -6780 15118 -6742
rect 15018 -6814 15034 -6780
rect 15102 -6814 15118 -6780
rect 15018 -6830 15118 -6814
rect 15176 -6780 15276 -6742
rect 15176 -6814 15192 -6780
rect 15260 -6814 15276 -6780
rect 15176 -6830 15276 -6814
rect 15334 -6780 15434 -6742
rect 15334 -6814 15350 -6780
rect 15418 -6814 15434 -6780
rect 15334 -6830 15434 -6814
rect 15492 -6780 15592 -6742
rect 15492 -6814 15508 -6780
rect 15576 -6814 15592 -6780
rect 15492 -6830 15592 -6814
rect 15650 -6780 15750 -6742
rect 15650 -6814 15666 -6780
rect 15734 -6814 15750 -6780
rect 15650 -6830 15750 -6814
rect 15808 -6780 15908 -6742
rect 15808 -6814 15824 -6780
rect 15892 -6814 15908 -6780
rect 15808 -6830 15908 -6814
rect 15966 -6780 16066 -6742
rect 15966 -6814 15982 -6780
rect 16050 -6814 16066 -6780
rect 15966 -6830 16066 -6814
rect 16124 -6780 16224 -6742
rect 16124 -6814 16140 -6780
rect 16208 -6814 16224 -6780
rect 16124 -6830 16224 -6814
rect 16282 -6780 16382 -6742
rect 16282 -6814 16298 -6780
rect 16366 -6814 16382 -6780
rect 16282 -6830 16382 -6814
rect 16440 -6780 16540 -6742
rect 16440 -6814 16456 -6780
rect 16524 -6814 16540 -6780
rect 16440 -6830 16540 -6814
rect 16598 -6780 16698 -6742
rect 16598 -6814 16614 -6780
rect 16682 -6814 16698 -6780
rect 16598 -6830 16698 -6814
rect 16756 -6780 16856 -6742
rect 16756 -6814 16772 -6780
rect 16840 -6814 16856 -6780
rect 16756 -6830 16856 -6814
rect 16914 -6780 17014 -6742
rect 16914 -6814 16930 -6780
rect 16998 -6814 17014 -6780
rect 16914 -6830 17014 -6814
rect 17072 -6780 17172 -6742
rect 17072 -6814 17088 -6780
rect 17156 -6814 17172 -6780
rect 17072 -6830 17172 -6814
rect 17230 -6780 17330 -6742
rect 17230 -6814 17246 -6780
rect 17314 -6814 17330 -6780
rect 17230 -6830 17330 -6814
rect 17388 -6780 17488 -6742
rect 17388 -6814 17404 -6780
rect 17472 -6814 17488 -6780
rect 17388 -6830 17488 -6814
rect 17546 -6780 17646 -6742
rect 17546 -6814 17562 -6780
rect 17630 -6814 17646 -6780
rect 17546 -6830 17646 -6814
rect 17704 -6780 17804 -6742
rect 17704 -6814 17720 -6780
rect 17788 -6814 17804 -6780
rect 17704 -6830 17804 -6814
rect 17862 -6780 17962 -6742
rect 17862 -6814 17878 -6780
rect 17946 -6814 17962 -6780
rect 17862 -6830 17962 -6814
rect 18020 -6780 18120 -6742
rect 18020 -6814 18036 -6780
rect 18104 -6814 18120 -6780
rect 18020 -6830 18120 -6814
rect 18178 -6780 18278 -6742
rect 18178 -6814 18194 -6780
rect 18262 -6814 18278 -6780
rect 18178 -6830 18278 -6814
rect 18336 -6780 18436 -6742
rect 18336 -6814 18352 -6780
rect 18420 -6814 18436 -6780
rect 18336 -6830 18436 -6814
rect 18494 -6780 18594 -6742
rect 18494 -6814 18510 -6780
rect 18578 -6814 18594 -6780
rect 18494 -6830 18594 -6814
rect 18652 -6780 18752 -6742
rect 18652 -6814 18668 -6780
rect 18736 -6814 18752 -6780
rect 18652 -6830 18752 -6814
rect 18810 -6780 18910 -6742
rect 18810 -6814 18826 -6780
rect 18894 -6814 18910 -6780
rect 18810 -6830 18910 -6814
rect 20528 -670 20628 -654
rect 20528 -704 20544 -670
rect 20612 -704 20628 -670
rect 20528 -742 20628 -704
rect 20686 -670 20786 -654
rect 20686 -704 20702 -670
rect 20770 -704 20786 -670
rect 20686 -742 20786 -704
rect 20844 -670 20944 -654
rect 20844 -704 20860 -670
rect 20928 -704 20944 -670
rect 20844 -742 20944 -704
rect 21002 -670 21102 -654
rect 21002 -704 21018 -670
rect 21086 -704 21102 -670
rect 21002 -742 21102 -704
rect 21160 -670 21260 -654
rect 21160 -704 21176 -670
rect 21244 -704 21260 -670
rect 21160 -742 21260 -704
rect 21318 -670 21418 -654
rect 21318 -704 21334 -670
rect 21402 -704 21418 -670
rect 21318 -742 21418 -704
rect 21476 -670 21576 -654
rect 21476 -704 21492 -670
rect 21560 -704 21576 -670
rect 21476 -742 21576 -704
rect 21634 -670 21734 -654
rect 21634 -704 21650 -670
rect 21718 -704 21734 -670
rect 21634 -742 21734 -704
rect 21792 -670 21892 -654
rect 21792 -704 21808 -670
rect 21876 -704 21892 -670
rect 21792 -742 21892 -704
rect 21950 -670 22050 -654
rect 21950 -704 21966 -670
rect 22034 -704 22050 -670
rect 21950 -742 22050 -704
rect 22108 -670 22208 -654
rect 22108 -704 22124 -670
rect 22192 -704 22208 -670
rect 22108 -742 22208 -704
rect 22266 -670 22366 -654
rect 22266 -704 22282 -670
rect 22350 -704 22366 -670
rect 22266 -742 22366 -704
rect 22424 -670 22524 -654
rect 22424 -704 22440 -670
rect 22508 -704 22524 -670
rect 22424 -742 22524 -704
rect 22582 -670 22682 -654
rect 22582 -704 22598 -670
rect 22666 -704 22682 -670
rect 22582 -742 22682 -704
rect 22740 -670 22840 -654
rect 22740 -704 22756 -670
rect 22824 -704 22840 -670
rect 22740 -742 22840 -704
rect 22898 -670 22998 -654
rect 22898 -704 22914 -670
rect 22982 -704 22998 -670
rect 22898 -742 22998 -704
rect 23056 -670 23156 -654
rect 23056 -704 23072 -670
rect 23140 -704 23156 -670
rect 23056 -742 23156 -704
rect 23214 -670 23314 -654
rect 23214 -704 23230 -670
rect 23298 -704 23314 -670
rect 23214 -742 23314 -704
rect 23372 -670 23472 -654
rect 23372 -704 23388 -670
rect 23456 -704 23472 -670
rect 23372 -742 23472 -704
rect 23530 -670 23630 -654
rect 23530 -704 23546 -670
rect 23614 -704 23630 -670
rect 23530 -742 23630 -704
rect 23688 -670 23788 -654
rect 23688 -704 23704 -670
rect 23772 -704 23788 -670
rect 23688 -742 23788 -704
rect 23846 -670 23946 -654
rect 23846 -704 23862 -670
rect 23930 -704 23946 -670
rect 23846 -742 23946 -704
rect 24004 -670 24104 -654
rect 24004 -704 24020 -670
rect 24088 -704 24104 -670
rect 24004 -742 24104 -704
rect 24162 -670 24262 -654
rect 24162 -704 24178 -670
rect 24246 -704 24262 -670
rect 24162 -742 24262 -704
rect 24320 -670 24420 -654
rect 24320 -704 24336 -670
rect 24404 -704 24420 -670
rect 24320 -742 24420 -704
rect 24478 -670 24578 -654
rect 24478 -704 24494 -670
rect 24562 -704 24578 -670
rect 24478 -742 24578 -704
rect 24636 -670 24736 -654
rect 24636 -704 24652 -670
rect 24720 -704 24736 -670
rect 24636 -742 24736 -704
rect 24794 -670 24894 -654
rect 24794 -704 24810 -670
rect 24878 -704 24894 -670
rect 24794 -742 24894 -704
rect 24952 -670 25052 -654
rect 24952 -704 24968 -670
rect 25036 -704 25052 -670
rect 24952 -742 25052 -704
rect 25110 -670 25210 -654
rect 25110 -704 25126 -670
rect 25194 -704 25210 -670
rect 25110 -742 25210 -704
rect 20528 -6780 20628 -6742
rect 20528 -6814 20544 -6780
rect 20612 -6814 20628 -6780
rect 20528 -6830 20628 -6814
rect 20686 -6780 20786 -6742
rect 20686 -6814 20702 -6780
rect 20770 -6814 20786 -6780
rect 20686 -6830 20786 -6814
rect 20844 -6780 20944 -6742
rect 20844 -6814 20860 -6780
rect 20928 -6814 20944 -6780
rect 20844 -6830 20944 -6814
rect 21002 -6780 21102 -6742
rect 21002 -6814 21018 -6780
rect 21086 -6814 21102 -6780
rect 21002 -6830 21102 -6814
rect 21160 -6780 21260 -6742
rect 21160 -6814 21176 -6780
rect 21244 -6814 21260 -6780
rect 21160 -6830 21260 -6814
rect 21318 -6780 21418 -6742
rect 21318 -6814 21334 -6780
rect 21402 -6814 21418 -6780
rect 21318 -6830 21418 -6814
rect 21476 -6780 21576 -6742
rect 21476 -6814 21492 -6780
rect 21560 -6814 21576 -6780
rect 21476 -6830 21576 -6814
rect 21634 -6780 21734 -6742
rect 21634 -6814 21650 -6780
rect 21718 -6814 21734 -6780
rect 21634 -6830 21734 -6814
rect 21792 -6780 21892 -6742
rect 21792 -6814 21808 -6780
rect 21876 -6814 21892 -6780
rect 21792 -6830 21892 -6814
rect 21950 -6780 22050 -6742
rect 21950 -6814 21966 -6780
rect 22034 -6814 22050 -6780
rect 21950 -6830 22050 -6814
rect 22108 -6780 22208 -6742
rect 22108 -6814 22124 -6780
rect 22192 -6814 22208 -6780
rect 22108 -6830 22208 -6814
rect 22266 -6780 22366 -6742
rect 22266 -6814 22282 -6780
rect 22350 -6814 22366 -6780
rect 22266 -6830 22366 -6814
rect 22424 -6780 22524 -6742
rect 22424 -6814 22440 -6780
rect 22508 -6814 22524 -6780
rect 22424 -6830 22524 -6814
rect 22582 -6780 22682 -6742
rect 22582 -6814 22598 -6780
rect 22666 -6814 22682 -6780
rect 22582 -6830 22682 -6814
rect 22740 -6780 22840 -6742
rect 22740 -6814 22756 -6780
rect 22824 -6814 22840 -6780
rect 22740 -6830 22840 -6814
rect 22898 -6780 22998 -6742
rect 22898 -6814 22914 -6780
rect 22982 -6814 22998 -6780
rect 22898 -6830 22998 -6814
rect 23056 -6780 23156 -6742
rect 23056 -6814 23072 -6780
rect 23140 -6814 23156 -6780
rect 23056 -6830 23156 -6814
rect 23214 -6780 23314 -6742
rect 23214 -6814 23230 -6780
rect 23298 -6814 23314 -6780
rect 23214 -6830 23314 -6814
rect 23372 -6780 23472 -6742
rect 23372 -6814 23388 -6780
rect 23456 -6814 23472 -6780
rect 23372 -6830 23472 -6814
rect 23530 -6780 23630 -6742
rect 23530 -6814 23546 -6780
rect 23614 -6814 23630 -6780
rect 23530 -6830 23630 -6814
rect 23688 -6780 23788 -6742
rect 23688 -6814 23704 -6780
rect 23772 -6814 23788 -6780
rect 23688 -6830 23788 -6814
rect 23846 -6780 23946 -6742
rect 23846 -6814 23862 -6780
rect 23930 -6814 23946 -6780
rect 23846 -6830 23946 -6814
rect 24004 -6780 24104 -6742
rect 24004 -6814 24020 -6780
rect 24088 -6814 24104 -6780
rect 24004 -6830 24104 -6814
rect 24162 -6780 24262 -6742
rect 24162 -6814 24178 -6780
rect 24246 -6814 24262 -6780
rect 24162 -6830 24262 -6814
rect 24320 -6780 24420 -6742
rect 24320 -6814 24336 -6780
rect 24404 -6814 24420 -6780
rect 24320 -6830 24420 -6814
rect 24478 -6780 24578 -6742
rect 24478 -6814 24494 -6780
rect 24562 -6814 24578 -6780
rect 24478 -6830 24578 -6814
rect 24636 -6780 24736 -6742
rect 24636 -6814 24652 -6780
rect 24720 -6814 24736 -6780
rect 24636 -6830 24736 -6814
rect 24794 -6780 24894 -6742
rect 24794 -6814 24810 -6780
rect 24878 -6814 24894 -6780
rect 24794 -6830 24894 -6814
rect 24952 -6780 25052 -6742
rect 24952 -6814 24968 -6780
rect 25036 -6814 25052 -6780
rect 24952 -6830 25052 -6814
rect 25110 -6780 25210 -6742
rect 25110 -6814 25126 -6780
rect 25194 -6814 25210 -6780
rect 25110 -6830 25210 -6814
<< polycont >>
rect 1644 6296 1712 6330
rect 1802 6296 1870 6330
rect 1960 6296 2028 6330
rect 2118 6296 2186 6330
rect 2276 6296 2344 6330
rect 2434 6296 2502 6330
rect 2592 6296 2660 6330
rect 2750 6296 2818 6330
rect 2908 6296 2976 6330
rect 3066 6296 3134 6330
rect 3224 6296 3292 6330
rect 3382 6296 3450 6330
rect 3540 6296 3608 6330
rect 3698 6296 3766 6330
rect 3856 6296 3924 6330
rect 4014 6296 4082 6330
rect 4172 6296 4240 6330
rect 4330 6296 4398 6330
rect 4488 6296 4556 6330
rect 4646 6296 4714 6330
rect 4804 6296 4872 6330
rect 4962 6296 5030 6330
rect 5120 6296 5188 6330
rect 5278 6296 5346 6330
rect 5436 6296 5504 6330
rect 5594 6296 5662 6330
rect 5752 6296 5820 6330
rect 5910 6296 5978 6330
rect 6068 6296 6136 6330
rect 6226 6296 6294 6330
rect 1644 186 1712 220
rect 1802 186 1870 220
rect 1960 186 2028 220
rect 2118 186 2186 220
rect 2276 186 2344 220
rect 2434 186 2502 220
rect 2592 186 2660 220
rect 2750 186 2818 220
rect 2908 186 2976 220
rect 3066 186 3134 220
rect 3224 186 3292 220
rect 3382 186 3450 220
rect 3540 186 3608 220
rect 3698 186 3766 220
rect 3856 186 3924 220
rect 4014 186 4082 220
rect 4172 186 4240 220
rect 4330 186 4398 220
rect 4488 186 4556 220
rect 4646 186 4714 220
rect 4804 186 4872 220
rect 4962 186 5030 220
rect 5120 186 5188 220
rect 5278 186 5346 220
rect 5436 186 5504 220
rect 5594 186 5662 220
rect 5752 186 5820 220
rect 5910 186 5978 220
rect 6068 186 6136 220
rect 6226 186 6294 220
rect 7944 6296 8012 6330
rect 8102 6296 8170 6330
rect 8260 6296 8328 6330
rect 8418 6296 8486 6330
rect 8576 6296 8644 6330
rect 8734 6296 8802 6330
rect 8892 6296 8960 6330
rect 9050 6296 9118 6330
rect 9208 6296 9276 6330
rect 9366 6296 9434 6330
rect 9524 6296 9592 6330
rect 9682 6296 9750 6330
rect 9840 6296 9908 6330
rect 9998 6296 10066 6330
rect 10156 6296 10224 6330
rect 10314 6296 10382 6330
rect 10472 6296 10540 6330
rect 10630 6296 10698 6330
rect 10788 6296 10856 6330
rect 10946 6296 11014 6330
rect 11104 6296 11172 6330
rect 11262 6296 11330 6330
rect 11420 6296 11488 6330
rect 11578 6296 11646 6330
rect 11736 6296 11804 6330
rect 11894 6296 11962 6330
rect 12052 6296 12120 6330
rect 12210 6296 12278 6330
rect 12368 6296 12436 6330
rect 12526 6296 12594 6330
rect 7944 186 8012 220
rect 8102 186 8170 220
rect 8260 186 8328 220
rect 8418 186 8486 220
rect 8576 186 8644 220
rect 8734 186 8802 220
rect 8892 186 8960 220
rect 9050 186 9118 220
rect 9208 186 9276 220
rect 9366 186 9434 220
rect 9524 186 9592 220
rect 9682 186 9750 220
rect 9840 186 9908 220
rect 9998 186 10066 220
rect 10156 186 10224 220
rect 10314 186 10382 220
rect 10472 186 10540 220
rect 10630 186 10698 220
rect 10788 186 10856 220
rect 10946 186 11014 220
rect 11104 186 11172 220
rect 11262 186 11330 220
rect 11420 186 11488 220
rect 11578 186 11646 220
rect 11736 186 11804 220
rect 11894 186 11962 220
rect 12052 186 12120 220
rect 12210 186 12278 220
rect 12368 186 12436 220
rect 12526 186 12594 220
rect 14244 6296 14312 6330
rect 14402 6296 14470 6330
rect 14560 6296 14628 6330
rect 14718 6296 14786 6330
rect 14876 6296 14944 6330
rect 15034 6296 15102 6330
rect 15192 6296 15260 6330
rect 15350 6296 15418 6330
rect 15508 6296 15576 6330
rect 15666 6296 15734 6330
rect 15824 6296 15892 6330
rect 15982 6296 16050 6330
rect 16140 6296 16208 6330
rect 16298 6296 16366 6330
rect 16456 6296 16524 6330
rect 16614 6296 16682 6330
rect 16772 6296 16840 6330
rect 16930 6296 16998 6330
rect 17088 6296 17156 6330
rect 17246 6296 17314 6330
rect 17404 6296 17472 6330
rect 17562 6296 17630 6330
rect 17720 6296 17788 6330
rect 17878 6296 17946 6330
rect 18036 6296 18104 6330
rect 18194 6296 18262 6330
rect 18352 6296 18420 6330
rect 18510 6296 18578 6330
rect 18668 6296 18736 6330
rect 18826 6296 18894 6330
rect 14244 186 14312 220
rect 14402 186 14470 220
rect 14560 186 14628 220
rect 14718 186 14786 220
rect 14876 186 14944 220
rect 15034 186 15102 220
rect 15192 186 15260 220
rect 15350 186 15418 220
rect 15508 186 15576 220
rect 15666 186 15734 220
rect 15824 186 15892 220
rect 15982 186 16050 220
rect 16140 186 16208 220
rect 16298 186 16366 220
rect 16456 186 16524 220
rect 16614 186 16682 220
rect 16772 186 16840 220
rect 16930 186 16998 220
rect 17088 186 17156 220
rect 17246 186 17314 220
rect 17404 186 17472 220
rect 17562 186 17630 220
rect 17720 186 17788 220
rect 17878 186 17946 220
rect 18036 186 18104 220
rect 18194 186 18262 220
rect 18352 186 18420 220
rect 18510 186 18578 220
rect 18668 186 18736 220
rect 18826 186 18894 220
rect 20544 6296 20612 6330
rect 20702 6296 20770 6330
rect 20860 6296 20928 6330
rect 21018 6296 21086 6330
rect 21176 6296 21244 6330
rect 21334 6296 21402 6330
rect 21492 6296 21560 6330
rect 21650 6296 21718 6330
rect 21808 6296 21876 6330
rect 21966 6296 22034 6330
rect 22124 6296 22192 6330
rect 22282 6296 22350 6330
rect 22440 6296 22508 6330
rect 22598 6296 22666 6330
rect 22756 6296 22824 6330
rect 22914 6296 22982 6330
rect 23072 6296 23140 6330
rect 23230 6296 23298 6330
rect 23388 6296 23456 6330
rect 23546 6296 23614 6330
rect 23704 6296 23772 6330
rect 23862 6296 23930 6330
rect 24020 6296 24088 6330
rect 24178 6296 24246 6330
rect 24336 6296 24404 6330
rect 24494 6296 24562 6330
rect 24652 6296 24720 6330
rect 24810 6296 24878 6330
rect 24968 6296 25036 6330
rect 25126 6296 25194 6330
rect 20544 186 20612 220
rect 20702 186 20770 220
rect 20860 186 20928 220
rect 21018 186 21086 220
rect 21176 186 21244 220
rect 21334 186 21402 220
rect 21492 186 21560 220
rect 21650 186 21718 220
rect 21808 186 21876 220
rect 21966 186 22034 220
rect 22124 186 22192 220
rect 22282 186 22350 220
rect 22440 186 22508 220
rect 22598 186 22666 220
rect 22756 186 22824 220
rect 22914 186 22982 220
rect 23072 186 23140 220
rect 23230 186 23298 220
rect 23388 186 23456 220
rect 23546 186 23614 220
rect 23704 186 23772 220
rect 23862 186 23930 220
rect 24020 186 24088 220
rect 24178 186 24246 220
rect 24336 186 24404 220
rect 24494 186 24562 220
rect 24652 186 24720 220
rect 24810 186 24878 220
rect 24968 186 25036 220
rect 25126 186 25194 220
rect 1644 -704 1712 -670
rect 1802 -704 1870 -670
rect 1960 -704 2028 -670
rect 2118 -704 2186 -670
rect 2276 -704 2344 -670
rect 2434 -704 2502 -670
rect 2592 -704 2660 -670
rect 2750 -704 2818 -670
rect 2908 -704 2976 -670
rect 3066 -704 3134 -670
rect 3224 -704 3292 -670
rect 3382 -704 3450 -670
rect 3540 -704 3608 -670
rect 3698 -704 3766 -670
rect 3856 -704 3924 -670
rect 4014 -704 4082 -670
rect 4172 -704 4240 -670
rect 4330 -704 4398 -670
rect 4488 -704 4556 -670
rect 4646 -704 4714 -670
rect 4804 -704 4872 -670
rect 4962 -704 5030 -670
rect 5120 -704 5188 -670
rect 5278 -704 5346 -670
rect 5436 -704 5504 -670
rect 5594 -704 5662 -670
rect 5752 -704 5820 -670
rect 5910 -704 5978 -670
rect 6068 -704 6136 -670
rect 6226 -704 6294 -670
rect 1644 -6814 1712 -6780
rect 1802 -6814 1870 -6780
rect 1960 -6814 2028 -6780
rect 2118 -6814 2186 -6780
rect 2276 -6814 2344 -6780
rect 2434 -6814 2502 -6780
rect 2592 -6814 2660 -6780
rect 2750 -6814 2818 -6780
rect 2908 -6814 2976 -6780
rect 3066 -6814 3134 -6780
rect 3224 -6814 3292 -6780
rect 3382 -6814 3450 -6780
rect 3540 -6814 3608 -6780
rect 3698 -6814 3766 -6780
rect 3856 -6814 3924 -6780
rect 4014 -6814 4082 -6780
rect 4172 -6814 4240 -6780
rect 4330 -6814 4398 -6780
rect 4488 -6814 4556 -6780
rect 4646 -6814 4714 -6780
rect 4804 -6814 4872 -6780
rect 4962 -6814 5030 -6780
rect 5120 -6814 5188 -6780
rect 5278 -6814 5346 -6780
rect 5436 -6814 5504 -6780
rect 5594 -6814 5662 -6780
rect 5752 -6814 5820 -6780
rect 5910 -6814 5978 -6780
rect 6068 -6814 6136 -6780
rect 6226 -6814 6294 -6780
rect 7944 -704 8012 -670
rect 8102 -704 8170 -670
rect 8260 -704 8328 -670
rect 8418 -704 8486 -670
rect 8576 -704 8644 -670
rect 8734 -704 8802 -670
rect 8892 -704 8960 -670
rect 9050 -704 9118 -670
rect 9208 -704 9276 -670
rect 9366 -704 9434 -670
rect 9524 -704 9592 -670
rect 9682 -704 9750 -670
rect 9840 -704 9908 -670
rect 9998 -704 10066 -670
rect 10156 -704 10224 -670
rect 10314 -704 10382 -670
rect 10472 -704 10540 -670
rect 10630 -704 10698 -670
rect 10788 -704 10856 -670
rect 10946 -704 11014 -670
rect 11104 -704 11172 -670
rect 11262 -704 11330 -670
rect 11420 -704 11488 -670
rect 11578 -704 11646 -670
rect 11736 -704 11804 -670
rect 11894 -704 11962 -670
rect 12052 -704 12120 -670
rect 12210 -704 12278 -670
rect 12368 -704 12436 -670
rect 12526 -704 12594 -670
rect 7944 -6814 8012 -6780
rect 8102 -6814 8170 -6780
rect 8260 -6814 8328 -6780
rect 8418 -6814 8486 -6780
rect 8576 -6814 8644 -6780
rect 8734 -6814 8802 -6780
rect 8892 -6814 8960 -6780
rect 9050 -6814 9118 -6780
rect 9208 -6814 9276 -6780
rect 9366 -6814 9434 -6780
rect 9524 -6814 9592 -6780
rect 9682 -6814 9750 -6780
rect 9840 -6814 9908 -6780
rect 9998 -6814 10066 -6780
rect 10156 -6814 10224 -6780
rect 10314 -6814 10382 -6780
rect 10472 -6814 10540 -6780
rect 10630 -6814 10698 -6780
rect 10788 -6814 10856 -6780
rect 10946 -6814 11014 -6780
rect 11104 -6814 11172 -6780
rect 11262 -6814 11330 -6780
rect 11420 -6814 11488 -6780
rect 11578 -6814 11646 -6780
rect 11736 -6814 11804 -6780
rect 11894 -6814 11962 -6780
rect 12052 -6814 12120 -6780
rect 12210 -6814 12278 -6780
rect 12368 -6814 12436 -6780
rect 12526 -6814 12594 -6780
rect 14244 -704 14312 -670
rect 14402 -704 14470 -670
rect 14560 -704 14628 -670
rect 14718 -704 14786 -670
rect 14876 -704 14944 -670
rect 15034 -704 15102 -670
rect 15192 -704 15260 -670
rect 15350 -704 15418 -670
rect 15508 -704 15576 -670
rect 15666 -704 15734 -670
rect 15824 -704 15892 -670
rect 15982 -704 16050 -670
rect 16140 -704 16208 -670
rect 16298 -704 16366 -670
rect 16456 -704 16524 -670
rect 16614 -704 16682 -670
rect 16772 -704 16840 -670
rect 16930 -704 16998 -670
rect 17088 -704 17156 -670
rect 17246 -704 17314 -670
rect 17404 -704 17472 -670
rect 17562 -704 17630 -670
rect 17720 -704 17788 -670
rect 17878 -704 17946 -670
rect 18036 -704 18104 -670
rect 18194 -704 18262 -670
rect 18352 -704 18420 -670
rect 18510 -704 18578 -670
rect 18668 -704 18736 -670
rect 18826 -704 18894 -670
rect 14244 -6814 14312 -6780
rect 14402 -6814 14470 -6780
rect 14560 -6814 14628 -6780
rect 14718 -6814 14786 -6780
rect 14876 -6814 14944 -6780
rect 15034 -6814 15102 -6780
rect 15192 -6814 15260 -6780
rect 15350 -6814 15418 -6780
rect 15508 -6814 15576 -6780
rect 15666 -6814 15734 -6780
rect 15824 -6814 15892 -6780
rect 15982 -6814 16050 -6780
rect 16140 -6814 16208 -6780
rect 16298 -6814 16366 -6780
rect 16456 -6814 16524 -6780
rect 16614 -6814 16682 -6780
rect 16772 -6814 16840 -6780
rect 16930 -6814 16998 -6780
rect 17088 -6814 17156 -6780
rect 17246 -6814 17314 -6780
rect 17404 -6814 17472 -6780
rect 17562 -6814 17630 -6780
rect 17720 -6814 17788 -6780
rect 17878 -6814 17946 -6780
rect 18036 -6814 18104 -6780
rect 18194 -6814 18262 -6780
rect 18352 -6814 18420 -6780
rect 18510 -6814 18578 -6780
rect 18668 -6814 18736 -6780
rect 18826 -6814 18894 -6780
rect 20544 -704 20612 -670
rect 20702 -704 20770 -670
rect 20860 -704 20928 -670
rect 21018 -704 21086 -670
rect 21176 -704 21244 -670
rect 21334 -704 21402 -670
rect 21492 -704 21560 -670
rect 21650 -704 21718 -670
rect 21808 -704 21876 -670
rect 21966 -704 22034 -670
rect 22124 -704 22192 -670
rect 22282 -704 22350 -670
rect 22440 -704 22508 -670
rect 22598 -704 22666 -670
rect 22756 -704 22824 -670
rect 22914 -704 22982 -670
rect 23072 -704 23140 -670
rect 23230 -704 23298 -670
rect 23388 -704 23456 -670
rect 23546 -704 23614 -670
rect 23704 -704 23772 -670
rect 23862 -704 23930 -670
rect 24020 -704 24088 -670
rect 24178 -704 24246 -670
rect 24336 -704 24404 -670
rect 24494 -704 24562 -670
rect 24652 -704 24720 -670
rect 24810 -704 24878 -670
rect 24968 -704 25036 -670
rect 25126 -704 25194 -670
rect 20544 -6814 20612 -6780
rect 20702 -6814 20770 -6780
rect 20860 -6814 20928 -6780
rect 21018 -6814 21086 -6780
rect 21176 -6814 21244 -6780
rect 21334 -6814 21402 -6780
rect 21492 -6814 21560 -6780
rect 21650 -6814 21718 -6780
rect 21808 -6814 21876 -6780
rect 21966 -6814 22034 -6780
rect 22124 -6814 22192 -6780
rect 22282 -6814 22350 -6780
rect 22440 -6814 22508 -6780
rect 22598 -6814 22666 -6780
rect 22756 -6814 22824 -6780
rect 22914 -6814 22982 -6780
rect 23072 -6814 23140 -6780
rect 23230 -6814 23298 -6780
rect 23388 -6814 23456 -6780
rect 23546 -6814 23614 -6780
rect 23704 -6814 23772 -6780
rect 23862 -6814 23930 -6780
rect 24020 -6814 24088 -6780
rect 24178 -6814 24246 -6780
rect 24336 -6814 24404 -6780
rect 24494 -6814 24562 -6780
rect 24652 -6814 24720 -6780
rect 24810 -6814 24878 -6780
rect 24968 -6814 25036 -6780
rect 25126 -6814 25194 -6780
<< locali >>
rect 1448 6434 1544 6468
rect 6394 6434 6490 6468
rect 1448 6372 1482 6434
rect 6456 6372 6490 6434
rect 1628 6296 1644 6330
rect 1712 6296 1728 6330
rect 1786 6296 1802 6330
rect 1870 6296 1886 6330
rect 1944 6296 1960 6330
rect 2028 6296 2044 6330
rect 2102 6296 2118 6330
rect 2186 6296 2202 6330
rect 2260 6296 2276 6330
rect 2344 6296 2360 6330
rect 2418 6296 2434 6330
rect 2502 6296 2518 6330
rect 2576 6296 2592 6330
rect 2660 6296 2676 6330
rect 2734 6296 2750 6330
rect 2818 6296 2834 6330
rect 2892 6296 2908 6330
rect 2976 6296 2992 6330
rect 3050 6296 3066 6330
rect 3134 6296 3150 6330
rect 3208 6296 3224 6330
rect 3292 6296 3308 6330
rect 3366 6296 3382 6330
rect 3450 6296 3466 6330
rect 3524 6296 3540 6330
rect 3608 6296 3624 6330
rect 3682 6296 3698 6330
rect 3766 6296 3782 6330
rect 3840 6296 3856 6330
rect 3924 6296 3940 6330
rect 3998 6296 4014 6330
rect 4082 6296 4098 6330
rect 4156 6296 4172 6330
rect 4240 6296 4256 6330
rect 4314 6296 4330 6330
rect 4398 6296 4414 6330
rect 4472 6296 4488 6330
rect 4556 6296 4572 6330
rect 4630 6296 4646 6330
rect 4714 6296 4730 6330
rect 4788 6296 4804 6330
rect 4872 6296 4888 6330
rect 4946 6296 4962 6330
rect 5030 6296 5046 6330
rect 5104 6296 5120 6330
rect 5188 6296 5204 6330
rect 5262 6296 5278 6330
rect 5346 6296 5362 6330
rect 5420 6296 5436 6330
rect 5504 6296 5520 6330
rect 5578 6296 5594 6330
rect 5662 6296 5678 6330
rect 5736 6296 5752 6330
rect 5820 6296 5836 6330
rect 5894 6296 5910 6330
rect 5978 6296 5994 6330
rect 6052 6296 6068 6330
rect 6136 6296 6152 6330
rect 6210 6296 6226 6330
rect 6294 6296 6310 6330
rect 7748 6434 7844 6468
rect 12694 6434 12790 6468
rect 7748 6372 7782 6434
rect 12756 6372 12790 6434
rect 7928 6296 7944 6330
rect 8012 6296 8028 6330
rect 8086 6296 8102 6330
rect 8170 6296 8186 6330
rect 8244 6296 8260 6330
rect 8328 6296 8344 6330
rect 8402 6296 8418 6330
rect 8486 6296 8502 6330
rect 8560 6296 8576 6330
rect 8644 6296 8660 6330
rect 8718 6296 8734 6330
rect 8802 6296 8818 6330
rect 8876 6296 8892 6330
rect 8960 6296 8976 6330
rect 9034 6296 9050 6330
rect 9118 6296 9134 6330
rect 9192 6296 9208 6330
rect 9276 6296 9292 6330
rect 9350 6296 9366 6330
rect 9434 6296 9450 6330
rect 9508 6296 9524 6330
rect 9592 6296 9608 6330
rect 9666 6296 9682 6330
rect 9750 6296 9766 6330
rect 9824 6296 9840 6330
rect 9908 6296 9924 6330
rect 9982 6296 9998 6330
rect 10066 6296 10082 6330
rect 10140 6296 10156 6330
rect 10224 6296 10240 6330
rect 10298 6296 10314 6330
rect 10382 6296 10398 6330
rect 10456 6296 10472 6330
rect 10540 6296 10556 6330
rect 10614 6296 10630 6330
rect 10698 6296 10714 6330
rect 10772 6296 10788 6330
rect 10856 6296 10872 6330
rect 10930 6296 10946 6330
rect 11014 6296 11030 6330
rect 11088 6296 11104 6330
rect 11172 6296 11188 6330
rect 11246 6296 11262 6330
rect 11330 6296 11346 6330
rect 11404 6296 11420 6330
rect 11488 6296 11504 6330
rect 11562 6296 11578 6330
rect 11646 6296 11662 6330
rect 11720 6296 11736 6330
rect 11804 6296 11820 6330
rect 11878 6296 11894 6330
rect 11962 6296 11978 6330
rect 12036 6296 12052 6330
rect 12120 6296 12136 6330
rect 12194 6296 12210 6330
rect 12278 6296 12294 6330
rect 12352 6296 12368 6330
rect 12436 6296 12452 6330
rect 12510 6296 12526 6330
rect 12594 6296 12610 6330
rect 14048 6434 14144 6468
rect 18994 6434 19090 6468
rect 14048 6372 14082 6434
rect 19056 6372 19090 6434
rect 14228 6296 14244 6330
rect 14312 6296 14328 6330
rect 14386 6296 14402 6330
rect 14470 6296 14486 6330
rect 14544 6296 14560 6330
rect 14628 6296 14644 6330
rect 14702 6296 14718 6330
rect 14786 6296 14802 6330
rect 14860 6296 14876 6330
rect 14944 6296 14960 6330
rect 15018 6296 15034 6330
rect 15102 6296 15118 6330
rect 15176 6296 15192 6330
rect 15260 6296 15276 6330
rect 15334 6296 15350 6330
rect 15418 6296 15434 6330
rect 15492 6296 15508 6330
rect 15576 6296 15592 6330
rect 15650 6296 15666 6330
rect 15734 6296 15750 6330
rect 15808 6296 15824 6330
rect 15892 6296 15908 6330
rect 15966 6296 15982 6330
rect 16050 6296 16066 6330
rect 16124 6296 16140 6330
rect 16208 6296 16224 6330
rect 16282 6296 16298 6330
rect 16366 6296 16382 6330
rect 16440 6296 16456 6330
rect 16524 6296 16540 6330
rect 16598 6296 16614 6330
rect 16682 6296 16698 6330
rect 16756 6296 16772 6330
rect 16840 6296 16856 6330
rect 16914 6296 16930 6330
rect 16998 6296 17014 6330
rect 17072 6296 17088 6330
rect 17156 6296 17172 6330
rect 17230 6296 17246 6330
rect 17314 6296 17330 6330
rect 17388 6296 17404 6330
rect 17472 6296 17488 6330
rect 17546 6296 17562 6330
rect 17630 6296 17646 6330
rect 17704 6296 17720 6330
rect 17788 6296 17804 6330
rect 17862 6296 17878 6330
rect 17946 6296 17962 6330
rect 18020 6296 18036 6330
rect 18104 6296 18120 6330
rect 18178 6296 18194 6330
rect 18262 6296 18278 6330
rect 18336 6296 18352 6330
rect 18420 6296 18436 6330
rect 18494 6296 18510 6330
rect 18578 6296 18594 6330
rect 18652 6296 18668 6330
rect 18736 6296 18752 6330
rect 18810 6296 18826 6330
rect 18894 6296 18910 6330
rect 20348 6434 20444 6468
rect 25294 6434 25390 6468
rect 20348 6372 20382 6434
rect 25356 6372 25390 6434
rect 20528 6296 20544 6330
rect 20612 6296 20628 6330
rect 20686 6296 20702 6330
rect 20770 6296 20786 6330
rect 20844 6296 20860 6330
rect 20928 6296 20944 6330
rect 21002 6296 21018 6330
rect 21086 6296 21102 6330
rect 21160 6296 21176 6330
rect 21244 6296 21260 6330
rect 21318 6296 21334 6330
rect 21402 6296 21418 6330
rect 21476 6296 21492 6330
rect 21560 6296 21576 6330
rect 21634 6296 21650 6330
rect 21718 6296 21734 6330
rect 21792 6296 21808 6330
rect 21876 6296 21892 6330
rect 21950 6296 21966 6330
rect 22034 6296 22050 6330
rect 22108 6296 22124 6330
rect 22192 6296 22208 6330
rect 22266 6296 22282 6330
rect 22350 6296 22366 6330
rect 22424 6296 22440 6330
rect 22508 6296 22524 6330
rect 22582 6296 22598 6330
rect 22666 6296 22682 6330
rect 22740 6296 22756 6330
rect 22824 6296 22840 6330
rect 22898 6296 22914 6330
rect 22982 6296 22998 6330
rect 23056 6296 23072 6330
rect 23140 6296 23156 6330
rect 23214 6296 23230 6330
rect 23298 6296 23314 6330
rect 23372 6296 23388 6330
rect 23456 6296 23472 6330
rect 23530 6296 23546 6330
rect 23614 6296 23630 6330
rect 23688 6296 23704 6330
rect 23772 6296 23788 6330
rect 23846 6296 23862 6330
rect 23930 6296 23946 6330
rect 24004 6296 24020 6330
rect 24088 6296 24104 6330
rect 24162 6296 24178 6330
rect 24246 6296 24262 6330
rect 24320 6296 24336 6330
rect 24404 6296 24420 6330
rect 24478 6296 24494 6330
rect 24562 6296 24578 6330
rect 24636 6296 24652 6330
rect 24720 6296 24736 6330
rect 24794 6296 24810 6330
rect 24878 6296 24894 6330
rect 24952 6296 24968 6330
rect 25036 6296 25052 6330
rect 25110 6296 25126 6330
rect 25194 6296 25210 6330
rect 1582 6246 1616 6262
rect 1582 254 1616 270
rect 1740 6246 1774 6262
rect 1740 254 1774 270
rect 1898 6246 1932 6262
rect 1898 254 1932 270
rect 2056 6246 2090 6262
rect 2056 254 2090 270
rect 2214 6246 2248 6262
rect 2214 254 2248 270
rect 2372 6246 2406 6262
rect 2372 254 2406 270
rect 2530 6246 2564 6262
rect 2530 254 2564 270
rect 2688 6246 2722 6262
rect 2688 254 2722 270
rect 2846 6246 2880 6262
rect 2846 254 2880 270
rect 3004 6246 3038 6262
rect 3004 254 3038 270
rect 3162 6246 3196 6262
rect 3162 254 3196 270
rect 3320 6246 3354 6262
rect 3320 254 3354 270
rect 3478 6246 3512 6262
rect 3478 254 3512 270
rect 3636 6246 3670 6262
rect 3636 254 3670 270
rect 3794 6246 3828 6262
rect 3794 254 3828 270
rect 3952 6246 3986 6262
rect 3952 254 3986 270
rect 4110 6246 4144 6262
rect 4110 254 4144 270
rect 4268 6246 4302 6262
rect 4268 254 4302 270
rect 4426 6246 4460 6262
rect 4426 254 4460 270
rect 4584 6246 4618 6262
rect 4584 254 4618 270
rect 4742 6246 4776 6262
rect 4742 254 4776 270
rect 4900 6246 4934 6262
rect 4900 254 4934 270
rect 5058 6246 5092 6262
rect 5058 254 5092 270
rect 5216 6246 5250 6262
rect 5216 254 5250 270
rect 5374 6246 5408 6262
rect 5374 254 5408 270
rect 5532 6246 5566 6262
rect 5532 254 5566 270
rect 5690 6246 5724 6262
rect 5690 254 5724 270
rect 5848 6246 5882 6262
rect 5848 254 5882 270
rect 6006 6246 6040 6262
rect 6006 254 6040 270
rect 6164 6246 6198 6262
rect 6164 254 6198 270
rect 6322 6246 6356 6262
rect 6322 254 6356 270
rect 7882 6246 7916 6262
rect 7882 254 7916 270
rect 8040 6246 8074 6262
rect 8040 254 8074 270
rect 8198 6246 8232 6262
rect 8198 254 8232 270
rect 8356 6246 8390 6262
rect 8356 254 8390 270
rect 8514 6246 8548 6262
rect 8514 254 8548 270
rect 8672 6246 8706 6262
rect 8672 254 8706 270
rect 8830 6246 8864 6262
rect 8830 254 8864 270
rect 8988 6246 9022 6262
rect 8988 254 9022 270
rect 9146 6246 9180 6262
rect 9146 254 9180 270
rect 9304 6246 9338 6262
rect 9304 254 9338 270
rect 9462 6246 9496 6262
rect 9462 254 9496 270
rect 9620 6246 9654 6262
rect 9620 254 9654 270
rect 9778 6246 9812 6262
rect 9778 254 9812 270
rect 9936 6246 9970 6262
rect 9936 254 9970 270
rect 10094 6246 10128 6262
rect 10094 254 10128 270
rect 10252 6246 10286 6262
rect 10252 254 10286 270
rect 10410 6246 10444 6262
rect 10410 254 10444 270
rect 10568 6246 10602 6262
rect 10568 254 10602 270
rect 10726 6246 10760 6262
rect 10726 254 10760 270
rect 10884 6246 10918 6262
rect 10884 254 10918 270
rect 11042 6246 11076 6262
rect 11042 254 11076 270
rect 11200 6246 11234 6262
rect 11200 254 11234 270
rect 11358 6246 11392 6262
rect 11358 254 11392 270
rect 11516 6246 11550 6262
rect 11516 254 11550 270
rect 11674 6246 11708 6262
rect 11674 254 11708 270
rect 11832 6246 11866 6262
rect 11832 254 11866 270
rect 11990 6246 12024 6262
rect 11990 254 12024 270
rect 12148 6246 12182 6262
rect 12148 254 12182 270
rect 12306 6246 12340 6262
rect 12306 254 12340 270
rect 12464 6246 12498 6262
rect 12464 254 12498 270
rect 12622 6246 12656 6262
rect 12622 254 12656 270
rect 14182 6246 14216 6262
rect 14182 254 14216 270
rect 14340 6246 14374 6262
rect 14340 254 14374 270
rect 14498 6246 14532 6262
rect 14498 254 14532 270
rect 14656 6246 14690 6262
rect 14656 254 14690 270
rect 14814 6246 14848 6262
rect 14814 254 14848 270
rect 14972 6246 15006 6262
rect 14972 254 15006 270
rect 15130 6246 15164 6262
rect 15130 254 15164 270
rect 15288 6246 15322 6262
rect 15288 254 15322 270
rect 15446 6246 15480 6262
rect 15446 254 15480 270
rect 15604 6246 15638 6262
rect 15604 254 15638 270
rect 15762 6246 15796 6262
rect 15762 254 15796 270
rect 15920 6246 15954 6262
rect 15920 254 15954 270
rect 16078 6246 16112 6262
rect 16078 254 16112 270
rect 16236 6246 16270 6262
rect 16236 254 16270 270
rect 16394 6246 16428 6262
rect 16394 254 16428 270
rect 16552 6246 16586 6262
rect 16552 254 16586 270
rect 16710 6246 16744 6262
rect 16710 254 16744 270
rect 16868 6246 16902 6262
rect 16868 254 16902 270
rect 17026 6246 17060 6262
rect 17026 254 17060 270
rect 17184 6246 17218 6262
rect 17184 254 17218 270
rect 17342 6246 17376 6262
rect 17342 254 17376 270
rect 17500 6246 17534 6262
rect 17500 254 17534 270
rect 17658 6246 17692 6262
rect 17658 254 17692 270
rect 17816 6246 17850 6262
rect 17816 254 17850 270
rect 17974 6246 18008 6262
rect 17974 254 18008 270
rect 18132 6246 18166 6262
rect 18132 254 18166 270
rect 18290 6246 18324 6262
rect 18290 254 18324 270
rect 18448 6246 18482 6262
rect 18448 254 18482 270
rect 18606 6246 18640 6262
rect 18606 254 18640 270
rect 18764 6246 18798 6262
rect 18764 254 18798 270
rect 18922 6246 18956 6262
rect 18922 254 18956 270
rect 20482 6246 20516 6262
rect 20482 254 20516 270
rect 20640 6246 20674 6262
rect 20640 254 20674 270
rect 20798 6246 20832 6262
rect 20798 254 20832 270
rect 20956 6246 20990 6262
rect 20956 254 20990 270
rect 21114 6246 21148 6262
rect 21114 254 21148 270
rect 21272 6246 21306 6262
rect 21272 254 21306 270
rect 21430 6246 21464 6262
rect 21430 254 21464 270
rect 21588 6246 21622 6262
rect 21588 254 21622 270
rect 21746 6246 21780 6262
rect 21746 254 21780 270
rect 21904 6246 21938 6262
rect 21904 254 21938 270
rect 22062 6246 22096 6262
rect 22062 254 22096 270
rect 22220 6246 22254 6262
rect 22220 254 22254 270
rect 22378 6246 22412 6262
rect 22378 254 22412 270
rect 22536 6246 22570 6262
rect 22536 254 22570 270
rect 22694 6246 22728 6262
rect 22694 254 22728 270
rect 22852 6246 22886 6262
rect 22852 254 22886 270
rect 23010 6246 23044 6262
rect 23010 254 23044 270
rect 23168 6246 23202 6262
rect 23168 254 23202 270
rect 23326 6246 23360 6262
rect 23326 254 23360 270
rect 23484 6246 23518 6262
rect 23484 254 23518 270
rect 23642 6246 23676 6262
rect 23642 254 23676 270
rect 23800 6246 23834 6262
rect 23800 254 23834 270
rect 23958 6246 23992 6262
rect 23958 254 23992 270
rect 24116 6246 24150 6262
rect 24116 254 24150 270
rect 24274 6246 24308 6262
rect 24274 254 24308 270
rect 24432 6246 24466 6262
rect 24432 254 24466 270
rect 24590 6246 24624 6262
rect 24590 254 24624 270
rect 24748 6246 24782 6262
rect 24748 254 24782 270
rect 24906 6246 24940 6262
rect 24906 254 24940 270
rect 25064 6246 25098 6262
rect 25064 254 25098 270
rect 25222 6246 25256 6262
rect 25222 254 25256 270
rect 1628 186 1644 220
rect 1712 186 1728 220
rect 1786 186 1802 220
rect 1870 186 1886 220
rect 1944 186 1960 220
rect 2028 186 2044 220
rect 2102 186 2118 220
rect 2186 186 2202 220
rect 2260 186 2276 220
rect 2344 186 2360 220
rect 2418 186 2434 220
rect 2502 186 2518 220
rect 2576 186 2592 220
rect 2660 186 2676 220
rect 2734 186 2750 220
rect 2818 186 2834 220
rect 2892 186 2908 220
rect 2976 186 2992 220
rect 3050 186 3066 220
rect 3134 186 3150 220
rect 3208 186 3224 220
rect 3292 186 3308 220
rect 3366 186 3382 220
rect 3450 186 3466 220
rect 3524 186 3540 220
rect 3608 186 3624 220
rect 3682 186 3698 220
rect 3766 186 3782 220
rect 3840 186 3856 220
rect 3924 186 3940 220
rect 3998 186 4014 220
rect 4082 186 4098 220
rect 4156 186 4172 220
rect 4240 186 4256 220
rect 4314 186 4330 220
rect 4398 186 4414 220
rect 4472 186 4488 220
rect 4556 186 4572 220
rect 4630 186 4646 220
rect 4714 186 4730 220
rect 4788 186 4804 220
rect 4872 186 4888 220
rect 4946 186 4962 220
rect 5030 186 5046 220
rect 5104 186 5120 220
rect 5188 186 5204 220
rect 5262 186 5278 220
rect 5346 186 5362 220
rect 5420 186 5436 220
rect 5504 186 5520 220
rect 5578 186 5594 220
rect 5662 186 5678 220
rect 5736 186 5752 220
rect 5820 186 5836 220
rect 5894 186 5910 220
rect 5978 186 5994 220
rect 6052 186 6068 220
rect 6136 186 6152 220
rect 6210 186 6226 220
rect 6294 186 6310 220
rect 1448 82 1482 144
rect 6456 82 6490 144
rect 1448 48 1544 82
rect 6394 48 6490 82
rect 7928 186 7944 220
rect 8012 186 8028 220
rect 8086 186 8102 220
rect 8170 186 8186 220
rect 8244 186 8260 220
rect 8328 186 8344 220
rect 8402 186 8418 220
rect 8486 186 8502 220
rect 8560 186 8576 220
rect 8644 186 8660 220
rect 8718 186 8734 220
rect 8802 186 8818 220
rect 8876 186 8892 220
rect 8960 186 8976 220
rect 9034 186 9050 220
rect 9118 186 9134 220
rect 9192 186 9208 220
rect 9276 186 9292 220
rect 9350 186 9366 220
rect 9434 186 9450 220
rect 9508 186 9524 220
rect 9592 186 9608 220
rect 9666 186 9682 220
rect 9750 186 9766 220
rect 9824 186 9840 220
rect 9908 186 9924 220
rect 9982 186 9998 220
rect 10066 186 10082 220
rect 10140 186 10156 220
rect 10224 186 10240 220
rect 10298 186 10314 220
rect 10382 186 10398 220
rect 10456 186 10472 220
rect 10540 186 10556 220
rect 10614 186 10630 220
rect 10698 186 10714 220
rect 10772 186 10788 220
rect 10856 186 10872 220
rect 10930 186 10946 220
rect 11014 186 11030 220
rect 11088 186 11104 220
rect 11172 186 11188 220
rect 11246 186 11262 220
rect 11330 186 11346 220
rect 11404 186 11420 220
rect 11488 186 11504 220
rect 11562 186 11578 220
rect 11646 186 11662 220
rect 11720 186 11736 220
rect 11804 186 11820 220
rect 11878 186 11894 220
rect 11962 186 11978 220
rect 12036 186 12052 220
rect 12120 186 12136 220
rect 12194 186 12210 220
rect 12278 186 12294 220
rect 12352 186 12368 220
rect 12436 186 12452 220
rect 12510 186 12526 220
rect 12594 186 12610 220
rect 7748 82 7782 144
rect 12756 82 12790 144
rect 7748 48 7844 82
rect 12694 48 12790 82
rect 14228 186 14244 220
rect 14312 186 14328 220
rect 14386 186 14402 220
rect 14470 186 14486 220
rect 14544 186 14560 220
rect 14628 186 14644 220
rect 14702 186 14718 220
rect 14786 186 14802 220
rect 14860 186 14876 220
rect 14944 186 14960 220
rect 15018 186 15034 220
rect 15102 186 15118 220
rect 15176 186 15192 220
rect 15260 186 15276 220
rect 15334 186 15350 220
rect 15418 186 15434 220
rect 15492 186 15508 220
rect 15576 186 15592 220
rect 15650 186 15666 220
rect 15734 186 15750 220
rect 15808 186 15824 220
rect 15892 186 15908 220
rect 15966 186 15982 220
rect 16050 186 16066 220
rect 16124 186 16140 220
rect 16208 186 16224 220
rect 16282 186 16298 220
rect 16366 186 16382 220
rect 16440 186 16456 220
rect 16524 186 16540 220
rect 16598 186 16614 220
rect 16682 186 16698 220
rect 16756 186 16772 220
rect 16840 186 16856 220
rect 16914 186 16930 220
rect 16998 186 17014 220
rect 17072 186 17088 220
rect 17156 186 17172 220
rect 17230 186 17246 220
rect 17314 186 17330 220
rect 17388 186 17404 220
rect 17472 186 17488 220
rect 17546 186 17562 220
rect 17630 186 17646 220
rect 17704 186 17720 220
rect 17788 186 17804 220
rect 17862 186 17878 220
rect 17946 186 17962 220
rect 18020 186 18036 220
rect 18104 186 18120 220
rect 18178 186 18194 220
rect 18262 186 18278 220
rect 18336 186 18352 220
rect 18420 186 18436 220
rect 18494 186 18510 220
rect 18578 186 18594 220
rect 18652 186 18668 220
rect 18736 186 18752 220
rect 18810 186 18826 220
rect 18894 186 18910 220
rect 14048 82 14082 144
rect 19056 82 19090 144
rect 14048 48 14144 82
rect 18994 48 19090 82
rect 20528 186 20544 220
rect 20612 186 20628 220
rect 20686 186 20702 220
rect 20770 186 20786 220
rect 20844 186 20860 220
rect 20928 186 20944 220
rect 21002 186 21018 220
rect 21086 186 21102 220
rect 21160 186 21176 220
rect 21244 186 21260 220
rect 21318 186 21334 220
rect 21402 186 21418 220
rect 21476 186 21492 220
rect 21560 186 21576 220
rect 21634 186 21650 220
rect 21718 186 21734 220
rect 21792 186 21808 220
rect 21876 186 21892 220
rect 21950 186 21966 220
rect 22034 186 22050 220
rect 22108 186 22124 220
rect 22192 186 22208 220
rect 22266 186 22282 220
rect 22350 186 22366 220
rect 22424 186 22440 220
rect 22508 186 22524 220
rect 22582 186 22598 220
rect 22666 186 22682 220
rect 22740 186 22756 220
rect 22824 186 22840 220
rect 22898 186 22914 220
rect 22982 186 22998 220
rect 23056 186 23072 220
rect 23140 186 23156 220
rect 23214 186 23230 220
rect 23298 186 23314 220
rect 23372 186 23388 220
rect 23456 186 23472 220
rect 23530 186 23546 220
rect 23614 186 23630 220
rect 23688 186 23704 220
rect 23772 186 23788 220
rect 23846 186 23862 220
rect 23930 186 23946 220
rect 24004 186 24020 220
rect 24088 186 24104 220
rect 24162 186 24178 220
rect 24246 186 24262 220
rect 24320 186 24336 220
rect 24404 186 24420 220
rect 24478 186 24494 220
rect 24562 186 24578 220
rect 24636 186 24652 220
rect 24720 186 24736 220
rect 24794 186 24810 220
rect 24878 186 24894 220
rect 24952 186 24968 220
rect 25036 186 25052 220
rect 25110 186 25126 220
rect 25194 186 25210 220
rect 20348 82 20382 144
rect 25356 82 25390 144
rect 20348 48 20444 82
rect 25294 48 25390 82
rect 1448 -566 1544 -532
rect 6394 -566 6490 -532
rect 1448 -628 1482 -566
rect 6456 -628 6490 -566
rect 1628 -704 1644 -670
rect 1712 -704 1728 -670
rect 1786 -704 1802 -670
rect 1870 -704 1886 -670
rect 1944 -704 1960 -670
rect 2028 -704 2044 -670
rect 2102 -704 2118 -670
rect 2186 -704 2202 -670
rect 2260 -704 2276 -670
rect 2344 -704 2360 -670
rect 2418 -704 2434 -670
rect 2502 -704 2518 -670
rect 2576 -704 2592 -670
rect 2660 -704 2676 -670
rect 2734 -704 2750 -670
rect 2818 -704 2834 -670
rect 2892 -704 2908 -670
rect 2976 -704 2992 -670
rect 3050 -704 3066 -670
rect 3134 -704 3150 -670
rect 3208 -704 3224 -670
rect 3292 -704 3308 -670
rect 3366 -704 3382 -670
rect 3450 -704 3466 -670
rect 3524 -704 3540 -670
rect 3608 -704 3624 -670
rect 3682 -704 3698 -670
rect 3766 -704 3782 -670
rect 3840 -704 3856 -670
rect 3924 -704 3940 -670
rect 3998 -704 4014 -670
rect 4082 -704 4098 -670
rect 4156 -704 4172 -670
rect 4240 -704 4256 -670
rect 4314 -704 4330 -670
rect 4398 -704 4414 -670
rect 4472 -704 4488 -670
rect 4556 -704 4572 -670
rect 4630 -704 4646 -670
rect 4714 -704 4730 -670
rect 4788 -704 4804 -670
rect 4872 -704 4888 -670
rect 4946 -704 4962 -670
rect 5030 -704 5046 -670
rect 5104 -704 5120 -670
rect 5188 -704 5204 -670
rect 5262 -704 5278 -670
rect 5346 -704 5362 -670
rect 5420 -704 5436 -670
rect 5504 -704 5520 -670
rect 5578 -704 5594 -670
rect 5662 -704 5678 -670
rect 5736 -704 5752 -670
rect 5820 -704 5836 -670
rect 5894 -704 5910 -670
rect 5978 -704 5994 -670
rect 6052 -704 6068 -670
rect 6136 -704 6152 -670
rect 6210 -704 6226 -670
rect 6294 -704 6310 -670
rect 7748 -566 7844 -532
rect 12694 -566 12790 -532
rect 7748 -628 7782 -566
rect 12756 -628 12790 -566
rect 7928 -704 7944 -670
rect 8012 -704 8028 -670
rect 8086 -704 8102 -670
rect 8170 -704 8186 -670
rect 8244 -704 8260 -670
rect 8328 -704 8344 -670
rect 8402 -704 8418 -670
rect 8486 -704 8502 -670
rect 8560 -704 8576 -670
rect 8644 -704 8660 -670
rect 8718 -704 8734 -670
rect 8802 -704 8818 -670
rect 8876 -704 8892 -670
rect 8960 -704 8976 -670
rect 9034 -704 9050 -670
rect 9118 -704 9134 -670
rect 9192 -704 9208 -670
rect 9276 -704 9292 -670
rect 9350 -704 9366 -670
rect 9434 -704 9450 -670
rect 9508 -704 9524 -670
rect 9592 -704 9608 -670
rect 9666 -704 9682 -670
rect 9750 -704 9766 -670
rect 9824 -704 9840 -670
rect 9908 -704 9924 -670
rect 9982 -704 9998 -670
rect 10066 -704 10082 -670
rect 10140 -704 10156 -670
rect 10224 -704 10240 -670
rect 10298 -704 10314 -670
rect 10382 -704 10398 -670
rect 10456 -704 10472 -670
rect 10540 -704 10556 -670
rect 10614 -704 10630 -670
rect 10698 -704 10714 -670
rect 10772 -704 10788 -670
rect 10856 -704 10872 -670
rect 10930 -704 10946 -670
rect 11014 -704 11030 -670
rect 11088 -704 11104 -670
rect 11172 -704 11188 -670
rect 11246 -704 11262 -670
rect 11330 -704 11346 -670
rect 11404 -704 11420 -670
rect 11488 -704 11504 -670
rect 11562 -704 11578 -670
rect 11646 -704 11662 -670
rect 11720 -704 11736 -670
rect 11804 -704 11820 -670
rect 11878 -704 11894 -670
rect 11962 -704 11978 -670
rect 12036 -704 12052 -670
rect 12120 -704 12136 -670
rect 12194 -704 12210 -670
rect 12278 -704 12294 -670
rect 12352 -704 12368 -670
rect 12436 -704 12452 -670
rect 12510 -704 12526 -670
rect 12594 -704 12610 -670
rect 14048 -566 14144 -532
rect 18994 -566 19090 -532
rect 14048 -628 14082 -566
rect 19056 -628 19090 -566
rect 14228 -704 14244 -670
rect 14312 -704 14328 -670
rect 14386 -704 14402 -670
rect 14470 -704 14486 -670
rect 14544 -704 14560 -670
rect 14628 -704 14644 -670
rect 14702 -704 14718 -670
rect 14786 -704 14802 -670
rect 14860 -704 14876 -670
rect 14944 -704 14960 -670
rect 15018 -704 15034 -670
rect 15102 -704 15118 -670
rect 15176 -704 15192 -670
rect 15260 -704 15276 -670
rect 15334 -704 15350 -670
rect 15418 -704 15434 -670
rect 15492 -704 15508 -670
rect 15576 -704 15592 -670
rect 15650 -704 15666 -670
rect 15734 -704 15750 -670
rect 15808 -704 15824 -670
rect 15892 -704 15908 -670
rect 15966 -704 15982 -670
rect 16050 -704 16066 -670
rect 16124 -704 16140 -670
rect 16208 -704 16224 -670
rect 16282 -704 16298 -670
rect 16366 -704 16382 -670
rect 16440 -704 16456 -670
rect 16524 -704 16540 -670
rect 16598 -704 16614 -670
rect 16682 -704 16698 -670
rect 16756 -704 16772 -670
rect 16840 -704 16856 -670
rect 16914 -704 16930 -670
rect 16998 -704 17014 -670
rect 17072 -704 17088 -670
rect 17156 -704 17172 -670
rect 17230 -704 17246 -670
rect 17314 -704 17330 -670
rect 17388 -704 17404 -670
rect 17472 -704 17488 -670
rect 17546 -704 17562 -670
rect 17630 -704 17646 -670
rect 17704 -704 17720 -670
rect 17788 -704 17804 -670
rect 17862 -704 17878 -670
rect 17946 -704 17962 -670
rect 18020 -704 18036 -670
rect 18104 -704 18120 -670
rect 18178 -704 18194 -670
rect 18262 -704 18278 -670
rect 18336 -704 18352 -670
rect 18420 -704 18436 -670
rect 18494 -704 18510 -670
rect 18578 -704 18594 -670
rect 18652 -704 18668 -670
rect 18736 -704 18752 -670
rect 18810 -704 18826 -670
rect 18894 -704 18910 -670
rect 20348 -566 20444 -532
rect 25294 -566 25390 -532
rect 20348 -628 20382 -566
rect 25356 -628 25390 -566
rect 20528 -704 20544 -670
rect 20612 -704 20628 -670
rect 20686 -704 20702 -670
rect 20770 -704 20786 -670
rect 20844 -704 20860 -670
rect 20928 -704 20944 -670
rect 21002 -704 21018 -670
rect 21086 -704 21102 -670
rect 21160 -704 21176 -670
rect 21244 -704 21260 -670
rect 21318 -704 21334 -670
rect 21402 -704 21418 -670
rect 21476 -704 21492 -670
rect 21560 -704 21576 -670
rect 21634 -704 21650 -670
rect 21718 -704 21734 -670
rect 21792 -704 21808 -670
rect 21876 -704 21892 -670
rect 21950 -704 21966 -670
rect 22034 -704 22050 -670
rect 22108 -704 22124 -670
rect 22192 -704 22208 -670
rect 22266 -704 22282 -670
rect 22350 -704 22366 -670
rect 22424 -704 22440 -670
rect 22508 -704 22524 -670
rect 22582 -704 22598 -670
rect 22666 -704 22682 -670
rect 22740 -704 22756 -670
rect 22824 -704 22840 -670
rect 22898 -704 22914 -670
rect 22982 -704 22998 -670
rect 23056 -704 23072 -670
rect 23140 -704 23156 -670
rect 23214 -704 23230 -670
rect 23298 -704 23314 -670
rect 23372 -704 23388 -670
rect 23456 -704 23472 -670
rect 23530 -704 23546 -670
rect 23614 -704 23630 -670
rect 23688 -704 23704 -670
rect 23772 -704 23788 -670
rect 23846 -704 23862 -670
rect 23930 -704 23946 -670
rect 24004 -704 24020 -670
rect 24088 -704 24104 -670
rect 24162 -704 24178 -670
rect 24246 -704 24262 -670
rect 24320 -704 24336 -670
rect 24404 -704 24420 -670
rect 24478 -704 24494 -670
rect 24562 -704 24578 -670
rect 24636 -704 24652 -670
rect 24720 -704 24736 -670
rect 24794 -704 24810 -670
rect 24878 -704 24894 -670
rect 24952 -704 24968 -670
rect 25036 -704 25052 -670
rect 25110 -704 25126 -670
rect 25194 -704 25210 -670
rect 1582 -754 1616 -738
rect 1582 -6746 1616 -6730
rect 1740 -754 1774 -738
rect 1740 -6746 1774 -6730
rect 1898 -754 1932 -738
rect 1898 -6746 1932 -6730
rect 2056 -754 2090 -738
rect 2056 -6746 2090 -6730
rect 2214 -754 2248 -738
rect 2214 -6746 2248 -6730
rect 2372 -754 2406 -738
rect 2372 -6746 2406 -6730
rect 2530 -754 2564 -738
rect 2530 -6746 2564 -6730
rect 2688 -754 2722 -738
rect 2688 -6746 2722 -6730
rect 2846 -754 2880 -738
rect 2846 -6746 2880 -6730
rect 3004 -754 3038 -738
rect 3004 -6746 3038 -6730
rect 3162 -754 3196 -738
rect 3162 -6746 3196 -6730
rect 3320 -754 3354 -738
rect 3320 -6746 3354 -6730
rect 3478 -754 3512 -738
rect 3478 -6746 3512 -6730
rect 3636 -754 3670 -738
rect 3636 -6746 3670 -6730
rect 3794 -754 3828 -738
rect 3794 -6746 3828 -6730
rect 3952 -754 3986 -738
rect 3952 -6746 3986 -6730
rect 4110 -754 4144 -738
rect 4110 -6746 4144 -6730
rect 4268 -754 4302 -738
rect 4268 -6746 4302 -6730
rect 4426 -754 4460 -738
rect 4426 -6746 4460 -6730
rect 4584 -754 4618 -738
rect 4584 -6746 4618 -6730
rect 4742 -754 4776 -738
rect 4742 -6746 4776 -6730
rect 4900 -754 4934 -738
rect 4900 -6746 4934 -6730
rect 5058 -754 5092 -738
rect 5058 -6746 5092 -6730
rect 5216 -754 5250 -738
rect 5216 -6746 5250 -6730
rect 5374 -754 5408 -738
rect 5374 -6746 5408 -6730
rect 5532 -754 5566 -738
rect 5532 -6746 5566 -6730
rect 5690 -754 5724 -738
rect 5690 -6746 5724 -6730
rect 5848 -754 5882 -738
rect 5848 -6746 5882 -6730
rect 6006 -754 6040 -738
rect 6006 -6746 6040 -6730
rect 6164 -754 6198 -738
rect 6164 -6746 6198 -6730
rect 6322 -754 6356 -738
rect 6322 -6746 6356 -6730
rect 7882 -754 7916 -738
rect 7882 -6746 7916 -6730
rect 8040 -754 8074 -738
rect 8040 -6746 8074 -6730
rect 8198 -754 8232 -738
rect 8198 -6746 8232 -6730
rect 8356 -754 8390 -738
rect 8356 -6746 8390 -6730
rect 8514 -754 8548 -738
rect 8514 -6746 8548 -6730
rect 8672 -754 8706 -738
rect 8672 -6746 8706 -6730
rect 8830 -754 8864 -738
rect 8830 -6746 8864 -6730
rect 8988 -754 9022 -738
rect 8988 -6746 9022 -6730
rect 9146 -754 9180 -738
rect 9146 -6746 9180 -6730
rect 9304 -754 9338 -738
rect 9304 -6746 9338 -6730
rect 9462 -754 9496 -738
rect 9462 -6746 9496 -6730
rect 9620 -754 9654 -738
rect 9620 -6746 9654 -6730
rect 9778 -754 9812 -738
rect 9778 -6746 9812 -6730
rect 9936 -754 9970 -738
rect 9936 -6746 9970 -6730
rect 10094 -754 10128 -738
rect 10094 -6746 10128 -6730
rect 10252 -754 10286 -738
rect 10252 -6746 10286 -6730
rect 10410 -754 10444 -738
rect 10410 -6746 10444 -6730
rect 10568 -754 10602 -738
rect 10568 -6746 10602 -6730
rect 10726 -754 10760 -738
rect 10726 -6746 10760 -6730
rect 10884 -754 10918 -738
rect 10884 -6746 10918 -6730
rect 11042 -754 11076 -738
rect 11042 -6746 11076 -6730
rect 11200 -754 11234 -738
rect 11200 -6746 11234 -6730
rect 11358 -754 11392 -738
rect 11358 -6746 11392 -6730
rect 11516 -754 11550 -738
rect 11516 -6746 11550 -6730
rect 11674 -754 11708 -738
rect 11674 -6746 11708 -6730
rect 11832 -754 11866 -738
rect 11832 -6746 11866 -6730
rect 11990 -754 12024 -738
rect 11990 -6746 12024 -6730
rect 12148 -754 12182 -738
rect 12148 -6746 12182 -6730
rect 12306 -754 12340 -738
rect 12306 -6746 12340 -6730
rect 12464 -754 12498 -738
rect 12464 -6746 12498 -6730
rect 12622 -754 12656 -738
rect 12622 -6746 12656 -6730
rect 14182 -754 14216 -738
rect 14182 -6746 14216 -6730
rect 14340 -754 14374 -738
rect 14340 -6746 14374 -6730
rect 14498 -754 14532 -738
rect 14498 -6746 14532 -6730
rect 14656 -754 14690 -738
rect 14656 -6746 14690 -6730
rect 14814 -754 14848 -738
rect 14814 -6746 14848 -6730
rect 14972 -754 15006 -738
rect 14972 -6746 15006 -6730
rect 15130 -754 15164 -738
rect 15130 -6746 15164 -6730
rect 15288 -754 15322 -738
rect 15288 -6746 15322 -6730
rect 15446 -754 15480 -738
rect 15446 -6746 15480 -6730
rect 15604 -754 15638 -738
rect 15604 -6746 15638 -6730
rect 15762 -754 15796 -738
rect 15762 -6746 15796 -6730
rect 15920 -754 15954 -738
rect 15920 -6746 15954 -6730
rect 16078 -754 16112 -738
rect 16078 -6746 16112 -6730
rect 16236 -754 16270 -738
rect 16236 -6746 16270 -6730
rect 16394 -754 16428 -738
rect 16394 -6746 16428 -6730
rect 16552 -754 16586 -738
rect 16552 -6746 16586 -6730
rect 16710 -754 16744 -738
rect 16710 -6746 16744 -6730
rect 16868 -754 16902 -738
rect 16868 -6746 16902 -6730
rect 17026 -754 17060 -738
rect 17026 -6746 17060 -6730
rect 17184 -754 17218 -738
rect 17184 -6746 17218 -6730
rect 17342 -754 17376 -738
rect 17342 -6746 17376 -6730
rect 17500 -754 17534 -738
rect 17500 -6746 17534 -6730
rect 17658 -754 17692 -738
rect 17658 -6746 17692 -6730
rect 17816 -754 17850 -738
rect 17816 -6746 17850 -6730
rect 17974 -754 18008 -738
rect 17974 -6746 18008 -6730
rect 18132 -754 18166 -738
rect 18132 -6746 18166 -6730
rect 18290 -754 18324 -738
rect 18290 -6746 18324 -6730
rect 18448 -754 18482 -738
rect 18448 -6746 18482 -6730
rect 18606 -754 18640 -738
rect 18606 -6746 18640 -6730
rect 18764 -754 18798 -738
rect 18764 -6746 18798 -6730
rect 18922 -754 18956 -738
rect 18922 -6746 18956 -6730
rect 20482 -754 20516 -738
rect 20482 -6746 20516 -6730
rect 20640 -754 20674 -738
rect 20640 -6746 20674 -6730
rect 20798 -754 20832 -738
rect 20798 -6746 20832 -6730
rect 20956 -754 20990 -738
rect 20956 -6746 20990 -6730
rect 21114 -754 21148 -738
rect 21114 -6746 21148 -6730
rect 21272 -754 21306 -738
rect 21272 -6746 21306 -6730
rect 21430 -754 21464 -738
rect 21430 -6746 21464 -6730
rect 21588 -754 21622 -738
rect 21588 -6746 21622 -6730
rect 21746 -754 21780 -738
rect 21746 -6746 21780 -6730
rect 21904 -754 21938 -738
rect 21904 -6746 21938 -6730
rect 22062 -754 22096 -738
rect 22062 -6746 22096 -6730
rect 22220 -754 22254 -738
rect 22220 -6746 22254 -6730
rect 22378 -754 22412 -738
rect 22378 -6746 22412 -6730
rect 22536 -754 22570 -738
rect 22536 -6746 22570 -6730
rect 22694 -754 22728 -738
rect 22694 -6746 22728 -6730
rect 22852 -754 22886 -738
rect 22852 -6746 22886 -6730
rect 23010 -754 23044 -738
rect 23010 -6746 23044 -6730
rect 23168 -754 23202 -738
rect 23168 -6746 23202 -6730
rect 23326 -754 23360 -738
rect 23326 -6746 23360 -6730
rect 23484 -754 23518 -738
rect 23484 -6746 23518 -6730
rect 23642 -754 23676 -738
rect 23642 -6746 23676 -6730
rect 23800 -754 23834 -738
rect 23800 -6746 23834 -6730
rect 23958 -754 23992 -738
rect 23958 -6746 23992 -6730
rect 24116 -754 24150 -738
rect 24116 -6746 24150 -6730
rect 24274 -754 24308 -738
rect 24274 -6746 24308 -6730
rect 24432 -754 24466 -738
rect 24432 -6746 24466 -6730
rect 24590 -754 24624 -738
rect 24590 -6746 24624 -6730
rect 24748 -754 24782 -738
rect 24748 -6746 24782 -6730
rect 24906 -754 24940 -738
rect 24906 -6746 24940 -6730
rect 25064 -754 25098 -738
rect 25064 -6746 25098 -6730
rect 25222 -754 25256 -738
rect 25222 -6746 25256 -6730
rect 1628 -6814 1644 -6780
rect 1712 -6814 1728 -6780
rect 1786 -6814 1802 -6780
rect 1870 -6814 1886 -6780
rect 1944 -6814 1960 -6780
rect 2028 -6814 2044 -6780
rect 2102 -6814 2118 -6780
rect 2186 -6814 2202 -6780
rect 2260 -6814 2276 -6780
rect 2344 -6814 2360 -6780
rect 2418 -6814 2434 -6780
rect 2502 -6814 2518 -6780
rect 2576 -6814 2592 -6780
rect 2660 -6814 2676 -6780
rect 2734 -6814 2750 -6780
rect 2818 -6814 2834 -6780
rect 2892 -6814 2908 -6780
rect 2976 -6814 2992 -6780
rect 3050 -6814 3066 -6780
rect 3134 -6814 3150 -6780
rect 3208 -6814 3224 -6780
rect 3292 -6814 3308 -6780
rect 3366 -6814 3382 -6780
rect 3450 -6814 3466 -6780
rect 3524 -6814 3540 -6780
rect 3608 -6814 3624 -6780
rect 3682 -6814 3698 -6780
rect 3766 -6814 3782 -6780
rect 3840 -6814 3856 -6780
rect 3924 -6814 3940 -6780
rect 3998 -6814 4014 -6780
rect 4082 -6814 4098 -6780
rect 4156 -6814 4172 -6780
rect 4240 -6814 4256 -6780
rect 4314 -6814 4330 -6780
rect 4398 -6814 4414 -6780
rect 4472 -6814 4488 -6780
rect 4556 -6814 4572 -6780
rect 4630 -6814 4646 -6780
rect 4714 -6814 4730 -6780
rect 4788 -6814 4804 -6780
rect 4872 -6814 4888 -6780
rect 4946 -6814 4962 -6780
rect 5030 -6814 5046 -6780
rect 5104 -6814 5120 -6780
rect 5188 -6814 5204 -6780
rect 5262 -6814 5278 -6780
rect 5346 -6814 5362 -6780
rect 5420 -6814 5436 -6780
rect 5504 -6814 5520 -6780
rect 5578 -6814 5594 -6780
rect 5662 -6814 5678 -6780
rect 5736 -6814 5752 -6780
rect 5820 -6814 5836 -6780
rect 5894 -6814 5910 -6780
rect 5978 -6814 5994 -6780
rect 6052 -6814 6068 -6780
rect 6136 -6814 6152 -6780
rect 6210 -6814 6226 -6780
rect 6294 -6814 6310 -6780
rect 1448 -6918 1482 -6856
rect 6456 -6918 6490 -6856
rect 1448 -6952 1544 -6918
rect 6394 -6952 6490 -6918
rect 7928 -6814 7944 -6780
rect 8012 -6814 8028 -6780
rect 8086 -6814 8102 -6780
rect 8170 -6814 8186 -6780
rect 8244 -6814 8260 -6780
rect 8328 -6814 8344 -6780
rect 8402 -6814 8418 -6780
rect 8486 -6814 8502 -6780
rect 8560 -6814 8576 -6780
rect 8644 -6814 8660 -6780
rect 8718 -6814 8734 -6780
rect 8802 -6814 8818 -6780
rect 8876 -6814 8892 -6780
rect 8960 -6814 8976 -6780
rect 9034 -6814 9050 -6780
rect 9118 -6814 9134 -6780
rect 9192 -6814 9208 -6780
rect 9276 -6814 9292 -6780
rect 9350 -6814 9366 -6780
rect 9434 -6814 9450 -6780
rect 9508 -6814 9524 -6780
rect 9592 -6814 9608 -6780
rect 9666 -6814 9682 -6780
rect 9750 -6814 9766 -6780
rect 9824 -6814 9840 -6780
rect 9908 -6814 9924 -6780
rect 9982 -6814 9998 -6780
rect 10066 -6814 10082 -6780
rect 10140 -6814 10156 -6780
rect 10224 -6814 10240 -6780
rect 10298 -6814 10314 -6780
rect 10382 -6814 10398 -6780
rect 10456 -6814 10472 -6780
rect 10540 -6814 10556 -6780
rect 10614 -6814 10630 -6780
rect 10698 -6814 10714 -6780
rect 10772 -6814 10788 -6780
rect 10856 -6814 10872 -6780
rect 10930 -6814 10946 -6780
rect 11014 -6814 11030 -6780
rect 11088 -6814 11104 -6780
rect 11172 -6814 11188 -6780
rect 11246 -6814 11262 -6780
rect 11330 -6814 11346 -6780
rect 11404 -6814 11420 -6780
rect 11488 -6814 11504 -6780
rect 11562 -6814 11578 -6780
rect 11646 -6814 11662 -6780
rect 11720 -6814 11736 -6780
rect 11804 -6814 11820 -6780
rect 11878 -6814 11894 -6780
rect 11962 -6814 11978 -6780
rect 12036 -6814 12052 -6780
rect 12120 -6814 12136 -6780
rect 12194 -6814 12210 -6780
rect 12278 -6814 12294 -6780
rect 12352 -6814 12368 -6780
rect 12436 -6814 12452 -6780
rect 12510 -6814 12526 -6780
rect 12594 -6814 12610 -6780
rect 7748 -6918 7782 -6856
rect 12756 -6918 12790 -6856
rect 7748 -6952 7844 -6918
rect 12694 -6952 12790 -6918
rect 14228 -6814 14244 -6780
rect 14312 -6814 14328 -6780
rect 14386 -6814 14402 -6780
rect 14470 -6814 14486 -6780
rect 14544 -6814 14560 -6780
rect 14628 -6814 14644 -6780
rect 14702 -6814 14718 -6780
rect 14786 -6814 14802 -6780
rect 14860 -6814 14876 -6780
rect 14944 -6814 14960 -6780
rect 15018 -6814 15034 -6780
rect 15102 -6814 15118 -6780
rect 15176 -6814 15192 -6780
rect 15260 -6814 15276 -6780
rect 15334 -6814 15350 -6780
rect 15418 -6814 15434 -6780
rect 15492 -6814 15508 -6780
rect 15576 -6814 15592 -6780
rect 15650 -6814 15666 -6780
rect 15734 -6814 15750 -6780
rect 15808 -6814 15824 -6780
rect 15892 -6814 15908 -6780
rect 15966 -6814 15982 -6780
rect 16050 -6814 16066 -6780
rect 16124 -6814 16140 -6780
rect 16208 -6814 16224 -6780
rect 16282 -6814 16298 -6780
rect 16366 -6814 16382 -6780
rect 16440 -6814 16456 -6780
rect 16524 -6814 16540 -6780
rect 16598 -6814 16614 -6780
rect 16682 -6814 16698 -6780
rect 16756 -6814 16772 -6780
rect 16840 -6814 16856 -6780
rect 16914 -6814 16930 -6780
rect 16998 -6814 17014 -6780
rect 17072 -6814 17088 -6780
rect 17156 -6814 17172 -6780
rect 17230 -6814 17246 -6780
rect 17314 -6814 17330 -6780
rect 17388 -6814 17404 -6780
rect 17472 -6814 17488 -6780
rect 17546 -6814 17562 -6780
rect 17630 -6814 17646 -6780
rect 17704 -6814 17720 -6780
rect 17788 -6814 17804 -6780
rect 17862 -6814 17878 -6780
rect 17946 -6814 17962 -6780
rect 18020 -6814 18036 -6780
rect 18104 -6814 18120 -6780
rect 18178 -6814 18194 -6780
rect 18262 -6814 18278 -6780
rect 18336 -6814 18352 -6780
rect 18420 -6814 18436 -6780
rect 18494 -6814 18510 -6780
rect 18578 -6814 18594 -6780
rect 18652 -6814 18668 -6780
rect 18736 -6814 18752 -6780
rect 18810 -6814 18826 -6780
rect 18894 -6814 18910 -6780
rect 14048 -6918 14082 -6856
rect 19056 -6918 19090 -6856
rect 14048 -6952 14144 -6918
rect 18994 -6952 19090 -6918
rect 20528 -6814 20544 -6780
rect 20612 -6814 20628 -6780
rect 20686 -6814 20702 -6780
rect 20770 -6814 20786 -6780
rect 20844 -6814 20860 -6780
rect 20928 -6814 20944 -6780
rect 21002 -6814 21018 -6780
rect 21086 -6814 21102 -6780
rect 21160 -6814 21176 -6780
rect 21244 -6814 21260 -6780
rect 21318 -6814 21334 -6780
rect 21402 -6814 21418 -6780
rect 21476 -6814 21492 -6780
rect 21560 -6814 21576 -6780
rect 21634 -6814 21650 -6780
rect 21718 -6814 21734 -6780
rect 21792 -6814 21808 -6780
rect 21876 -6814 21892 -6780
rect 21950 -6814 21966 -6780
rect 22034 -6814 22050 -6780
rect 22108 -6814 22124 -6780
rect 22192 -6814 22208 -6780
rect 22266 -6814 22282 -6780
rect 22350 -6814 22366 -6780
rect 22424 -6814 22440 -6780
rect 22508 -6814 22524 -6780
rect 22582 -6814 22598 -6780
rect 22666 -6814 22682 -6780
rect 22740 -6814 22756 -6780
rect 22824 -6814 22840 -6780
rect 22898 -6814 22914 -6780
rect 22982 -6814 22998 -6780
rect 23056 -6814 23072 -6780
rect 23140 -6814 23156 -6780
rect 23214 -6814 23230 -6780
rect 23298 -6814 23314 -6780
rect 23372 -6814 23388 -6780
rect 23456 -6814 23472 -6780
rect 23530 -6814 23546 -6780
rect 23614 -6814 23630 -6780
rect 23688 -6814 23704 -6780
rect 23772 -6814 23788 -6780
rect 23846 -6814 23862 -6780
rect 23930 -6814 23946 -6780
rect 24004 -6814 24020 -6780
rect 24088 -6814 24104 -6780
rect 24162 -6814 24178 -6780
rect 24246 -6814 24262 -6780
rect 24320 -6814 24336 -6780
rect 24404 -6814 24420 -6780
rect 24478 -6814 24494 -6780
rect 24562 -6814 24578 -6780
rect 24636 -6814 24652 -6780
rect 24720 -6814 24736 -6780
rect 24794 -6814 24810 -6780
rect 24878 -6814 24894 -6780
rect 24952 -6814 24968 -6780
rect 25036 -6814 25052 -6780
rect 25110 -6814 25126 -6780
rect 25194 -6814 25210 -6780
rect 20348 -6918 20382 -6856
rect 25356 -6918 25390 -6856
rect 20348 -6952 20444 -6918
rect 25294 -6952 25390 -6918
<< viali >>
rect 1636 6468 6359 6470
rect 7936 6468 12659 6470
rect 14236 6468 18959 6470
rect 20536 6468 25259 6470
rect 1636 6434 6359 6468
rect 1636 6432 6359 6434
rect 1644 6296 1712 6330
rect 1802 6296 1870 6330
rect 1960 6296 2028 6330
rect 2118 6296 2186 6330
rect 2276 6296 2344 6330
rect 2434 6296 2502 6330
rect 2592 6296 2660 6330
rect 2750 6296 2818 6330
rect 2908 6296 2976 6330
rect 3066 6296 3134 6330
rect 3224 6296 3292 6330
rect 3382 6296 3450 6330
rect 3540 6296 3608 6330
rect 3698 6296 3766 6330
rect 3856 6296 3924 6330
rect 4014 6296 4082 6330
rect 4172 6296 4240 6330
rect 4330 6296 4398 6330
rect 4488 6296 4556 6330
rect 4646 6296 4714 6330
rect 4804 6296 4872 6330
rect 4962 6296 5030 6330
rect 5120 6296 5188 6330
rect 5278 6296 5346 6330
rect 5436 6296 5504 6330
rect 5594 6296 5662 6330
rect 5752 6296 5820 6330
rect 5910 6296 5978 6330
rect 6068 6296 6136 6330
rect 6226 6296 6294 6330
rect 7936 6434 12659 6468
rect 7936 6432 12659 6434
rect 7944 6296 8012 6330
rect 8102 6296 8170 6330
rect 8260 6296 8328 6330
rect 8418 6296 8486 6330
rect 8576 6296 8644 6330
rect 8734 6296 8802 6330
rect 8892 6296 8960 6330
rect 9050 6296 9118 6330
rect 9208 6296 9276 6330
rect 9366 6296 9434 6330
rect 9524 6296 9592 6330
rect 9682 6296 9750 6330
rect 9840 6296 9908 6330
rect 9998 6296 10066 6330
rect 10156 6296 10224 6330
rect 10314 6296 10382 6330
rect 10472 6296 10540 6330
rect 10630 6296 10698 6330
rect 10788 6296 10856 6330
rect 10946 6296 11014 6330
rect 11104 6296 11172 6330
rect 11262 6296 11330 6330
rect 11420 6296 11488 6330
rect 11578 6296 11646 6330
rect 11736 6296 11804 6330
rect 11894 6296 11962 6330
rect 12052 6296 12120 6330
rect 12210 6296 12278 6330
rect 12368 6296 12436 6330
rect 12526 6296 12594 6330
rect 14236 6434 18959 6468
rect 14236 6432 18959 6434
rect 14244 6296 14312 6330
rect 14402 6296 14470 6330
rect 14560 6296 14628 6330
rect 14718 6296 14786 6330
rect 14876 6296 14944 6330
rect 15034 6296 15102 6330
rect 15192 6296 15260 6330
rect 15350 6296 15418 6330
rect 15508 6296 15576 6330
rect 15666 6296 15734 6330
rect 15824 6296 15892 6330
rect 15982 6296 16050 6330
rect 16140 6296 16208 6330
rect 16298 6296 16366 6330
rect 16456 6296 16524 6330
rect 16614 6296 16682 6330
rect 16772 6296 16840 6330
rect 16930 6296 16998 6330
rect 17088 6296 17156 6330
rect 17246 6296 17314 6330
rect 17404 6296 17472 6330
rect 17562 6296 17630 6330
rect 17720 6296 17788 6330
rect 17878 6296 17946 6330
rect 18036 6296 18104 6330
rect 18194 6296 18262 6330
rect 18352 6296 18420 6330
rect 18510 6296 18578 6330
rect 18668 6296 18736 6330
rect 18826 6296 18894 6330
rect 20536 6434 25259 6468
rect 20536 6432 25259 6434
rect 20544 6296 20612 6330
rect 20702 6296 20770 6330
rect 20860 6296 20928 6330
rect 21018 6296 21086 6330
rect 21176 6296 21244 6330
rect 21334 6296 21402 6330
rect 21492 6296 21560 6330
rect 21650 6296 21718 6330
rect 21808 6296 21876 6330
rect 21966 6296 22034 6330
rect 22124 6296 22192 6330
rect 22282 6296 22350 6330
rect 22440 6296 22508 6330
rect 22598 6296 22666 6330
rect 22756 6296 22824 6330
rect 22914 6296 22982 6330
rect 23072 6296 23140 6330
rect 23230 6296 23298 6330
rect 23388 6296 23456 6330
rect 23546 6296 23614 6330
rect 23704 6296 23772 6330
rect 23862 6296 23930 6330
rect 24020 6296 24088 6330
rect 24178 6296 24246 6330
rect 24336 6296 24404 6330
rect 24494 6296 24562 6330
rect 24652 6296 24720 6330
rect 24810 6296 24878 6330
rect 24968 6296 25036 6330
rect 25126 6296 25194 6330
rect 1446 236 1448 6280
rect 1448 236 1482 6280
rect 1482 236 1484 6280
rect 1582 270 1616 6246
rect 1740 270 1774 6246
rect 1898 270 1932 6246
rect 2056 270 2090 6246
rect 2214 270 2248 6246
rect 2372 270 2406 6246
rect 2530 270 2564 6246
rect 2688 270 2722 6246
rect 2846 270 2880 6246
rect 3004 270 3038 6246
rect 3162 270 3196 6246
rect 3320 270 3354 6246
rect 3478 270 3512 6246
rect 3636 270 3670 6246
rect 3794 270 3828 6246
rect 3952 270 3986 6246
rect 4110 270 4144 6246
rect 4268 270 4302 6246
rect 4426 270 4460 6246
rect 4584 270 4618 6246
rect 4742 270 4776 6246
rect 4900 270 4934 6246
rect 5058 270 5092 6246
rect 5216 270 5250 6246
rect 5374 270 5408 6246
rect 5532 270 5566 6246
rect 5690 270 5724 6246
rect 5848 270 5882 6246
rect 6006 270 6040 6246
rect 6164 270 6198 6246
rect 6322 270 6356 6246
rect 6454 236 6456 6280
rect 6456 236 6490 6280
rect 6490 236 6492 6280
rect 7746 236 7748 6280
rect 7748 236 7782 6280
rect 7782 236 7784 6280
rect 7882 270 7916 6246
rect 8040 270 8074 6246
rect 8198 270 8232 6246
rect 8356 270 8390 6246
rect 8514 270 8548 6246
rect 8672 270 8706 6246
rect 8830 270 8864 6246
rect 8988 270 9022 6246
rect 9146 270 9180 6246
rect 9304 270 9338 6246
rect 9462 270 9496 6246
rect 9620 270 9654 6246
rect 9778 270 9812 6246
rect 9936 270 9970 6246
rect 10094 270 10128 6246
rect 10252 270 10286 6246
rect 10410 270 10444 6246
rect 10568 270 10602 6246
rect 10726 270 10760 6246
rect 10884 270 10918 6246
rect 11042 270 11076 6246
rect 11200 270 11234 6246
rect 11358 270 11392 6246
rect 11516 270 11550 6246
rect 11674 270 11708 6246
rect 11832 270 11866 6246
rect 11990 270 12024 6246
rect 12148 270 12182 6246
rect 12306 270 12340 6246
rect 12464 270 12498 6246
rect 12622 270 12656 6246
rect 12754 236 12756 6280
rect 12756 236 12790 6280
rect 12790 236 12792 6280
rect 14046 236 14048 6280
rect 14048 236 14082 6280
rect 14082 236 14084 6280
rect 14182 270 14216 6246
rect 14340 270 14374 6246
rect 14498 270 14532 6246
rect 14656 270 14690 6246
rect 14814 270 14848 6246
rect 14972 270 15006 6246
rect 15130 270 15164 6246
rect 15288 270 15322 6246
rect 15446 270 15480 6246
rect 15604 270 15638 6246
rect 15762 270 15796 6246
rect 15920 270 15954 6246
rect 16078 270 16112 6246
rect 16236 270 16270 6246
rect 16394 270 16428 6246
rect 16552 270 16586 6246
rect 16710 270 16744 6246
rect 16868 270 16902 6246
rect 17026 270 17060 6246
rect 17184 270 17218 6246
rect 17342 270 17376 6246
rect 17500 270 17534 6246
rect 17658 270 17692 6246
rect 17816 270 17850 6246
rect 17974 270 18008 6246
rect 18132 270 18166 6246
rect 18290 270 18324 6246
rect 18448 270 18482 6246
rect 18606 270 18640 6246
rect 18764 270 18798 6246
rect 18922 270 18956 6246
rect 19054 236 19056 6280
rect 19056 236 19090 6280
rect 19090 236 19092 6280
rect 20346 236 20348 6280
rect 20348 236 20382 6280
rect 20382 236 20384 6280
rect 20482 270 20516 6246
rect 20640 270 20674 6246
rect 20798 270 20832 6246
rect 20956 270 20990 6246
rect 21114 270 21148 6246
rect 21272 270 21306 6246
rect 21430 270 21464 6246
rect 21588 270 21622 6246
rect 21746 270 21780 6246
rect 21904 270 21938 6246
rect 22062 270 22096 6246
rect 22220 270 22254 6246
rect 22378 270 22412 6246
rect 22536 270 22570 6246
rect 22694 270 22728 6246
rect 22852 270 22886 6246
rect 23010 270 23044 6246
rect 23168 270 23202 6246
rect 23326 270 23360 6246
rect 23484 270 23518 6246
rect 23642 270 23676 6246
rect 23800 270 23834 6246
rect 23958 270 23992 6246
rect 24116 270 24150 6246
rect 24274 270 24308 6246
rect 24432 270 24466 6246
rect 24590 270 24624 6246
rect 24748 270 24782 6246
rect 24906 270 24940 6246
rect 25064 270 25098 6246
rect 25222 270 25256 6246
rect 25354 236 25356 6280
rect 25356 236 25390 6280
rect 25390 236 25392 6280
rect 1644 186 1712 220
rect 1802 186 1870 220
rect 1960 186 2028 220
rect 2118 186 2186 220
rect 2276 186 2344 220
rect 2434 186 2502 220
rect 2592 186 2660 220
rect 2750 186 2818 220
rect 2908 186 2976 220
rect 3066 186 3134 220
rect 3224 186 3292 220
rect 3382 186 3450 220
rect 3540 186 3608 220
rect 3698 186 3766 220
rect 3856 186 3924 220
rect 4014 186 4082 220
rect 4172 186 4240 220
rect 4330 186 4398 220
rect 4488 186 4556 220
rect 4646 186 4714 220
rect 4804 186 4872 220
rect 4962 186 5030 220
rect 5120 186 5188 220
rect 5278 186 5346 220
rect 5436 186 5504 220
rect 5594 186 5662 220
rect 5752 186 5820 220
rect 5910 186 5978 220
rect 6068 186 6136 220
rect 6226 186 6294 220
rect 1636 82 6302 84
rect 1636 48 6302 82
rect 7944 186 8012 220
rect 8102 186 8170 220
rect 8260 186 8328 220
rect 8418 186 8486 220
rect 8576 186 8644 220
rect 8734 186 8802 220
rect 8892 186 8960 220
rect 9050 186 9118 220
rect 9208 186 9276 220
rect 9366 186 9434 220
rect 9524 186 9592 220
rect 9682 186 9750 220
rect 9840 186 9908 220
rect 9998 186 10066 220
rect 10156 186 10224 220
rect 10314 186 10382 220
rect 10472 186 10540 220
rect 10630 186 10698 220
rect 10788 186 10856 220
rect 10946 186 11014 220
rect 11104 186 11172 220
rect 11262 186 11330 220
rect 11420 186 11488 220
rect 11578 186 11646 220
rect 11736 186 11804 220
rect 11894 186 11962 220
rect 12052 186 12120 220
rect 12210 186 12278 220
rect 12368 186 12436 220
rect 12526 186 12594 220
rect 7936 82 12602 84
rect 7936 48 12602 82
rect 14244 186 14312 220
rect 14402 186 14470 220
rect 14560 186 14628 220
rect 14718 186 14786 220
rect 14876 186 14944 220
rect 15034 186 15102 220
rect 15192 186 15260 220
rect 15350 186 15418 220
rect 15508 186 15576 220
rect 15666 186 15734 220
rect 15824 186 15892 220
rect 15982 186 16050 220
rect 16140 186 16208 220
rect 16298 186 16366 220
rect 16456 186 16524 220
rect 16614 186 16682 220
rect 16772 186 16840 220
rect 16930 186 16998 220
rect 17088 186 17156 220
rect 17246 186 17314 220
rect 17404 186 17472 220
rect 17562 186 17630 220
rect 17720 186 17788 220
rect 17878 186 17946 220
rect 18036 186 18104 220
rect 18194 186 18262 220
rect 18352 186 18420 220
rect 18510 186 18578 220
rect 18668 186 18736 220
rect 18826 186 18894 220
rect 14236 82 18902 84
rect 14236 48 18902 82
rect 20544 186 20612 220
rect 20702 186 20770 220
rect 20860 186 20928 220
rect 21018 186 21086 220
rect 21176 186 21244 220
rect 21334 186 21402 220
rect 21492 186 21560 220
rect 21650 186 21718 220
rect 21808 186 21876 220
rect 21966 186 22034 220
rect 22124 186 22192 220
rect 22282 186 22350 220
rect 22440 186 22508 220
rect 22598 186 22666 220
rect 22756 186 22824 220
rect 22914 186 22982 220
rect 23072 186 23140 220
rect 23230 186 23298 220
rect 23388 186 23456 220
rect 23546 186 23614 220
rect 23704 186 23772 220
rect 23862 186 23930 220
rect 24020 186 24088 220
rect 24178 186 24246 220
rect 24336 186 24404 220
rect 24494 186 24562 220
rect 24652 186 24720 220
rect 24810 186 24878 220
rect 24968 186 25036 220
rect 25126 186 25194 220
rect 20536 82 25202 84
rect 20536 48 25202 82
rect 1636 46 6302 48
rect 7936 46 12602 48
rect 14236 46 18902 48
rect 20536 46 25202 48
rect 1636 -532 6359 -530
rect 7936 -532 12659 -530
rect 14236 -532 18959 -530
rect 20536 -532 25259 -530
rect 1636 -566 6359 -532
rect 1636 -568 6359 -566
rect 1644 -704 1712 -670
rect 1802 -704 1870 -670
rect 1960 -704 2028 -670
rect 2118 -704 2186 -670
rect 2276 -704 2344 -670
rect 2434 -704 2502 -670
rect 2592 -704 2660 -670
rect 2750 -704 2818 -670
rect 2908 -704 2976 -670
rect 3066 -704 3134 -670
rect 3224 -704 3292 -670
rect 3382 -704 3450 -670
rect 3540 -704 3608 -670
rect 3698 -704 3766 -670
rect 3856 -704 3924 -670
rect 4014 -704 4082 -670
rect 4172 -704 4240 -670
rect 4330 -704 4398 -670
rect 4488 -704 4556 -670
rect 4646 -704 4714 -670
rect 4804 -704 4872 -670
rect 4962 -704 5030 -670
rect 5120 -704 5188 -670
rect 5278 -704 5346 -670
rect 5436 -704 5504 -670
rect 5594 -704 5662 -670
rect 5752 -704 5820 -670
rect 5910 -704 5978 -670
rect 6068 -704 6136 -670
rect 6226 -704 6294 -670
rect 7936 -566 12659 -532
rect 7936 -568 12659 -566
rect 7944 -704 8012 -670
rect 8102 -704 8170 -670
rect 8260 -704 8328 -670
rect 8418 -704 8486 -670
rect 8576 -704 8644 -670
rect 8734 -704 8802 -670
rect 8892 -704 8960 -670
rect 9050 -704 9118 -670
rect 9208 -704 9276 -670
rect 9366 -704 9434 -670
rect 9524 -704 9592 -670
rect 9682 -704 9750 -670
rect 9840 -704 9908 -670
rect 9998 -704 10066 -670
rect 10156 -704 10224 -670
rect 10314 -704 10382 -670
rect 10472 -704 10540 -670
rect 10630 -704 10698 -670
rect 10788 -704 10856 -670
rect 10946 -704 11014 -670
rect 11104 -704 11172 -670
rect 11262 -704 11330 -670
rect 11420 -704 11488 -670
rect 11578 -704 11646 -670
rect 11736 -704 11804 -670
rect 11894 -704 11962 -670
rect 12052 -704 12120 -670
rect 12210 -704 12278 -670
rect 12368 -704 12436 -670
rect 12526 -704 12594 -670
rect 14236 -566 18959 -532
rect 14236 -568 18959 -566
rect 14244 -704 14312 -670
rect 14402 -704 14470 -670
rect 14560 -704 14628 -670
rect 14718 -704 14786 -670
rect 14876 -704 14944 -670
rect 15034 -704 15102 -670
rect 15192 -704 15260 -670
rect 15350 -704 15418 -670
rect 15508 -704 15576 -670
rect 15666 -704 15734 -670
rect 15824 -704 15892 -670
rect 15982 -704 16050 -670
rect 16140 -704 16208 -670
rect 16298 -704 16366 -670
rect 16456 -704 16524 -670
rect 16614 -704 16682 -670
rect 16772 -704 16840 -670
rect 16930 -704 16998 -670
rect 17088 -704 17156 -670
rect 17246 -704 17314 -670
rect 17404 -704 17472 -670
rect 17562 -704 17630 -670
rect 17720 -704 17788 -670
rect 17878 -704 17946 -670
rect 18036 -704 18104 -670
rect 18194 -704 18262 -670
rect 18352 -704 18420 -670
rect 18510 -704 18578 -670
rect 18668 -704 18736 -670
rect 18826 -704 18894 -670
rect 20536 -566 25259 -532
rect 20536 -568 25259 -566
rect 20544 -704 20612 -670
rect 20702 -704 20770 -670
rect 20860 -704 20928 -670
rect 21018 -704 21086 -670
rect 21176 -704 21244 -670
rect 21334 -704 21402 -670
rect 21492 -704 21560 -670
rect 21650 -704 21718 -670
rect 21808 -704 21876 -670
rect 21966 -704 22034 -670
rect 22124 -704 22192 -670
rect 22282 -704 22350 -670
rect 22440 -704 22508 -670
rect 22598 -704 22666 -670
rect 22756 -704 22824 -670
rect 22914 -704 22982 -670
rect 23072 -704 23140 -670
rect 23230 -704 23298 -670
rect 23388 -704 23456 -670
rect 23546 -704 23614 -670
rect 23704 -704 23772 -670
rect 23862 -704 23930 -670
rect 24020 -704 24088 -670
rect 24178 -704 24246 -670
rect 24336 -704 24404 -670
rect 24494 -704 24562 -670
rect 24652 -704 24720 -670
rect 24810 -704 24878 -670
rect 24968 -704 25036 -670
rect 25126 -704 25194 -670
rect 1446 -6764 1448 -720
rect 1448 -6764 1482 -720
rect 1482 -6764 1484 -720
rect 1582 -6730 1616 -754
rect 1740 -6730 1774 -754
rect 1898 -6730 1932 -754
rect 2056 -6730 2090 -754
rect 2214 -6730 2248 -754
rect 2372 -6730 2406 -754
rect 2530 -6730 2564 -754
rect 2688 -6730 2722 -754
rect 2846 -6730 2880 -754
rect 3004 -6730 3038 -754
rect 3162 -6730 3196 -754
rect 3320 -6730 3354 -754
rect 3478 -6730 3512 -754
rect 3636 -6730 3670 -754
rect 3794 -6730 3828 -754
rect 3952 -6730 3986 -754
rect 4110 -6730 4144 -754
rect 4268 -6730 4302 -754
rect 4426 -6730 4460 -754
rect 4584 -6730 4618 -754
rect 4742 -6730 4776 -754
rect 4900 -6730 4934 -754
rect 5058 -6730 5092 -754
rect 5216 -6730 5250 -754
rect 5374 -6730 5408 -754
rect 5532 -6730 5566 -754
rect 5690 -6730 5724 -754
rect 5848 -6730 5882 -754
rect 6006 -6730 6040 -754
rect 6164 -6730 6198 -754
rect 6322 -6730 6356 -754
rect 6454 -6764 6456 -720
rect 6456 -6764 6490 -720
rect 6490 -6764 6492 -720
rect 7746 -6764 7748 -720
rect 7748 -6764 7782 -720
rect 7782 -6764 7784 -720
rect 7882 -6730 7916 -754
rect 8040 -6730 8074 -754
rect 8198 -6730 8232 -754
rect 8356 -6730 8390 -754
rect 8514 -6730 8548 -754
rect 8672 -6730 8706 -754
rect 8830 -6730 8864 -754
rect 8988 -6730 9022 -754
rect 9146 -6730 9180 -754
rect 9304 -6730 9338 -754
rect 9462 -6730 9496 -754
rect 9620 -6730 9654 -754
rect 9778 -6730 9812 -754
rect 9936 -6730 9970 -754
rect 10094 -6730 10128 -754
rect 10252 -6730 10286 -754
rect 10410 -6730 10444 -754
rect 10568 -6730 10602 -754
rect 10726 -6730 10760 -754
rect 10884 -6730 10918 -754
rect 11042 -6730 11076 -754
rect 11200 -6730 11234 -754
rect 11358 -6730 11392 -754
rect 11516 -6730 11550 -754
rect 11674 -6730 11708 -754
rect 11832 -6730 11866 -754
rect 11990 -6730 12024 -754
rect 12148 -6730 12182 -754
rect 12306 -6730 12340 -754
rect 12464 -6730 12498 -754
rect 12622 -6730 12656 -754
rect 12754 -6764 12756 -720
rect 12756 -6764 12790 -720
rect 12790 -6764 12792 -720
rect 14046 -6764 14048 -720
rect 14048 -6764 14082 -720
rect 14082 -6764 14084 -720
rect 14182 -6730 14216 -754
rect 14340 -6730 14374 -754
rect 14498 -6730 14532 -754
rect 14656 -6730 14690 -754
rect 14814 -6730 14848 -754
rect 14972 -6730 15006 -754
rect 15130 -6730 15164 -754
rect 15288 -6730 15322 -754
rect 15446 -6730 15480 -754
rect 15604 -6730 15638 -754
rect 15762 -6730 15796 -754
rect 15920 -6730 15954 -754
rect 16078 -6730 16112 -754
rect 16236 -6730 16270 -754
rect 16394 -6730 16428 -754
rect 16552 -6730 16586 -754
rect 16710 -6730 16744 -754
rect 16868 -6730 16902 -754
rect 17026 -6730 17060 -754
rect 17184 -6730 17218 -754
rect 17342 -6730 17376 -754
rect 17500 -6730 17534 -754
rect 17658 -6730 17692 -754
rect 17816 -6730 17850 -754
rect 17974 -6730 18008 -754
rect 18132 -6730 18166 -754
rect 18290 -6730 18324 -754
rect 18448 -6730 18482 -754
rect 18606 -6730 18640 -754
rect 18764 -6730 18798 -754
rect 18922 -6730 18956 -754
rect 19054 -6764 19056 -720
rect 19056 -6764 19090 -720
rect 19090 -6764 19092 -720
rect 20346 -6764 20348 -720
rect 20348 -6764 20382 -720
rect 20382 -6764 20384 -720
rect 20482 -6730 20516 -754
rect 20640 -6730 20674 -754
rect 20798 -6730 20832 -754
rect 20956 -6730 20990 -754
rect 21114 -6730 21148 -754
rect 21272 -6730 21306 -754
rect 21430 -6730 21464 -754
rect 21588 -6730 21622 -754
rect 21746 -6730 21780 -754
rect 21904 -6730 21938 -754
rect 22062 -6730 22096 -754
rect 22220 -6730 22254 -754
rect 22378 -6730 22412 -754
rect 22536 -6730 22570 -754
rect 22694 -6730 22728 -754
rect 22852 -6730 22886 -754
rect 23010 -6730 23044 -754
rect 23168 -6730 23202 -754
rect 23326 -6730 23360 -754
rect 23484 -6730 23518 -754
rect 23642 -6730 23676 -754
rect 23800 -6730 23834 -754
rect 23958 -6730 23992 -754
rect 24116 -6730 24150 -754
rect 24274 -6730 24308 -754
rect 24432 -6730 24466 -754
rect 24590 -6730 24624 -754
rect 24748 -6730 24782 -754
rect 24906 -6730 24940 -754
rect 25064 -6730 25098 -754
rect 25222 -6730 25256 -754
rect 25354 -6764 25356 -720
rect 25356 -6764 25390 -720
rect 25390 -6764 25392 -720
rect 1644 -6814 1712 -6780
rect 1802 -6814 1870 -6780
rect 1960 -6814 2028 -6780
rect 2118 -6814 2186 -6780
rect 2276 -6814 2344 -6780
rect 2434 -6814 2502 -6780
rect 2592 -6814 2660 -6780
rect 2750 -6814 2818 -6780
rect 2908 -6814 2976 -6780
rect 3066 -6814 3134 -6780
rect 3224 -6814 3292 -6780
rect 3382 -6814 3450 -6780
rect 3540 -6814 3608 -6780
rect 3698 -6814 3766 -6780
rect 3856 -6814 3924 -6780
rect 4014 -6814 4082 -6780
rect 4172 -6814 4240 -6780
rect 4330 -6814 4398 -6780
rect 4488 -6814 4556 -6780
rect 4646 -6814 4714 -6780
rect 4804 -6814 4872 -6780
rect 4962 -6814 5030 -6780
rect 5120 -6814 5188 -6780
rect 5278 -6814 5346 -6780
rect 5436 -6814 5504 -6780
rect 5594 -6814 5662 -6780
rect 5752 -6814 5820 -6780
rect 5910 -6814 5978 -6780
rect 6068 -6814 6136 -6780
rect 6226 -6814 6294 -6780
rect 1636 -6918 6302 -6916
rect 1636 -6952 6302 -6918
rect 7944 -6814 8012 -6780
rect 8102 -6814 8170 -6780
rect 8260 -6814 8328 -6780
rect 8418 -6814 8486 -6780
rect 8576 -6814 8644 -6780
rect 8734 -6814 8802 -6780
rect 8892 -6814 8960 -6780
rect 9050 -6814 9118 -6780
rect 9208 -6814 9276 -6780
rect 9366 -6814 9434 -6780
rect 9524 -6814 9592 -6780
rect 9682 -6814 9750 -6780
rect 9840 -6814 9908 -6780
rect 9998 -6814 10066 -6780
rect 10156 -6814 10224 -6780
rect 10314 -6814 10382 -6780
rect 10472 -6814 10540 -6780
rect 10630 -6814 10698 -6780
rect 10788 -6814 10856 -6780
rect 10946 -6814 11014 -6780
rect 11104 -6814 11172 -6780
rect 11262 -6814 11330 -6780
rect 11420 -6814 11488 -6780
rect 11578 -6814 11646 -6780
rect 11736 -6814 11804 -6780
rect 11894 -6814 11962 -6780
rect 12052 -6814 12120 -6780
rect 12210 -6814 12278 -6780
rect 12368 -6814 12436 -6780
rect 12526 -6814 12594 -6780
rect 7936 -6918 12602 -6916
rect 7936 -6952 12602 -6918
rect 14244 -6814 14312 -6780
rect 14402 -6814 14470 -6780
rect 14560 -6814 14628 -6780
rect 14718 -6814 14786 -6780
rect 14876 -6814 14944 -6780
rect 15034 -6814 15102 -6780
rect 15192 -6814 15260 -6780
rect 15350 -6814 15418 -6780
rect 15508 -6814 15576 -6780
rect 15666 -6814 15734 -6780
rect 15824 -6814 15892 -6780
rect 15982 -6814 16050 -6780
rect 16140 -6814 16208 -6780
rect 16298 -6814 16366 -6780
rect 16456 -6814 16524 -6780
rect 16614 -6814 16682 -6780
rect 16772 -6814 16840 -6780
rect 16930 -6814 16998 -6780
rect 17088 -6814 17156 -6780
rect 17246 -6814 17314 -6780
rect 17404 -6814 17472 -6780
rect 17562 -6814 17630 -6780
rect 17720 -6814 17788 -6780
rect 17878 -6814 17946 -6780
rect 18036 -6814 18104 -6780
rect 18194 -6814 18262 -6780
rect 18352 -6814 18420 -6780
rect 18510 -6814 18578 -6780
rect 18668 -6814 18736 -6780
rect 18826 -6814 18894 -6780
rect 14236 -6918 18902 -6916
rect 14236 -6952 18902 -6918
rect 20544 -6814 20612 -6780
rect 20702 -6814 20770 -6780
rect 20860 -6814 20928 -6780
rect 21018 -6814 21086 -6780
rect 21176 -6814 21244 -6780
rect 21334 -6814 21402 -6780
rect 21492 -6814 21560 -6780
rect 21650 -6814 21718 -6780
rect 21808 -6814 21876 -6780
rect 21966 -6814 22034 -6780
rect 22124 -6814 22192 -6780
rect 22282 -6814 22350 -6780
rect 22440 -6814 22508 -6780
rect 22598 -6814 22666 -6780
rect 22756 -6814 22824 -6780
rect 22914 -6814 22982 -6780
rect 23072 -6814 23140 -6780
rect 23230 -6814 23298 -6780
rect 23388 -6814 23456 -6780
rect 23546 -6814 23614 -6780
rect 23704 -6814 23772 -6780
rect 23862 -6814 23930 -6780
rect 24020 -6814 24088 -6780
rect 24178 -6814 24246 -6780
rect 24336 -6814 24404 -6780
rect 24494 -6814 24562 -6780
rect 24652 -6814 24720 -6780
rect 24810 -6814 24878 -6780
rect 24968 -6814 25036 -6780
rect 25126 -6814 25194 -6780
rect 20536 -6918 25202 -6916
rect 20536 -6952 25202 -6918
rect 1636 -6954 6302 -6952
rect 7936 -6954 12602 -6952
rect 14236 -6954 18902 -6952
rect 20536 -6954 25202 -6952
<< metal1 >>
rect 1430 6470 6510 6480
rect 1430 6432 1636 6470
rect 6359 6432 6510 6470
rect 1430 6422 6510 6432
rect 1430 6420 1500 6422
rect 6440 6420 6510 6422
rect 1632 6330 1652 6390
rect 6286 6330 6306 6390
rect 1632 6296 1644 6330
rect 6294 6296 6306 6330
rect 1632 6290 1652 6296
rect 6286 6290 6306 6296
rect 1565 6246 1631 6258
rect 1565 6238 1582 6246
rect 1616 6238 1631 6246
rect 1565 270 1582 278
rect 1616 270 1631 278
rect 1565 258 1631 270
rect 1723 6246 1789 6258
rect 1723 6238 1740 6246
rect 1774 6238 1789 6246
rect 1723 270 1740 278
rect 1774 270 1789 278
rect 1723 258 1789 270
rect 1881 6246 1947 6258
rect 1881 6238 1898 6246
rect 1932 6238 1947 6246
rect 1881 270 1898 278
rect 1932 270 1947 278
rect 1881 258 1947 270
rect 2039 6246 2105 6258
rect 2039 6238 2056 6246
rect 2090 6238 2105 6246
rect 2039 270 2056 278
rect 2090 270 2105 278
rect 2039 258 2105 270
rect 2197 6246 2263 6258
rect 2197 6238 2214 6246
rect 2248 6238 2263 6246
rect 2197 270 2214 278
rect 2248 270 2263 278
rect 2197 258 2263 270
rect 2355 6246 2421 6258
rect 2355 6238 2372 6246
rect 2406 6238 2421 6246
rect 2355 270 2372 278
rect 2406 270 2421 278
rect 2355 258 2421 270
rect 2513 6246 2579 6258
rect 2513 6238 2530 6246
rect 2564 6238 2579 6246
rect 2513 270 2530 278
rect 2564 270 2579 278
rect 2513 258 2579 270
rect 2671 6246 2737 6258
rect 2671 6238 2688 6246
rect 2722 6238 2737 6246
rect 2671 270 2688 278
rect 2722 270 2737 278
rect 2671 258 2737 270
rect 2829 6246 2895 6258
rect 2829 6238 2846 6246
rect 2880 6238 2895 6246
rect 2829 270 2846 278
rect 2880 270 2895 278
rect 2829 258 2895 270
rect 2987 6246 3053 6258
rect 2987 6238 3004 6246
rect 3038 6238 3053 6246
rect 2987 270 3004 278
rect 3038 270 3053 278
rect 2987 258 3053 270
rect 3145 6246 3211 6258
rect 3145 6238 3162 6246
rect 3196 6238 3211 6246
rect 3145 270 3162 278
rect 3196 270 3211 278
rect 3145 258 3211 270
rect 3303 6246 3369 6258
rect 3303 6238 3320 6246
rect 3354 6238 3369 6246
rect 3303 270 3320 278
rect 3354 270 3369 278
rect 3303 258 3369 270
rect 3461 6246 3527 6258
rect 3461 6238 3478 6246
rect 3512 6238 3527 6246
rect 3461 270 3478 278
rect 3512 270 3527 278
rect 3461 258 3527 270
rect 3619 6246 3685 6258
rect 3619 6238 3636 6246
rect 3670 6238 3685 6246
rect 3619 270 3636 278
rect 3670 270 3685 278
rect 3619 258 3685 270
rect 3777 6246 3843 6258
rect 3777 6238 3794 6246
rect 3828 6238 3843 6246
rect 3777 270 3794 278
rect 3828 270 3843 278
rect 3777 258 3843 270
rect 3935 6246 4001 6258
rect 3935 6238 3952 6246
rect 3986 6238 4001 6246
rect 3935 270 3952 278
rect 3986 270 4001 278
rect 3935 258 4001 270
rect 4093 6246 4159 6258
rect 4093 6238 4110 6246
rect 4144 6238 4159 6246
rect 4093 270 4110 278
rect 4144 270 4159 278
rect 4093 258 4159 270
rect 4251 6246 4317 6258
rect 4251 6238 4268 6246
rect 4302 6238 4317 6246
rect 4251 270 4268 278
rect 4302 270 4317 278
rect 4251 258 4317 270
rect 4409 6246 4475 6258
rect 4409 6238 4426 6246
rect 4460 6238 4475 6246
rect 4409 270 4426 278
rect 4460 270 4475 278
rect 4409 258 4475 270
rect 4567 6246 4633 6258
rect 4567 6238 4584 6246
rect 4618 6238 4633 6246
rect 4567 270 4584 278
rect 4618 270 4633 278
rect 4567 258 4633 270
rect 4725 6246 4791 6258
rect 4725 6238 4742 6246
rect 4776 6238 4791 6246
rect 4725 270 4742 278
rect 4776 270 4791 278
rect 4725 258 4791 270
rect 4883 6246 4949 6258
rect 4883 6238 4900 6246
rect 4934 6238 4949 6246
rect 4883 270 4900 278
rect 4934 270 4949 278
rect 4883 258 4949 270
rect 5041 6246 5107 6258
rect 5041 6238 5058 6246
rect 5092 6238 5107 6246
rect 5041 270 5058 278
rect 5092 270 5107 278
rect 5041 258 5107 270
rect 5199 6246 5265 6258
rect 5199 6238 5216 6246
rect 5250 6238 5265 6246
rect 5199 270 5216 278
rect 5250 270 5265 278
rect 5199 258 5265 270
rect 5357 6246 5423 6258
rect 5357 6238 5374 6246
rect 5408 6238 5423 6246
rect 5357 270 5374 278
rect 5408 270 5423 278
rect 5357 258 5423 270
rect 5515 6246 5581 6258
rect 5515 6238 5532 6246
rect 5566 6238 5581 6246
rect 5515 270 5532 278
rect 5566 270 5581 278
rect 5515 258 5581 270
rect 5673 6246 5739 6258
rect 5673 6238 5690 6246
rect 5724 6238 5739 6246
rect 5673 270 5690 278
rect 5724 270 5739 278
rect 5673 258 5739 270
rect 5831 6246 5897 6258
rect 5831 6238 5848 6246
rect 5882 6238 5897 6246
rect 5831 270 5848 278
rect 5882 270 5897 278
rect 5831 258 5897 270
rect 5989 6246 6055 6258
rect 5989 6238 6006 6246
rect 6040 6238 6055 6246
rect 5989 270 6006 278
rect 6040 270 6055 278
rect 5989 258 6055 270
rect 6147 6246 6213 6258
rect 6147 6238 6164 6246
rect 6198 6238 6213 6246
rect 6147 270 6164 278
rect 6198 270 6213 278
rect 6147 258 6213 270
rect 6305 6246 6371 6258
rect 6305 6238 6322 6246
rect 6356 6238 6371 6246
rect 6305 270 6322 278
rect 6356 270 6371 278
rect 6305 258 6371 270
rect 1632 220 1652 226
rect 6286 220 6306 226
rect 1632 186 1644 220
rect 6294 186 6306 220
rect 1632 126 1652 186
rect 6286 126 6306 186
rect 1430 94 1500 100
rect 6440 94 6510 100
rect 1430 84 6510 94
rect 1430 46 1636 84
rect 6302 46 6510 84
rect 1430 30 6510 46
rect 7730 6470 12810 6480
rect 7730 6432 7936 6470
rect 12659 6432 12810 6470
rect 7730 6422 12810 6432
rect 7730 6420 7800 6422
rect 12740 6420 12810 6422
rect 7932 6330 7952 6390
rect 12586 6330 12606 6390
rect 7932 6296 7944 6330
rect 12594 6296 12606 6330
rect 7932 6290 7952 6296
rect 12586 6290 12606 6296
rect 7865 6246 7931 6258
rect 7865 6238 7882 6246
rect 7916 6238 7931 6246
rect 7865 270 7882 278
rect 7916 270 7931 278
rect 7865 258 7931 270
rect 8023 6246 8089 6258
rect 8023 6238 8040 6246
rect 8074 6238 8089 6246
rect 8023 270 8040 278
rect 8074 270 8089 278
rect 8023 258 8089 270
rect 8181 6246 8247 6258
rect 8181 6238 8198 6246
rect 8232 6238 8247 6246
rect 8181 270 8198 278
rect 8232 270 8247 278
rect 8181 258 8247 270
rect 8339 6246 8405 6258
rect 8339 6238 8356 6246
rect 8390 6238 8405 6246
rect 8339 270 8356 278
rect 8390 270 8405 278
rect 8339 258 8405 270
rect 8497 6246 8563 6258
rect 8497 6238 8514 6246
rect 8548 6238 8563 6246
rect 8497 270 8514 278
rect 8548 270 8563 278
rect 8497 258 8563 270
rect 8655 6246 8721 6258
rect 8655 6238 8672 6246
rect 8706 6238 8721 6246
rect 8655 270 8672 278
rect 8706 270 8721 278
rect 8655 258 8721 270
rect 8813 6246 8879 6258
rect 8813 6238 8830 6246
rect 8864 6238 8879 6246
rect 8813 270 8830 278
rect 8864 270 8879 278
rect 8813 258 8879 270
rect 8971 6246 9037 6258
rect 8971 6238 8988 6246
rect 9022 6238 9037 6246
rect 8971 270 8988 278
rect 9022 270 9037 278
rect 8971 258 9037 270
rect 9129 6246 9195 6258
rect 9129 6238 9146 6246
rect 9180 6238 9195 6246
rect 9129 270 9146 278
rect 9180 270 9195 278
rect 9129 258 9195 270
rect 9287 6246 9353 6258
rect 9287 6238 9304 6246
rect 9338 6238 9353 6246
rect 9287 270 9304 278
rect 9338 270 9353 278
rect 9287 258 9353 270
rect 9445 6246 9511 6258
rect 9445 6238 9462 6246
rect 9496 6238 9511 6246
rect 9445 270 9462 278
rect 9496 270 9511 278
rect 9445 258 9511 270
rect 9603 6246 9669 6258
rect 9603 6238 9620 6246
rect 9654 6238 9669 6246
rect 9603 270 9620 278
rect 9654 270 9669 278
rect 9603 258 9669 270
rect 9761 6246 9827 6258
rect 9761 6238 9778 6246
rect 9812 6238 9827 6246
rect 9761 270 9778 278
rect 9812 270 9827 278
rect 9761 258 9827 270
rect 9919 6246 9985 6258
rect 9919 6238 9936 6246
rect 9970 6238 9985 6246
rect 9919 270 9936 278
rect 9970 270 9985 278
rect 9919 258 9985 270
rect 10077 6246 10143 6258
rect 10077 6238 10094 6246
rect 10128 6238 10143 6246
rect 10077 270 10094 278
rect 10128 270 10143 278
rect 10077 258 10143 270
rect 10235 6246 10301 6258
rect 10235 6238 10252 6246
rect 10286 6238 10301 6246
rect 10235 270 10252 278
rect 10286 270 10301 278
rect 10235 258 10301 270
rect 10393 6246 10459 6258
rect 10393 6238 10410 6246
rect 10444 6238 10459 6246
rect 10393 270 10410 278
rect 10444 270 10459 278
rect 10393 258 10459 270
rect 10551 6246 10617 6258
rect 10551 6238 10568 6246
rect 10602 6238 10617 6246
rect 10551 270 10568 278
rect 10602 270 10617 278
rect 10551 258 10617 270
rect 10709 6246 10775 6258
rect 10709 6238 10726 6246
rect 10760 6238 10775 6246
rect 10709 270 10726 278
rect 10760 270 10775 278
rect 10709 258 10775 270
rect 10867 6246 10933 6258
rect 10867 6238 10884 6246
rect 10918 6238 10933 6246
rect 10867 270 10884 278
rect 10918 270 10933 278
rect 10867 258 10933 270
rect 11025 6246 11091 6258
rect 11025 6238 11042 6246
rect 11076 6238 11091 6246
rect 11025 270 11042 278
rect 11076 270 11091 278
rect 11025 258 11091 270
rect 11183 6246 11249 6258
rect 11183 6238 11200 6246
rect 11234 6238 11249 6246
rect 11183 270 11200 278
rect 11234 270 11249 278
rect 11183 258 11249 270
rect 11341 6246 11407 6258
rect 11341 6238 11358 6246
rect 11392 6238 11407 6246
rect 11341 270 11358 278
rect 11392 270 11407 278
rect 11341 258 11407 270
rect 11499 6246 11565 6258
rect 11499 6238 11516 6246
rect 11550 6238 11565 6246
rect 11499 270 11516 278
rect 11550 270 11565 278
rect 11499 258 11565 270
rect 11657 6246 11723 6258
rect 11657 6238 11674 6246
rect 11708 6238 11723 6246
rect 11657 270 11674 278
rect 11708 270 11723 278
rect 11657 258 11723 270
rect 11815 6246 11881 6258
rect 11815 6238 11832 6246
rect 11866 6238 11881 6246
rect 11815 270 11832 278
rect 11866 270 11881 278
rect 11815 258 11881 270
rect 11973 6246 12039 6258
rect 11973 6238 11990 6246
rect 12024 6238 12039 6246
rect 11973 270 11990 278
rect 12024 270 12039 278
rect 11973 258 12039 270
rect 12131 6246 12197 6258
rect 12131 6238 12148 6246
rect 12182 6238 12197 6246
rect 12131 270 12148 278
rect 12182 270 12197 278
rect 12131 258 12197 270
rect 12289 6246 12355 6258
rect 12289 6238 12306 6246
rect 12340 6238 12355 6246
rect 12289 270 12306 278
rect 12340 270 12355 278
rect 12289 258 12355 270
rect 12447 6246 12513 6258
rect 12447 6238 12464 6246
rect 12498 6238 12513 6246
rect 12447 270 12464 278
rect 12498 270 12513 278
rect 12447 258 12513 270
rect 12605 6246 12671 6258
rect 12605 6238 12622 6246
rect 12656 6238 12671 6246
rect 12605 270 12622 278
rect 12656 270 12671 278
rect 12605 258 12671 270
rect 7932 220 7952 226
rect 12586 220 12606 226
rect 7932 186 7944 220
rect 12594 186 12606 220
rect 7932 126 7952 186
rect 12586 126 12606 186
rect 7730 94 7800 100
rect 12740 94 12810 100
rect 7730 84 12810 94
rect 7730 46 7936 84
rect 12602 46 12810 84
rect 7730 30 12810 46
rect 14030 6470 19110 6480
rect 14030 6432 14236 6470
rect 18959 6432 19110 6470
rect 14030 6422 19110 6432
rect 14030 6420 14100 6422
rect 19040 6420 19110 6422
rect 14232 6330 14252 6390
rect 18886 6330 18906 6390
rect 14232 6296 14244 6330
rect 18894 6296 18906 6330
rect 14232 6290 14252 6296
rect 18886 6290 18906 6296
rect 14165 6246 14231 6258
rect 14165 6238 14182 6246
rect 14216 6238 14231 6246
rect 14165 270 14182 278
rect 14216 270 14231 278
rect 14165 258 14231 270
rect 14323 6246 14389 6258
rect 14323 6238 14340 6246
rect 14374 6238 14389 6246
rect 14323 270 14340 278
rect 14374 270 14389 278
rect 14323 258 14389 270
rect 14481 6246 14547 6258
rect 14481 6238 14498 6246
rect 14532 6238 14547 6246
rect 14481 270 14498 278
rect 14532 270 14547 278
rect 14481 258 14547 270
rect 14639 6246 14705 6258
rect 14639 6238 14656 6246
rect 14690 6238 14705 6246
rect 14639 270 14656 278
rect 14690 270 14705 278
rect 14639 258 14705 270
rect 14797 6246 14863 6258
rect 14797 6238 14814 6246
rect 14848 6238 14863 6246
rect 14797 270 14814 278
rect 14848 270 14863 278
rect 14797 258 14863 270
rect 14955 6246 15021 6258
rect 14955 6238 14972 6246
rect 15006 6238 15021 6246
rect 14955 270 14972 278
rect 15006 270 15021 278
rect 14955 258 15021 270
rect 15113 6246 15179 6258
rect 15113 6238 15130 6246
rect 15164 6238 15179 6246
rect 15113 270 15130 278
rect 15164 270 15179 278
rect 15113 258 15179 270
rect 15271 6246 15337 6258
rect 15271 6238 15288 6246
rect 15322 6238 15337 6246
rect 15271 270 15288 278
rect 15322 270 15337 278
rect 15271 258 15337 270
rect 15429 6246 15495 6258
rect 15429 6238 15446 6246
rect 15480 6238 15495 6246
rect 15429 270 15446 278
rect 15480 270 15495 278
rect 15429 258 15495 270
rect 15587 6246 15653 6258
rect 15587 6238 15604 6246
rect 15638 6238 15653 6246
rect 15587 270 15604 278
rect 15638 270 15653 278
rect 15587 258 15653 270
rect 15745 6246 15811 6258
rect 15745 6238 15762 6246
rect 15796 6238 15811 6246
rect 15745 270 15762 278
rect 15796 270 15811 278
rect 15745 258 15811 270
rect 15903 6246 15969 6258
rect 15903 6238 15920 6246
rect 15954 6238 15969 6246
rect 15903 270 15920 278
rect 15954 270 15969 278
rect 15903 258 15969 270
rect 16061 6246 16127 6258
rect 16061 6238 16078 6246
rect 16112 6238 16127 6246
rect 16061 270 16078 278
rect 16112 270 16127 278
rect 16061 258 16127 270
rect 16219 6246 16285 6258
rect 16219 6238 16236 6246
rect 16270 6238 16285 6246
rect 16219 270 16236 278
rect 16270 270 16285 278
rect 16219 258 16285 270
rect 16377 6246 16443 6258
rect 16377 6238 16394 6246
rect 16428 6238 16443 6246
rect 16377 270 16394 278
rect 16428 270 16443 278
rect 16377 258 16443 270
rect 16535 6246 16601 6258
rect 16535 6238 16552 6246
rect 16586 6238 16601 6246
rect 16535 270 16552 278
rect 16586 270 16601 278
rect 16535 258 16601 270
rect 16693 6246 16759 6258
rect 16693 6238 16710 6246
rect 16744 6238 16759 6246
rect 16693 270 16710 278
rect 16744 270 16759 278
rect 16693 258 16759 270
rect 16851 6246 16917 6258
rect 16851 6238 16868 6246
rect 16902 6238 16917 6246
rect 16851 270 16868 278
rect 16902 270 16917 278
rect 16851 258 16917 270
rect 17009 6246 17075 6258
rect 17009 6238 17026 6246
rect 17060 6238 17075 6246
rect 17009 270 17026 278
rect 17060 270 17075 278
rect 17009 258 17075 270
rect 17167 6246 17233 6258
rect 17167 6238 17184 6246
rect 17218 6238 17233 6246
rect 17167 270 17184 278
rect 17218 270 17233 278
rect 17167 258 17233 270
rect 17325 6246 17391 6258
rect 17325 6238 17342 6246
rect 17376 6238 17391 6246
rect 17325 270 17342 278
rect 17376 270 17391 278
rect 17325 258 17391 270
rect 17483 6246 17549 6258
rect 17483 6238 17500 6246
rect 17534 6238 17549 6246
rect 17483 270 17500 278
rect 17534 270 17549 278
rect 17483 258 17549 270
rect 17641 6246 17707 6258
rect 17641 6238 17658 6246
rect 17692 6238 17707 6246
rect 17641 270 17658 278
rect 17692 270 17707 278
rect 17641 258 17707 270
rect 17799 6246 17865 6258
rect 17799 6238 17816 6246
rect 17850 6238 17865 6246
rect 17799 270 17816 278
rect 17850 270 17865 278
rect 17799 258 17865 270
rect 17957 6246 18023 6258
rect 17957 6238 17974 6246
rect 18008 6238 18023 6246
rect 17957 270 17974 278
rect 18008 270 18023 278
rect 17957 258 18023 270
rect 18115 6246 18181 6258
rect 18115 6238 18132 6246
rect 18166 6238 18181 6246
rect 18115 270 18132 278
rect 18166 270 18181 278
rect 18115 258 18181 270
rect 18273 6246 18339 6258
rect 18273 6238 18290 6246
rect 18324 6238 18339 6246
rect 18273 270 18290 278
rect 18324 270 18339 278
rect 18273 258 18339 270
rect 18431 6246 18497 6258
rect 18431 6238 18448 6246
rect 18482 6238 18497 6246
rect 18431 270 18448 278
rect 18482 270 18497 278
rect 18431 258 18497 270
rect 18589 6246 18655 6258
rect 18589 6238 18606 6246
rect 18640 6238 18655 6246
rect 18589 270 18606 278
rect 18640 270 18655 278
rect 18589 258 18655 270
rect 18747 6246 18813 6258
rect 18747 6238 18764 6246
rect 18798 6238 18813 6246
rect 18747 270 18764 278
rect 18798 270 18813 278
rect 18747 258 18813 270
rect 18905 6246 18971 6258
rect 18905 6238 18922 6246
rect 18956 6238 18971 6246
rect 18905 270 18922 278
rect 18956 270 18971 278
rect 18905 258 18971 270
rect 14232 220 14252 226
rect 18886 220 18906 226
rect 14232 186 14244 220
rect 18894 186 18906 220
rect 14232 126 14252 186
rect 18886 126 18906 186
rect 14030 94 14100 100
rect 19040 94 19110 100
rect 14030 84 19110 94
rect 14030 46 14236 84
rect 18902 46 19110 84
rect 14030 30 19110 46
rect 20330 6470 25410 6480
rect 20330 6432 20536 6470
rect 25259 6432 25410 6470
rect 20330 6422 25410 6432
rect 20330 6420 20400 6422
rect 25340 6420 25410 6422
rect 20532 6330 20552 6390
rect 25186 6330 25206 6390
rect 20532 6296 20544 6330
rect 25194 6296 25206 6330
rect 20532 6290 20552 6296
rect 25186 6290 25206 6296
rect 20465 6246 20531 6258
rect 20465 6238 20482 6246
rect 20516 6238 20531 6246
rect 20465 270 20482 278
rect 20516 270 20531 278
rect 20465 258 20531 270
rect 20623 6246 20689 6258
rect 20623 6238 20640 6246
rect 20674 6238 20689 6246
rect 20623 270 20640 278
rect 20674 270 20689 278
rect 20623 258 20689 270
rect 20781 6246 20847 6258
rect 20781 6238 20798 6246
rect 20832 6238 20847 6246
rect 20781 270 20798 278
rect 20832 270 20847 278
rect 20781 258 20847 270
rect 20939 6246 21005 6258
rect 20939 6238 20956 6246
rect 20990 6238 21005 6246
rect 20939 270 20956 278
rect 20990 270 21005 278
rect 20939 258 21005 270
rect 21097 6246 21163 6258
rect 21097 6238 21114 6246
rect 21148 6238 21163 6246
rect 21097 270 21114 278
rect 21148 270 21163 278
rect 21097 258 21163 270
rect 21255 6246 21321 6258
rect 21255 6238 21272 6246
rect 21306 6238 21321 6246
rect 21255 270 21272 278
rect 21306 270 21321 278
rect 21255 258 21321 270
rect 21413 6246 21479 6258
rect 21413 6238 21430 6246
rect 21464 6238 21479 6246
rect 21413 270 21430 278
rect 21464 270 21479 278
rect 21413 258 21479 270
rect 21571 6246 21637 6258
rect 21571 6238 21588 6246
rect 21622 6238 21637 6246
rect 21571 270 21588 278
rect 21622 270 21637 278
rect 21571 258 21637 270
rect 21729 6246 21795 6258
rect 21729 6238 21746 6246
rect 21780 6238 21795 6246
rect 21729 270 21746 278
rect 21780 270 21795 278
rect 21729 258 21795 270
rect 21887 6246 21953 6258
rect 21887 6238 21904 6246
rect 21938 6238 21953 6246
rect 21887 270 21904 278
rect 21938 270 21953 278
rect 21887 258 21953 270
rect 22045 6246 22111 6258
rect 22045 6238 22062 6246
rect 22096 6238 22111 6246
rect 22045 270 22062 278
rect 22096 270 22111 278
rect 22045 258 22111 270
rect 22203 6246 22269 6258
rect 22203 6238 22220 6246
rect 22254 6238 22269 6246
rect 22203 270 22220 278
rect 22254 270 22269 278
rect 22203 258 22269 270
rect 22361 6246 22427 6258
rect 22361 6238 22378 6246
rect 22412 6238 22427 6246
rect 22361 270 22378 278
rect 22412 270 22427 278
rect 22361 258 22427 270
rect 22519 6246 22585 6258
rect 22519 6238 22536 6246
rect 22570 6238 22585 6246
rect 22519 270 22536 278
rect 22570 270 22585 278
rect 22519 258 22585 270
rect 22677 6246 22743 6258
rect 22677 6238 22694 6246
rect 22728 6238 22743 6246
rect 22677 270 22694 278
rect 22728 270 22743 278
rect 22677 258 22743 270
rect 22835 6246 22901 6258
rect 22835 6238 22852 6246
rect 22886 6238 22901 6246
rect 22835 270 22852 278
rect 22886 270 22901 278
rect 22835 258 22901 270
rect 22993 6246 23059 6258
rect 22993 6238 23010 6246
rect 23044 6238 23059 6246
rect 22993 270 23010 278
rect 23044 270 23059 278
rect 22993 258 23059 270
rect 23151 6246 23217 6258
rect 23151 6238 23168 6246
rect 23202 6238 23217 6246
rect 23151 270 23168 278
rect 23202 270 23217 278
rect 23151 258 23217 270
rect 23309 6246 23375 6258
rect 23309 6238 23326 6246
rect 23360 6238 23375 6246
rect 23309 270 23326 278
rect 23360 270 23375 278
rect 23309 258 23375 270
rect 23467 6246 23533 6258
rect 23467 6238 23484 6246
rect 23518 6238 23533 6246
rect 23467 270 23484 278
rect 23518 270 23533 278
rect 23467 258 23533 270
rect 23625 6246 23691 6258
rect 23625 6238 23642 6246
rect 23676 6238 23691 6246
rect 23625 270 23642 278
rect 23676 270 23691 278
rect 23625 258 23691 270
rect 23783 6246 23849 6258
rect 23783 6238 23800 6246
rect 23834 6238 23849 6246
rect 23783 270 23800 278
rect 23834 270 23849 278
rect 23783 258 23849 270
rect 23941 6246 24007 6258
rect 23941 6238 23958 6246
rect 23992 6238 24007 6246
rect 23941 270 23958 278
rect 23992 270 24007 278
rect 23941 258 24007 270
rect 24099 6246 24165 6258
rect 24099 6238 24116 6246
rect 24150 6238 24165 6246
rect 24099 270 24116 278
rect 24150 270 24165 278
rect 24099 258 24165 270
rect 24257 6246 24323 6258
rect 24257 6238 24274 6246
rect 24308 6238 24323 6246
rect 24257 270 24274 278
rect 24308 270 24323 278
rect 24257 258 24323 270
rect 24415 6246 24481 6258
rect 24415 6238 24432 6246
rect 24466 6238 24481 6246
rect 24415 270 24432 278
rect 24466 270 24481 278
rect 24415 258 24481 270
rect 24573 6246 24639 6258
rect 24573 6238 24590 6246
rect 24624 6238 24639 6246
rect 24573 270 24590 278
rect 24624 270 24639 278
rect 24573 258 24639 270
rect 24731 6246 24797 6258
rect 24731 6238 24748 6246
rect 24782 6238 24797 6246
rect 24731 270 24748 278
rect 24782 270 24797 278
rect 24731 258 24797 270
rect 24889 6246 24955 6258
rect 24889 6238 24906 6246
rect 24940 6238 24955 6246
rect 24889 270 24906 278
rect 24940 270 24955 278
rect 24889 258 24955 270
rect 25047 6246 25113 6258
rect 25047 6238 25064 6246
rect 25098 6238 25113 6246
rect 25047 270 25064 278
rect 25098 270 25113 278
rect 25047 258 25113 270
rect 25205 6246 25271 6258
rect 25205 6238 25222 6246
rect 25256 6238 25271 6246
rect 25205 270 25222 278
rect 25256 270 25271 278
rect 25205 258 25271 270
rect 20532 220 20552 226
rect 25186 220 25206 226
rect 20532 186 20544 220
rect 25194 186 25206 220
rect 20532 126 20552 186
rect 25186 126 25206 186
rect 20330 94 20400 100
rect 25340 94 25410 100
rect 20330 84 25410 94
rect 20330 46 20536 84
rect 25202 46 25410 84
rect 20330 30 25410 46
rect 1430 -530 6510 -520
rect 1430 -568 1636 -530
rect 6359 -568 6510 -530
rect 1430 -578 6510 -568
rect 1430 -580 1500 -578
rect 6440 -580 6510 -578
rect 1632 -670 1652 -610
rect 6286 -670 6306 -610
rect 1632 -704 1644 -670
rect 6294 -704 6306 -670
rect 1632 -710 1652 -704
rect 6286 -710 6306 -704
rect 1565 -754 1631 -742
rect 1565 -762 1582 -754
rect 1616 -762 1631 -754
rect 1565 -6730 1582 -6722
rect 1616 -6730 1631 -6722
rect 1565 -6742 1631 -6730
rect 1723 -754 1789 -742
rect 1723 -762 1740 -754
rect 1774 -762 1789 -754
rect 1723 -6730 1740 -6722
rect 1774 -6730 1789 -6722
rect 1723 -6742 1789 -6730
rect 1881 -754 1947 -742
rect 1881 -762 1898 -754
rect 1932 -762 1947 -754
rect 1881 -6730 1898 -6722
rect 1932 -6730 1947 -6722
rect 1881 -6742 1947 -6730
rect 2039 -754 2105 -742
rect 2039 -762 2056 -754
rect 2090 -762 2105 -754
rect 2039 -6730 2056 -6722
rect 2090 -6730 2105 -6722
rect 2039 -6742 2105 -6730
rect 2197 -754 2263 -742
rect 2197 -762 2214 -754
rect 2248 -762 2263 -754
rect 2197 -6730 2214 -6722
rect 2248 -6730 2263 -6722
rect 2197 -6742 2263 -6730
rect 2355 -754 2421 -742
rect 2355 -762 2372 -754
rect 2406 -762 2421 -754
rect 2355 -6730 2372 -6722
rect 2406 -6730 2421 -6722
rect 2355 -6742 2421 -6730
rect 2513 -754 2579 -742
rect 2513 -762 2530 -754
rect 2564 -762 2579 -754
rect 2513 -6730 2530 -6722
rect 2564 -6730 2579 -6722
rect 2513 -6742 2579 -6730
rect 2671 -754 2737 -742
rect 2671 -762 2688 -754
rect 2722 -762 2737 -754
rect 2671 -6730 2688 -6722
rect 2722 -6730 2737 -6722
rect 2671 -6742 2737 -6730
rect 2829 -754 2895 -742
rect 2829 -762 2846 -754
rect 2880 -762 2895 -754
rect 2829 -6730 2846 -6722
rect 2880 -6730 2895 -6722
rect 2829 -6742 2895 -6730
rect 2987 -754 3053 -742
rect 2987 -762 3004 -754
rect 3038 -762 3053 -754
rect 2987 -6730 3004 -6722
rect 3038 -6730 3053 -6722
rect 2987 -6742 3053 -6730
rect 3145 -754 3211 -742
rect 3145 -762 3162 -754
rect 3196 -762 3211 -754
rect 3145 -6730 3162 -6722
rect 3196 -6730 3211 -6722
rect 3145 -6742 3211 -6730
rect 3303 -754 3369 -742
rect 3303 -762 3320 -754
rect 3354 -762 3369 -754
rect 3303 -6730 3320 -6722
rect 3354 -6730 3369 -6722
rect 3303 -6742 3369 -6730
rect 3461 -754 3527 -742
rect 3461 -762 3478 -754
rect 3512 -762 3527 -754
rect 3461 -6730 3478 -6722
rect 3512 -6730 3527 -6722
rect 3461 -6742 3527 -6730
rect 3619 -754 3685 -742
rect 3619 -762 3636 -754
rect 3670 -762 3685 -754
rect 3619 -6730 3636 -6722
rect 3670 -6730 3685 -6722
rect 3619 -6742 3685 -6730
rect 3777 -754 3843 -742
rect 3777 -762 3794 -754
rect 3828 -762 3843 -754
rect 3777 -6730 3794 -6722
rect 3828 -6730 3843 -6722
rect 3777 -6742 3843 -6730
rect 3935 -754 4001 -742
rect 3935 -762 3952 -754
rect 3986 -762 4001 -754
rect 3935 -6730 3952 -6722
rect 3986 -6730 4001 -6722
rect 3935 -6742 4001 -6730
rect 4093 -754 4159 -742
rect 4093 -762 4110 -754
rect 4144 -762 4159 -754
rect 4093 -6730 4110 -6722
rect 4144 -6730 4159 -6722
rect 4093 -6742 4159 -6730
rect 4251 -754 4317 -742
rect 4251 -762 4268 -754
rect 4302 -762 4317 -754
rect 4251 -6730 4268 -6722
rect 4302 -6730 4317 -6722
rect 4251 -6742 4317 -6730
rect 4409 -754 4475 -742
rect 4409 -762 4426 -754
rect 4460 -762 4475 -754
rect 4409 -6730 4426 -6722
rect 4460 -6730 4475 -6722
rect 4409 -6742 4475 -6730
rect 4567 -754 4633 -742
rect 4567 -762 4584 -754
rect 4618 -762 4633 -754
rect 4567 -6730 4584 -6722
rect 4618 -6730 4633 -6722
rect 4567 -6742 4633 -6730
rect 4725 -754 4791 -742
rect 4725 -762 4742 -754
rect 4776 -762 4791 -754
rect 4725 -6730 4742 -6722
rect 4776 -6730 4791 -6722
rect 4725 -6742 4791 -6730
rect 4883 -754 4949 -742
rect 4883 -762 4900 -754
rect 4934 -762 4949 -754
rect 4883 -6730 4900 -6722
rect 4934 -6730 4949 -6722
rect 4883 -6742 4949 -6730
rect 5041 -754 5107 -742
rect 5041 -762 5058 -754
rect 5092 -762 5107 -754
rect 5041 -6730 5058 -6722
rect 5092 -6730 5107 -6722
rect 5041 -6742 5107 -6730
rect 5199 -754 5265 -742
rect 5199 -762 5216 -754
rect 5250 -762 5265 -754
rect 5199 -6730 5216 -6722
rect 5250 -6730 5265 -6722
rect 5199 -6742 5265 -6730
rect 5357 -754 5423 -742
rect 5357 -762 5374 -754
rect 5408 -762 5423 -754
rect 5357 -6730 5374 -6722
rect 5408 -6730 5423 -6722
rect 5357 -6742 5423 -6730
rect 5515 -754 5581 -742
rect 5515 -762 5532 -754
rect 5566 -762 5581 -754
rect 5515 -6730 5532 -6722
rect 5566 -6730 5581 -6722
rect 5515 -6742 5581 -6730
rect 5673 -754 5739 -742
rect 5673 -762 5690 -754
rect 5724 -762 5739 -754
rect 5673 -6730 5690 -6722
rect 5724 -6730 5739 -6722
rect 5673 -6742 5739 -6730
rect 5831 -754 5897 -742
rect 5831 -762 5848 -754
rect 5882 -762 5897 -754
rect 5831 -6730 5848 -6722
rect 5882 -6730 5897 -6722
rect 5831 -6742 5897 -6730
rect 5989 -754 6055 -742
rect 5989 -762 6006 -754
rect 6040 -762 6055 -754
rect 5989 -6730 6006 -6722
rect 6040 -6730 6055 -6722
rect 5989 -6742 6055 -6730
rect 6147 -754 6213 -742
rect 6147 -762 6164 -754
rect 6198 -762 6213 -754
rect 6147 -6730 6164 -6722
rect 6198 -6730 6213 -6722
rect 6147 -6742 6213 -6730
rect 6305 -754 6371 -742
rect 6305 -762 6322 -754
rect 6356 -762 6371 -754
rect 6305 -6730 6322 -6722
rect 6356 -6730 6371 -6722
rect 6305 -6742 6371 -6730
rect 1632 -6780 1652 -6774
rect 6286 -6780 6306 -6774
rect 1632 -6814 1644 -6780
rect 6294 -6814 6306 -6780
rect 1632 -6874 1652 -6814
rect 6286 -6874 6306 -6814
rect 1430 -6906 1500 -6900
rect 6440 -6906 6510 -6900
rect 1430 -6916 6510 -6906
rect 1430 -6954 1636 -6916
rect 6302 -6954 6510 -6916
rect 1430 -6970 6510 -6954
rect 7730 -530 12810 -520
rect 7730 -568 7936 -530
rect 12659 -568 12810 -530
rect 7730 -578 12810 -568
rect 7730 -580 7800 -578
rect 12740 -580 12810 -578
rect 7932 -670 7952 -610
rect 12586 -670 12606 -610
rect 7932 -704 7944 -670
rect 12594 -704 12606 -670
rect 7932 -710 7952 -704
rect 12586 -710 12606 -704
rect 7865 -754 7931 -742
rect 7865 -762 7882 -754
rect 7916 -762 7931 -754
rect 7865 -6730 7882 -6722
rect 7916 -6730 7931 -6722
rect 7865 -6742 7931 -6730
rect 8023 -754 8089 -742
rect 8023 -762 8040 -754
rect 8074 -762 8089 -754
rect 8023 -6730 8040 -6722
rect 8074 -6730 8089 -6722
rect 8023 -6742 8089 -6730
rect 8181 -754 8247 -742
rect 8181 -762 8198 -754
rect 8232 -762 8247 -754
rect 8181 -6730 8198 -6722
rect 8232 -6730 8247 -6722
rect 8181 -6742 8247 -6730
rect 8339 -754 8405 -742
rect 8339 -762 8356 -754
rect 8390 -762 8405 -754
rect 8339 -6730 8356 -6722
rect 8390 -6730 8405 -6722
rect 8339 -6742 8405 -6730
rect 8497 -754 8563 -742
rect 8497 -762 8514 -754
rect 8548 -762 8563 -754
rect 8497 -6730 8514 -6722
rect 8548 -6730 8563 -6722
rect 8497 -6742 8563 -6730
rect 8655 -754 8721 -742
rect 8655 -762 8672 -754
rect 8706 -762 8721 -754
rect 8655 -6730 8672 -6722
rect 8706 -6730 8721 -6722
rect 8655 -6742 8721 -6730
rect 8813 -754 8879 -742
rect 8813 -762 8830 -754
rect 8864 -762 8879 -754
rect 8813 -6730 8830 -6722
rect 8864 -6730 8879 -6722
rect 8813 -6742 8879 -6730
rect 8971 -754 9037 -742
rect 8971 -762 8988 -754
rect 9022 -762 9037 -754
rect 8971 -6730 8988 -6722
rect 9022 -6730 9037 -6722
rect 8971 -6742 9037 -6730
rect 9129 -754 9195 -742
rect 9129 -762 9146 -754
rect 9180 -762 9195 -754
rect 9129 -6730 9146 -6722
rect 9180 -6730 9195 -6722
rect 9129 -6742 9195 -6730
rect 9287 -754 9353 -742
rect 9287 -762 9304 -754
rect 9338 -762 9353 -754
rect 9287 -6730 9304 -6722
rect 9338 -6730 9353 -6722
rect 9287 -6742 9353 -6730
rect 9445 -754 9511 -742
rect 9445 -762 9462 -754
rect 9496 -762 9511 -754
rect 9445 -6730 9462 -6722
rect 9496 -6730 9511 -6722
rect 9445 -6742 9511 -6730
rect 9603 -754 9669 -742
rect 9603 -762 9620 -754
rect 9654 -762 9669 -754
rect 9603 -6730 9620 -6722
rect 9654 -6730 9669 -6722
rect 9603 -6742 9669 -6730
rect 9761 -754 9827 -742
rect 9761 -762 9778 -754
rect 9812 -762 9827 -754
rect 9761 -6730 9778 -6722
rect 9812 -6730 9827 -6722
rect 9761 -6742 9827 -6730
rect 9919 -754 9985 -742
rect 9919 -762 9936 -754
rect 9970 -762 9985 -754
rect 9919 -6730 9936 -6722
rect 9970 -6730 9985 -6722
rect 9919 -6742 9985 -6730
rect 10077 -754 10143 -742
rect 10077 -762 10094 -754
rect 10128 -762 10143 -754
rect 10077 -6730 10094 -6722
rect 10128 -6730 10143 -6722
rect 10077 -6742 10143 -6730
rect 10235 -754 10301 -742
rect 10235 -762 10252 -754
rect 10286 -762 10301 -754
rect 10235 -6730 10252 -6722
rect 10286 -6730 10301 -6722
rect 10235 -6742 10301 -6730
rect 10393 -754 10459 -742
rect 10393 -762 10410 -754
rect 10444 -762 10459 -754
rect 10393 -6730 10410 -6722
rect 10444 -6730 10459 -6722
rect 10393 -6742 10459 -6730
rect 10551 -754 10617 -742
rect 10551 -762 10568 -754
rect 10602 -762 10617 -754
rect 10551 -6730 10568 -6722
rect 10602 -6730 10617 -6722
rect 10551 -6742 10617 -6730
rect 10709 -754 10775 -742
rect 10709 -762 10726 -754
rect 10760 -762 10775 -754
rect 10709 -6730 10726 -6722
rect 10760 -6730 10775 -6722
rect 10709 -6742 10775 -6730
rect 10867 -754 10933 -742
rect 10867 -762 10884 -754
rect 10918 -762 10933 -754
rect 10867 -6730 10884 -6722
rect 10918 -6730 10933 -6722
rect 10867 -6742 10933 -6730
rect 11025 -754 11091 -742
rect 11025 -762 11042 -754
rect 11076 -762 11091 -754
rect 11025 -6730 11042 -6722
rect 11076 -6730 11091 -6722
rect 11025 -6742 11091 -6730
rect 11183 -754 11249 -742
rect 11183 -762 11200 -754
rect 11234 -762 11249 -754
rect 11183 -6730 11200 -6722
rect 11234 -6730 11249 -6722
rect 11183 -6742 11249 -6730
rect 11341 -754 11407 -742
rect 11341 -762 11358 -754
rect 11392 -762 11407 -754
rect 11341 -6730 11358 -6722
rect 11392 -6730 11407 -6722
rect 11341 -6742 11407 -6730
rect 11499 -754 11565 -742
rect 11499 -762 11516 -754
rect 11550 -762 11565 -754
rect 11499 -6730 11516 -6722
rect 11550 -6730 11565 -6722
rect 11499 -6742 11565 -6730
rect 11657 -754 11723 -742
rect 11657 -762 11674 -754
rect 11708 -762 11723 -754
rect 11657 -6730 11674 -6722
rect 11708 -6730 11723 -6722
rect 11657 -6742 11723 -6730
rect 11815 -754 11881 -742
rect 11815 -762 11832 -754
rect 11866 -762 11881 -754
rect 11815 -6730 11832 -6722
rect 11866 -6730 11881 -6722
rect 11815 -6742 11881 -6730
rect 11973 -754 12039 -742
rect 11973 -762 11990 -754
rect 12024 -762 12039 -754
rect 11973 -6730 11990 -6722
rect 12024 -6730 12039 -6722
rect 11973 -6742 12039 -6730
rect 12131 -754 12197 -742
rect 12131 -762 12148 -754
rect 12182 -762 12197 -754
rect 12131 -6730 12148 -6722
rect 12182 -6730 12197 -6722
rect 12131 -6742 12197 -6730
rect 12289 -754 12355 -742
rect 12289 -762 12306 -754
rect 12340 -762 12355 -754
rect 12289 -6730 12306 -6722
rect 12340 -6730 12355 -6722
rect 12289 -6742 12355 -6730
rect 12447 -754 12513 -742
rect 12447 -762 12464 -754
rect 12498 -762 12513 -754
rect 12447 -6730 12464 -6722
rect 12498 -6730 12513 -6722
rect 12447 -6742 12513 -6730
rect 12605 -754 12671 -742
rect 12605 -762 12622 -754
rect 12656 -762 12671 -754
rect 12605 -6730 12622 -6722
rect 12656 -6730 12671 -6722
rect 12605 -6742 12671 -6730
rect 7932 -6780 7952 -6774
rect 12586 -6780 12606 -6774
rect 7932 -6814 7944 -6780
rect 12594 -6814 12606 -6780
rect 7932 -6874 7952 -6814
rect 12586 -6874 12606 -6814
rect 7730 -6906 7800 -6900
rect 12740 -6906 12810 -6900
rect 7730 -6916 12810 -6906
rect 7730 -6954 7936 -6916
rect 12602 -6954 12810 -6916
rect 7730 -6970 12810 -6954
rect 14030 -530 19110 -520
rect 14030 -568 14236 -530
rect 18959 -568 19110 -530
rect 14030 -578 19110 -568
rect 14030 -580 14100 -578
rect 19040 -580 19110 -578
rect 14232 -670 14252 -610
rect 18886 -670 18906 -610
rect 14232 -704 14244 -670
rect 18894 -704 18906 -670
rect 14232 -710 14252 -704
rect 18886 -710 18906 -704
rect 14165 -754 14231 -742
rect 14165 -762 14182 -754
rect 14216 -762 14231 -754
rect 14165 -6730 14182 -6722
rect 14216 -6730 14231 -6722
rect 14165 -6742 14231 -6730
rect 14323 -754 14389 -742
rect 14323 -762 14340 -754
rect 14374 -762 14389 -754
rect 14323 -6730 14340 -6722
rect 14374 -6730 14389 -6722
rect 14323 -6742 14389 -6730
rect 14481 -754 14547 -742
rect 14481 -762 14498 -754
rect 14532 -762 14547 -754
rect 14481 -6730 14498 -6722
rect 14532 -6730 14547 -6722
rect 14481 -6742 14547 -6730
rect 14639 -754 14705 -742
rect 14639 -762 14656 -754
rect 14690 -762 14705 -754
rect 14639 -6730 14656 -6722
rect 14690 -6730 14705 -6722
rect 14639 -6742 14705 -6730
rect 14797 -754 14863 -742
rect 14797 -762 14814 -754
rect 14848 -762 14863 -754
rect 14797 -6730 14814 -6722
rect 14848 -6730 14863 -6722
rect 14797 -6742 14863 -6730
rect 14955 -754 15021 -742
rect 14955 -762 14972 -754
rect 15006 -762 15021 -754
rect 14955 -6730 14972 -6722
rect 15006 -6730 15021 -6722
rect 14955 -6742 15021 -6730
rect 15113 -754 15179 -742
rect 15113 -762 15130 -754
rect 15164 -762 15179 -754
rect 15113 -6730 15130 -6722
rect 15164 -6730 15179 -6722
rect 15113 -6742 15179 -6730
rect 15271 -754 15337 -742
rect 15271 -762 15288 -754
rect 15322 -762 15337 -754
rect 15271 -6730 15288 -6722
rect 15322 -6730 15337 -6722
rect 15271 -6742 15337 -6730
rect 15429 -754 15495 -742
rect 15429 -762 15446 -754
rect 15480 -762 15495 -754
rect 15429 -6730 15446 -6722
rect 15480 -6730 15495 -6722
rect 15429 -6742 15495 -6730
rect 15587 -754 15653 -742
rect 15587 -762 15604 -754
rect 15638 -762 15653 -754
rect 15587 -6730 15604 -6722
rect 15638 -6730 15653 -6722
rect 15587 -6742 15653 -6730
rect 15745 -754 15811 -742
rect 15745 -762 15762 -754
rect 15796 -762 15811 -754
rect 15745 -6730 15762 -6722
rect 15796 -6730 15811 -6722
rect 15745 -6742 15811 -6730
rect 15903 -754 15969 -742
rect 15903 -762 15920 -754
rect 15954 -762 15969 -754
rect 15903 -6730 15920 -6722
rect 15954 -6730 15969 -6722
rect 15903 -6742 15969 -6730
rect 16061 -754 16127 -742
rect 16061 -762 16078 -754
rect 16112 -762 16127 -754
rect 16061 -6730 16078 -6722
rect 16112 -6730 16127 -6722
rect 16061 -6742 16127 -6730
rect 16219 -754 16285 -742
rect 16219 -762 16236 -754
rect 16270 -762 16285 -754
rect 16219 -6730 16236 -6722
rect 16270 -6730 16285 -6722
rect 16219 -6742 16285 -6730
rect 16377 -754 16443 -742
rect 16377 -762 16394 -754
rect 16428 -762 16443 -754
rect 16377 -6730 16394 -6722
rect 16428 -6730 16443 -6722
rect 16377 -6742 16443 -6730
rect 16535 -754 16601 -742
rect 16535 -762 16552 -754
rect 16586 -762 16601 -754
rect 16535 -6730 16552 -6722
rect 16586 -6730 16601 -6722
rect 16535 -6742 16601 -6730
rect 16693 -754 16759 -742
rect 16693 -762 16710 -754
rect 16744 -762 16759 -754
rect 16693 -6730 16710 -6722
rect 16744 -6730 16759 -6722
rect 16693 -6742 16759 -6730
rect 16851 -754 16917 -742
rect 16851 -762 16868 -754
rect 16902 -762 16917 -754
rect 16851 -6730 16868 -6722
rect 16902 -6730 16917 -6722
rect 16851 -6742 16917 -6730
rect 17009 -754 17075 -742
rect 17009 -762 17026 -754
rect 17060 -762 17075 -754
rect 17009 -6730 17026 -6722
rect 17060 -6730 17075 -6722
rect 17009 -6742 17075 -6730
rect 17167 -754 17233 -742
rect 17167 -762 17184 -754
rect 17218 -762 17233 -754
rect 17167 -6730 17184 -6722
rect 17218 -6730 17233 -6722
rect 17167 -6742 17233 -6730
rect 17325 -754 17391 -742
rect 17325 -762 17342 -754
rect 17376 -762 17391 -754
rect 17325 -6730 17342 -6722
rect 17376 -6730 17391 -6722
rect 17325 -6742 17391 -6730
rect 17483 -754 17549 -742
rect 17483 -762 17500 -754
rect 17534 -762 17549 -754
rect 17483 -6730 17500 -6722
rect 17534 -6730 17549 -6722
rect 17483 -6742 17549 -6730
rect 17641 -754 17707 -742
rect 17641 -762 17658 -754
rect 17692 -762 17707 -754
rect 17641 -6730 17658 -6722
rect 17692 -6730 17707 -6722
rect 17641 -6742 17707 -6730
rect 17799 -754 17865 -742
rect 17799 -762 17816 -754
rect 17850 -762 17865 -754
rect 17799 -6730 17816 -6722
rect 17850 -6730 17865 -6722
rect 17799 -6742 17865 -6730
rect 17957 -754 18023 -742
rect 17957 -762 17974 -754
rect 18008 -762 18023 -754
rect 17957 -6730 17974 -6722
rect 18008 -6730 18023 -6722
rect 17957 -6742 18023 -6730
rect 18115 -754 18181 -742
rect 18115 -762 18132 -754
rect 18166 -762 18181 -754
rect 18115 -6730 18132 -6722
rect 18166 -6730 18181 -6722
rect 18115 -6742 18181 -6730
rect 18273 -754 18339 -742
rect 18273 -762 18290 -754
rect 18324 -762 18339 -754
rect 18273 -6730 18290 -6722
rect 18324 -6730 18339 -6722
rect 18273 -6742 18339 -6730
rect 18431 -754 18497 -742
rect 18431 -762 18448 -754
rect 18482 -762 18497 -754
rect 18431 -6730 18448 -6722
rect 18482 -6730 18497 -6722
rect 18431 -6742 18497 -6730
rect 18589 -754 18655 -742
rect 18589 -762 18606 -754
rect 18640 -762 18655 -754
rect 18589 -6730 18606 -6722
rect 18640 -6730 18655 -6722
rect 18589 -6742 18655 -6730
rect 18747 -754 18813 -742
rect 18747 -762 18764 -754
rect 18798 -762 18813 -754
rect 18747 -6730 18764 -6722
rect 18798 -6730 18813 -6722
rect 18747 -6742 18813 -6730
rect 18905 -754 18971 -742
rect 18905 -762 18922 -754
rect 18956 -762 18971 -754
rect 18905 -6730 18922 -6722
rect 18956 -6730 18971 -6722
rect 18905 -6742 18971 -6730
rect 14232 -6780 14252 -6774
rect 18886 -6780 18906 -6774
rect 14232 -6814 14244 -6780
rect 18894 -6814 18906 -6780
rect 14232 -6874 14252 -6814
rect 18886 -6874 18906 -6814
rect 14030 -6906 14100 -6900
rect 19040 -6906 19110 -6900
rect 14030 -6916 19110 -6906
rect 14030 -6954 14236 -6916
rect 18902 -6954 19110 -6916
rect 14030 -6970 19110 -6954
rect 20330 -530 25410 -520
rect 20330 -568 20536 -530
rect 25259 -568 25410 -530
rect 20330 -578 25410 -568
rect 20330 -580 20400 -578
rect 25340 -580 25410 -578
rect 20532 -670 20552 -610
rect 25186 -670 25206 -610
rect 20532 -704 20544 -670
rect 25194 -704 25206 -670
rect 20532 -710 20552 -704
rect 25186 -710 25206 -704
rect 20465 -754 20531 -742
rect 20465 -762 20482 -754
rect 20516 -762 20531 -754
rect 20465 -6730 20482 -6722
rect 20516 -6730 20531 -6722
rect 20465 -6742 20531 -6730
rect 20623 -754 20689 -742
rect 20623 -762 20640 -754
rect 20674 -762 20689 -754
rect 20623 -6730 20640 -6722
rect 20674 -6730 20689 -6722
rect 20623 -6742 20689 -6730
rect 20781 -754 20847 -742
rect 20781 -762 20798 -754
rect 20832 -762 20847 -754
rect 20781 -6730 20798 -6722
rect 20832 -6730 20847 -6722
rect 20781 -6742 20847 -6730
rect 20939 -754 21005 -742
rect 20939 -762 20956 -754
rect 20990 -762 21005 -754
rect 20939 -6730 20956 -6722
rect 20990 -6730 21005 -6722
rect 20939 -6742 21005 -6730
rect 21097 -754 21163 -742
rect 21097 -762 21114 -754
rect 21148 -762 21163 -754
rect 21097 -6730 21114 -6722
rect 21148 -6730 21163 -6722
rect 21097 -6742 21163 -6730
rect 21255 -754 21321 -742
rect 21255 -762 21272 -754
rect 21306 -762 21321 -754
rect 21255 -6730 21272 -6722
rect 21306 -6730 21321 -6722
rect 21255 -6742 21321 -6730
rect 21413 -754 21479 -742
rect 21413 -762 21430 -754
rect 21464 -762 21479 -754
rect 21413 -6730 21430 -6722
rect 21464 -6730 21479 -6722
rect 21413 -6742 21479 -6730
rect 21571 -754 21637 -742
rect 21571 -762 21588 -754
rect 21622 -762 21637 -754
rect 21571 -6730 21588 -6722
rect 21622 -6730 21637 -6722
rect 21571 -6742 21637 -6730
rect 21729 -754 21795 -742
rect 21729 -762 21746 -754
rect 21780 -762 21795 -754
rect 21729 -6730 21746 -6722
rect 21780 -6730 21795 -6722
rect 21729 -6742 21795 -6730
rect 21887 -754 21953 -742
rect 21887 -762 21904 -754
rect 21938 -762 21953 -754
rect 21887 -6730 21904 -6722
rect 21938 -6730 21953 -6722
rect 21887 -6742 21953 -6730
rect 22045 -754 22111 -742
rect 22045 -762 22062 -754
rect 22096 -762 22111 -754
rect 22045 -6730 22062 -6722
rect 22096 -6730 22111 -6722
rect 22045 -6742 22111 -6730
rect 22203 -754 22269 -742
rect 22203 -762 22220 -754
rect 22254 -762 22269 -754
rect 22203 -6730 22220 -6722
rect 22254 -6730 22269 -6722
rect 22203 -6742 22269 -6730
rect 22361 -754 22427 -742
rect 22361 -762 22378 -754
rect 22412 -762 22427 -754
rect 22361 -6730 22378 -6722
rect 22412 -6730 22427 -6722
rect 22361 -6742 22427 -6730
rect 22519 -754 22585 -742
rect 22519 -762 22536 -754
rect 22570 -762 22585 -754
rect 22519 -6730 22536 -6722
rect 22570 -6730 22585 -6722
rect 22519 -6742 22585 -6730
rect 22677 -754 22743 -742
rect 22677 -762 22694 -754
rect 22728 -762 22743 -754
rect 22677 -6730 22694 -6722
rect 22728 -6730 22743 -6722
rect 22677 -6742 22743 -6730
rect 22835 -754 22901 -742
rect 22835 -762 22852 -754
rect 22886 -762 22901 -754
rect 22835 -6730 22852 -6722
rect 22886 -6730 22901 -6722
rect 22835 -6742 22901 -6730
rect 22993 -754 23059 -742
rect 22993 -762 23010 -754
rect 23044 -762 23059 -754
rect 22993 -6730 23010 -6722
rect 23044 -6730 23059 -6722
rect 22993 -6742 23059 -6730
rect 23151 -754 23217 -742
rect 23151 -762 23168 -754
rect 23202 -762 23217 -754
rect 23151 -6730 23168 -6722
rect 23202 -6730 23217 -6722
rect 23151 -6742 23217 -6730
rect 23309 -754 23375 -742
rect 23309 -762 23326 -754
rect 23360 -762 23375 -754
rect 23309 -6730 23326 -6722
rect 23360 -6730 23375 -6722
rect 23309 -6742 23375 -6730
rect 23467 -754 23533 -742
rect 23467 -762 23484 -754
rect 23518 -762 23533 -754
rect 23467 -6730 23484 -6722
rect 23518 -6730 23533 -6722
rect 23467 -6742 23533 -6730
rect 23625 -754 23691 -742
rect 23625 -762 23642 -754
rect 23676 -762 23691 -754
rect 23625 -6730 23642 -6722
rect 23676 -6730 23691 -6722
rect 23625 -6742 23691 -6730
rect 23783 -754 23849 -742
rect 23783 -762 23800 -754
rect 23834 -762 23849 -754
rect 23783 -6730 23800 -6722
rect 23834 -6730 23849 -6722
rect 23783 -6742 23849 -6730
rect 23941 -754 24007 -742
rect 23941 -762 23958 -754
rect 23992 -762 24007 -754
rect 23941 -6730 23958 -6722
rect 23992 -6730 24007 -6722
rect 23941 -6742 24007 -6730
rect 24099 -754 24165 -742
rect 24099 -762 24116 -754
rect 24150 -762 24165 -754
rect 24099 -6730 24116 -6722
rect 24150 -6730 24165 -6722
rect 24099 -6742 24165 -6730
rect 24257 -754 24323 -742
rect 24257 -762 24274 -754
rect 24308 -762 24323 -754
rect 24257 -6730 24274 -6722
rect 24308 -6730 24323 -6722
rect 24257 -6742 24323 -6730
rect 24415 -754 24481 -742
rect 24415 -762 24432 -754
rect 24466 -762 24481 -754
rect 24415 -6730 24432 -6722
rect 24466 -6730 24481 -6722
rect 24415 -6742 24481 -6730
rect 24573 -754 24639 -742
rect 24573 -762 24590 -754
rect 24624 -762 24639 -754
rect 24573 -6730 24590 -6722
rect 24624 -6730 24639 -6722
rect 24573 -6742 24639 -6730
rect 24731 -754 24797 -742
rect 24731 -762 24748 -754
rect 24782 -762 24797 -754
rect 24731 -6730 24748 -6722
rect 24782 -6730 24797 -6722
rect 24731 -6742 24797 -6730
rect 24889 -754 24955 -742
rect 24889 -762 24906 -754
rect 24940 -762 24955 -754
rect 24889 -6730 24906 -6722
rect 24940 -6730 24955 -6722
rect 24889 -6742 24955 -6730
rect 25047 -754 25113 -742
rect 25047 -762 25064 -754
rect 25098 -762 25113 -754
rect 25047 -6730 25064 -6722
rect 25098 -6730 25113 -6722
rect 25047 -6742 25113 -6730
rect 25205 -754 25271 -742
rect 25205 -762 25222 -754
rect 25256 -762 25271 -754
rect 25205 -6730 25222 -6722
rect 25256 -6730 25271 -6722
rect 25205 -6742 25271 -6730
rect 20532 -6780 20552 -6774
rect 25186 -6780 25206 -6774
rect 20532 -6814 20544 -6780
rect 25194 -6814 25206 -6780
rect 20532 -6874 20552 -6814
rect 25186 -6874 25206 -6814
rect 20330 -6906 20400 -6900
rect 25340 -6906 25410 -6900
rect 20330 -6916 25410 -6906
rect 20330 -6954 20536 -6916
rect 25202 -6954 25410 -6916
rect 20330 -6970 25410 -6954
<< via1 >>
rect 1430 6280 1500 6420
rect 1652 6330 6286 6390
rect 1652 6296 1712 6330
rect 1712 6296 1802 6330
rect 1802 6296 1870 6330
rect 1870 6296 1960 6330
rect 1960 6296 2028 6330
rect 2028 6296 2118 6330
rect 2118 6296 2186 6330
rect 2186 6296 2276 6330
rect 2276 6296 2344 6330
rect 2344 6296 2434 6330
rect 2434 6296 2502 6330
rect 2502 6296 2592 6330
rect 2592 6296 2660 6330
rect 2660 6296 2750 6330
rect 2750 6296 2818 6330
rect 2818 6296 2908 6330
rect 2908 6296 2976 6330
rect 2976 6296 3066 6330
rect 3066 6296 3134 6330
rect 3134 6296 3224 6330
rect 3224 6296 3292 6330
rect 3292 6296 3382 6330
rect 3382 6296 3450 6330
rect 3450 6296 3540 6330
rect 3540 6296 3608 6330
rect 3608 6296 3698 6330
rect 3698 6296 3766 6330
rect 3766 6296 3856 6330
rect 3856 6296 3924 6330
rect 3924 6296 4014 6330
rect 4014 6296 4082 6330
rect 4082 6296 4172 6330
rect 4172 6296 4240 6330
rect 4240 6296 4330 6330
rect 4330 6296 4398 6330
rect 4398 6296 4488 6330
rect 4488 6296 4556 6330
rect 4556 6296 4646 6330
rect 4646 6296 4714 6330
rect 4714 6296 4804 6330
rect 4804 6296 4872 6330
rect 4872 6296 4962 6330
rect 4962 6296 5030 6330
rect 5030 6296 5120 6330
rect 5120 6296 5188 6330
rect 5188 6296 5278 6330
rect 5278 6296 5346 6330
rect 5346 6296 5436 6330
rect 5436 6296 5504 6330
rect 5504 6296 5594 6330
rect 5594 6296 5662 6330
rect 5662 6296 5752 6330
rect 5752 6296 5820 6330
rect 5820 6296 5910 6330
rect 5910 6296 5978 6330
rect 5978 6296 6068 6330
rect 6068 6296 6136 6330
rect 6136 6296 6226 6330
rect 6226 6296 6286 6330
rect 1652 6290 6286 6296
rect 1430 236 1446 6280
rect 1446 236 1484 6280
rect 1484 236 1500 6280
rect 6440 6280 6510 6420
rect 1565 278 1582 6238
rect 1582 278 1616 6238
rect 1616 278 1631 6238
rect 1723 278 1740 6238
rect 1740 278 1774 6238
rect 1774 278 1789 6238
rect 1881 278 1898 6238
rect 1898 278 1932 6238
rect 1932 278 1947 6238
rect 2039 278 2056 6238
rect 2056 278 2090 6238
rect 2090 278 2105 6238
rect 2197 278 2214 6238
rect 2214 278 2248 6238
rect 2248 278 2263 6238
rect 2355 278 2372 6238
rect 2372 278 2406 6238
rect 2406 278 2421 6238
rect 2513 278 2530 6238
rect 2530 278 2564 6238
rect 2564 278 2579 6238
rect 2671 278 2688 6238
rect 2688 278 2722 6238
rect 2722 278 2737 6238
rect 2829 278 2846 6238
rect 2846 278 2880 6238
rect 2880 278 2895 6238
rect 2987 278 3004 6238
rect 3004 278 3038 6238
rect 3038 278 3053 6238
rect 3145 278 3162 6238
rect 3162 278 3196 6238
rect 3196 278 3211 6238
rect 3303 278 3320 6238
rect 3320 278 3354 6238
rect 3354 278 3369 6238
rect 3461 278 3478 6238
rect 3478 278 3512 6238
rect 3512 278 3527 6238
rect 3619 278 3636 6238
rect 3636 278 3670 6238
rect 3670 278 3685 6238
rect 3777 278 3794 6238
rect 3794 278 3828 6238
rect 3828 278 3843 6238
rect 3935 278 3952 6238
rect 3952 278 3986 6238
rect 3986 278 4001 6238
rect 4093 278 4110 6238
rect 4110 278 4144 6238
rect 4144 278 4159 6238
rect 4251 278 4268 6238
rect 4268 278 4302 6238
rect 4302 278 4317 6238
rect 4409 278 4426 6238
rect 4426 278 4460 6238
rect 4460 278 4475 6238
rect 4567 278 4584 6238
rect 4584 278 4618 6238
rect 4618 278 4633 6238
rect 4725 278 4742 6238
rect 4742 278 4776 6238
rect 4776 278 4791 6238
rect 4883 278 4900 6238
rect 4900 278 4934 6238
rect 4934 278 4949 6238
rect 5041 278 5058 6238
rect 5058 278 5092 6238
rect 5092 278 5107 6238
rect 5199 278 5216 6238
rect 5216 278 5250 6238
rect 5250 278 5265 6238
rect 5357 278 5374 6238
rect 5374 278 5408 6238
rect 5408 278 5423 6238
rect 5515 278 5532 6238
rect 5532 278 5566 6238
rect 5566 278 5581 6238
rect 5673 278 5690 6238
rect 5690 278 5724 6238
rect 5724 278 5739 6238
rect 5831 278 5848 6238
rect 5848 278 5882 6238
rect 5882 278 5897 6238
rect 5989 278 6006 6238
rect 6006 278 6040 6238
rect 6040 278 6055 6238
rect 6147 278 6164 6238
rect 6164 278 6198 6238
rect 6198 278 6213 6238
rect 6305 278 6322 6238
rect 6322 278 6356 6238
rect 6356 278 6371 6238
rect 1430 100 1500 236
rect 6440 236 6454 6280
rect 6454 236 6492 6280
rect 6492 236 6510 6280
rect 1652 220 6286 226
rect 1652 186 1712 220
rect 1712 186 1802 220
rect 1802 186 1870 220
rect 1870 186 1960 220
rect 1960 186 2028 220
rect 2028 186 2118 220
rect 2118 186 2186 220
rect 2186 186 2276 220
rect 2276 186 2344 220
rect 2344 186 2434 220
rect 2434 186 2502 220
rect 2502 186 2592 220
rect 2592 186 2660 220
rect 2660 186 2750 220
rect 2750 186 2818 220
rect 2818 186 2908 220
rect 2908 186 2976 220
rect 2976 186 3066 220
rect 3066 186 3134 220
rect 3134 186 3224 220
rect 3224 186 3292 220
rect 3292 186 3382 220
rect 3382 186 3450 220
rect 3450 186 3540 220
rect 3540 186 3608 220
rect 3608 186 3698 220
rect 3698 186 3766 220
rect 3766 186 3856 220
rect 3856 186 3924 220
rect 3924 186 4014 220
rect 4014 186 4082 220
rect 4082 186 4172 220
rect 4172 186 4240 220
rect 4240 186 4330 220
rect 4330 186 4398 220
rect 4398 186 4488 220
rect 4488 186 4556 220
rect 4556 186 4646 220
rect 4646 186 4714 220
rect 4714 186 4804 220
rect 4804 186 4872 220
rect 4872 186 4962 220
rect 4962 186 5030 220
rect 5030 186 5120 220
rect 5120 186 5188 220
rect 5188 186 5278 220
rect 5278 186 5346 220
rect 5346 186 5436 220
rect 5436 186 5504 220
rect 5504 186 5594 220
rect 5594 186 5662 220
rect 5662 186 5752 220
rect 5752 186 5820 220
rect 5820 186 5910 220
rect 5910 186 5978 220
rect 5978 186 6068 220
rect 6068 186 6136 220
rect 6136 186 6226 220
rect 6226 186 6286 220
rect 1652 126 6286 186
rect 6440 100 6510 236
rect 7730 6280 7800 6420
rect 7952 6330 12586 6390
rect 7952 6296 8012 6330
rect 8012 6296 8102 6330
rect 8102 6296 8170 6330
rect 8170 6296 8260 6330
rect 8260 6296 8328 6330
rect 8328 6296 8418 6330
rect 8418 6296 8486 6330
rect 8486 6296 8576 6330
rect 8576 6296 8644 6330
rect 8644 6296 8734 6330
rect 8734 6296 8802 6330
rect 8802 6296 8892 6330
rect 8892 6296 8960 6330
rect 8960 6296 9050 6330
rect 9050 6296 9118 6330
rect 9118 6296 9208 6330
rect 9208 6296 9276 6330
rect 9276 6296 9366 6330
rect 9366 6296 9434 6330
rect 9434 6296 9524 6330
rect 9524 6296 9592 6330
rect 9592 6296 9682 6330
rect 9682 6296 9750 6330
rect 9750 6296 9840 6330
rect 9840 6296 9908 6330
rect 9908 6296 9998 6330
rect 9998 6296 10066 6330
rect 10066 6296 10156 6330
rect 10156 6296 10224 6330
rect 10224 6296 10314 6330
rect 10314 6296 10382 6330
rect 10382 6296 10472 6330
rect 10472 6296 10540 6330
rect 10540 6296 10630 6330
rect 10630 6296 10698 6330
rect 10698 6296 10788 6330
rect 10788 6296 10856 6330
rect 10856 6296 10946 6330
rect 10946 6296 11014 6330
rect 11014 6296 11104 6330
rect 11104 6296 11172 6330
rect 11172 6296 11262 6330
rect 11262 6296 11330 6330
rect 11330 6296 11420 6330
rect 11420 6296 11488 6330
rect 11488 6296 11578 6330
rect 11578 6296 11646 6330
rect 11646 6296 11736 6330
rect 11736 6296 11804 6330
rect 11804 6296 11894 6330
rect 11894 6296 11962 6330
rect 11962 6296 12052 6330
rect 12052 6296 12120 6330
rect 12120 6296 12210 6330
rect 12210 6296 12278 6330
rect 12278 6296 12368 6330
rect 12368 6296 12436 6330
rect 12436 6296 12526 6330
rect 12526 6296 12586 6330
rect 7952 6290 12586 6296
rect 7730 236 7746 6280
rect 7746 236 7784 6280
rect 7784 236 7800 6280
rect 12740 6280 12810 6420
rect 7865 278 7882 6238
rect 7882 278 7916 6238
rect 7916 278 7931 6238
rect 8023 278 8040 6238
rect 8040 278 8074 6238
rect 8074 278 8089 6238
rect 8181 278 8198 6238
rect 8198 278 8232 6238
rect 8232 278 8247 6238
rect 8339 278 8356 6238
rect 8356 278 8390 6238
rect 8390 278 8405 6238
rect 8497 278 8514 6238
rect 8514 278 8548 6238
rect 8548 278 8563 6238
rect 8655 278 8672 6238
rect 8672 278 8706 6238
rect 8706 278 8721 6238
rect 8813 278 8830 6238
rect 8830 278 8864 6238
rect 8864 278 8879 6238
rect 8971 278 8988 6238
rect 8988 278 9022 6238
rect 9022 278 9037 6238
rect 9129 278 9146 6238
rect 9146 278 9180 6238
rect 9180 278 9195 6238
rect 9287 278 9304 6238
rect 9304 278 9338 6238
rect 9338 278 9353 6238
rect 9445 278 9462 6238
rect 9462 278 9496 6238
rect 9496 278 9511 6238
rect 9603 278 9620 6238
rect 9620 278 9654 6238
rect 9654 278 9669 6238
rect 9761 278 9778 6238
rect 9778 278 9812 6238
rect 9812 278 9827 6238
rect 9919 278 9936 6238
rect 9936 278 9970 6238
rect 9970 278 9985 6238
rect 10077 278 10094 6238
rect 10094 278 10128 6238
rect 10128 278 10143 6238
rect 10235 278 10252 6238
rect 10252 278 10286 6238
rect 10286 278 10301 6238
rect 10393 278 10410 6238
rect 10410 278 10444 6238
rect 10444 278 10459 6238
rect 10551 278 10568 6238
rect 10568 278 10602 6238
rect 10602 278 10617 6238
rect 10709 278 10726 6238
rect 10726 278 10760 6238
rect 10760 278 10775 6238
rect 10867 278 10884 6238
rect 10884 278 10918 6238
rect 10918 278 10933 6238
rect 11025 278 11042 6238
rect 11042 278 11076 6238
rect 11076 278 11091 6238
rect 11183 278 11200 6238
rect 11200 278 11234 6238
rect 11234 278 11249 6238
rect 11341 278 11358 6238
rect 11358 278 11392 6238
rect 11392 278 11407 6238
rect 11499 278 11516 6238
rect 11516 278 11550 6238
rect 11550 278 11565 6238
rect 11657 278 11674 6238
rect 11674 278 11708 6238
rect 11708 278 11723 6238
rect 11815 278 11832 6238
rect 11832 278 11866 6238
rect 11866 278 11881 6238
rect 11973 278 11990 6238
rect 11990 278 12024 6238
rect 12024 278 12039 6238
rect 12131 278 12148 6238
rect 12148 278 12182 6238
rect 12182 278 12197 6238
rect 12289 278 12306 6238
rect 12306 278 12340 6238
rect 12340 278 12355 6238
rect 12447 278 12464 6238
rect 12464 278 12498 6238
rect 12498 278 12513 6238
rect 12605 278 12622 6238
rect 12622 278 12656 6238
rect 12656 278 12671 6238
rect 7730 100 7800 236
rect 12740 236 12754 6280
rect 12754 236 12792 6280
rect 12792 236 12810 6280
rect 7952 220 12586 226
rect 7952 186 8012 220
rect 8012 186 8102 220
rect 8102 186 8170 220
rect 8170 186 8260 220
rect 8260 186 8328 220
rect 8328 186 8418 220
rect 8418 186 8486 220
rect 8486 186 8576 220
rect 8576 186 8644 220
rect 8644 186 8734 220
rect 8734 186 8802 220
rect 8802 186 8892 220
rect 8892 186 8960 220
rect 8960 186 9050 220
rect 9050 186 9118 220
rect 9118 186 9208 220
rect 9208 186 9276 220
rect 9276 186 9366 220
rect 9366 186 9434 220
rect 9434 186 9524 220
rect 9524 186 9592 220
rect 9592 186 9682 220
rect 9682 186 9750 220
rect 9750 186 9840 220
rect 9840 186 9908 220
rect 9908 186 9998 220
rect 9998 186 10066 220
rect 10066 186 10156 220
rect 10156 186 10224 220
rect 10224 186 10314 220
rect 10314 186 10382 220
rect 10382 186 10472 220
rect 10472 186 10540 220
rect 10540 186 10630 220
rect 10630 186 10698 220
rect 10698 186 10788 220
rect 10788 186 10856 220
rect 10856 186 10946 220
rect 10946 186 11014 220
rect 11014 186 11104 220
rect 11104 186 11172 220
rect 11172 186 11262 220
rect 11262 186 11330 220
rect 11330 186 11420 220
rect 11420 186 11488 220
rect 11488 186 11578 220
rect 11578 186 11646 220
rect 11646 186 11736 220
rect 11736 186 11804 220
rect 11804 186 11894 220
rect 11894 186 11962 220
rect 11962 186 12052 220
rect 12052 186 12120 220
rect 12120 186 12210 220
rect 12210 186 12278 220
rect 12278 186 12368 220
rect 12368 186 12436 220
rect 12436 186 12526 220
rect 12526 186 12586 220
rect 7952 126 12586 186
rect 12740 100 12810 236
rect 14030 6280 14100 6420
rect 14252 6330 18886 6390
rect 14252 6296 14312 6330
rect 14312 6296 14402 6330
rect 14402 6296 14470 6330
rect 14470 6296 14560 6330
rect 14560 6296 14628 6330
rect 14628 6296 14718 6330
rect 14718 6296 14786 6330
rect 14786 6296 14876 6330
rect 14876 6296 14944 6330
rect 14944 6296 15034 6330
rect 15034 6296 15102 6330
rect 15102 6296 15192 6330
rect 15192 6296 15260 6330
rect 15260 6296 15350 6330
rect 15350 6296 15418 6330
rect 15418 6296 15508 6330
rect 15508 6296 15576 6330
rect 15576 6296 15666 6330
rect 15666 6296 15734 6330
rect 15734 6296 15824 6330
rect 15824 6296 15892 6330
rect 15892 6296 15982 6330
rect 15982 6296 16050 6330
rect 16050 6296 16140 6330
rect 16140 6296 16208 6330
rect 16208 6296 16298 6330
rect 16298 6296 16366 6330
rect 16366 6296 16456 6330
rect 16456 6296 16524 6330
rect 16524 6296 16614 6330
rect 16614 6296 16682 6330
rect 16682 6296 16772 6330
rect 16772 6296 16840 6330
rect 16840 6296 16930 6330
rect 16930 6296 16998 6330
rect 16998 6296 17088 6330
rect 17088 6296 17156 6330
rect 17156 6296 17246 6330
rect 17246 6296 17314 6330
rect 17314 6296 17404 6330
rect 17404 6296 17472 6330
rect 17472 6296 17562 6330
rect 17562 6296 17630 6330
rect 17630 6296 17720 6330
rect 17720 6296 17788 6330
rect 17788 6296 17878 6330
rect 17878 6296 17946 6330
rect 17946 6296 18036 6330
rect 18036 6296 18104 6330
rect 18104 6296 18194 6330
rect 18194 6296 18262 6330
rect 18262 6296 18352 6330
rect 18352 6296 18420 6330
rect 18420 6296 18510 6330
rect 18510 6296 18578 6330
rect 18578 6296 18668 6330
rect 18668 6296 18736 6330
rect 18736 6296 18826 6330
rect 18826 6296 18886 6330
rect 14252 6290 18886 6296
rect 14030 236 14046 6280
rect 14046 236 14084 6280
rect 14084 236 14100 6280
rect 19040 6280 19110 6420
rect 14165 278 14182 6238
rect 14182 278 14216 6238
rect 14216 278 14231 6238
rect 14323 278 14340 6238
rect 14340 278 14374 6238
rect 14374 278 14389 6238
rect 14481 278 14498 6238
rect 14498 278 14532 6238
rect 14532 278 14547 6238
rect 14639 278 14656 6238
rect 14656 278 14690 6238
rect 14690 278 14705 6238
rect 14797 278 14814 6238
rect 14814 278 14848 6238
rect 14848 278 14863 6238
rect 14955 278 14972 6238
rect 14972 278 15006 6238
rect 15006 278 15021 6238
rect 15113 278 15130 6238
rect 15130 278 15164 6238
rect 15164 278 15179 6238
rect 15271 278 15288 6238
rect 15288 278 15322 6238
rect 15322 278 15337 6238
rect 15429 278 15446 6238
rect 15446 278 15480 6238
rect 15480 278 15495 6238
rect 15587 278 15604 6238
rect 15604 278 15638 6238
rect 15638 278 15653 6238
rect 15745 278 15762 6238
rect 15762 278 15796 6238
rect 15796 278 15811 6238
rect 15903 278 15920 6238
rect 15920 278 15954 6238
rect 15954 278 15969 6238
rect 16061 278 16078 6238
rect 16078 278 16112 6238
rect 16112 278 16127 6238
rect 16219 278 16236 6238
rect 16236 278 16270 6238
rect 16270 278 16285 6238
rect 16377 278 16394 6238
rect 16394 278 16428 6238
rect 16428 278 16443 6238
rect 16535 278 16552 6238
rect 16552 278 16586 6238
rect 16586 278 16601 6238
rect 16693 278 16710 6238
rect 16710 278 16744 6238
rect 16744 278 16759 6238
rect 16851 278 16868 6238
rect 16868 278 16902 6238
rect 16902 278 16917 6238
rect 17009 278 17026 6238
rect 17026 278 17060 6238
rect 17060 278 17075 6238
rect 17167 278 17184 6238
rect 17184 278 17218 6238
rect 17218 278 17233 6238
rect 17325 278 17342 6238
rect 17342 278 17376 6238
rect 17376 278 17391 6238
rect 17483 278 17500 6238
rect 17500 278 17534 6238
rect 17534 278 17549 6238
rect 17641 278 17658 6238
rect 17658 278 17692 6238
rect 17692 278 17707 6238
rect 17799 278 17816 6238
rect 17816 278 17850 6238
rect 17850 278 17865 6238
rect 17957 278 17974 6238
rect 17974 278 18008 6238
rect 18008 278 18023 6238
rect 18115 278 18132 6238
rect 18132 278 18166 6238
rect 18166 278 18181 6238
rect 18273 278 18290 6238
rect 18290 278 18324 6238
rect 18324 278 18339 6238
rect 18431 278 18448 6238
rect 18448 278 18482 6238
rect 18482 278 18497 6238
rect 18589 278 18606 6238
rect 18606 278 18640 6238
rect 18640 278 18655 6238
rect 18747 278 18764 6238
rect 18764 278 18798 6238
rect 18798 278 18813 6238
rect 18905 278 18922 6238
rect 18922 278 18956 6238
rect 18956 278 18971 6238
rect 14030 100 14100 236
rect 19040 236 19054 6280
rect 19054 236 19092 6280
rect 19092 236 19110 6280
rect 14252 220 18886 226
rect 14252 186 14312 220
rect 14312 186 14402 220
rect 14402 186 14470 220
rect 14470 186 14560 220
rect 14560 186 14628 220
rect 14628 186 14718 220
rect 14718 186 14786 220
rect 14786 186 14876 220
rect 14876 186 14944 220
rect 14944 186 15034 220
rect 15034 186 15102 220
rect 15102 186 15192 220
rect 15192 186 15260 220
rect 15260 186 15350 220
rect 15350 186 15418 220
rect 15418 186 15508 220
rect 15508 186 15576 220
rect 15576 186 15666 220
rect 15666 186 15734 220
rect 15734 186 15824 220
rect 15824 186 15892 220
rect 15892 186 15982 220
rect 15982 186 16050 220
rect 16050 186 16140 220
rect 16140 186 16208 220
rect 16208 186 16298 220
rect 16298 186 16366 220
rect 16366 186 16456 220
rect 16456 186 16524 220
rect 16524 186 16614 220
rect 16614 186 16682 220
rect 16682 186 16772 220
rect 16772 186 16840 220
rect 16840 186 16930 220
rect 16930 186 16998 220
rect 16998 186 17088 220
rect 17088 186 17156 220
rect 17156 186 17246 220
rect 17246 186 17314 220
rect 17314 186 17404 220
rect 17404 186 17472 220
rect 17472 186 17562 220
rect 17562 186 17630 220
rect 17630 186 17720 220
rect 17720 186 17788 220
rect 17788 186 17878 220
rect 17878 186 17946 220
rect 17946 186 18036 220
rect 18036 186 18104 220
rect 18104 186 18194 220
rect 18194 186 18262 220
rect 18262 186 18352 220
rect 18352 186 18420 220
rect 18420 186 18510 220
rect 18510 186 18578 220
rect 18578 186 18668 220
rect 18668 186 18736 220
rect 18736 186 18826 220
rect 18826 186 18886 220
rect 14252 126 18886 186
rect 19040 100 19110 236
rect 20330 6280 20400 6420
rect 20552 6330 25186 6390
rect 20552 6296 20612 6330
rect 20612 6296 20702 6330
rect 20702 6296 20770 6330
rect 20770 6296 20860 6330
rect 20860 6296 20928 6330
rect 20928 6296 21018 6330
rect 21018 6296 21086 6330
rect 21086 6296 21176 6330
rect 21176 6296 21244 6330
rect 21244 6296 21334 6330
rect 21334 6296 21402 6330
rect 21402 6296 21492 6330
rect 21492 6296 21560 6330
rect 21560 6296 21650 6330
rect 21650 6296 21718 6330
rect 21718 6296 21808 6330
rect 21808 6296 21876 6330
rect 21876 6296 21966 6330
rect 21966 6296 22034 6330
rect 22034 6296 22124 6330
rect 22124 6296 22192 6330
rect 22192 6296 22282 6330
rect 22282 6296 22350 6330
rect 22350 6296 22440 6330
rect 22440 6296 22508 6330
rect 22508 6296 22598 6330
rect 22598 6296 22666 6330
rect 22666 6296 22756 6330
rect 22756 6296 22824 6330
rect 22824 6296 22914 6330
rect 22914 6296 22982 6330
rect 22982 6296 23072 6330
rect 23072 6296 23140 6330
rect 23140 6296 23230 6330
rect 23230 6296 23298 6330
rect 23298 6296 23388 6330
rect 23388 6296 23456 6330
rect 23456 6296 23546 6330
rect 23546 6296 23614 6330
rect 23614 6296 23704 6330
rect 23704 6296 23772 6330
rect 23772 6296 23862 6330
rect 23862 6296 23930 6330
rect 23930 6296 24020 6330
rect 24020 6296 24088 6330
rect 24088 6296 24178 6330
rect 24178 6296 24246 6330
rect 24246 6296 24336 6330
rect 24336 6296 24404 6330
rect 24404 6296 24494 6330
rect 24494 6296 24562 6330
rect 24562 6296 24652 6330
rect 24652 6296 24720 6330
rect 24720 6296 24810 6330
rect 24810 6296 24878 6330
rect 24878 6296 24968 6330
rect 24968 6296 25036 6330
rect 25036 6296 25126 6330
rect 25126 6296 25186 6330
rect 20552 6290 25186 6296
rect 20330 236 20346 6280
rect 20346 236 20384 6280
rect 20384 236 20400 6280
rect 25340 6280 25410 6420
rect 20465 278 20482 6238
rect 20482 278 20516 6238
rect 20516 278 20531 6238
rect 20623 278 20640 6238
rect 20640 278 20674 6238
rect 20674 278 20689 6238
rect 20781 278 20798 6238
rect 20798 278 20832 6238
rect 20832 278 20847 6238
rect 20939 278 20956 6238
rect 20956 278 20990 6238
rect 20990 278 21005 6238
rect 21097 278 21114 6238
rect 21114 278 21148 6238
rect 21148 278 21163 6238
rect 21255 278 21272 6238
rect 21272 278 21306 6238
rect 21306 278 21321 6238
rect 21413 278 21430 6238
rect 21430 278 21464 6238
rect 21464 278 21479 6238
rect 21571 278 21588 6238
rect 21588 278 21622 6238
rect 21622 278 21637 6238
rect 21729 278 21746 6238
rect 21746 278 21780 6238
rect 21780 278 21795 6238
rect 21887 278 21904 6238
rect 21904 278 21938 6238
rect 21938 278 21953 6238
rect 22045 278 22062 6238
rect 22062 278 22096 6238
rect 22096 278 22111 6238
rect 22203 278 22220 6238
rect 22220 278 22254 6238
rect 22254 278 22269 6238
rect 22361 278 22378 6238
rect 22378 278 22412 6238
rect 22412 278 22427 6238
rect 22519 278 22536 6238
rect 22536 278 22570 6238
rect 22570 278 22585 6238
rect 22677 278 22694 6238
rect 22694 278 22728 6238
rect 22728 278 22743 6238
rect 22835 278 22852 6238
rect 22852 278 22886 6238
rect 22886 278 22901 6238
rect 22993 278 23010 6238
rect 23010 278 23044 6238
rect 23044 278 23059 6238
rect 23151 278 23168 6238
rect 23168 278 23202 6238
rect 23202 278 23217 6238
rect 23309 278 23326 6238
rect 23326 278 23360 6238
rect 23360 278 23375 6238
rect 23467 278 23484 6238
rect 23484 278 23518 6238
rect 23518 278 23533 6238
rect 23625 278 23642 6238
rect 23642 278 23676 6238
rect 23676 278 23691 6238
rect 23783 278 23800 6238
rect 23800 278 23834 6238
rect 23834 278 23849 6238
rect 23941 278 23958 6238
rect 23958 278 23992 6238
rect 23992 278 24007 6238
rect 24099 278 24116 6238
rect 24116 278 24150 6238
rect 24150 278 24165 6238
rect 24257 278 24274 6238
rect 24274 278 24308 6238
rect 24308 278 24323 6238
rect 24415 278 24432 6238
rect 24432 278 24466 6238
rect 24466 278 24481 6238
rect 24573 278 24590 6238
rect 24590 278 24624 6238
rect 24624 278 24639 6238
rect 24731 278 24748 6238
rect 24748 278 24782 6238
rect 24782 278 24797 6238
rect 24889 278 24906 6238
rect 24906 278 24940 6238
rect 24940 278 24955 6238
rect 25047 278 25064 6238
rect 25064 278 25098 6238
rect 25098 278 25113 6238
rect 25205 278 25222 6238
rect 25222 278 25256 6238
rect 25256 278 25271 6238
rect 20330 100 20400 236
rect 25340 236 25354 6280
rect 25354 236 25392 6280
rect 25392 236 25410 6280
rect 20552 220 25186 226
rect 20552 186 20612 220
rect 20612 186 20702 220
rect 20702 186 20770 220
rect 20770 186 20860 220
rect 20860 186 20928 220
rect 20928 186 21018 220
rect 21018 186 21086 220
rect 21086 186 21176 220
rect 21176 186 21244 220
rect 21244 186 21334 220
rect 21334 186 21402 220
rect 21402 186 21492 220
rect 21492 186 21560 220
rect 21560 186 21650 220
rect 21650 186 21718 220
rect 21718 186 21808 220
rect 21808 186 21876 220
rect 21876 186 21966 220
rect 21966 186 22034 220
rect 22034 186 22124 220
rect 22124 186 22192 220
rect 22192 186 22282 220
rect 22282 186 22350 220
rect 22350 186 22440 220
rect 22440 186 22508 220
rect 22508 186 22598 220
rect 22598 186 22666 220
rect 22666 186 22756 220
rect 22756 186 22824 220
rect 22824 186 22914 220
rect 22914 186 22982 220
rect 22982 186 23072 220
rect 23072 186 23140 220
rect 23140 186 23230 220
rect 23230 186 23298 220
rect 23298 186 23388 220
rect 23388 186 23456 220
rect 23456 186 23546 220
rect 23546 186 23614 220
rect 23614 186 23704 220
rect 23704 186 23772 220
rect 23772 186 23862 220
rect 23862 186 23930 220
rect 23930 186 24020 220
rect 24020 186 24088 220
rect 24088 186 24178 220
rect 24178 186 24246 220
rect 24246 186 24336 220
rect 24336 186 24404 220
rect 24404 186 24494 220
rect 24494 186 24562 220
rect 24562 186 24652 220
rect 24652 186 24720 220
rect 24720 186 24810 220
rect 24810 186 24878 220
rect 24878 186 24968 220
rect 24968 186 25036 220
rect 25036 186 25126 220
rect 25126 186 25186 220
rect 20552 126 25186 186
rect 25340 100 25410 236
rect 1430 -720 1500 -580
rect 1652 -670 6286 -610
rect 1652 -704 1712 -670
rect 1712 -704 1802 -670
rect 1802 -704 1870 -670
rect 1870 -704 1960 -670
rect 1960 -704 2028 -670
rect 2028 -704 2118 -670
rect 2118 -704 2186 -670
rect 2186 -704 2276 -670
rect 2276 -704 2344 -670
rect 2344 -704 2434 -670
rect 2434 -704 2502 -670
rect 2502 -704 2592 -670
rect 2592 -704 2660 -670
rect 2660 -704 2750 -670
rect 2750 -704 2818 -670
rect 2818 -704 2908 -670
rect 2908 -704 2976 -670
rect 2976 -704 3066 -670
rect 3066 -704 3134 -670
rect 3134 -704 3224 -670
rect 3224 -704 3292 -670
rect 3292 -704 3382 -670
rect 3382 -704 3450 -670
rect 3450 -704 3540 -670
rect 3540 -704 3608 -670
rect 3608 -704 3698 -670
rect 3698 -704 3766 -670
rect 3766 -704 3856 -670
rect 3856 -704 3924 -670
rect 3924 -704 4014 -670
rect 4014 -704 4082 -670
rect 4082 -704 4172 -670
rect 4172 -704 4240 -670
rect 4240 -704 4330 -670
rect 4330 -704 4398 -670
rect 4398 -704 4488 -670
rect 4488 -704 4556 -670
rect 4556 -704 4646 -670
rect 4646 -704 4714 -670
rect 4714 -704 4804 -670
rect 4804 -704 4872 -670
rect 4872 -704 4962 -670
rect 4962 -704 5030 -670
rect 5030 -704 5120 -670
rect 5120 -704 5188 -670
rect 5188 -704 5278 -670
rect 5278 -704 5346 -670
rect 5346 -704 5436 -670
rect 5436 -704 5504 -670
rect 5504 -704 5594 -670
rect 5594 -704 5662 -670
rect 5662 -704 5752 -670
rect 5752 -704 5820 -670
rect 5820 -704 5910 -670
rect 5910 -704 5978 -670
rect 5978 -704 6068 -670
rect 6068 -704 6136 -670
rect 6136 -704 6226 -670
rect 6226 -704 6286 -670
rect 1652 -710 6286 -704
rect 1430 -6764 1446 -720
rect 1446 -6764 1484 -720
rect 1484 -6764 1500 -720
rect 6440 -720 6510 -580
rect 1565 -6722 1582 -762
rect 1582 -6722 1616 -762
rect 1616 -6722 1631 -762
rect 1723 -6722 1740 -762
rect 1740 -6722 1774 -762
rect 1774 -6722 1789 -762
rect 1881 -6722 1898 -762
rect 1898 -6722 1932 -762
rect 1932 -6722 1947 -762
rect 2039 -6722 2056 -762
rect 2056 -6722 2090 -762
rect 2090 -6722 2105 -762
rect 2197 -6722 2214 -762
rect 2214 -6722 2248 -762
rect 2248 -6722 2263 -762
rect 2355 -6722 2372 -762
rect 2372 -6722 2406 -762
rect 2406 -6722 2421 -762
rect 2513 -6722 2530 -762
rect 2530 -6722 2564 -762
rect 2564 -6722 2579 -762
rect 2671 -6722 2688 -762
rect 2688 -6722 2722 -762
rect 2722 -6722 2737 -762
rect 2829 -6722 2846 -762
rect 2846 -6722 2880 -762
rect 2880 -6722 2895 -762
rect 2987 -6722 3004 -762
rect 3004 -6722 3038 -762
rect 3038 -6722 3053 -762
rect 3145 -6722 3162 -762
rect 3162 -6722 3196 -762
rect 3196 -6722 3211 -762
rect 3303 -6722 3320 -762
rect 3320 -6722 3354 -762
rect 3354 -6722 3369 -762
rect 3461 -6722 3478 -762
rect 3478 -6722 3512 -762
rect 3512 -6722 3527 -762
rect 3619 -6722 3636 -762
rect 3636 -6722 3670 -762
rect 3670 -6722 3685 -762
rect 3777 -6722 3794 -762
rect 3794 -6722 3828 -762
rect 3828 -6722 3843 -762
rect 3935 -6722 3952 -762
rect 3952 -6722 3986 -762
rect 3986 -6722 4001 -762
rect 4093 -6722 4110 -762
rect 4110 -6722 4144 -762
rect 4144 -6722 4159 -762
rect 4251 -6722 4268 -762
rect 4268 -6722 4302 -762
rect 4302 -6722 4317 -762
rect 4409 -6722 4426 -762
rect 4426 -6722 4460 -762
rect 4460 -6722 4475 -762
rect 4567 -6722 4584 -762
rect 4584 -6722 4618 -762
rect 4618 -6722 4633 -762
rect 4725 -6722 4742 -762
rect 4742 -6722 4776 -762
rect 4776 -6722 4791 -762
rect 4883 -6722 4900 -762
rect 4900 -6722 4934 -762
rect 4934 -6722 4949 -762
rect 5041 -6722 5058 -762
rect 5058 -6722 5092 -762
rect 5092 -6722 5107 -762
rect 5199 -6722 5216 -762
rect 5216 -6722 5250 -762
rect 5250 -6722 5265 -762
rect 5357 -6722 5374 -762
rect 5374 -6722 5408 -762
rect 5408 -6722 5423 -762
rect 5515 -6722 5532 -762
rect 5532 -6722 5566 -762
rect 5566 -6722 5581 -762
rect 5673 -6722 5690 -762
rect 5690 -6722 5724 -762
rect 5724 -6722 5739 -762
rect 5831 -6722 5848 -762
rect 5848 -6722 5882 -762
rect 5882 -6722 5897 -762
rect 5989 -6722 6006 -762
rect 6006 -6722 6040 -762
rect 6040 -6722 6055 -762
rect 6147 -6722 6164 -762
rect 6164 -6722 6198 -762
rect 6198 -6722 6213 -762
rect 6305 -6722 6322 -762
rect 6322 -6722 6356 -762
rect 6356 -6722 6371 -762
rect 1430 -6900 1500 -6764
rect 6440 -6764 6454 -720
rect 6454 -6764 6492 -720
rect 6492 -6764 6510 -720
rect 1652 -6780 6286 -6774
rect 1652 -6814 1712 -6780
rect 1712 -6814 1802 -6780
rect 1802 -6814 1870 -6780
rect 1870 -6814 1960 -6780
rect 1960 -6814 2028 -6780
rect 2028 -6814 2118 -6780
rect 2118 -6814 2186 -6780
rect 2186 -6814 2276 -6780
rect 2276 -6814 2344 -6780
rect 2344 -6814 2434 -6780
rect 2434 -6814 2502 -6780
rect 2502 -6814 2592 -6780
rect 2592 -6814 2660 -6780
rect 2660 -6814 2750 -6780
rect 2750 -6814 2818 -6780
rect 2818 -6814 2908 -6780
rect 2908 -6814 2976 -6780
rect 2976 -6814 3066 -6780
rect 3066 -6814 3134 -6780
rect 3134 -6814 3224 -6780
rect 3224 -6814 3292 -6780
rect 3292 -6814 3382 -6780
rect 3382 -6814 3450 -6780
rect 3450 -6814 3540 -6780
rect 3540 -6814 3608 -6780
rect 3608 -6814 3698 -6780
rect 3698 -6814 3766 -6780
rect 3766 -6814 3856 -6780
rect 3856 -6814 3924 -6780
rect 3924 -6814 4014 -6780
rect 4014 -6814 4082 -6780
rect 4082 -6814 4172 -6780
rect 4172 -6814 4240 -6780
rect 4240 -6814 4330 -6780
rect 4330 -6814 4398 -6780
rect 4398 -6814 4488 -6780
rect 4488 -6814 4556 -6780
rect 4556 -6814 4646 -6780
rect 4646 -6814 4714 -6780
rect 4714 -6814 4804 -6780
rect 4804 -6814 4872 -6780
rect 4872 -6814 4962 -6780
rect 4962 -6814 5030 -6780
rect 5030 -6814 5120 -6780
rect 5120 -6814 5188 -6780
rect 5188 -6814 5278 -6780
rect 5278 -6814 5346 -6780
rect 5346 -6814 5436 -6780
rect 5436 -6814 5504 -6780
rect 5504 -6814 5594 -6780
rect 5594 -6814 5662 -6780
rect 5662 -6814 5752 -6780
rect 5752 -6814 5820 -6780
rect 5820 -6814 5910 -6780
rect 5910 -6814 5978 -6780
rect 5978 -6814 6068 -6780
rect 6068 -6814 6136 -6780
rect 6136 -6814 6226 -6780
rect 6226 -6814 6286 -6780
rect 1652 -6874 6286 -6814
rect 6440 -6900 6510 -6764
rect 7730 -720 7800 -580
rect 7952 -670 12586 -610
rect 7952 -704 8012 -670
rect 8012 -704 8102 -670
rect 8102 -704 8170 -670
rect 8170 -704 8260 -670
rect 8260 -704 8328 -670
rect 8328 -704 8418 -670
rect 8418 -704 8486 -670
rect 8486 -704 8576 -670
rect 8576 -704 8644 -670
rect 8644 -704 8734 -670
rect 8734 -704 8802 -670
rect 8802 -704 8892 -670
rect 8892 -704 8960 -670
rect 8960 -704 9050 -670
rect 9050 -704 9118 -670
rect 9118 -704 9208 -670
rect 9208 -704 9276 -670
rect 9276 -704 9366 -670
rect 9366 -704 9434 -670
rect 9434 -704 9524 -670
rect 9524 -704 9592 -670
rect 9592 -704 9682 -670
rect 9682 -704 9750 -670
rect 9750 -704 9840 -670
rect 9840 -704 9908 -670
rect 9908 -704 9998 -670
rect 9998 -704 10066 -670
rect 10066 -704 10156 -670
rect 10156 -704 10224 -670
rect 10224 -704 10314 -670
rect 10314 -704 10382 -670
rect 10382 -704 10472 -670
rect 10472 -704 10540 -670
rect 10540 -704 10630 -670
rect 10630 -704 10698 -670
rect 10698 -704 10788 -670
rect 10788 -704 10856 -670
rect 10856 -704 10946 -670
rect 10946 -704 11014 -670
rect 11014 -704 11104 -670
rect 11104 -704 11172 -670
rect 11172 -704 11262 -670
rect 11262 -704 11330 -670
rect 11330 -704 11420 -670
rect 11420 -704 11488 -670
rect 11488 -704 11578 -670
rect 11578 -704 11646 -670
rect 11646 -704 11736 -670
rect 11736 -704 11804 -670
rect 11804 -704 11894 -670
rect 11894 -704 11962 -670
rect 11962 -704 12052 -670
rect 12052 -704 12120 -670
rect 12120 -704 12210 -670
rect 12210 -704 12278 -670
rect 12278 -704 12368 -670
rect 12368 -704 12436 -670
rect 12436 -704 12526 -670
rect 12526 -704 12586 -670
rect 7952 -710 12586 -704
rect 7730 -6764 7746 -720
rect 7746 -6764 7784 -720
rect 7784 -6764 7800 -720
rect 12740 -720 12810 -580
rect 7865 -6722 7882 -762
rect 7882 -6722 7916 -762
rect 7916 -6722 7931 -762
rect 8023 -6722 8040 -762
rect 8040 -6722 8074 -762
rect 8074 -6722 8089 -762
rect 8181 -6722 8198 -762
rect 8198 -6722 8232 -762
rect 8232 -6722 8247 -762
rect 8339 -6722 8356 -762
rect 8356 -6722 8390 -762
rect 8390 -6722 8405 -762
rect 8497 -6722 8514 -762
rect 8514 -6722 8548 -762
rect 8548 -6722 8563 -762
rect 8655 -6722 8672 -762
rect 8672 -6722 8706 -762
rect 8706 -6722 8721 -762
rect 8813 -6722 8830 -762
rect 8830 -6722 8864 -762
rect 8864 -6722 8879 -762
rect 8971 -6722 8988 -762
rect 8988 -6722 9022 -762
rect 9022 -6722 9037 -762
rect 9129 -6722 9146 -762
rect 9146 -6722 9180 -762
rect 9180 -6722 9195 -762
rect 9287 -6722 9304 -762
rect 9304 -6722 9338 -762
rect 9338 -6722 9353 -762
rect 9445 -6722 9462 -762
rect 9462 -6722 9496 -762
rect 9496 -6722 9511 -762
rect 9603 -6722 9620 -762
rect 9620 -6722 9654 -762
rect 9654 -6722 9669 -762
rect 9761 -6722 9778 -762
rect 9778 -6722 9812 -762
rect 9812 -6722 9827 -762
rect 9919 -6722 9936 -762
rect 9936 -6722 9970 -762
rect 9970 -6722 9985 -762
rect 10077 -6722 10094 -762
rect 10094 -6722 10128 -762
rect 10128 -6722 10143 -762
rect 10235 -6722 10252 -762
rect 10252 -6722 10286 -762
rect 10286 -6722 10301 -762
rect 10393 -6722 10410 -762
rect 10410 -6722 10444 -762
rect 10444 -6722 10459 -762
rect 10551 -6722 10568 -762
rect 10568 -6722 10602 -762
rect 10602 -6722 10617 -762
rect 10709 -6722 10726 -762
rect 10726 -6722 10760 -762
rect 10760 -6722 10775 -762
rect 10867 -6722 10884 -762
rect 10884 -6722 10918 -762
rect 10918 -6722 10933 -762
rect 11025 -6722 11042 -762
rect 11042 -6722 11076 -762
rect 11076 -6722 11091 -762
rect 11183 -6722 11200 -762
rect 11200 -6722 11234 -762
rect 11234 -6722 11249 -762
rect 11341 -6722 11358 -762
rect 11358 -6722 11392 -762
rect 11392 -6722 11407 -762
rect 11499 -6722 11516 -762
rect 11516 -6722 11550 -762
rect 11550 -6722 11565 -762
rect 11657 -6722 11674 -762
rect 11674 -6722 11708 -762
rect 11708 -6722 11723 -762
rect 11815 -6722 11832 -762
rect 11832 -6722 11866 -762
rect 11866 -6722 11881 -762
rect 11973 -6722 11990 -762
rect 11990 -6722 12024 -762
rect 12024 -6722 12039 -762
rect 12131 -6722 12148 -762
rect 12148 -6722 12182 -762
rect 12182 -6722 12197 -762
rect 12289 -6722 12306 -762
rect 12306 -6722 12340 -762
rect 12340 -6722 12355 -762
rect 12447 -6722 12464 -762
rect 12464 -6722 12498 -762
rect 12498 -6722 12513 -762
rect 12605 -6722 12622 -762
rect 12622 -6722 12656 -762
rect 12656 -6722 12671 -762
rect 7730 -6900 7800 -6764
rect 12740 -6764 12754 -720
rect 12754 -6764 12792 -720
rect 12792 -6764 12810 -720
rect 7952 -6780 12586 -6774
rect 7952 -6814 8012 -6780
rect 8012 -6814 8102 -6780
rect 8102 -6814 8170 -6780
rect 8170 -6814 8260 -6780
rect 8260 -6814 8328 -6780
rect 8328 -6814 8418 -6780
rect 8418 -6814 8486 -6780
rect 8486 -6814 8576 -6780
rect 8576 -6814 8644 -6780
rect 8644 -6814 8734 -6780
rect 8734 -6814 8802 -6780
rect 8802 -6814 8892 -6780
rect 8892 -6814 8960 -6780
rect 8960 -6814 9050 -6780
rect 9050 -6814 9118 -6780
rect 9118 -6814 9208 -6780
rect 9208 -6814 9276 -6780
rect 9276 -6814 9366 -6780
rect 9366 -6814 9434 -6780
rect 9434 -6814 9524 -6780
rect 9524 -6814 9592 -6780
rect 9592 -6814 9682 -6780
rect 9682 -6814 9750 -6780
rect 9750 -6814 9840 -6780
rect 9840 -6814 9908 -6780
rect 9908 -6814 9998 -6780
rect 9998 -6814 10066 -6780
rect 10066 -6814 10156 -6780
rect 10156 -6814 10224 -6780
rect 10224 -6814 10314 -6780
rect 10314 -6814 10382 -6780
rect 10382 -6814 10472 -6780
rect 10472 -6814 10540 -6780
rect 10540 -6814 10630 -6780
rect 10630 -6814 10698 -6780
rect 10698 -6814 10788 -6780
rect 10788 -6814 10856 -6780
rect 10856 -6814 10946 -6780
rect 10946 -6814 11014 -6780
rect 11014 -6814 11104 -6780
rect 11104 -6814 11172 -6780
rect 11172 -6814 11262 -6780
rect 11262 -6814 11330 -6780
rect 11330 -6814 11420 -6780
rect 11420 -6814 11488 -6780
rect 11488 -6814 11578 -6780
rect 11578 -6814 11646 -6780
rect 11646 -6814 11736 -6780
rect 11736 -6814 11804 -6780
rect 11804 -6814 11894 -6780
rect 11894 -6814 11962 -6780
rect 11962 -6814 12052 -6780
rect 12052 -6814 12120 -6780
rect 12120 -6814 12210 -6780
rect 12210 -6814 12278 -6780
rect 12278 -6814 12368 -6780
rect 12368 -6814 12436 -6780
rect 12436 -6814 12526 -6780
rect 12526 -6814 12586 -6780
rect 7952 -6874 12586 -6814
rect 12740 -6900 12810 -6764
rect 14030 -720 14100 -580
rect 14252 -670 18886 -610
rect 14252 -704 14312 -670
rect 14312 -704 14402 -670
rect 14402 -704 14470 -670
rect 14470 -704 14560 -670
rect 14560 -704 14628 -670
rect 14628 -704 14718 -670
rect 14718 -704 14786 -670
rect 14786 -704 14876 -670
rect 14876 -704 14944 -670
rect 14944 -704 15034 -670
rect 15034 -704 15102 -670
rect 15102 -704 15192 -670
rect 15192 -704 15260 -670
rect 15260 -704 15350 -670
rect 15350 -704 15418 -670
rect 15418 -704 15508 -670
rect 15508 -704 15576 -670
rect 15576 -704 15666 -670
rect 15666 -704 15734 -670
rect 15734 -704 15824 -670
rect 15824 -704 15892 -670
rect 15892 -704 15982 -670
rect 15982 -704 16050 -670
rect 16050 -704 16140 -670
rect 16140 -704 16208 -670
rect 16208 -704 16298 -670
rect 16298 -704 16366 -670
rect 16366 -704 16456 -670
rect 16456 -704 16524 -670
rect 16524 -704 16614 -670
rect 16614 -704 16682 -670
rect 16682 -704 16772 -670
rect 16772 -704 16840 -670
rect 16840 -704 16930 -670
rect 16930 -704 16998 -670
rect 16998 -704 17088 -670
rect 17088 -704 17156 -670
rect 17156 -704 17246 -670
rect 17246 -704 17314 -670
rect 17314 -704 17404 -670
rect 17404 -704 17472 -670
rect 17472 -704 17562 -670
rect 17562 -704 17630 -670
rect 17630 -704 17720 -670
rect 17720 -704 17788 -670
rect 17788 -704 17878 -670
rect 17878 -704 17946 -670
rect 17946 -704 18036 -670
rect 18036 -704 18104 -670
rect 18104 -704 18194 -670
rect 18194 -704 18262 -670
rect 18262 -704 18352 -670
rect 18352 -704 18420 -670
rect 18420 -704 18510 -670
rect 18510 -704 18578 -670
rect 18578 -704 18668 -670
rect 18668 -704 18736 -670
rect 18736 -704 18826 -670
rect 18826 -704 18886 -670
rect 14252 -710 18886 -704
rect 14030 -6764 14046 -720
rect 14046 -6764 14084 -720
rect 14084 -6764 14100 -720
rect 19040 -720 19110 -580
rect 14165 -6722 14182 -762
rect 14182 -6722 14216 -762
rect 14216 -6722 14231 -762
rect 14323 -6722 14340 -762
rect 14340 -6722 14374 -762
rect 14374 -6722 14389 -762
rect 14481 -6722 14498 -762
rect 14498 -6722 14532 -762
rect 14532 -6722 14547 -762
rect 14639 -6722 14656 -762
rect 14656 -6722 14690 -762
rect 14690 -6722 14705 -762
rect 14797 -6722 14814 -762
rect 14814 -6722 14848 -762
rect 14848 -6722 14863 -762
rect 14955 -6722 14972 -762
rect 14972 -6722 15006 -762
rect 15006 -6722 15021 -762
rect 15113 -6722 15130 -762
rect 15130 -6722 15164 -762
rect 15164 -6722 15179 -762
rect 15271 -6722 15288 -762
rect 15288 -6722 15322 -762
rect 15322 -6722 15337 -762
rect 15429 -6722 15446 -762
rect 15446 -6722 15480 -762
rect 15480 -6722 15495 -762
rect 15587 -6722 15604 -762
rect 15604 -6722 15638 -762
rect 15638 -6722 15653 -762
rect 15745 -6722 15762 -762
rect 15762 -6722 15796 -762
rect 15796 -6722 15811 -762
rect 15903 -6722 15920 -762
rect 15920 -6722 15954 -762
rect 15954 -6722 15969 -762
rect 16061 -6722 16078 -762
rect 16078 -6722 16112 -762
rect 16112 -6722 16127 -762
rect 16219 -6722 16236 -762
rect 16236 -6722 16270 -762
rect 16270 -6722 16285 -762
rect 16377 -6722 16394 -762
rect 16394 -6722 16428 -762
rect 16428 -6722 16443 -762
rect 16535 -6722 16552 -762
rect 16552 -6722 16586 -762
rect 16586 -6722 16601 -762
rect 16693 -6722 16710 -762
rect 16710 -6722 16744 -762
rect 16744 -6722 16759 -762
rect 16851 -6722 16868 -762
rect 16868 -6722 16902 -762
rect 16902 -6722 16917 -762
rect 17009 -6722 17026 -762
rect 17026 -6722 17060 -762
rect 17060 -6722 17075 -762
rect 17167 -6722 17184 -762
rect 17184 -6722 17218 -762
rect 17218 -6722 17233 -762
rect 17325 -6722 17342 -762
rect 17342 -6722 17376 -762
rect 17376 -6722 17391 -762
rect 17483 -6722 17500 -762
rect 17500 -6722 17534 -762
rect 17534 -6722 17549 -762
rect 17641 -6722 17658 -762
rect 17658 -6722 17692 -762
rect 17692 -6722 17707 -762
rect 17799 -6722 17816 -762
rect 17816 -6722 17850 -762
rect 17850 -6722 17865 -762
rect 17957 -6722 17974 -762
rect 17974 -6722 18008 -762
rect 18008 -6722 18023 -762
rect 18115 -6722 18132 -762
rect 18132 -6722 18166 -762
rect 18166 -6722 18181 -762
rect 18273 -6722 18290 -762
rect 18290 -6722 18324 -762
rect 18324 -6722 18339 -762
rect 18431 -6722 18448 -762
rect 18448 -6722 18482 -762
rect 18482 -6722 18497 -762
rect 18589 -6722 18606 -762
rect 18606 -6722 18640 -762
rect 18640 -6722 18655 -762
rect 18747 -6722 18764 -762
rect 18764 -6722 18798 -762
rect 18798 -6722 18813 -762
rect 18905 -6722 18922 -762
rect 18922 -6722 18956 -762
rect 18956 -6722 18971 -762
rect 14030 -6900 14100 -6764
rect 19040 -6764 19054 -720
rect 19054 -6764 19092 -720
rect 19092 -6764 19110 -720
rect 14252 -6780 18886 -6774
rect 14252 -6814 14312 -6780
rect 14312 -6814 14402 -6780
rect 14402 -6814 14470 -6780
rect 14470 -6814 14560 -6780
rect 14560 -6814 14628 -6780
rect 14628 -6814 14718 -6780
rect 14718 -6814 14786 -6780
rect 14786 -6814 14876 -6780
rect 14876 -6814 14944 -6780
rect 14944 -6814 15034 -6780
rect 15034 -6814 15102 -6780
rect 15102 -6814 15192 -6780
rect 15192 -6814 15260 -6780
rect 15260 -6814 15350 -6780
rect 15350 -6814 15418 -6780
rect 15418 -6814 15508 -6780
rect 15508 -6814 15576 -6780
rect 15576 -6814 15666 -6780
rect 15666 -6814 15734 -6780
rect 15734 -6814 15824 -6780
rect 15824 -6814 15892 -6780
rect 15892 -6814 15982 -6780
rect 15982 -6814 16050 -6780
rect 16050 -6814 16140 -6780
rect 16140 -6814 16208 -6780
rect 16208 -6814 16298 -6780
rect 16298 -6814 16366 -6780
rect 16366 -6814 16456 -6780
rect 16456 -6814 16524 -6780
rect 16524 -6814 16614 -6780
rect 16614 -6814 16682 -6780
rect 16682 -6814 16772 -6780
rect 16772 -6814 16840 -6780
rect 16840 -6814 16930 -6780
rect 16930 -6814 16998 -6780
rect 16998 -6814 17088 -6780
rect 17088 -6814 17156 -6780
rect 17156 -6814 17246 -6780
rect 17246 -6814 17314 -6780
rect 17314 -6814 17404 -6780
rect 17404 -6814 17472 -6780
rect 17472 -6814 17562 -6780
rect 17562 -6814 17630 -6780
rect 17630 -6814 17720 -6780
rect 17720 -6814 17788 -6780
rect 17788 -6814 17878 -6780
rect 17878 -6814 17946 -6780
rect 17946 -6814 18036 -6780
rect 18036 -6814 18104 -6780
rect 18104 -6814 18194 -6780
rect 18194 -6814 18262 -6780
rect 18262 -6814 18352 -6780
rect 18352 -6814 18420 -6780
rect 18420 -6814 18510 -6780
rect 18510 -6814 18578 -6780
rect 18578 -6814 18668 -6780
rect 18668 -6814 18736 -6780
rect 18736 -6814 18826 -6780
rect 18826 -6814 18886 -6780
rect 14252 -6874 18886 -6814
rect 19040 -6900 19110 -6764
rect 20330 -720 20400 -580
rect 20552 -670 25186 -610
rect 20552 -704 20612 -670
rect 20612 -704 20702 -670
rect 20702 -704 20770 -670
rect 20770 -704 20860 -670
rect 20860 -704 20928 -670
rect 20928 -704 21018 -670
rect 21018 -704 21086 -670
rect 21086 -704 21176 -670
rect 21176 -704 21244 -670
rect 21244 -704 21334 -670
rect 21334 -704 21402 -670
rect 21402 -704 21492 -670
rect 21492 -704 21560 -670
rect 21560 -704 21650 -670
rect 21650 -704 21718 -670
rect 21718 -704 21808 -670
rect 21808 -704 21876 -670
rect 21876 -704 21966 -670
rect 21966 -704 22034 -670
rect 22034 -704 22124 -670
rect 22124 -704 22192 -670
rect 22192 -704 22282 -670
rect 22282 -704 22350 -670
rect 22350 -704 22440 -670
rect 22440 -704 22508 -670
rect 22508 -704 22598 -670
rect 22598 -704 22666 -670
rect 22666 -704 22756 -670
rect 22756 -704 22824 -670
rect 22824 -704 22914 -670
rect 22914 -704 22982 -670
rect 22982 -704 23072 -670
rect 23072 -704 23140 -670
rect 23140 -704 23230 -670
rect 23230 -704 23298 -670
rect 23298 -704 23388 -670
rect 23388 -704 23456 -670
rect 23456 -704 23546 -670
rect 23546 -704 23614 -670
rect 23614 -704 23704 -670
rect 23704 -704 23772 -670
rect 23772 -704 23862 -670
rect 23862 -704 23930 -670
rect 23930 -704 24020 -670
rect 24020 -704 24088 -670
rect 24088 -704 24178 -670
rect 24178 -704 24246 -670
rect 24246 -704 24336 -670
rect 24336 -704 24404 -670
rect 24404 -704 24494 -670
rect 24494 -704 24562 -670
rect 24562 -704 24652 -670
rect 24652 -704 24720 -670
rect 24720 -704 24810 -670
rect 24810 -704 24878 -670
rect 24878 -704 24968 -670
rect 24968 -704 25036 -670
rect 25036 -704 25126 -670
rect 25126 -704 25186 -670
rect 20552 -710 25186 -704
rect 20330 -6764 20346 -720
rect 20346 -6764 20384 -720
rect 20384 -6764 20400 -720
rect 25340 -720 25410 -580
rect 20465 -6722 20482 -762
rect 20482 -6722 20516 -762
rect 20516 -6722 20531 -762
rect 20623 -6722 20640 -762
rect 20640 -6722 20674 -762
rect 20674 -6722 20689 -762
rect 20781 -6722 20798 -762
rect 20798 -6722 20832 -762
rect 20832 -6722 20847 -762
rect 20939 -6722 20956 -762
rect 20956 -6722 20990 -762
rect 20990 -6722 21005 -762
rect 21097 -6722 21114 -762
rect 21114 -6722 21148 -762
rect 21148 -6722 21163 -762
rect 21255 -6722 21272 -762
rect 21272 -6722 21306 -762
rect 21306 -6722 21321 -762
rect 21413 -6722 21430 -762
rect 21430 -6722 21464 -762
rect 21464 -6722 21479 -762
rect 21571 -6722 21588 -762
rect 21588 -6722 21622 -762
rect 21622 -6722 21637 -762
rect 21729 -6722 21746 -762
rect 21746 -6722 21780 -762
rect 21780 -6722 21795 -762
rect 21887 -6722 21904 -762
rect 21904 -6722 21938 -762
rect 21938 -6722 21953 -762
rect 22045 -6722 22062 -762
rect 22062 -6722 22096 -762
rect 22096 -6722 22111 -762
rect 22203 -6722 22220 -762
rect 22220 -6722 22254 -762
rect 22254 -6722 22269 -762
rect 22361 -6722 22378 -762
rect 22378 -6722 22412 -762
rect 22412 -6722 22427 -762
rect 22519 -6722 22536 -762
rect 22536 -6722 22570 -762
rect 22570 -6722 22585 -762
rect 22677 -6722 22694 -762
rect 22694 -6722 22728 -762
rect 22728 -6722 22743 -762
rect 22835 -6722 22852 -762
rect 22852 -6722 22886 -762
rect 22886 -6722 22901 -762
rect 22993 -6722 23010 -762
rect 23010 -6722 23044 -762
rect 23044 -6722 23059 -762
rect 23151 -6722 23168 -762
rect 23168 -6722 23202 -762
rect 23202 -6722 23217 -762
rect 23309 -6722 23326 -762
rect 23326 -6722 23360 -762
rect 23360 -6722 23375 -762
rect 23467 -6722 23484 -762
rect 23484 -6722 23518 -762
rect 23518 -6722 23533 -762
rect 23625 -6722 23642 -762
rect 23642 -6722 23676 -762
rect 23676 -6722 23691 -762
rect 23783 -6722 23800 -762
rect 23800 -6722 23834 -762
rect 23834 -6722 23849 -762
rect 23941 -6722 23958 -762
rect 23958 -6722 23992 -762
rect 23992 -6722 24007 -762
rect 24099 -6722 24116 -762
rect 24116 -6722 24150 -762
rect 24150 -6722 24165 -762
rect 24257 -6722 24274 -762
rect 24274 -6722 24308 -762
rect 24308 -6722 24323 -762
rect 24415 -6722 24432 -762
rect 24432 -6722 24466 -762
rect 24466 -6722 24481 -762
rect 24573 -6722 24590 -762
rect 24590 -6722 24624 -762
rect 24624 -6722 24639 -762
rect 24731 -6722 24748 -762
rect 24748 -6722 24782 -762
rect 24782 -6722 24797 -762
rect 24889 -6722 24906 -762
rect 24906 -6722 24940 -762
rect 24940 -6722 24955 -762
rect 25047 -6722 25064 -762
rect 25064 -6722 25098 -762
rect 25098 -6722 25113 -762
rect 25205 -6722 25222 -762
rect 25222 -6722 25256 -762
rect 25256 -6722 25271 -762
rect 20330 -6900 20400 -6764
rect 25340 -6764 25354 -720
rect 25354 -6764 25392 -720
rect 25392 -6764 25410 -720
rect 20552 -6780 25186 -6774
rect 20552 -6814 20612 -6780
rect 20612 -6814 20702 -6780
rect 20702 -6814 20770 -6780
rect 20770 -6814 20860 -6780
rect 20860 -6814 20928 -6780
rect 20928 -6814 21018 -6780
rect 21018 -6814 21086 -6780
rect 21086 -6814 21176 -6780
rect 21176 -6814 21244 -6780
rect 21244 -6814 21334 -6780
rect 21334 -6814 21402 -6780
rect 21402 -6814 21492 -6780
rect 21492 -6814 21560 -6780
rect 21560 -6814 21650 -6780
rect 21650 -6814 21718 -6780
rect 21718 -6814 21808 -6780
rect 21808 -6814 21876 -6780
rect 21876 -6814 21966 -6780
rect 21966 -6814 22034 -6780
rect 22034 -6814 22124 -6780
rect 22124 -6814 22192 -6780
rect 22192 -6814 22282 -6780
rect 22282 -6814 22350 -6780
rect 22350 -6814 22440 -6780
rect 22440 -6814 22508 -6780
rect 22508 -6814 22598 -6780
rect 22598 -6814 22666 -6780
rect 22666 -6814 22756 -6780
rect 22756 -6814 22824 -6780
rect 22824 -6814 22914 -6780
rect 22914 -6814 22982 -6780
rect 22982 -6814 23072 -6780
rect 23072 -6814 23140 -6780
rect 23140 -6814 23230 -6780
rect 23230 -6814 23298 -6780
rect 23298 -6814 23388 -6780
rect 23388 -6814 23456 -6780
rect 23456 -6814 23546 -6780
rect 23546 -6814 23614 -6780
rect 23614 -6814 23704 -6780
rect 23704 -6814 23772 -6780
rect 23772 -6814 23862 -6780
rect 23862 -6814 23930 -6780
rect 23930 -6814 24020 -6780
rect 24020 -6814 24088 -6780
rect 24088 -6814 24178 -6780
rect 24178 -6814 24246 -6780
rect 24246 -6814 24336 -6780
rect 24336 -6814 24404 -6780
rect 24404 -6814 24494 -6780
rect 24494 -6814 24562 -6780
rect 24562 -6814 24652 -6780
rect 24652 -6814 24720 -6780
rect 24720 -6814 24810 -6780
rect 24810 -6814 24878 -6780
rect 24878 -6814 24968 -6780
rect 24968 -6814 25036 -6780
rect 25036 -6814 25126 -6780
rect 25126 -6814 25186 -6780
rect 20552 -6874 25186 -6814
rect 25340 -6900 25410 -6764
<< metal2 >>
rect 6500 6480 7800 6500
rect 12800 6480 14100 6600
rect 19100 6480 20400 6500
rect 1430 6420 1500 6480
rect 6440 6420 7800 6480
rect 1632 6380 1652 6390
rect 6286 6380 6306 6390
rect 1632 6310 1640 6380
rect 6300 6310 6306 6380
rect 1632 6290 1652 6310
rect 6286 6290 6306 6310
rect 1565 6238 1631 6258
rect 1565 258 1631 278
rect 1723 6238 1789 6258
rect 1723 258 1789 278
rect 1881 6238 1947 6258
rect 1881 258 1947 278
rect 2039 6238 2105 6258
rect 2039 258 2105 278
rect 2197 6238 2263 6258
rect 2197 258 2263 278
rect 2355 6238 2421 6258
rect 2355 258 2421 278
rect 2513 6238 2579 6258
rect 2513 258 2579 278
rect 2671 6238 2737 6258
rect 2671 258 2737 278
rect 2829 6238 2895 6258
rect 2829 258 2895 278
rect 2987 6238 3053 6258
rect 2987 258 3053 278
rect 3145 6238 3211 6258
rect 3145 258 3211 278
rect 3303 6238 3369 6258
rect 3303 258 3369 278
rect 3461 6238 3527 6258
rect 3461 258 3527 278
rect 3619 6238 3685 6258
rect 3619 258 3685 278
rect 3777 6238 3843 6258
rect 3777 258 3843 278
rect 3935 6238 4001 6258
rect 3935 258 4001 278
rect 4093 6238 4159 6258
rect 4093 258 4159 278
rect 4251 6238 4317 6258
rect 4251 258 4317 278
rect 4409 6238 4475 6258
rect 4409 258 4475 278
rect 4567 6238 4633 6258
rect 4567 258 4633 278
rect 4725 6238 4791 6258
rect 4725 258 4791 278
rect 4883 6238 4949 6258
rect 4883 258 4949 278
rect 5041 6238 5107 6258
rect 5041 258 5107 278
rect 5199 6238 5265 6258
rect 5199 258 5265 278
rect 5357 6238 5423 6258
rect 5357 258 5423 278
rect 5515 6238 5581 6258
rect 5515 258 5581 278
rect 5673 6238 5739 6258
rect 5673 258 5739 278
rect 5831 6238 5897 6258
rect 5831 258 5897 278
rect 5989 6238 6055 6258
rect 5989 258 6055 278
rect 6147 6238 6213 6258
rect 6147 258 6213 278
rect 6305 6238 6371 6258
rect 6305 258 6371 278
rect 1632 210 1652 226
rect 6286 210 6306 226
rect 1632 140 1640 210
rect 6290 140 6306 210
rect 1632 126 1652 140
rect 6286 126 6306 140
rect 1430 30 1500 100
rect 6510 6100 7730 6420
rect 6510 5500 7730 5900
rect 6510 4900 7730 5300
rect 6510 4300 7730 4700
rect 6510 3700 7730 4100
rect 6510 3100 7730 3500
rect 6510 2500 7730 2900
rect 6510 1900 7730 2300
rect 6510 1300 7730 1700
rect 6510 700 7730 1100
rect 6510 100 7730 500
rect 12740 6420 14100 6480
rect 7932 6380 7952 6390
rect 12586 6380 12606 6390
rect 7932 6310 7940 6380
rect 12600 6310 12606 6380
rect 7932 6290 7952 6310
rect 12586 6290 12606 6310
rect 7865 6238 7931 6258
rect 7865 258 7931 278
rect 8023 6238 8089 6258
rect 8023 258 8089 278
rect 8181 6238 8247 6258
rect 8181 258 8247 278
rect 8339 6238 8405 6258
rect 8339 258 8405 278
rect 8497 6238 8563 6258
rect 8497 258 8563 278
rect 8655 6238 8721 6258
rect 8655 258 8721 278
rect 8813 6238 8879 6258
rect 8813 258 8879 278
rect 8971 6238 9037 6258
rect 8971 258 9037 278
rect 9129 6238 9195 6258
rect 9129 258 9195 278
rect 9287 6238 9353 6258
rect 9287 258 9353 278
rect 9445 6238 9511 6258
rect 9445 258 9511 278
rect 9603 6238 9669 6258
rect 9603 258 9669 278
rect 9761 6238 9827 6258
rect 9761 258 9827 278
rect 9919 6238 9985 6258
rect 9919 258 9985 278
rect 10077 6238 10143 6258
rect 10077 258 10143 278
rect 10235 6238 10301 6258
rect 10235 258 10301 278
rect 10393 6238 10459 6258
rect 10393 258 10459 278
rect 10551 6238 10617 6258
rect 10551 258 10617 278
rect 10709 6238 10775 6258
rect 10709 258 10775 278
rect 10867 6238 10933 6258
rect 10867 258 10933 278
rect 11025 6238 11091 6258
rect 11025 258 11091 278
rect 11183 6238 11249 6258
rect 11183 258 11249 278
rect 11341 6238 11407 6258
rect 11341 258 11407 278
rect 11499 6238 11565 6258
rect 11499 258 11565 278
rect 11657 6238 11723 6258
rect 11657 258 11723 278
rect 11815 6238 11881 6258
rect 11815 258 11881 278
rect 11973 6238 12039 6258
rect 11973 258 12039 278
rect 12131 6238 12197 6258
rect 12131 258 12197 278
rect 12289 6238 12355 6258
rect 12289 258 12355 278
rect 12447 6238 12513 6258
rect 12447 258 12513 278
rect 12605 6238 12671 6258
rect 12605 258 12671 278
rect 7932 210 7952 226
rect 12586 210 12606 226
rect 7932 140 7940 210
rect 12590 140 12606 210
rect 7932 126 7952 140
rect 12586 126 12606 140
rect 6440 30 6510 100
rect 6900 -500 7400 100
rect 7730 30 7800 100
rect 12810 6200 14030 6420
rect 12810 5600 14030 6000
rect 12810 5000 14030 5400
rect 12810 4400 14030 4800
rect 12810 3800 14030 4200
rect 12810 3200 14030 3600
rect 12810 2600 14030 3000
rect 12810 2000 14030 2400
rect 12810 1400 14030 1800
rect 12810 800 14030 1200
rect 12810 200 14030 600
rect 12740 30 12810 100
rect 13200 -500 13700 200
rect 19040 6420 20400 6480
rect 14232 6380 14252 6390
rect 18886 6380 18906 6390
rect 14232 6310 14240 6380
rect 18900 6310 18906 6380
rect 14232 6290 14252 6310
rect 18886 6290 18906 6310
rect 14165 6238 14231 6258
rect 14165 258 14231 278
rect 14323 6238 14389 6258
rect 14323 258 14389 278
rect 14481 6238 14547 6258
rect 14481 258 14547 278
rect 14639 6238 14705 6258
rect 14639 258 14705 278
rect 14797 6238 14863 6258
rect 14797 258 14863 278
rect 14955 6238 15021 6258
rect 14955 258 15021 278
rect 15113 6238 15179 6258
rect 15113 258 15179 278
rect 15271 6238 15337 6258
rect 15271 258 15337 278
rect 15429 6238 15495 6258
rect 15429 258 15495 278
rect 15587 6238 15653 6258
rect 15587 258 15653 278
rect 15745 6238 15811 6258
rect 15745 258 15811 278
rect 15903 6238 15969 6258
rect 15903 258 15969 278
rect 16061 6238 16127 6258
rect 16061 258 16127 278
rect 16219 6238 16285 6258
rect 16219 258 16285 278
rect 16377 6238 16443 6258
rect 16377 258 16443 278
rect 16535 6238 16601 6258
rect 16535 258 16601 278
rect 16693 6238 16759 6258
rect 16693 258 16759 278
rect 16851 6238 16917 6258
rect 16851 258 16917 278
rect 17009 6238 17075 6258
rect 17009 258 17075 278
rect 17167 6238 17233 6258
rect 17167 258 17233 278
rect 17325 6238 17391 6258
rect 17325 258 17391 278
rect 17483 6238 17549 6258
rect 17483 258 17549 278
rect 17641 6238 17707 6258
rect 17641 258 17707 278
rect 17799 6238 17865 6258
rect 17799 258 17865 278
rect 17957 6238 18023 6258
rect 17957 258 18023 278
rect 18115 6238 18181 6258
rect 18115 258 18181 278
rect 18273 6238 18339 6258
rect 18273 258 18339 278
rect 18431 6238 18497 6258
rect 18431 258 18497 278
rect 18589 6238 18655 6258
rect 18589 258 18655 278
rect 18747 6238 18813 6258
rect 18747 258 18813 278
rect 18905 6238 18971 6258
rect 18905 258 18971 278
rect 14232 210 14252 226
rect 18886 210 18906 226
rect 14232 140 14240 210
rect 18890 140 18906 210
rect 14232 126 14252 140
rect 18886 126 18906 140
rect 14030 30 14100 100
rect 19110 6100 20330 6420
rect 19110 5500 20330 5900
rect 19110 4900 20330 5300
rect 19110 4300 20330 4700
rect 19110 3700 20330 4100
rect 19110 3100 20330 3500
rect 19110 2500 20330 2900
rect 19110 1900 20330 2300
rect 19110 1300 20330 1700
rect 19110 700 20330 1100
rect 19110 100 20330 500
rect 25340 6420 25410 6480
rect 20532 6380 20552 6390
rect 25186 6380 25206 6390
rect 20532 6310 20540 6380
rect 25200 6310 25206 6380
rect 20532 6290 20552 6310
rect 25186 6290 25206 6310
rect 20465 6238 20531 6258
rect 20465 258 20531 278
rect 20623 6238 20689 6258
rect 20623 258 20689 278
rect 20781 6238 20847 6258
rect 20781 258 20847 278
rect 20939 6238 21005 6258
rect 20939 258 21005 278
rect 21097 6238 21163 6258
rect 21097 258 21163 278
rect 21255 6238 21321 6258
rect 21255 258 21321 278
rect 21413 6238 21479 6258
rect 21413 258 21479 278
rect 21571 6238 21637 6258
rect 21571 258 21637 278
rect 21729 6238 21795 6258
rect 21729 258 21795 278
rect 21887 6238 21953 6258
rect 21887 258 21953 278
rect 22045 6238 22111 6258
rect 22045 258 22111 278
rect 22203 6238 22269 6258
rect 22203 258 22269 278
rect 22361 6238 22427 6258
rect 22361 258 22427 278
rect 22519 6238 22585 6258
rect 22519 258 22585 278
rect 22677 6238 22743 6258
rect 22677 258 22743 278
rect 22835 6238 22901 6258
rect 22835 258 22901 278
rect 22993 6238 23059 6258
rect 22993 258 23059 278
rect 23151 6238 23217 6258
rect 23151 258 23217 278
rect 23309 6238 23375 6258
rect 23309 258 23375 278
rect 23467 6238 23533 6258
rect 23467 258 23533 278
rect 23625 6238 23691 6258
rect 23625 258 23691 278
rect 23783 6238 23849 6258
rect 23783 258 23849 278
rect 23941 6238 24007 6258
rect 23941 258 24007 278
rect 24099 6238 24165 6258
rect 24099 258 24165 278
rect 24257 6238 24323 6258
rect 24257 258 24323 278
rect 24415 6238 24481 6258
rect 24415 258 24481 278
rect 24573 6238 24639 6258
rect 24573 258 24639 278
rect 24731 6238 24797 6258
rect 24731 258 24797 278
rect 24889 6238 24955 6258
rect 24889 258 24955 278
rect 25047 6238 25113 6258
rect 25047 258 25113 278
rect 25205 6238 25271 6258
rect 25205 258 25271 278
rect 20532 210 20552 226
rect 25186 210 25206 226
rect 20532 140 20540 210
rect 25190 140 25206 210
rect 20532 126 20552 140
rect 25186 126 25206 140
rect 19040 30 19110 100
rect 19500 -500 20000 100
rect 20330 30 20400 100
rect 25340 30 25410 100
rect 6500 -520 7800 -500
rect 12800 -520 14100 -500
rect 19100 -520 20400 -500
rect 1430 -580 1500 -520
rect 6440 -580 7800 -520
rect 1632 -620 1652 -610
rect 6286 -620 6306 -610
rect 1632 -690 1640 -620
rect 6300 -690 6306 -620
rect 1632 -710 1652 -690
rect 6286 -710 6306 -690
rect 1565 -762 1631 -742
rect 1565 -6742 1631 -6722
rect 1723 -762 1789 -742
rect 1723 -6742 1789 -6722
rect 1881 -762 1947 -742
rect 1881 -6742 1947 -6722
rect 2039 -762 2105 -742
rect 2039 -6742 2105 -6722
rect 2197 -762 2263 -742
rect 2197 -6742 2263 -6722
rect 2355 -762 2421 -742
rect 2355 -6742 2421 -6722
rect 2513 -762 2579 -742
rect 2513 -6742 2579 -6722
rect 2671 -762 2737 -742
rect 2671 -6742 2737 -6722
rect 2829 -762 2895 -742
rect 2829 -6742 2895 -6722
rect 2987 -762 3053 -742
rect 2987 -6742 3053 -6722
rect 3145 -762 3211 -742
rect 3145 -6742 3211 -6722
rect 3303 -762 3369 -742
rect 3303 -6742 3369 -6722
rect 3461 -762 3527 -742
rect 3461 -6742 3527 -6722
rect 3619 -762 3685 -742
rect 3619 -6742 3685 -6722
rect 3777 -762 3843 -742
rect 3777 -6742 3843 -6722
rect 3935 -762 4001 -742
rect 3935 -6742 4001 -6722
rect 4093 -762 4159 -742
rect 4093 -6742 4159 -6722
rect 4251 -762 4317 -742
rect 4251 -6742 4317 -6722
rect 4409 -762 4475 -742
rect 4409 -6742 4475 -6722
rect 4567 -762 4633 -742
rect 4567 -6742 4633 -6722
rect 4725 -762 4791 -742
rect 4725 -6742 4791 -6722
rect 4883 -762 4949 -742
rect 4883 -6742 4949 -6722
rect 5041 -762 5107 -742
rect 5041 -6742 5107 -6722
rect 5199 -762 5265 -742
rect 5199 -6742 5265 -6722
rect 5357 -762 5423 -742
rect 5357 -6742 5423 -6722
rect 5515 -762 5581 -742
rect 5515 -6742 5581 -6722
rect 5673 -762 5739 -742
rect 5673 -6742 5739 -6722
rect 5831 -762 5897 -742
rect 5831 -6742 5897 -6722
rect 5989 -762 6055 -742
rect 5989 -6742 6055 -6722
rect 6147 -762 6213 -742
rect 6147 -6742 6213 -6722
rect 6305 -762 6371 -742
rect 6305 -6742 6371 -6722
rect 1632 -6790 1652 -6774
rect 6286 -6790 6306 -6774
rect 1632 -6860 1640 -6790
rect 6290 -6860 6306 -6790
rect 1632 -6874 1652 -6860
rect 6286 -6874 6306 -6860
rect 1430 -6970 1500 -6900
rect 6510 -900 7730 -580
rect 6510 -1500 7730 -1100
rect 6510 -2100 7730 -1700
rect 6510 -2700 7730 -2300
rect 6510 -3300 7730 -2900
rect 6510 -3900 7730 -3500
rect 6510 -4500 7730 -4100
rect 6510 -5100 7730 -4700
rect 6510 -5700 7730 -5300
rect 6510 -6300 7730 -5900
rect 6510 -6900 7730 -6500
rect 12740 -580 14100 -520
rect 7932 -620 7952 -610
rect 12586 -620 12606 -610
rect 7932 -690 7940 -620
rect 12600 -690 12606 -620
rect 7932 -710 7952 -690
rect 12586 -710 12606 -690
rect 7865 -762 7931 -742
rect 7865 -6742 7931 -6722
rect 8023 -762 8089 -742
rect 8023 -6742 8089 -6722
rect 8181 -762 8247 -742
rect 8181 -6742 8247 -6722
rect 8339 -762 8405 -742
rect 8339 -6742 8405 -6722
rect 8497 -762 8563 -742
rect 8497 -6742 8563 -6722
rect 8655 -762 8721 -742
rect 8655 -6742 8721 -6722
rect 8813 -762 8879 -742
rect 8813 -6742 8879 -6722
rect 8971 -762 9037 -742
rect 8971 -6742 9037 -6722
rect 9129 -762 9195 -742
rect 9129 -6742 9195 -6722
rect 9287 -762 9353 -742
rect 9287 -6742 9353 -6722
rect 9445 -762 9511 -742
rect 9445 -6742 9511 -6722
rect 9603 -762 9669 -742
rect 9603 -6742 9669 -6722
rect 9761 -762 9827 -742
rect 9761 -6742 9827 -6722
rect 9919 -762 9985 -742
rect 9919 -6742 9985 -6722
rect 10077 -762 10143 -742
rect 10077 -6742 10143 -6722
rect 10235 -762 10301 -742
rect 10235 -6742 10301 -6722
rect 10393 -762 10459 -742
rect 10393 -6742 10459 -6722
rect 10551 -762 10617 -742
rect 10551 -6742 10617 -6722
rect 10709 -762 10775 -742
rect 10709 -6742 10775 -6722
rect 10867 -762 10933 -742
rect 10867 -6742 10933 -6722
rect 11025 -762 11091 -742
rect 11025 -6742 11091 -6722
rect 11183 -762 11249 -742
rect 11183 -6742 11249 -6722
rect 11341 -762 11407 -742
rect 11341 -6742 11407 -6722
rect 11499 -762 11565 -742
rect 11499 -6742 11565 -6722
rect 11657 -762 11723 -742
rect 11657 -6742 11723 -6722
rect 11815 -762 11881 -742
rect 11815 -6742 11881 -6722
rect 11973 -762 12039 -742
rect 11973 -6742 12039 -6722
rect 12131 -762 12197 -742
rect 12131 -6742 12197 -6722
rect 12289 -762 12355 -742
rect 12289 -6742 12355 -6722
rect 12447 -762 12513 -742
rect 12447 -6742 12513 -6722
rect 12605 -762 12671 -742
rect 12605 -6742 12671 -6722
rect 7932 -6790 7952 -6774
rect 12586 -6790 12606 -6774
rect 7932 -6860 7940 -6790
rect 12590 -6860 12606 -6790
rect 7932 -6874 7952 -6860
rect 12586 -6874 12606 -6860
rect 6440 -6970 6510 -6900
rect 7730 -6970 7800 -6900
rect 12810 -900 14030 -580
rect 12810 -1500 14030 -1100
rect 12810 -2100 14030 -1700
rect 12810 -2700 14030 -2300
rect 12810 -3300 14030 -2900
rect 12810 -3900 14030 -3500
rect 12810 -4500 14030 -4100
rect 12810 -5100 14030 -4700
rect 12810 -5700 14030 -5300
rect 12810 -6300 14030 -5900
rect 12810 -6900 14030 -6500
rect 19040 -580 20400 -520
rect 14232 -620 14252 -610
rect 18886 -620 18906 -610
rect 14232 -690 14240 -620
rect 18900 -690 18906 -620
rect 14232 -710 14252 -690
rect 18886 -710 18906 -690
rect 14165 -762 14231 -742
rect 14165 -6742 14231 -6722
rect 14323 -762 14389 -742
rect 14323 -6742 14389 -6722
rect 14481 -762 14547 -742
rect 14481 -6742 14547 -6722
rect 14639 -762 14705 -742
rect 14639 -6742 14705 -6722
rect 14797 -762 14863 -742
rect 14797 -6742 14863 -6722
rect 14955 -762 15021 -742
rect 14955 -6742 15021 -6722
rect 15113 -762 15179 -742
rect 15113 -6742 15179 -6722
rect 15271 -762 15337 -742
rect 15271 -6742 15337 -6722
rect 15429 -762 15495 -742
rect 15429 -6742 15495 -6722
rect 15587 -762 15653 -742
rect 15587 -6742 15653 -6722
rect 15745 -762 15811 -742
rect 15745 -6742 15811 -6722
rect 15903 -762 15969 -742
rect 15903 -6742 15969 -6722
rect 16061 -762 16127 -742
rect 16061 -6742 16127 -6722
rect 16219 -762 16285 -742
rect 16219 -6742 16285 -6722
rect 16377 -762 16443 -742
rect 16377 -6742 16443 -6722
rect 16535 -762 16601 -742
rect 16535 -6742 16601 -6722
rect 16693 -762 16759 -742
rect 16693 -6742 16759 -6722
rect 16851 -762 16917 -742
rect 16851 -6742 16917 -6722
rect 17009 -762 17075 -742
rect 17009 -6742 17075 -6722
rect 17167 -762 17233 -742
rect 17167 -6742 17233 -6722
rect 17325 -762 17391 -742
rect 17325 -6742 17391 -6722
rect 17483 -762 17549 -742
rect 17483 -6742 17549 -6722
rect 17641 -762 17707 -742
rect 17641 -6742 17707 -6722
rect 17799 -762 17865 -742
rect 17799 -6742 17865 -6722
rect 17957 -762 18023 -742
rect 17957 -6742 18023 -6722
rect 18115 -762 18181 -742
rect 18115 -6742 18181 -6722
rect 18273 -762 18339 -742
rect 18273 -6742 18339 -6722
rect 18431 -762 18497 -742
rect 18431 -6742 18497 -6722
rect 18589 -762 18655 -742
rect 18589 -6742 18655 -6722
rect 18747 -762 18813 -742
rect 18747 -6742 18813 -6722
rect 18905 -762 18971 -742
rect 18905 -6742 18971 -6722
rect 14232 -6790 14252 -6774
rect 18886 -6790 18906 -6774
rect 14232 -6860 14240 -6790
rect 18890 -6860 18906 -6790
rect 14232 -6874 14252 -6860
rect 18886 -6874 18906 -6860
rect 12740 -6970 12810 -6900
rect 14030 -6970 14100 -6900
rect 19110 -900 20330 -580
rect 19110 -1500 20330 -1100
rect 19110 -2100 20330 -1700
rect 19110 -2700 20330 -2300
rect 19110 -3300 20330 -2900
rect 19110 -3900 20330 -3500
rect 19110 -4500 20330 -4100
rect 19110 -5100 20330 -4700
rect 19110 -5700 20330 -5300
rect 19110 -6300 20330 -5900
rect 19110 -6900 20330 -6500
rect 25340 -580 25410 -520
rect 20532 -620 20552 -610
rect 25186 -620 25206 -610
rect 20532 -690 20540 -620
rect 25200 -690 25206 -620
rect 20532 -710 20552 -690
rect 25186 -710 25206 -690
rect 20465 -762 20531 -742
rect 20465 -6742 20531 -6722
rect 20623 -762 20689 -742
rect 20623 -6742 20689 -6722
rect 20781 -762 20847 -742
rect 20781 -6742 20847 -6722
rect 20939 -762 21005 -742
rect 20939 -6742 21005 -6722
rect 21097 -762 21163 -742
rect 21097 -6742 21163 -6722
rect 21255 -762 21321 -742
rect 21255 -6742 21321 -6722
rect 21413 -762 21479 -742
rect 21413 -6742 21479 -6722
rect 21571 -762 21637 -742
rect 21571 -6742 21637 -6722
rect 21729 -762 21795 -742
rect 21729 -6742 21795 -6722
rect 21887 -762 21953 -742
rect 21887 -6742 21953 -6722
rect 22045 -762 22111 -742
rect 22045 -6742 22111 -6722
rect 22203 -762 22269 -742
rect 22203 -6742 22269 -6722
rect 22361 -762 22427 -742
rect 22361 -6742 22427 -6722
rect 22519 -762 22585 -742
rect 22519 -6742 22585 -6722
rect 22677 -762 22743 -742
rect 22677 -6742 22743 -6722
rect 22835 -762 22901 -742
rect 22835 -6742 22901 -6722
rect 22993 -762 23059 -742
rect 22993 -6742 23059 -6722
rect 23151 -762 23217 -742
rect 23151 -6742 23217 -6722
rect 23309 -762 23375 -742
rect 23309 -6742 23375 -6722
rect 23467 -762 23533 -742
rect 23467 -6742 23533 -6722
rect 23625 -762 23691 -742
rect 23625 -6742 23691 -6722
rect 23783 -762 23849 -742
rect 23783 -6742 23849 -6722
rect 23941 -762 24007 -742
rect 23941 -6742 24007 -6722
rect 24099 -762 24165 -742
rect 24099 -6742 24165 -6722
rect 24257 -762 24323 -742
rect 24257 -6742 24323 -6722
rect 24415 -762 24481 -742
rect 24415 -6742 24481 -6722
rect 24573 -762 24639 -742
rect 24573 -6742 24639 -6722
rect 24731 -762 24797 -742
rect 24731 -6742 24797 -6722
rect 24889 -762 24955 -742
rect 24889 -6742 24955 -6722
rect 25047 -762 25113 -742
rect 25047 -6742 25113 -6722
rect 25205 -762 25271 -742
rect 25205 -6742 25271 -6722
rect 20532 -6790 20552 -6774
rect 25186 -6790 25206 -6774
rect 20532 -6860 20540 -6790
rect 25190 -6860 25206 -6790
rect 20532 -6874 20552 -6860
rect 25186 -6874 25206 -6860
rect 19040 -6970 19110 -6900
rect 20330 -6970 20400 -6900
rect 25340 -6970 25410 -6900
<< via2 >>
rect 1640 6310 1652 6380
rect 1652 6310 6286 6380
rect 6286 6310 6300 6380
rect 1565 885 1631 2645
rect 1723 3885 1789 5645
rect 1881 885 1947 2645
rect 2039 3885 2105 5645
rect 2197 885 2263 2645
rect 2355 3885 2421 5645
rect 2513 885 2579 2645
rect 2671 3885 2737 5645
rect 2829 885 2895 2645
rect 2987 3885 3053 5645
rect 3145 885 3211 2645
rect 3303 3885 3369 5645
rect 3461 885 3527 2645
rect 3619 3885 3685 5645
rect 3777 885 3843 2645
rect 3935 3885 4001 5645
rect 4093 885 4159 2645
rect 4251 3885 4317 5645
rect 4409 885 4475 2645
rect 4567 3885 4633 5645
rect 4725 885 4791 2645
rect 4883 3885 4949 5645
rect 5041 885 5107 2645
rect 5199 3885 5265 5645
rect 5357 885 5423 2645
rect 5515 3885 5581 5645
rect 5673 885 5739 2645
rect 5831 3885 5897 5645
rect 5989 885 6055 2645
rect 6147 3885 6213 5645
rect 6305 885 6371 2645
rect 1640 140 1652 210
rect 1652 140 6286 210
rect 6286 140 6290 210
rect 7940 6310 7952 6380
rect 7952 6310 12586 6380
rect 12586 6310 12600 6380
rect 7865 885 7931 2645
rect 8023 3885 8089 5645
rect 8181 885 8247 2645
rect 8339 3885 8405 5645
rect 8497 885 8563 2645
rect 8655 3885 8721 5645
rect 8813 885 8879 2645
rect 8971 3885 9037 5645
rect 9129 885 9195 2645
rect 9287 3885 9353 5645
rect 9445 885 9511 2645
rect 9603 3885 9669 5645
rect 9761 885 9827 2645
rect 9919 3885 9985 5645
rect 10077 885 10143 2645
rect 10235 3885 10301 5645
rect 10393 885 10459 2645
rect 10551 3885 10617 5645
rect 10709 885 10775 2645
rect 10867 3885 10933 5645
rect 11025 885 11091 2645
rect 11183 3885 11249 5645
rect 11341 885 11407 2645
rect 11499 3885 11565 5645
rect 11657 885 11723 2645
rect 11815 3885 11881 5645
rect 11973 885 12039 2645
rect 12131 3885 12197 5645
rect 12289 885 12355 2645
rect 12447 3885 12513 5645
rect 12605 885 12671 2645
rect 7940 140 7952 210
rect 7952 140 12586 210
rect 12586 140 12590 210
rect 14240 6310 14252 6380
rect 14252 6310 18886 6380
rect 18886 6310 18900 6380
rect 14165 885 14231 2645
rect 14323 3885 14389 5645
rect 14481 885 14547 2645
rect 14639 3885 14705 5645
rect 14797 885 14863 2645
rect 14955 3885 15021 5645
rect 15113 885 15179 2645
rect 15271 3885 15337 5645
rect 15429 885 15495 2645
rect 15587 3885 15653 5645
rect 15745 885 15811 2645
rect 15903 3885 15969 5645
rect 16061 885 16127 2645
rect 16219 3885 16285 5645
rect 16377 885 16443 2645
rect 16535 3885 16601 5645
rect 16693 885 16759 2645
rect 16851 3885 16917 5645
rect 17009 885 17075 2645
rect 17167 3885 17233 5645
rect 17325 885 17391 2645
rect 17483 3885 17549 5645
rect 17641 885 17707 2645
rect 17799 3885 17865 5645
rect 17957 885 18023 2645
rect 18115 3885 18181 5645
rect 18273 885 18339 2645
rect 18431 3885 18497 5645
rect 18589 885 18655 2645
rect 18747 3885 18813 5645
rect 18905 885 18971 2645
rect 14240 140 14252 210
rect 14252 140 18886 210
rect 18886 140 18890 210
rect 20540 6310 20552 6380
rect 20552 6310 25186 6380
rect 25186 6310 25200 6380
rect 20465 885 20531 2645
rect 20623 3885 20689 5645
rect 20781 885 20847 2645
rect 20939 3885 21005 5645
rect 21097 885 21163 2645
rect 21255 3885 21321 5645
rect 21413 885 21479 2645
rect 21571 3885 21637 5645
rect 21729 885 21795 2645
rect 21887 3885 21953 5645
rect 22045 885 22111 2645
rect 22203 3885 22269 5645
rect 22361 885 22427 2645
rect 22519 3885 22585 5645
rect 22677 885 22743 2645
rect 22835 3885 22901 5645
rect 22993 885 23059 2645
rect 23151 3885 23217 5645
rect 23309 885 23375 2645
rect 23467 3885 23533 5645
rect 23625 885 23691 2645
rect 23783 3885 23849 5645
rect 23941 885 24007 2645
rect 24099 3885 24165 5645
rect 24257 885 24323 2645
rect 24415 3885 24481 5645
rect 24573 885 24639 2645
rect 24731 3885 24797 5645
rect 24889 885 24955 2645
rect 25047 3885 25113 5645
rect 25205 885 25271 2645
rect 20540 140 20552 210
rect 20552 140 25186 210
rect 25186 140 25190 210
rect 1640 -690 1652 -620
rect 1652 -690 6286 -620
rect 6286 -690 6300 -620
rect 1565 -6115 1631 -4355
rect 1723 -3115 1789 -1355
rect 1881 -6115 1947 -4355
rect 2039 -3115 2105 -1355
rect 2197 -6115 2263 -4355
rect 2355 -3115 2421 -1355
rect 2513 -6115 2579 -4355
rect 2671 -3115 2737 -1355
rect 2829 -6115 2895 -4355
rect 2987 -3115 3053 -1355
rect 3145 -6115 3211 -4355
rect 3303 -3115 3369 -1355
rect 3461 -6115 3527 -4355
rect 3619 -3115 3685 -1355
rect 3777 -6115 3843 -4355
rect 3935 -3115 4001 -1355
rect 4093 -6115 4159 -4355
rect 4251 -3115 4317 -1355
rect 4409 -6115 4475 -4355
rect 4567 -3115 4633 -1355
rect 4725 -6115 4791 -4355
rect 4883 -3115 4949 -1355
rect 5041 -6115 5107 -4355
rect 5199 -3115 5265 -1355
rect 5357 -6115 5423 -4355
rect 5515 -3115 5581 -1355
rect 5673 -6115 5739 -4355
rect 5831 -3115 5897 -1355
rect 5989 -6115 6055 -4355
rect 6147 -3115 6213 -1355
rect 6305 -6115 6371 -4355
rect 1640 -6860 1652 -6790
rect 1652 -6860 6286 -6790
rect 6286 -6860 6290 -6790
rect 7940 -690 7952 -620
rect 7952 -690 12586 -620
rect 12586 -690 12600 -620
rect 7865 -6115 7931 -4355
rect 8023 -3115 8089 -1355
rect 8181 -6115 8247 -4355
rect 8339 -3115 8405 -1355
rect 8497 -6115 8563 -4355
rect 8655 -3115 8721 -1355
rect 8813 -6115 8879 -4355
rect 8971 -3115 9037 -1355
rect 9129 -6115 9195 -4355
rect 9287 -3115 9353 -1355
rect 9445 -6115 9511 -4355
rect 9603 -3115 9669 -1355
rect 9761 -6115 9827 -4355
rect 9919 -3115 9985 -1355
rect 10077 -6115 10143 -4355
rect 10235 -3115 10301 -1355
rect 10393 -6115 10459 -4355
rect 10551 -3115 10617 -1355
rect 10709 -6115 10775 -4355
rect 10867 -3115 10933 -1355
rect 11025 -6115 11091 -4355
rect 11183 -3115 11249 -1355
rect 11341 -6115 11407 -4355
rect 11499 -3115 11565 -1355
rect 11657 -6115 11723 -4355
rect 11815 -3115 11881 -1355
rect 11973 -6115 12039 -4355
rect 12131 -3115 12197 -1355
rect 12289 -6115 12355 -4355
rect 12447 -3115 12513 -1355
rect 12605 -6115 12671 -4355
rect 7940 -6860 7952 -6790
rect 7952 -6860 12586 -6790
rect 12586 -6860 12590 -6790
rect 14240 -690 14252 -620
rect 14252 -690 18886 -620
rect 18886 -690 18900 -620
rect 14165 -6115 14231 -4355
rect 14323 -3115 14389 -1355
rect 14481 -6115 14547 -4355
rect 14639 -3115 14705 -1355
rect 14797 -6115 14863 -4355
rect 14955 -3115 15021 -1355
rect 15113 -6115 15179 -4355
rect 15271 -3115 15337 -1355
rect 15429 -6115 15495 -4355
rect 15587 -3115 15653 -1355
rect 15745 -6115 15811 -4355
rect 15903 -3115 15969 -1355
rect 16061 -6115 16127 -4355
rect 16219 -3115 16285 -1355
rect 16377 -6115 16443 -4355
rect 16535 -3115 16601 -1355
rect 16693 -6115 16759 -4355
rect 16851 -3115 16917 -1355
rect 17009 -6115 17075 -4355
rect 17167 -3115 17233 -1355
rect 17325 -6115 17391 -4355
rect 17483 -3115 17549 -1355
rect 17641 -6115 17707 -4355
rect 17799 -3115 17865 -1355
rect 17957 -6115 18023 -4355
rect 18115 -3115 18181 -1355
rect 18273 -6115 18339 -4355
rect 18431 -3115 18497 -1355
rect 18589 -6115 18655 -4355
rect 18747 -3115 18813 -1355
rect 18905 -6115 18971 -4355
rect 14240 -6860 14252 -6790
rect 14252 -6860 18886 -6790
rect 18886 -6860 18890 -6790
rect 20540 -690 20552 -620
rect 20552 -690 25186 -620
rect 25186 -690 25200 -620
rect 20465 -6115 20531 -4355
rect 20623 -3115 20689 -1355
rect 20781 -6115 20847 -4355
rect 20939 -3115 21005 -1355
rect 21097 -6115 21163 -4355
rect 21255 -3115 21321 -1355
rect 21413 -6115 21479 -4355
rect 21571 -3115 21637 -1355
rect 21729 -6115 21795 -4355
rect 21887 -3115 21953 -1355
rect 22045 -6115 22111 -4355
rect 22203 -3115 22269 -1355
rect 22361 -6115 22427 -4355
rect 22519 -3115 22585 -1355
rect 22677 -6115 22743 -4355
rect 22835 -3115 22901 -1355
rect 22993 -6115 23059 -4355
rect 23151 -3115 23217 -1355
rect 23309 -6115 23375 -4355
rect 23467 -3115 23533 -1355
rect 23625 -6115 23691 -4355
rect 23783 -3115 23849 -1355
rect 23941 -6115 24007 -4355
rect 24099 -3115 24165 -1355
rect 24257 -6115 24323 -4355
rect 24415 -3115 24481 -1355
rect 24573 -6115 24639 -4355
rect 24731 -3115 24797 -1355
rect 24889 -6115 24955 -4355
rect 25047 -3115 25113 -1355
rect 25205 -6115 25271 -4355
rect 20540 -6860 20552 -6790
rect 20552 -6860 25186 -6790
rect 25186 -6860 25190 -6790
<< metal3 >>
rect 1500 6380 6500 6500
rect 1500 6310 1640 6380
rect 6300 6310 6500 6380
rect 1500 6300 6500 6310
rect 7800 6380 12800 6500
rect 7800 6310 7940 6380
rect 12600 6310 12800 6380
rect 7800 6300 12800 6310
rect 14100 6380 19100 6500
rect 14100 6310 14240 6380
rect 18900 6310 19100 6380
rect 14100 6300 19100 6310
rect 20400 6380 25400 6500
rect 20400 6310 20540 6380
rect 25200 6310 25400 6380
rect 20400 6300 25400 6310
rect 1400 5700 6510 5800
rect 1400 3900 1500 5700
rect 2800 5645 6510 5700
rect 2800 3900 2987 5645
rect 1400 3885 1723 3900
rect 1789 3885 2039 3900
rect 2105 3885 2355 3900
rect 2421 3885 2671 3900
rect 2737 3885 2987 3900
rect 3053 3885 3303 5645
rect 3369 3885 3619 5645
rect 3685 3885 3935 5645
rect 4001 3885 4251 5645
rect 4317 3885 4567 5645
rect 4633 3885 4883 5645
rect 4949 3885 5199 5645
rect 5265 3885 5515 5645
rect 5581 3885 5831 5645
rect 5897 3885 6147 5645
rect 6213 3885 6510 5645
rect 1400 3800 6510 3885
rect 7700 5700 12810 5800
rect 7700 3900 7800 5700
rect 9000 5645 12810 5700
rect 7700 3885 8023 3900
rect 8089 3885 8339 3900
rect 8405 3885 8655 3900
rect 8721 3885 8971 3900
rect 9037 3885 9287 5645
rect 9353 3885 9603 5645
rect 9669 3885 9919 5645
rect 9985 3885 10235 5645
rect 10301 3885 10551 5645
rect 10617 3885 10867 5645
rect 10933 3885 11183 5645
rect 11249 3885 11499 5645
rect 11565 3885 11815 5645
rect 11881 3885 12131 5645
rect 12197 3885 12447 5645
rect 12513 3885 12810 5645
rect 7700 3800 12810 3885
rect 14000 5700 19110 5800
rect 14000 3900 14100 5700
rect 15400 5645 19110 5700
rect 15400 3900 15587 5645
rect 14000 3885 14323 3900
rect 14389 3885 14639 3900
rect 14705 3885 14955 3900
rect 15021 3885 15271 3900
rect 15337 3885 15587 3900
rect 15653 3885 15903 5645
rect 15969 3885 16219 5645
rect 16285 3885 16535 5645
rect 16601 3885 16851 5645
rect 16917 3885 17167 5645
rect 17233 3885 17483 5645
rect 17549 3885 17799 5645
rect 17865 3885 18115 5645
rect 18181 3885 18431 5645
rect 18497 3885 18747 5645
rect 18813 3885 19110 5645
rect 14000 3800 19110 3885
rect 20300 5700 25410 5800
rect 20300 3900 20400 5700
rect 21600 5645 25410 5700
rect 20300 3885 20623 3900
rect 20689 3885 20939 3900
rect 21005 3885 21255 3900
rect 21321 3885 21571 3900
rect 21637 3885 21887 5645
rect 21953 3885 22203 5645
rect 22269 3885 22519 5645
rect 22585 3885 22835 5645
rect 22901 3885 23151 5645
rect 23217 3885 23467 5645
rect 23533 3885 23783 5645
rect 23849 3885 24099 5645
rect 24165 3885 24415 5645
rect 24481 3885 24731 5645
rect 24797 3885 25047 5645
rect 25113 3885 25410 5645
rect 20300 3800 25410 3885
rect 1400 2700 6510 2800
rect 1400 900 1500 2700
rect 2800 2645 6510 2700
rect 2800 900 2829 2645
rect 1400 885 1565 900
rect 1631 885 1881 900
rect 1947 885 2197 900
rect 2263 885 2513 900
rect 2579 885 2829 900
rect 2895 885 3145 2645
rect 3211 885 3461 2645
rect 3527 885 3777 2645
rect 3843 885 4093 2645
rect 4159 885 4409 2645
rect 4475 885 4725 2645
rect 4791 885 5041 2645
rect 5107 885 5357 2645
rect 5423 885 5673 2645
rect 5739 885 5989 2645
rect 6055 885 6305 2645
rect 6371 885 6510 2645
rect 1400 800 6510 885
rect 7730 2700 13000 2800
rect 7730 2645 11600 2700
rect 7730 885 7865 2645
rect 7931 885 8181 2645
rect 8247 885 8497 2645
rect 8563 885 8813 2645
rect 8879 885 9129 2645
rect 9195 885 9445 2645
rect 9511 885 9761 2645
rect 9827 885 10077 2645
rect 10143 885 10393 2645
rect 10459 885 10709 2645
rect 10775 885 11025 2645
rect 11091 885 11341 2645
rect 11407 900 11600 2645
rect 12900 900 13000 2700
rect 11407 885 11657 900
rect 11723 885 11973 900
rect 12039 885 12289 900
rect 12355 885 12605 900
rect 12671 885 13000 900
rect 7730 800 13000 885
rect 14000 2700 19110 2800
rect 14000 900 14100 2700
rect 15400 2645 19110 2700
rect 15400 900 15429 2645
rect 14000 885 14165 900
rect 14231 885 14481 900
rect 14547 885 14797 900
rect 14863 885 15113 900
rect 15179 885 15429 900
rect 15495 885 15745 2645
rect 15811 885 16061 2645
rect 16127 885 16377 2645
rect 16443 885 16693 2645
rect 16759 885 17009 2645
rect 17075 885 17325 2645
rect 17391 885 17641 2645
rect 17707 885 17957 2645
rect 18023 885 18273 2645
rect 18339 885 18589 2645
rect 18655 885 18905 2645
rect 18971 885 19110 2645
rect 14000 800 19110 885
rect 20330 2700 25600 2800
rect 20330 2645 24200 2700
rect 20330 885 20465 2645
rect 20531 885 20781 2645
rect 20847 885 21097 2645
rect 21163 885 21413 2645
rect 21479 885 21729 2645
rect 21795 885 22045 2645
rect 22111 885 22361 2645
rect 22427 885 22677 2645
rect 22743 885 22993 2645
rect 23059 885 23309 2645
rect 23375 885 23625 2645
rect 23691 885 23941 2645
rect 24007 900 24200 2645
rect 25500 900 25600 2700
rect 24007 885 24257 900
rect 24323 885 24573 900
rect 24639 885 24889 900
rect 24955 885 25205 900
rect 25271 885 25600 900
rect 20330 800 25600 885
rect 3100 400 5000 500
rect 3100 300 3300 400
rect 1400 210 3300 300
rect 4800 300 5000 400
rect 15700 400 17600 500
rect 15700 300 15900 400
rect 4800 210 7400 300
rect 1400 140 1640 210
rect 6290 180 7400 210
rect 6290 140 7020 180
rect 1400 100 3300 140
rect 4800 100 7020 140
rect 1400 20 7020 100
rect 7380 20 7400 180
rect 1400 0 7400 20
rect 7600 210 13700 300
rect 7600 140 7940 210
rect 12590 180 13700 210
rect 12590 140 13320 180
rect 7600 20 13320 140
rect 13680 20 13700 180
rect 7600 0 13700 20
rect 13900 210 15900 300
rect 17400 300 17600 400
rect 17400 210 20000 300
rect 13900 140 14240 210
rect 18890 180 20000 210
rect 18890 140 19620 180
rect 13900 100 15900 140
rect 17400 100 19620 140
rect 13900 20 19620 100
rect 19980 20 20000 180
rect 13900 0 20000 20
rect 20200 210 25400 300
rect 20200 140 20540 210
rect 25190 140 25400 210
rect 20200 0 25400 140
rect 7600 -200 7900 0
rect 9400 -100 12000 0
rect 13900 -100 14100 0
rect 20200 -100 20500 0
rect 22000 -100 24600 0
rect 6500 -400 7900 -200
rect 12800 -300 14100 -100
rect 19100 -300 20500 -100
rect 3100 -500 5000 -400
rect 6500 -500 6800 -400
rect 9400 -500 12000 -400
rect 12800 -500 13100 -300
rect 15700 -500 17600 -400
rect 19100 -500 19400 -300
rect 22000 -500 24600 -400
rect 1400 -620 3300 -500
rect 4800 -620 6800 -500
rect 1400 -690 1640 -620
rect 6300 -690 6800 -620
rect 1400 -800 3300 -690
rect 4800 -800 6800 -690
rect 7000 -520 13100 -500
rect 7000 -680 7020 -520
rect 7380 -620 13100 -520
rect 7380 -680 7940 -620
rect 7000 -690 7940 -680
rect 12600 -690 13100 -620
rect 7000 -800 13100 -690
rect 13300 -520 15900 -500
rect 13300 -680 13320 -520
rect 13680 -620 15900 -520
rect 17400 -620 19400 -500
rect 13680 -680 14240 -620
rect 13300 -690 14240 -680
rect 18900 -690 19400 -620
rect 13300 -800 15900 -690
rect 17400 -800 19400 -690
rect 19600 -520 25400 -500
rect 19600 -680 19620 -520
rect 19980 -620 25400 -520
rect 19980 -680 20540 -620
rect 19600 -690 20540 -680
rect 25200 -690 25400 -620
rect 19600 -800 25400 -690
rect 3100 -900 5000 -800
rect 15700 -900 17600 -800
rect 1430 -1300 6510 -1200
rect 1430 -1355 3400 -1300
rect 4700 -1355 6510 -1300
rect 1430 -3115 1723 -1355
rect 1789 -3115 2039 -1355
rect 2105 -3115 2355 -1355
rect 2421 -3115 2671 -1355
rect 2737 -3115 2987 -1355
rect 3053 -3115 3303 -1355
rect 3369 -3100 3400 -1355
rect 4700 -3100 4883 -1355
rect 3369 -3115 3619 -3100
rect 3685 -3115 3935 -3100
rect 4001 -3115 4251 -3100
rect 4317 -3115 4567 -3100
rect 4633 -3115 4883 -3100
rect 4949 -3115 5199 -1355
rect 5265 -3115 5515 -1355
rect 5581 -3115 5831 -1355
rect 5897 -3115 6147 -1355
rect 6213 -3115 6510 -1355
rect 1430 -3200 6510 -3115
rect 7700 -1300 12810 -1200
rect 7700 -3100 7800 -1300
rect 9100 -1355 12810 -1300
rect 9100 -3100 9287 -1355
rect 7700 -3115 8023 -3100
rect 8089 -3115 8339 -3100
rect 8405 -3115 8655 -3100
rect 8721 -3115 8971 -3100
rect 9037 -3115 9287 -3100
rect 9353 -3115 9603 -1355
rect 9669 -3115 9919 -1355
rect 9985 -3115 10235 -1355
rect 10301 -3115 10551 -1355
rect 10617 -3115 10867 -1355
rect 10933 -3115 11183 -1355
rect 11249 -3115 11499 -1355
rect 11565 -3115 11815 -1355
rect 11881 -3115 12131 -1355
rect 12197 -3115 12447 -1355
rect 12513 -3115 12810 -1355
rect 7700 -3200 12810 -3115
rect 14030 -1300 19110 -1200
rect 14030 -1355 16000 -1300
rect 17300 -1355 19110 -1300
rect 14030 -3115 14323 -1355
rect 14389 -3115 14639 -1355
rect 14705 -3115 14955 -1355
rect 15021 -3115 15271 -1355
rect 15337 -3115 15587 -1355
rect 15653 -3115 15903 -1355
rect 15969 -3100 16000 -1355
rect 17300 -3100 17483 -1355
rect 15969 -3115 16219 -3100
rect 16285 -3115 16535 -3100
rect 16601 -3115 16851 -3100
rect 16917 -3115 17167 -3100
rect 17233 -3115 17483 -3100
rect 17549 -3115 17799 -1355
rect 17865 -3115 18115 -1355
rect 18181 -3115 18431 -1355
rect 18497 -3115 18747 -1355
rect 18813 -3115 19110 -1355
rect 14030 -3200 19110 -3115
rect 20300 -1300 25410 -1200
rect 20300 -3100 20400 -1300
rect 21700 -1355 25410 -1300
rect 21700 -3100 21887 -1355
rect 20300 -3115 20623 -3100
rect 20689 -3115 20939 -3100
rect 21005 -3115 21255 -3100
rect 21321 -3115 21571 -3100
rect 21637 -3115 21887 -3100
rect 21953 -3115 22203 -1355
rect 22269 -3115 22519 -1355
rect 22585 -3115 22835 -1355
rect 22901 -3115 23151 -1355
rect 23217 -3115 23467 -1355
rect 23533 -3115 23783 -1355
rect 23849 -3115 24099 -1355
rect 24165 -3115 24415 -1355
rect 24481 -3115 24731 -1355
rect 24797 -3115 25047 -1355
rect 25113 -3115 25410 -1355
rect 20300 -3200 25410 -3115
rect 1430 -4300 6700 -4200
rect 1430 -4355 5300 -4300
rect 1430 -6115 1565 -4355
rect 1631 -6115 1881 -4355
rect 1947 -6115 2197 -4355
rect 2263 -6115 2513 -4355
rect 2579 -6115 2829 -4355
rect 2895 -6115 3145 -4355
rect 3211 -6115 3461 -4355
rect 3527 -6115 3777 -4355
rect 3843 -6115 4093 -4355
rect 4159 -6115 4409 -4355
rect 4475 -6115 4725 -4355
rect 4791 -6115 5041 -4355
rect 5107 -6100 5300 -4355
rect 6600 -6100 6700 -4300
rect 5107 -6115 5357 -6100
rect 5423 -6115 5673 -6100
rect 5739 -6115 5989 -6100
rect 6055 -6115 6305 -6100
rect 6371 -6115 6700 -6100
rect 1430 -6200 6700 -6115
rect 7730 -4300 12810 -4200
rect 7730 -4355 9700 -4300
rect 11000 -4355 12810 -4300
rect 7730 -6115 7865 -4355
rect 7931 -6115 8181 -4355
rect 8247 -6115 8497 -4355
rect 8563 -6115 8813 -4355
rect 8879 -6115 9129 -4355
rect 9195 -6115 9445 -4355
rect 9511 -6100 9700 -4355
rect 11000 -6100 11025 -4355
rect 9511 -6115 9761 -6100
rect 9827 -6115 10077 -6100
rect 10143 -6115 10393 -6100
rect 10459 -6115 10709 -6100
rect 10775 -6115 11025 -6100
rect 11091 -6115 11341 -4355
rect 11407 -6115 11657 -4355
rect 11723 -6115 11973 -4355
rect 12039 -6115 12289 -4355
rect 12355 -6115 12605 -4355
rect 12671 -6115 12810 -4355
rect 7730 -6200 12810 -6115
rect 14030 -4300 19300 -4200
rect 14030 -4355 17900 -4300
rect 14030 -6115 14165 -4355
rect 14231 -6115 14481 -4355
rect 14547 -6115 14797 -4355
rect 14863 -6115 15113 -4355
rect 15179 -6115 15429 -4355
rect 15495 -6115 15745 -4355
rect 15811 -6115 16061 -4355
rect 16127 -6115 16377 -4355
rect 16443 -6115 16693 -4355
rect 16759 -6115 17009 -4355
rect 17075 -6115 17325 -4355
rect 17391 -6115 17641 -4355
rect 17707 -6100 17900 -4355
rect 19200 -6100 19300 -4300
rect 17707 -6115 17957 -6100
rect 18023 -6115 18273 -6100
rect 18339 -6115 18589 -6100
rect 18655 -6115 18905 -6100
rect 18971 -6115 19300 -6100
rect 14030 -6200 19300 -6115
rect 20300 -4300 25600 -4200
rect 20300 -4355 22300 -4300
rect 23600 -4355 25600 -4300
rect 20300 -6115 20465 -4355
rect 20531 -6115 20781 -4355
rect 20847 -6115 21097 -4355
rect 21163 -6115 21413 -4355
rect 21479 -6115 21729 -4355
rect 21795 -6115 22045 -4355
rect 22111 -6100 22300 -4355
rect 23600 -6100 23625 -4355
rect 22111 -6115 22361 -6100
rect 22427 -6115 22677 -6100
rect 22743 -6115 22993 -6100
rect 23059 -6115 23309 -6100
rect 23375 -6115 23625 -6100
rect 23691 -6115 23941 -4355
rect 24007 -6115 24257 -4355
rect 24323 -6115 24573 -4355
rect 24639 -6115 24889 -4355
rect 24955 -6115 25205 -4355
rect 25271 -6115 25600 -4355
rect 20300 -6200 25600 -6115
rect 1500 -6790 6500 -6770
rect 1500 -6860 1640 -6790
rect 6290 -6860 6500 -6790
rect 1500 -6970 6500 -6860
rect 7800 -6790 12800 -6770
rect 7800 -6860 7940 -6790
rect 12590 -6860 12800 -6790
rect 7800 -6970 12800 -6860
rect 14100 -6790 19100 -6770
rect 14100 -6860 14240 -6790
rect 18890 -6860 19100 -6790
rect 14100 -6970 19100 -6860
rect 20400 -6790 25400 -6770
rect 20400 -6860 20540 -6790
rect 25190 -6860 25400 -6790
rect 20400 -6970 25400 -6860
<< via3 >>
rect 1500 5645 2800 5700
rect 1500 3900 1723 5645
rect 1723 3900 1789 5645
rect 1789 3900 2039 5645
rect 2039 3900 2105 5645
rect 2105 3900 2355 5645
rect 2355 3900 2421 5645
rect 2421 3900 2671 5645
rect 2671 3900 2737 5645
rect 2737 3900 2800 5645
rect 7800 5645 9000 5700
rect 7800 3900 8023 5645
rect 8023 3900 8089 5645
rect 8089 3900 8339 5645
rect 8339 3900 8405 5645
rect 8405 3900 8655 5645
rect 8655 3900 8721 5645
rect 8721 3900 8971 5645
rect 8971 3900 9000 5645
rect 14100 5645 15400 5700
rect 14100 3900 14323 5645
rect 14323 3900 14389 5645
rect 14389 3900 14639 5645
rect 14639 3900 14705 5645
rect 14705 3900 14955 5645
rect 14955 3900 15021 5645
rect 15021 3900 15271 5645
rect 15271 3900 15337 5645
rect 15337 3900 15400 5645
rect 20400 5645 21600 5700
rect 20400 3900 20623 5645
rect 20623 3900 20689 5645
rect 20689 3900 20939 5645
rect 20939 3900 21005 5645
rect 21005 3900 21255 5645
rect 21255 3900 21321 5645
rect 21321 3900 21571 5645
rect 21571 3900 21600 5645
rect 1500 2645 2800 2700
rect 1500 900 1565 2645
rect 1565 900 1631 2645
rect 1631 900 1881 2645
rect 1881 900 1947 2645
rect 1947 900 2197 2645
rect 2197 900 2263 2645
rect 2263 900 2513 2645
rect 2513 900 2579 2645
rect 2579 900 2800 2645
rect 11600 2645 12900 2700
rect 11600 900 11657 2645
rect 11657 900 11723 2645
rect 11723 900 11973 2645
rect 11973 900 12039 2645
rect 12039 900 12289 2645
rect 12289 900 12355 2645
rect 12355 900 12605 2645
rect 12605 900 12671 2645
rect 12671 900 12900 2645
rect 14100 2645 15400 2700
rect 14100 900 14165 2645
rect 14165 900 14231 2645
rect 14231 900 14481 2645
rect 14481 900 14547 2645
rect 14547 900 14797 2645
rect 14797 900 14863 2645
rect 14863 900 15113 2645
rect 15113 900 15179 2645
rect 15179 900 15400 2645
rect 24200 2645 25500 2700
rect 24200 900 24257 2645
rect 24257 900 24323 2645
rect 24323 900 24573 2645
rect 24573 900 24639 2645
rect 24639 900 24889 2645
rect 24889 900 24955 2645
rect 24955 900 25205 2645
rect 25205 900 25271 2645
rect 25271 900 25500 2645
rect 3300 210 4800 400
rect 3300 140 4800 210
rect 3300 100 4800 140
rect 7020 20 7380 180
rect 13320 20 13680 180
rect 15900 210 17400 400
rect 15900 140 17400 210
rect 15900 100 17400 140
rect 19620 20 19980 180
rect 3300 -620 4800 -500
rect 3300 -690 4800 -620
rect 3300 -800 4800 -690
rect 7020 -680 7380 -520
rect 13320 -680 13680 -520
rect 15900 -620 17400 -500
rect 15900 -690 17400 -620
rect 15900 -800 17400 -690
rect 19620 -680 19980 -520
rect 3400 -1355 4700 -1300
rect 3400 -3100 3619 -1355
rect 3619 -3100 3685 -1355
rect 3685 -3100 3935 -1355
rect 3935 -3100 4001 -1355
rect 4001 -3100 4251 -1355
rect 4251 -3100 4317 -1355
rect 4317 -3100 4567 -1355
rect 4567 -3100 4633 -1355
rect 4633 -3100 4700 -1355
rect 7800 -1355 9100 -1300
rect 7800 -3100 8023 -1355
rect 8023 -3100 8089 -1355
rect 8089 -3100 8339 -1355
rect 8339 -3100 8405 -1355
rect 8405 -3100 8655 -1355
rect 8655 -3100 8721 -1355
rect 8721 -3100 8971 -1355
rect 8971 -3100 9037 -1355
rect 9037 -3100 9100 -1355
rect 16000 -1355 17300 -1300
rect 16000 -3100 16219 -1355
rect 16219 -3100 16285 -1355
rect 16285 -3100 16535 -1355
rect 16535 -3100 16601 -1355
rect 16601 -3100 16851 -1355
rect 16851 -3100 16917 -1355
rect 16917 -3100 17167 -1355
rect 17167 -3100 17233 -1355
rect 17233 -3100 17300 -1355
rect 20400 -1355 21700 -1300
rect 20400 -3100 20623 -1355
rect 20623 -3100 20689 -1355
rect 20689 -3100 20939 -1355
rect 20939 -3100 21005 -1355
rect 21005 -3100 21255 -1355
rect 21255 -3100 21321 -1355
rect 21321 -3100 21571 -1355
rect 21571 -3100 21637 -1355
rect 21637 -3100 21700 -1355
rect 5300 -4355 6600 -4300
rect 5300 -6100 5357 -4355
rect 5357 -6100 5423 -4355
rect 5423 -6100 5673 -4355
rect 5673 -6100 5739 -4355
rect 5739 -6100 5989 -4355
rect 5989 -6100 6055 -4355
rect 6055 -6100 6305 -4355
rect 6305 -6100 6371 -4355
rect 6371 -6100 6600 -4355
rect 9700 -4355 11000 -4300
rect 9700 -6100 9761 -4355
rect 9761 -6100 9827 -4355
rect 9827 -6100 10077 -4355
rect 10077 -6100 10143 -4355
rect 10143 -6100 10393 -4355
rect 10393 -6100 10459 -4355
rect 10459 -6100 10709 -4355
rect 10709 -6100 10775 -4355
rect 10775 -6100 11000 -4355
rect 17900 -4355 19200 -4300
rect 17900 -6100 17957 -4355
rect 17957 -6100 18023 -4355
rect 18023 -6100 18273 -4355
rect 18273 -6100 18339 -4355
rect 18339 -6100 18589 -4355
rect 18589 -6100 18655 -4355
rect 18655 -6100 18905 -4355
rect 18905 -6100 18971 -4355
rect 18971 -6100 19200 -4355
rect 22300 -4355 23600 -4300
rect 22300 -6100 22361 -4355
rect 22361 -6100 22427 -4355
rect 22427 -6100 22677 -4355
rect 22677 -6100 22743 -4355
rect 22743 -6100 22993 -4355
rect 22993 -6100 23059 -4355
rect 23059 -6100 23309 -4355
rect 23309 -6100 23375 -4355
rect 23375 -6100 23600 -4355
<< metal4 >>
rect 5200 11100 6700 11200
rect 5200 9500 5300 11100
rect 6600 9500 6700 11100
rect 1400 8000 2900 8200
rect 1400 6600 1600 8000
rect 2800 6600 2900 8000
rect 1400 5700 2900 6600
rect 1400 3900 1500 5700
rect 2800 3900 2900 5700
rect 1400 3800 2900 3900
rect 1400 2700 2900 2800
rect 1400 900 1500 2700
rect 2800 900 2900 2700
rect 1400 -9900 2900 900
rect 3200 400 4900 500
rect 3200 100 3300 400
rect 4800 100 4900 400
rect 3200 0 4900 100
rect 3200 -500 4900 -400
rect 3200 -800 3300 -500
rect 4800 -800 4900 -500
rect 3200 -900 4900 -800
rect 3300 -1300 4800 -1200
rect 3300 -3100 3400 -1300
rect 4700 -3100 4800 -1300
rect 3300 -6900 4800 -3100
rect 5200 -4300 6700 9500
rect 7700 11100 9200 11200
rect 7700 9500 7800 11100
rect 9100 9500 9200 11100
rect 7700 5700 9200 9500
rect 17800 11100 19300 11200
rect 17800 9500 17900 11100
rect 19200 9500 19300 11100
rect 7700 3900 7800 5700
rect 9000 3900 9200 5700
rect 7700 3800 9200 3900
rect 9600 8100 11100 8200
rect 9600 6500 9800 8100
rect 11000 6500 11100 8100
rect 7000 180 7400 200
rect 7000 20 7020 180
rect 7380 20 7400 180
rect 7000 -520 7400 20
rect 7000 -680 7020 -520
rect 7380 -680 7400 -520
rect 7000 -700 7400 -680
rect 5200 -6100 5300 -4300
rect 6600 -6100 6700 -4300
rect 5200 -6200 6700 -6100
rect 7700 -1300 9200 -1200
rect 7700 -3100 7800 -1300
rect 9100 -3100 9200 -1300
rect 3300 -8500 3400 -6900
rect 4700 -8500 4800 -6900
rect 3300 -8600 4800 -8500
rect 1400 -11500 1500 -9900
rect 2800 -11500 2900 -9900
rect 1400 -11600 2900 -11500
rect 7700 -9900 9200 -3100
rect 9600 -4300 11100 6500
rect 14000 8000 15500 8200
rect 14000 6600 14200 8000
rect 15400 6600 15500 8000
rect 14000 5700 15500 6600
rect 14000 3900 14100 5700
rect 15400 3900 15500 5700
rect 14000 3800 15500 3900
rect 9600 -6100 9700 -4300
rect 11000 -6100 11100 -4300
rect 9600 -6200 11100 -6100
rect 11500 2700 13000 2800
rect 11500 900 11600 2700
rect 12900 900 13000 2700
rect 11500 -6900 13000 900
rect 14000 2700 15500 2800
rect 14000 900 14100 2700
rect 15400 900 15500 2700
rect 13300 180 13700 200
rect 13300 20 13320 180
rect 13680 20 13700 180
rect 13300 -520 13700 20
rect 13300 -680 13320 -520
rect 13680 -680 13700 -520
rect 13300 -700 13700 -680
rect 11500 -8500 11600 -6900
rect 12900 -8500 13000 -6900
rect 11500 -8600 13000 -8500
rect 14000 -9900 15500 900
rect 15800 400 17500 500
rect 15800 100 15900 400
rect 17400 100 17500 400
rect 15800 0 17500 100
rect 15800 -500 17500 -400
rect 15800 -800 15900 -500
rect 17400 -800 17500 -500
rect 15800 -900 17500 -800
rect 15900 -1300 17400 -1200
rect 15900 -3100 16000 -1300
rect 17300 -3100 17400 -1300
rect 15900 -6900 17400 -3100
rect 17800 -4300 19300 9500
rect 20300 11100 21800 11200
rect 20300 9500 20400 11100
rect 21700 9500 21800 11100
rect 20300 8200 21800 9500
rect 20300 6600 21900 8200
rect 22200 8100 23700 8200
rect 20300 5700 21800 6600
rect 20300 3900 20400 5700
rect 21600 3900 21800 5700
rect 20300 3800 21800 3900
rect 22200 6500 22400 8100
rect 23600 6500 23700 8100
rect 19600 180 20000 200
rect 19600 20 19620 180
rect 19980 20 20000 180
rect 19600 -520 20000 20
rect 19600 -680 19620 -520
rect 19980 -680 20000 -520
rect 19600 -700 20000 -680
rect 17800 -6100 17900 -4300
rect 19200 -6100 19300 -4300
rect 17800 -6200 19300 -6100
rect 20300 -1300 21800 -1200
rect 20300 -3100 20400 -1300
rect 21700 -3100 21800 -1300
rect 15900 -8500 16000 -6900
rect 17300 -8500 17400 -6900
rect 15900 -8600 17400 -8500
rect 7700 -11500 7800 -9900
rect 9100 -11500 9200 -9900
rect 7700 -11600 9200 -11500
rect 11500 -11500 11600 -9900
rect 12800 -11500 13000 -9900
rect 11500 -11600 13000 -11500
rect 14000 -11500 14100 -9900
rect 15400 -11500 15500 -9900
rect 14000 -11600 15500 -11500
rect 20300 -9900 21800 -3100
rect 22200 -4300 23700 6500
rect 22200 -6100 22300 -4300
rect 23600 -6100 23700 -4300
rect 22200 -6200 23700 -6100
rect 24100 2700 25600 2800
rect 24100 900 24200 2700
rect 25500 900 25600 2700
rect 24100 -6900 25600 900
rect 24100 -8500 24200 -6900
rect 25500 -8500 25600 -6900
rect 24100 -8600 25600 -8500
rect 20300 -11500 20400 -9900
rect 21700 -11500 21800 -9900
rect 20300 -11600 21800 -11500
<< via4 >>
rect 5300 9500 6600 11100
rect 1600 6600 2800 8000
rect 3300 100 4800 400
rect 3300 -800 4800 -500
rect 7800 9500 9100 11100
rect 17900 9500 19200 11100
rect 9800 6500 11000 8100
rect 3400 -8500 4700 -6900
rect 1500 -11500 2800 -9900
rect 14200 6600 15400 8000
rect 11600 -8500 12900 -6900
rect 15900 100 17400 400
rect 15900 -800 17400 -500
rect 20400 9500 21700 11100
rect 22400 6500 23600 8100
rect 16000 -8500 17300 -6900
rect 7800 -11500 9100 -9900
rect 14100 -11500 15400 -9900
rect 24200 -8500 25500 -6900
rect 20400 -11500 21700 -9900
<< metal5 >>
rect 1400 8200 4200 11400
rect 22800 11200 25600 11400
rect 5200 11100 25600 11200
rect 5200 9500 5300 11100
rect 6600 9500 7800 11100
rect 9100 9500 17900 11100
rect 19200 9500 20400 11100
rect 21700 9500 25600 11100
rect 5200 9400 25600 9500
rect 1400 8100 23700 8200
rect 1400 8000 9800 8100
rect 1400 6600 1600 8000
rect 2800 6600 9800 8000
rect 1400 6500 9800 6600
rect 11000 8000 22400 8100
rect 11000 6600 14200 8000
rect 15400 6600 22400 8000
rect 11000 6500 22400 6600
rect 23600 6500 23700 8100
rect 1400 6400 23700 6500
rect 1300 400 25500 500
rect 1300 100 3300 400
rect 4800 100 15900 400
rect 17400 100 25500 400
rect 1300 0 25500 100
rect 1300 -500 25500 -400
rect 1300 -800 3300 -500
rect 4800 -800 15900 -500
rect 17400 -800 25500 -500
rect 1300 -900 25500 -800
rect 3300 -6900 25600 -6800
rect 3300 -8500 3400 -6900
rect 4700 -8500 11600 -6900
rect 12900 -8500 16000 -6900
rect 17300 -8500 24200 -6900
rect 25500 -8500 25600 -6900
rect 3300 -8600 25600 -8500
rect 1400 -9900 21800 -9800
rect 1400 -11500 1500 -9900
rect 2800 -11500 7800 -9900
rect 9100 -11500 14100 -9900
rect 15400 -11500 20400 -9900
rect 21700 -11500 21800 -9900
rect 1400 -11600 21800 -11500
rect 1400 -11800 4200 -11600
rect 22800 -11800 25600 -8600
<< labels >>
rlabel metal5 1300 0 1400 500 1 GL
rlabel metal5 1300 -900 1400 -400 1 GR
rlabel metal5 1400 -11800 4200 -11600 1 SD2L
rlabel metal5 22800 -11800 25600 -11600 1 SD2R
rlabel metal5 22800 11200 25600 11400 1 SD1R
rlabel metal5 1400 11200 4200 11400 1 SD1L
rlabel metal2 14030 -580 14100 -520 1 SUB
<< end >>
