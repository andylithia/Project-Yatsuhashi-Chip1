magic
tech sky130B
magscale 1 2
timestamp 1661127237
<< metal3 >>
rect 12000 23800 20000 24000
rect 12000 20400 12200 23800
rect 19800 20400 20000 23800
rect 12000 20200 20000 20400
rect 21000 23800 25000 24000
rect 21000 19200 21200 23800
rect 12800 14200 21200 19200
rect 24800 14200 25000 23800
rect 12800 14000 25000 14200
rect 12800 8000 20000 14000
<< via3 >>
rect 12200 20400 19800 23800
rect 21200 14200 24800 23800
rect -1400 2600 -600 6600
<< mimcap >>
rect 13000 18800 19800 19000
rect 13000 8400 13200 18800
rect 19600 8400 19800 18800
rect 13000 8200 19800 8400
<< mimcapcontact >>
rect 13200 8400 19600 18800
<< metal4 >>
rect 12000 23800 20000 24000
rect 12000 20400 12200 23800
rect 19800 20400 20000 23800
rect 12000 18800 20000 20400
rect 12000 14000 13200 18800
rect -5200 12000 -600 13200
rect 12800 8400 13200 14000
rect 19600 8400 20000 18800
rect 21000 23800 25000 24000
rect 21000 14200 21200 23800
rect 24800 14200 25000 23800
rect 21000 14000 25000 14200
rect 12800 8000 20000 8400
rect -1600 6600 -400 6800
rect -1600 2600 -1400 6600
rect -600 2600 -400 6600
rect -1600 2400 -400 2600
rect 13800 1200 18000 6000
rect 16000 1000 18000 1200
rect 16000 800 20000 1000
rect 16000 600 47400 800
rect 16000 -4000 33600 600
rect 20000 -4200 41000 -4000
rect 40800 -10800 41000 -4200
rect 47200 -10800 47400 600
rect 40800 -16800 47400 -10800
<< via4 >>
rect 21200 14200 24800 23800
rect -1400 2600 -600 6600
rect 33600 -4000 47200 600
rect 41000 -10800 47200 -4000
<< mimcap2 >>
rect 13000 18800 19800 19000
rect 13000 8400 13200 18800
rect 19600 8400 19800 18800
rect 13000 8200 19800 8400
<< mimcap2contact >>
rect 13200 8400 19600 18800
<< metal5 >>
rect 20600 24000 26000 25200
rect 20000 23800 54600 24000
rect 20000 19200 21200 23800
rect 12800 18800 21200 19200
rect 12800 8400 13200 18800
rect 19600 14200 21200 18800
rect 24800 20000 54600 23800
rect 24800 19000 30000 20000
rect 24800 18000 29000 19000
rect 24800 17000 28000 18000
rect 24800 16000 27000 17000
rect 24800 15000 26000 16000
rect 24800 14200 25000 15000
rect 19600 14000 25000 14200
rect 19600 13000 24000 14000
rect 19600 12000 23000 13000
rect 19600 8400 20000 12000
rect 12800 8000 20000 8400
rect -6600 6600 -400 6800
rect -6600 5800 -1400 6600
rect -1600 2600 -1400 5800
rect -600 2600 -400 6600
rect -1600 2400 -400 2600
rect 33400 600 47400 800
rect 33400 -4000 33600 600
rect 33400 -4200 41000 -4000
rect 40800 -10800 41000 -4200
rect 47200 -10800 47400 600
rect 40800 -16800 47400 -10800
use PA_complete_without_ind  PA_complete_without_ind_0
timestamp 1661126380
transform 1 0 1 0 1 0
box -9600 -4000 17800 12600
use octa_ind_3t_140_160_flat  octa_ind_3t_140_160_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1660524083
transform 0 -1 -24800 1 0 49100
box -39300 -34000 -5300 -6000
use octa_ind_thick_1p8n_flat_mod1  octa_ind_thick_1p8n_flat_mod1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1660790920
transform 0 1 65600 -1 0 -23300
box -47300 -45000 2700 5000
<< end >>
