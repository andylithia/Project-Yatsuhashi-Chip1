magic
tech sky130A
magscale 1 2
timestamp 1664821665
<< pwell >>
rect 30600 12500 31000 14016
<< psubdiff >>
rect 30634 13946 30730 13980
rect 30868 13946 30964 13980
rect 30634 13884 30668 13946
rect 30930 13884 30964 13946
rect 30634 12570 30668 12632
rect 30930 12570 30964 12632
rect 30634 12536 30730 12570
rect 30868 12536 30964 12570
<< psubdiffcont >>
rect 30730 13946 30868 13980
rect 30634 12632 30668 13884
rect 30930 12632 30964 13884
rect 30730 12536 30868 12570
<< xpolycontact >>
rect 30764 13418 30834 13850
rect 30764 12666 30834 13098
<< ppolyres >>
rect 30764 13098 30834 13418
<< locali >>
rect 30634 13946 30730 13980
rect 30868 13946 30964 13980
rect 30634 13884 30668 13946
rect 30930 13884 30964 13946
rect 30634 12570 30668 12632
rect 30930 12570 30964 12632
rect 30634 12536 30730 12570
rect 30868 12536 30964 12570
<< viali >>
rect 30780 13435 30818 13832
rect 30780 12684 30818 13081
<< metal1 >>
rect -1520 40090 -1280 40100
rect -1520 39910 -1510 40090
rect -1290 39910 -1280 40090
rect -1520 39900 -1280 39910
rect 20 40090 260 40100
rect 20 39910 30 40090
rect 250 39910 260 40090
rect 20 39900 260 39910
rect 26540 39190 26780 39200
rect 26540 39010 26550 39190
rect 26770 39010 26780 39190
rect 26540 39000 26780 39010
rect 28080 39190 28320 39200
rect 28080 39010 28090 39190
rect 28310 39010 28320 39190
rect 28080 39000 28320 39010
rect -4300 27250 -4100 27260
rect -4300 27030 -4290 27250
rect -4110 27030 -4100 27250
rect -4300 27020 -4100 27030
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect -4300 25710 -4100 25720
rect -4300 25490 -4290 25710
rect -4110 25490 -4100 25710
rect -4300 25480 -4100 25490
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect -4300 13900 -4100 13910
rect -4300 13420 -4290 13900
rect -4110 13420 -4100 13900
rect -4300 13410 -4100 13420
rect 30700 13900 30900 13910
rect 30700 13420 30710 13900
rect 30890 13420 30900 13900
rect 30700 13410 30900 13420
rect -4300 13090 -4100 13100
rect -4300 12610 -4290 13090
rect -4110 12610 -4100 13090
rect -4300 12600 -4100 12610
rect 30700 13090 30900 13100
rect 30700 12610 30710 13090
rect 30890 12610 30900 13090
rect 30700 12600 30900 12610
<< via1 >>
rect -1510 39910 -1290 40090
rect 30 39910 250 40090
rect 26550 39010 26770 39190
rect 28090 39010 28310 39190
rect -4290 27030 -4110 27250
rect 30910 27030 31090 27250
rect -4290 25490 -4110 25710
rect 30910 25490 31090 25710
rect -4290 13420 -4110 13900
rect 30710 13832 30890 13900
rect 30710 13435 30780 13832
rect 30780 13435 30818 13832
rect 30818 13435 30890 13832
rect 30710 13420 30890 13435
rect -4290 12610 -4110 13090
rect 30710 13081 30890 13090
rect 30710 12684 30780 13081
rect 30780 12684 30818 13081
rect 30818 12684 30890 13081
rect 30710 12610 30890 12684
<< metal2 >>
rect -1520 40090 -1280 40100
rect -1520 39910 -1510 40090
rect -1290 39910 -1280 40090
rect -1520 39900 -1280 39910
rect 20 40090 260 40100
rect 20 39910 30 40090
rect 250 39910 260 40090
rect 20 39900 260 39910
rect 26540 39190 26780 39200
rect 26540 39010 26550 39190
rect 26770 39010 26780 39190
rect 26540 39000 26780 39010
rect 28080 39190 28320 39200
rect 28080 39010 28090 39190
rect 28310 39010 28320 39190
rect 28080 39000 28320 39010
rect -4300 27250 -4100 27260
rect -4300 27030 -4290 27250
rect -4110 27030 -4100 27250
rect -4300 27020 -4100 27030
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect -4300 25710 -4100 25720
rect -4300 25490 -4290 25710
rect -4110 25490 -4100 25710
rect -4300 25480 -4100 25490
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect -4300 13900 -4100 13910
rect -4300 13420 -4290 13900
rect -4110 13420 -4100 13900
rect -4300 13410 -4100 13420
rect 30700 13900 30900 13910
rect 30700 13420 30710 13900
rect 30890 13420 30900 13900
rect 30700 13410 30900 13420
rect -4300 13090 -4100 13100
rect -4300 12610 -4290 13090
rect -4110 12610 -4100 13090
rect -4300 12600 -4100 12610
rect 30700 13090 30900 13100
rect 30700 12610 30710 13090
rect 30890 12610 30900 13090
rect 30700 12600 30900 12610
<< via2 >>
rect -1510 39910 -1290 40090
rect 30 39910 250 40090
rect 26550 39010 26770 39190
rect 28090 39010 28310 39190
rect -4290 27030 -4110 27250
rect 30910 27030 31090 27250
rect -4290 25490 -4110 25710
rect 30910 25490 31090 25710
rect -4290 13420 -4110 13900
rect 30710 13420 30890 13900
rect -4290 12610 -4110 13090
rect 30710 12610 30890 13090
<< metal3 >>
rect -1520 40190 -1280 40200
rect -1520 39810 -1510 40190
rect -1290 39810 -1280 40190
rect -1520 39800 -1280 39810
rect 0 40180 300 40200
rect 0 39820 20 40180
rect 280 39820 300 40180
rect 0 39800 300 39820
rect 26500 39280 26800 39300
rect 26500 38920 26520 39280
rect 26780 38920 26800 39280
rect 26500 38900 26800 38920
rect 28080 39290 28320 39300
rect 28080 38910 28090 39290
rect 28310 38910 28320 39290
rect 28080 38900 28320 38910
rect -4400 31700 2800 31800
rect -4400 31100 1400 31700
rect 2700 31100 2800 31700
rect -4400 31000 2800 31100
rect 24000 31700 31200 31800
rect 24000 31100 24100 31700
rect 25400 31100 31200 31700
rect 24000 31000 31200 31100
rect -4400 27250 -3900 31000
rect -4400 27030 -4290 27250
rect -4110 27030 -3900 27250
rect -4400 27000 -3900 27030
rect 30700 27250 31200 31000
rect 30700 27030 30910 27250
rect 31090 27030 31200 27250
rect 30700 27000 31200 27030
rect -4400 25710 -4000 25720
rect -4400 25490 -4390 25710
rect -4010 25490 -4000 25710
rect -4400 25480 -4000 25490
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25480 31200 25490
rect -4400 14000 -4000 14010
rect -4400 13420 -4390 14000
rect -4010 13420 -4000 14000
rect -4400 13410 -4000 13420
rect 30600 14000 31000 14010
rect 30600 13420 30610 14000
rect 30990 13420 31000 14000
rect 30600 13410 31000 13420
rect -4400 13090 -4000 13100
rect -4400 12510 -4390 13090
rect -4010 12510 -4000 13090
rect -4400 12500 -4000 12510
rect 30600 13090 31000 13100
rect 30600 12510 30610 13090
rect 30990 12510 31000 13090
rect 30600 12500 31000 12510
<< via3 >>
rect -1510 40090 -1290 40190
rect -1510 39910 -1290 40090
rect -1510 39810 -1290 39910
rect 20 40090 280 40180
rect 20 39910 30 40090
rect 30 39910 250 40090
rect 250 39910 280 40090
rect 20 39820 280 39910
rect 26520 39190 26780 39280
rect 26520 39010 26550 39190
rect 26550 39010 26770 39190
rect 26770 39010 26780 39190
rect 26520 38920 26780 39010
rect 28090 39190 28310 39290
rect 28090 39010 28310 39190
rect 28090 38910 28310 39010
rect 1400 31100 2700 31700
rect 24100 31100 25400 31700
rect -4390 25490 -4290 25710
rect -4290 25490 -4110 25710
rect -4110 25490 -4010 25710
rect 30810 25490 30910 25710
rect 30910 25490 31090 25710
rect 31090 25490 31190 25710
rect -4390 13900 -4010 14000
rect -4390 13420 -4290 13900
rect -4290 13420 -4110 13900
rect -4110 13420 -4010 13900
rect 30610 13900 30990 14000
rect 30610 13420 30710 13900
rect 30710 13420 30890 13900
rect 30890 13420 30990 13900
rect -4390 12610 -4290 13090
rect -4290 12610 -4110 13090
rect -4110 12610 -4010 13090
rect -4390 12510 -4010 12610
rect 30610 12610 30710 13090
rect 30710 12610 30890 13090
rect 30890 12610 30990 13090
rect 30610 12510 30990 12610
<< metal4 >>
rect -600 47500 800 47600
rect -600 46500 -500 47500
rect 700 46500 800 47500
rect -600 46400 800 46500
rect -1000 46000 800 46400
rect -3400 40800 800 46000
rect -1580 40190 -1280 40200
rect -1580 40170 -1510 40190
rect -1580 39830 -1550 40170
rect -1580 39810 -1510 39830
rect -1290 39810 -1280 40190
rect -1580 39800 -1280 39810
rect -1000 40180 800 40800
rect -1000 39820 20 40180
rect 280 39820 800 40180
rect -1000 39100 800 39820
rect -3400 38600 -1600 38700
rect -3400 37600 -2900 38600
rect -1700 37600 -1600 38600
rect -4400 25710 -4000 25720
rect -4400 25490 -4390 25710
rect -4010 25490 -4000 25710
rect -4400 25450 -4370 25490
rect -4030 25450 -4000 25490
rect -4400 25430 -4000 25450
rect -3400 24900 -1600 37600
rect -6100 14300 -1600 24900
rect -4400 14000 -4000 14010
rect -4400 13420 -4390 14000
rect -4010 13420 -4000 14000
rect -4400 13410 -4000 13420
rect -3400 13800 -1600 14300
rect -3400 13100 -3300 13800
rect -4400 13090 -3300 13100
rect -4400 12510 -4390 13090
rect -4010 12600 -3300 13090
rect -1700 12600 -1600 13800
rect -4010 12510 -1600 12600
rect -4400 12500 -1600 12510
rect -1000 25500 -600 39100
rect 700 25500 800 39100
rect 26000 47500 27400 47600
rect 26000 46500 26100 47500
rect 27300 46500 27400 47500
rect 26000 46400 27400 46500
rect 26000 46000 27800 46400
rect 26000 40800 30200 46000
rect 26000 39280 27800 40800
rect 26000 38920 26520 39280
rect 26780 38920 27800 39280
rect 26000 38200 27800 38920
rect 28080 39290 28380 39300
rect 28080 38910 28090 39290
rect 28310 39270 28380 39290
rect 28350 38930 28380 39270
rect 28310 38910 28380 38930
rect 28080 38900 28380 38910
rect -1000 23200 800 25500
rect -1000 18500 -600 23200
rect 700 18500 800 23200
rect -1000 12100 800 18500
rect -1000 8000 -600 12100
rect 700 10100 800 12100
rect 200 10000 800 10100
rect 26000 25500 26100 38200
rect 27400 25500 27800 38200
rect 26000 23200 27800 25500
rect 26000 16300 26100 23200
rect 27400 16300 27800 23200
rect 26000 11900 27800 16300
rect 28400 38600 30200 38700
rect 28400 37600 28500 38600
rect 29700 37600 30200 38600
rect 28400 24900 30200 37600
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25450 30830 25490
rect 31170 25450 31200 25490
rect 30800 25430 31200 25450
rect 28400 14300 32900 24900
rect 28400 13700 30200 14300
rect 28400 12600 28500 13700
rect 30100 13100 30200 13700
rect 30600 14000 31000 14010
rect 30600 13420 30610 14000
rect 30990 13420 31000 14000
rect 30600 13410 31000 13420
rect 30100 13090 31000 13100
rect 30100 12600 30610 13090
rect 28400 12510 30610 12600
rect 30990 12510 31000 13090
rect 28400 12500 31000 12510
rect 200 8000 300 10000
rect 26000 9200 26100 11900
rect 26000 9100 26600 9200
rect -1000 7900 300 8000
rect 26500 8000 26600 9100
rect 27400 8000 27800 11900
rect 26500 7900 27800 8000
rect -1000 7400 800 7900
rect -3400 2200 800 7400
rect 26000 7400 27800 7900
rect 26000 2200 30200 7400
<< via4 >>
rect -500 46500 700 47500
rect -1550 39830 -1510 40170
rect -1510 39830 -1310 40170
rect -2900 37600 -1700 38600
rect -4370 25490 -4030 25690
rect -4370 25450 -4030 25490
rect -4370 13440 -4030 13980
rect -3300 12600 -1700 13800
rect -600 25500 700 39100
rect 26100 46500 27300 47500
rect 28110 38930 28310 39270
rect 28310 38930 28350 39270
rect -600 18500 700 23200
rect -600 10100 700 12100
rect -600 8000 200 10100
rect 26100 25500 27400 38200
rect 26100 16300 27400 23200
rect 28500 37600 29700 38600
rect 30830 25490 31170 25690
rect 30830 25450 31170 25490
rect 28500 12600 30100 13700
rect 30630 13440 30970 13980
rect 26100 9200 27400 11900
rect 26600 8000 27400 9200
<< mimcap2 >>
rect -3300 45800 700 45900
rect -3300 41000 -3200 45800
rect 600 41000 700 45800
rect -3300 40900 700 41000
rect 26100 45800 30100 45900
rect 26100 41000 26200 45800
rect 30000 41000 30100 45800
rect 26100 40900 30100 41000
rect -3300 36900 -1700 37000
rect -3300 26700 -3200 36900
rect -1800 26700 -1700 36900
rect -3300 26600 -1700 26700
rect 28500 36900 30100 37000
rect 28500 26700 28600 36900
rect 30000 26700 30100 36900
rect 28500 26600 30100 26700
rect -6000 24700 -1700 24800
rect -6000 14500 -5900 24700
rect -1800 14500 -1700 24700
rect -6000 14400 -1700 14500
rect 28500 24700 32800 24800
rect 28500 14500 28600 24700
rect 32700 14500 32800 24700
rect 28500 14400 32800 14500
rect -3300 7200 700 7300
rect -3300 2400 -3200 7200
rect 600 2400 700 7200
rect -3300 2300 700 2400
rect 26100 7200 30100 7300
rect 26100 2400 26200 7200
rect 30000 2400 30100 7200
rect 26100 2300 30100 2400
<< mimcap2contact >>
rect -3200 41000 600 45800
rect 26200 41000 30000 45800
rect -3200 26700 -1800 36900
rect 28600 26700 30000 36900
rect -5900 14500 -1800 24700
rect 28600 14500 32700 24700
rect -3200 2400 600 7200
rect 26200 2400 30000 7200
<< metal5 >>
rect 1300 48100 2800 48500
rect 24000 48100 25500 48500
rect -600 47500 1300 47600
rect -600 46500 -500 47500
rect 700 46700 1300 47500
rect 25500 47500 27400 47600
rect 25500 46700 26100 47500
rect 700 46500 800 46700
rect -600 46400 800 46500
rect 26000 46500 26100 46700
rect 27300 46500 27400 47500
rect 26000 46400 27400 46500
rect -3400 45800 800 46000
rect -3400 41000 -3200 45800
rect 600 41000 800 45800
rect -3400 40800 800 41000
rect 26000 45800 30200 46000
rect 26000 41000 26200 45800
rect 30000 41000 30200 45800
rect 26000 40800 30200 41000
rect -3000 40170 1200 40200
rect -3000 39830 -1550 40170
rect -1310 39830 1200 40170
rect -3000 39700 1200 39830
rect -3000 38600 -1600 39700
rect 25400 39270 29800 39300
rect -3000 37600 -2900 38600
rect -1700 37600 -1600 38600
rect -3000 37500 -1600 37600
rect -700 39100 800 39200
rect -3400 36900 -1600 37100
rect -3400 26700 -3200 36900
rect -1800 26700 -1600 36900
rect -3400 26500 -1600 26700
rect -4400 25690 -4000 25720
rect -4400 25450 -4370 25690
rect -4030 25450 -4000 25690
rect -4400 24900 -4000 25450
rect -700 25500 -600 39100
rect 700 25500 800 39100
rect 25400 38930 28110 39270
rect 28350 38930 29800 39270
rect 25400 38800 29800 38930
rect 28400 38600 29800 38800
rect -700 25400 800 25500
rect 26000 38200 27500 38300
rect 26000 25500 26100 38200
rect 27400 25500 27500 38200
rect 28400 37600 28500 38600
rect 29700 37600 29800 38600
rect 28400 37500 29800 37600
rect 28400 36900 30200 37100
rect 28400 26700 28600 36900
rect 30000 26700 30200 36900
rect 28400 26500 30200 26700
rect 26000 25400 27500 25500
rect 30800 25690 31200 25720
rect 30800 25450 30830 25690
rect 31170 25450 31200 25690
rect 30800 24900 31200 25450
rect -6100 24700 1200 24900
rect 25400 24700 32900 24900
rect -6100 14500 -5900 24700
rect -1800 24000 2100 24700
rect 25400 24600 28600 24700
rect -1800 23800 1200 24000
rect 24500 23900 28600 24600
rect 25400 23800 28600 23900
rect -1800 14500 -1600 23800
rect 25400 23500 25600 23800
rect -700 23200 800 23300
rect -700 18500 -600 23200
rect 700 18500 800 23200
rect -700 18400 800 18500
rect 26000 23200 27500 23300
rect -6100 14300 -1600 14500
rect -1200 16500 1300 17900
rect -4400 13980 -4000 14300
rect -4400 13440 -4370 13980
rect -4030 13440 -4000 13980
rect -1200 13900 0 16500
rect 26000 16300 26100 23200
rect 27400 16300 27500 23200
rect 26000 16200 27500 16300
rect 25500 14300 28000 15700
rect 28400 14500 28600 23800
rect 32700 14500 32900 24700
rect 28400 14300 32900 14500
rect -4400 13410 -4000 13440
rect -3400 13800 0 13900
rect -3400 12600 -3300 13800
rect -1700 12600 0 13800
rect 26800 13800 28000 14300
rect 30600 13980 31000 14300
rect 26800 13700 30200 13800
rect 26800 12600 28500 13700
rect 30100 12600 30200 13700
rect 30600 13440 30630 13980
rect 30970 13440 31000 13980
rect 30600 13410 31000 13440
rect -3400 7400 -1600 12600
rect 26800 12500 30200 12600
rect -700 12100 800 12200
rect -700 8000 -600 12100
rect 700 10100 800 12100
rect 200 10000 800 10100
rect 26000 11900 27500 12000
rect 200 8000 300 10000
rect 700 9100 1200 9600
rect 26000 9200 26100 11900
rect 26000 9100 26600 9200
rect 25400 8200 26100 8700
rect -700 7900 300 8000
rect 26500 8000 26600 9100
rect 27400 8000 27500 11900
rect 26500 7900 27500 8000
rect 28400 7400 30200 12500
rect -3400 7200 800 7400
rect -3400 2400 -3200 7200
rect 600 3600 800 7200
rect 26000 7200 30200 7400
rect 26000 3600 26200 7200
rect 600 2400 1400 3600
rect -3400 2200 1400 2400
rect 24000 2400 26200 3600
rect 30000 2400 30200 7200
rect 24000 2200 30200 2400
rect 24000 1700 25500 2200
rect 1300 0 2800 400
rect 24000 0 25500 400
use cascode_1  cascode_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/CLASSE
timestamp 1664506494
transform 1 0 14700 0 1 -3700
box -14700 3700 10800 52200
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_0
timestamp 1664814488
transform -1 0 31001 0 1 26369
box -199 -889 199 889
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_1
timestamp 1664814488
transform 1 0 -4201 0 1 26369
box -199 -889 199 889
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_3
timestamp 1664814488
transform 0 1 -631 -1 0 40001
box -199 -889 199 889
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_4
timestamp 1664814488
transform 0 -1 27431 -1 0 39101
box -199 -889 199 889
use sky130_fd_pr__res_high_po_0p35_FFWWQH  sky130_fd_pr__res_high_po_0p35_FFWWQH_0
timestamp 1664805031
transform 1 0 -4199 0 1 13258
box -201 -758 201 758
use sky130_fd_pr__res_high_po_0p35_FFWWQH  sky130_fd_pr__res_high_po_0p35_FFWWQH_1
timestamp 1664805031
transform -1 0 30799 0 1 13258
box -201 -758 201 758
<< labels >>
rlabel metal5 25800 8200 26100 8700 1 VINP
rlabel metal5 700 9100 1000 9600 1 VINN
rlabel metal5 1300 0 2800 400 1 VSS
rlabel metal5 24000 0 25500 400 1 VSSH
rlabel metal5 1300 48100 2800 48500 1 VDN
rlabel metal5 24000 48100 25500 48500 1 VDP
rlabel metal5 900 39700 1200 40200 1 VGN
rlabel metal5 25600 38800 25900 39300 1 VGP
rlabel metal5 800 24400 1100 24900 1 N2
rlabel metal5 900 16500 1200 17900 1 N
rlabel metal5 25600 14300 25900 15700 1 P
<< end >>
