magic
tech sky130B
magscale 1 2
timestamp 1660448881
<< error_p >>
rect -29 13339 29 13345
rect -29 13305 -17 13339
rect -29 13299 29 13305
rect -29 13029 29 13035
rect -29 12995 -17 13029
rect -29 12989 29 12995
rect -29 12921 29 12927
rect -29 12887 -17 12921
rect -29 12881 29 12887
rect -29 12611 29 12617
rect -29 12577 -17 12611
rect -29 12571 29 12577
rect -29 12503 29 12509
rect -29 12469 -17 12503
rect -29 12463 29 12469
rect -29 12193 29 12199
rect -29 12159 -17 12193
rect -29 12153 29 12159
rect -29 12085 29 12091
rect -29 12051 -17 12085
rect -29 12045 29 12051
rect -29 11775 29 11781
rect -29 11741 -17 11775
rect -29 11735 29 11741
rect -29 11667 29 11673
rect -29 11633 -17 11667
rect -29 11627 29 11633
rect -29 11357 29 11363
rect -29 11323 -17 11357
rect -29 11317 29 11323
rect -29 11249 29 11255
rect -29 11215 -17 11249
rect -29 11209 29 11215
rect -29 10939 29 10945
rect -29 10905 -17 10939
rect -29 10899 29 10905
rect -29 10831 29 10837
rect -29 10797 -17 10831
rect -29 10791 29 10797
rect -29 10521 29 10527
rect -29 10487 -17 10521
rect -29 10481 29 10487
rect -29 10413 29 10419
rect -29 10379 -17 10413
rect -29 10373 29 10379
rect -29 10103 29 10109
rect -29 10069 -17 10103
rect -29 10063 29 10069
rect -29 9995 29 10001
rect -29 9961 -17 9995
rect -29 9955 29 9961
rect -29 9685 29 9691
rect -29 9651 -17 9685
rect -29 9645 29 9651
rect -29 9577 29 9583
rect -29 9543 -17 9577
rect -29 9537 29 9543
rect -29 9267 29 9273
rect -29 9233 -17 9267
rect -29 9227 29 9233
rect -29 9159 29 9165
rect -29 9125 -17 9159
rect -29 9119 29 9125
rect -29 8849 29 8855
rect -29 8815 -17 8849
rect -29 8809 29 8815
rect -29 8741 29 8747
rect -29 8707 -17 8741
rect -29 8701 29 8707
rect -29 8431 29 8437
rect -29 8397 -17 8431
rect -29 8391 29 8397
rect -29 8323 29 8329
rect -29 8289 -17 8323
rect -29 8283 29 8289
rect -29 8013 29 8019
rect -29 7979 -17 8013
rect -29 7973 29 7979
rect -29 7905 29 7911
rect -29 7871 -17 7905
rect -29 7865 29 7871
rect -29 7595 29 7601
rect -29 7561 -17 7595
rect -29 7555 29 7561
rect -29 7487 29 7493
rect -29 7453 -17 7487
rect -29 7447 29 7453
rect -29 7177 29 7183
rect -29 7143 -17 7177
rect -29 7137 29 7143
rect -29 7069 29 7075
rect -29 7035 -17 7069
rect -29 7029 29 7035
rect -29 6759 29 6765
rect -29 6725 -17 6759
rect -29 6719 29 6725
rect -29 6651 29 6657
rect -29 6617 -17 6651
rect -29 6611 29 6617
rect -29 6341 29 6347
rect -29 6307 -17 6341
rect -29 6301 29 6307
rect -29 6233 29 6239
rect -29 6199 -17 6233
rect -29 6193 29 6199
rect -29 5923 29 5929
rect -29 5889 -17 5923
rect -29 5883 29 5889
rect -29 5815 29 5821
rect -29 5781 -17 5815
rect -29 5775 29 5781
rect -29 5505 29 5511
rect -29 5471 -17 5505
rect -29 5465 29 5471
rect -29 5397 29 5403
rect -29 5363 -17 5397
rect -29 5357 29 5363
rect -29 5087 29 5093
rect -29 5053 -17 5087
rect -29 5047 29 5053
rect -29 4979 29 4985
rect -29 4945 -17 4979
rect -29 4939 29 4945
rect -29 4669 29 4675
rect -29 4635 -17 4669
rect -29 4629 29 4635
rect -29 4561 29 4567
rect -29 4527 -17 4561
rect -29 4521 29 4527
rect -29 4251 29 4257
rect -29 4217 -17 4251
rect -29 4211 29 4217
rect -29 4143 29 4149
rect -29 4109 -17 4143
rect -29 4103 29 4109
rect -29 3833 29 3839
rect -29 3799 -17 3833
rect -29 3793 29 3799
rect -29 3725 29 3731
rect -29 3691 -17 3725
rect -29 3685 29 3691
rect -29 3415 29 3421
rect -29 3381 -17 3415
rect -29 3375 29 3381
rect -29 3307 29 3313
rect -29 3273 -17 3307
rect -29 3267 29 3273
rect -29 2997 29 3003
rect -29 2963 -17 2997
rect -29 2957 29 2963
rect -29 2889 29 2895
rect -29 2855 -17 2889
rect -29 2849 29 2855
rect -29 2579 29 2585
rect -29 2545 -17 2579
rect -29 2539 29 2545
rect -29 2471 29 2477
rect -29 2437 -17 2471
rect -29 2431 29 2437
rect -29 2161 29 2167
rect -29 2127 -17 2161
rect -29 2121 29 2127
rect -29 2053 29 2059
rect -29 2019 -17 2053
rect -29 2013 29 2019
rect -29 1743 29 1749
rect -29 1709 -17 1743
rect -29 1703 29 1709
rect -29 1635 29 1641
rect -29 1601 -17 1635
rect -29 1595 29 1601
rect -29 1325 29 1331
rect -29 1291 -17 1325
rect -29 1285 29 1291
rect -29 1217 29 1223
rect -29 1183 -17 1217
rect -29 1177 29 1183
rect -29 907 29 913
rect -29 873 -17 907
rect -29 867 29 873
rect -29 799 29 805
rect -29 765 -17 799
rect -29 759 29 765
rect -29 489 29 495
rect -29 455 -17 489
rect -29 449 29 455
rect -29 381 29 387
rect -29 347 -17 381
rect -29 341 29 347
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect -29 -387 29 -381
rect -29 -455 29 -449
rect -29 -489 -17 -455
rect -29 -495 29 -489
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect -29 -805 29 -799
rect -29 -873 29 -867
rect -29 -907 -17 -873
rect -29 -913 29 -907
rect -29 -1183 29 -1177
rect -29 -1217 -17 -1183
rect -29 -1223 29 -1217
rect -29 -1291 29 -1285
rect -29 -1325 -17 -1291
rect -29 -1331 29 -1325
rect -29 -1601 29 -1595
rect -29 -1635 -17 -1601
rect -29 -1641 29 -1635
rect -29 -1709 29 -1703
rect -29 -1743 -17 -1709
rect -29 -1749 29 -1743
rect -29 -2019 29 -2013
rect -29 -2053 -17 -2019
rect -29 -2059 29 -2053
rect -29 -2127 29 -2121
rect -29 -2161 -17 -2127
rect -29 -2167 29 -2161
rect -29 -2437 29 -2431
rect -29 -2471 -17 -2437
rect -29 -2477 29 -2471
rect -29 -2545 29 -2539
rect -29 -2579 -17 -2545
rect -29 -2585 29 -2579
rect -29 -2855 29 -2849
rect -29 -2889 -17 -2855
rect -29 -2895 29 -2889
rect -29 -2963 29 -2957
rect -29 -2997 -17 -2963
rect -29 -3003 29 -2997
rect -29 -3273 29 -3267
rect -29 -3307 -17 -3273
rect -29 -3313 29 -3307
rect -29 -3381 29 -3375
rect -29 -3415 -17 -3381
rect -29 -3421 29 -3415
rect -29 -3691 29 -3685
rect -29 -3725 -17 -3691
rect -29 -3731 29 -3725
rect -29 -3799 29 -3793
rect -29 -3833 -17 -3799
rect -29 -3839 29 -3833
rect -29 -4109 29 -4103
rect -29 -4143 -17 -4109
rect -29 -4149 29 -4143
rect -29 -4217 29 -4211
rect -29 -4251 -17 -4217
rect -29 -4257 29 -4251
rect -29 -4527 29 -4521
rect -29 -4561 -17 -4527
rect -29 -4567 29 -4561
rect -29 -4635 29 -4629
rect -29 -4669 -17 -4635
rect -29 -4675 29 -4669
rect -29 -4945 29 -4939
rect -29 -4979 -17 -4945
rect -29 -4985 29 -4979
rect -29 -5053 29 -5047
rect -29 -5087 -17 -5053
rect -29 -5093 29 -5087
rect -29 -5363 29 -5357
rect -29 -5397 -17 -5363
rect -29 -5403 29 -5397
rect -29 -5471 29 -5465
rect -29 -5505 -17 -5471
rect -29 -5511 29 -5505
rect -29 -5781 29 -5775
rect -29 -5815 -17 -5781
rect -29 -5821 29 -5815
rect -29 -5889 29 -5883
rect -29 -5923 -17 -5889
rect -29 -5929 29 -5923
rect -29 -6199 29 -6193
rect -29 -6233 -17 -6199
rect -29 -6239 29 -6233
rect -29 -6307 29 -6301
rect -29 -6341 -17 -6307
rect -29 -6347 29 -6341
rect -29 -6617 29 -6611
rect -29 -6651 -17 -6617
rect -29 -6657 29 -6651
rect -29 -6725 29 -6719
rect -29 -6759 -17 -6725
rect -29 -6765 29 -6759
rect -29 -7035 29 -7029
rect -29 -7069 -17 -7035
rect -29 -7075 29 -7069
rect -29 -7143 29 -7137
rect -29 -7177 -17 -7143
rect -29 -7183 29 -7177
rect -29 -7453 29 -7447
rect -29 -7487 -17 -7453
rect -29 -7493 29 -7487
rect -29 -7561 29 -7555
rect -29 -7595 -17 -7561
rect -29 -7601 29 -7595
rect -29 -7871 29 -7865
rect -29 -7905 -17 -7871
rect -29 -7911 29 -7905
rect -29 -7979 29 -7973
rect -29 -8013 -17 -7979
rect -29 -8019 29 -8013
rect -29 -8289 29 -8283
rect -29 -8323 -17 -8289
rect -29 -8329 29 -8323
rect -29 -8397 29 -8391
rect -29 -8431 -17 -8397
rect -29 -8437 29 -8431
rect -29 -8707 29 -8701
rect -29 -8741 -17 -8707
rect -29 -8747 29 -8741
rect -29 -8815 29 -8809
rect -29 -8849 -17 -8815
rect -29 -8855 29 -8849
rect -29 -9125 29 -9119
rect -29 -9159 -17 -9125
rect -29 -9165 29 -9159
rect -29 -9233 29 -9227
rect -29 -9267 -17 -9233
rect -29 -9273 29 -9267
rect -29 -9543 29 -9537
rect -29 -9577 -17 -9543
rect -29 -9583 29 -9577
rect -29 -9651 29 -9645
rect -29 -9685 -17 -9651
rect -29 -9691 29 -9685
rect -29 -9961 29 -9955
rect -29 -9995 -17 -9961
rect -29 -10001 29 -9995
rect -29 -10069 29 -10063
rect -29 -10103 -17 -10069
rect -29 -10109 29 -10103
rect -29 -10379 29 -10373
rect -29 -10413 -17 -10379
rect -29 -10419 29 -10413
rect -29 -10487 29 -10481
rect -29 -10521 -17 -10487
rect -29 -10527 29 -10521
rect -29 -10797 29 -10791
rect -29 -10831 -17 -10797
rect -29 -10837 29 -10831
rect -29 -10905 29 -10899
rect -29 -10939 -17 -10905
rect -29 -10945 29 -10939
rect -29 -11215 29 -11209
rect -29 -11249 -17 -11215
rect -29 -11255 29 -11249
rect -29 -11323 29 -11317
rect -29 -11357 -17 -11323
rect -29 -11363 29 -11357
rect -29 -11633 29 -11627
rect -29 -11667 -17 -11633
rect -29 -11673 29 -11667
rect -29 -11741 29 -11735
rect -29 -11775 -17 -11741
rect -29 -11781 29 -11775
rect -29 -12051 29 -12045
rect -29 -12085 -17 -12051
rect -29 -12091 29 -12085
rect -29 -12159 29 -12153
rect -29 -12193 -17 -12159
rect -29 -12199 29 -12193
rect -29 -12469 29 -12463
rect -29 -12503 -17 -12469
rect -29 -12509 29 -12503
rect -29 -12577 29 -12571
rect -29 -12611 -17 -12577
rect -29 -12617 29 -12611
rect -29 -12887 29 -12881
rect -29 -12921 -17 -12887
rect -29 -12927 29 -12921
rect -29 -12995 29 -12989
rect -29 -13029 -17 -12995
rect -29 -13035 29 -13029
rect -29 -13305 29 -13299
rect -29 -13339 -17 -13305
rect -29 -13345 29 -13339
<< pwell >>
rect -211 -13477 211 13477
<< nmos >>
rect -15 13067 15 13267
rect -15 12649 15 12849
rect -15 12231 15 12431
rect -15 11813 15 12013
rect -15 11395 15 11595
rect -15 10977 15 11177
rect -15 10559 15 10759
rect -15 10141 15 10341
rect -15 9723 15 9923
rect -15 9305 15 9505
rect -15 8887 15 9087
rect -15 8469 15 8669
rect -15 8051 15 8251
rect -15 7633 15 7833
rect -15 7215 15 7415
rect -15 6797 15 6997
rect -15 6379 15 6579
rect -15 5961 15 6161
rect -15 5543 15 5743
rect -15 5125 15 5325
rect -15 4707 15 4907
rect -15 4289 15 4489
rect -15 3871 15 4071
rect -15 3453 15 3653
rect -15 3035 15 3235
rect -15 2617 15 2817
rect -15 2199 15 2399
rect -15 1781 15 1981
rect -15 1363 15 1563
rect -15 945 15 1145
rect -15 527 15 727
rect -15 109 15 309
rect -15 -309 15 -109
rect -15 -727 15 -527
rect -15 -1145 15 -945
rect -15 -1563 15 -1363
rect -15 -1981 15 -1781
rect -15 -2399 15 -2199
rect -15 -2817 15 -2617
rect -15 -3235 15 -3035
rect -15 -3653 15 -3453
rect -15 -4071 15 -3871
rect -15 -4489 15 -4289
rect -15 -4907 15 -4707
rect -15 -5325 15 -5125
rect -15 -5743 15 -5543
rect -15 -6161 15 -5961
rect -15 -6579 15 -6379
rect -15 -6997 15 -6797
rect -15 -7415 15 -7215
rect -15 -7833 15 -7633
rect -15 -8251 15 -8051
rect -15 -8669 15 -8469
rect -15 -9087 15 -8887
rect -15 -9505 15 -9305
rect -15 -9923 15 -9723
rect -15 -10341 15 -10141
rect -15 -10759 15 -10559
rect -15 -11177 15 -10977
rect -15 -11595 15 -11395
rect -15 -12013 15 -11813
rect -15 -12431 15 -12231
rect -15 -12849 15 -12649
rect -15 -13267 15 -13067
<< ndiff >>
rect -73 13255 -15 13267
rect -73 13079 -61 13255
rect -27 13079 -15 13255
rect -73 13067 -15 13079
rect 15 13255 73 13267
rect 15 13079 27 13255
rect 61 13079 73 13255
rect 15 13067 73 13079
rect -73 12837 -15 12849
rect -73 12661 -61 12837
rect -27 12661 -15 12837
rect -73 12649 -15 12661
rect 15 12837 73 12849
rect 15 12661 27 12837
rect 61 12661 73 12837
rect 15 12649 73 12661
rect -73 12419 -15 12431
rect -73 12243 -61 12419
rect -27 12243 -15 12419
rect -73 12231 -15 12243
rect 15 12419 73 12431
rect 15 12243 27 12419
rect 61 12243 73 12419
rect 15 12231 73 12243
rect -73 12001 -15 12013
rect -73 11825 -61 12001
rect -27 11825 -15 12001
rect -73 11813 -15 11825
rect 15 12001 73 12013
rect 15 11825 27 12001
rect 61 11825 73 12001
rect 15 11813 73 11825
rect -73 11583 -15 11595
rect -73 11407 -61 11583
rect -27 11407 -15 11583
rect -73 11395 -15 11407
rect 15 11583 73 11595
rect 15 11407 27 11583
rect 61 11407 73 11583
rect 15 11395 73 11407
rect -73 11165 -15 11177
rect -73 10989 -61 11165
rect -27 10989 -15 11165
rect -73 10977 -15 10989
rect 15 11165 73 11177
rect 15 10989 27 11165
rect 61 10989 73 11165
rect 15 10977 73 10989
rect -73 10747 -15 10759
rect -73 10571 -61 10747
rect -27 10571 -15 10747
rect -73 10559 -15 10571
rect 15 10747 73 10759
rect 15 10571 27 10747
rect 61 10571 73 10747
rect 15 10559 73 10571
rect -73 10329 -15 10341
rect -73 10153 -61 10329
rect -27 10153 -15 10329
rect -73 10141 -15 10153
rect 15 10329 73 10341
rect 15 10153 27 10329
rect 61 10153 73 10329
rect 15 10141 73 10153
rect -73 9911 -15 9923
rect -73 9735 -61 9911
rect -27 9735 -15 9911
rect -73 9723 -15 9735
rect 15 9911 73 9923
rect 15 9735 27 9911
rect 61 9735 73 9911
rect 15 9723 73 9735
rect -73 9493 -15 9505
rect -73 9317 -61 9493
rect -27 9317 -15 9493
rect -73 9305 -15 9317
rect 15 9493 73 9505
rect 15 9317 27 9493
rect 61 9317 73 9493
rect 15 9305 73 9317
rect -73 9075 -15 9087
rect -73 8899 -61 9075
rect -27 8899 -15 9075
rect -73 8887 -15 8899
rect 15 9075 73 9087
rect 15 8899 27 9075
rect 61 8899 73 9075
rect 15 8887 73 8899
rect -73 8657 -15 8669
rect -73 8481 -61 8657
rect -27 8481 -15 8657
rect -73 8469 -15 8481
rect 15 8657 73 8669
rect 15 8481 27 8657
rect 61 8481 73 8657
rect 15 8469 73 8481
rect -73 8239 -15 8251
rect -73 8063 -61 8239
rect -27 8063 -15 8239
rect -73 8051 -15 8063
rect 15 8239 73 8251
rect 15 8063 27 8239
rect 61 8063 73 8239
rect 15 8051 73 8063
rect -73 7821 -15 7833
rect -73 7645 -61 7821
rect -27 7645 -15 7821
rect -73 7633 -15 7645
rect 15 7821 73 7833
rect 15 7645 27 7821
rect 61 7645 73 7821
rect 15 7633 73 7645
rect -73 7403 -15 7415
rect -73 7227 -61 7403
rect -27 7227 -15 7403
rect -73 7215 -15 7227
rect 15 7403 73 7415
rect 15 7227 27 7403
rect 61 7227 73 7403
rect 15 7215 73 7227
rect -73 6985 -15 6997
rect -73 6809 -61 6985
rect -27 6809 -15 6985
rect -73 6797 -15 6809
rect 15 6985 73 6997
rect 15 6809 27 6985
rect 61 6809 73 6985
rect 15 6797 73 6809
rect -73 6567 -15 6579
rect -73 6391 -61 6567
rect -27 6391 -15 6567
rect -73 6379 -15 6391
rect 15 6567 73 6579
rect 15 6391 27 6567
rect 61 6391 73 6567
rect 15 6379 73 6391
rect -73 6149 -15 6161
rect -73 5973 -61 6149
rect -27 5973 -15 6149
rect -73 5961 -15 5973
rect 15 6149 73 6161
rect 15 5973 27 6149
rect 61 5973 73 6149
rect 15 5961 73 5973
rect -73 5731 -15 5743
rect -73 5555 -61 5731
rect -27 5555 -15 5731
rect -73 5543 -15 5555
rect 15 5731 73 5743
rect 15 5555 27 5731
rect 61 5555 73 5731
rect 15 5543 73 5555
rect -73 5313 -15 5325
rect -73 5137 -61 5313
rect -27 5137 -15 5313
rect -73 5125 -15 5137
rect 15 5313 73 5325
rect 15 5137 27 5313
rect 61 5137 73 5313
rect 15 5125 73 5137
rect -73 4895 -15 4907
rect -73 4719 -61 4895
rect -27 4719 -15 4895
rect -73 4707 -15 4719
rect 15 4895 73 4907
rect 15 4719 27 4895
rect 61 4719 73 4895
rect 15 4707 73 4719
rect -73 4477 -15 4489
rect -73 4301 -61 4477
rect -27 4301 -15 4477
rect -73 4289 -15 4301
rect 15 4477 73 4489
rect 15 4301 27 4477
rect 61 4301 73 4477
rect 15 4289 73 4301
rect -73 4059 -15 4071
rect -73 3883 -61 4059
rect -27 3883 -15 4059
rect -73 3871 -15 3883
rect 15 4059 73 4071
rect 15 3883 27 4059
rect 61 3883 73 4059
rect 15 3871 73 3883
rect -73 3641 -15 3653
rect -73 3465 -61 3641
rect -27 3465 -15 3641
rect -73 3453 -15 3465
rect 15 3641 73 3653
rect 15 3465 27 3641
rect 61 3465 73 3641
rect 15 3453 73 3465
rect -73 3223 -15 3235
rect -73 3047 -61 3223
rect -27 3047 -15 3223
rect -73 3035 -15 3047
rect 15 3223 73 3235
rect 15 3047 27 3223
rect 61 3047 73 3223
rect 15 3035 73 3047
rect -73 2805 -15 2817
rect -73 2629 -61 2805
rect -27 2629 -15 2805
rect -73 2617 -15 2629
rect 15 2805 73 2817
rect 15 2629 27 2805
rect 61 2629 73 2805
rect 15 2617 73 2629
rect -73 2387 -15 2399
rect -73 2211 -61 2387
rect -27 2211 -15 2387
rect -73 2199 -15 2211
rect 15 2387 73 2399
rect 15 2211 27 2387
rect 61 2211 73 2387
rect 15 2199 73 2211
rect -73 1969 -15 1981
rect -73 1793 -61 1969
rect -27 1793 -15 1969
rect -73 1781 -15 1793
rect 15 1969 73 1981
rect 15 1793 27 1969
rect 61 1793 73 1969
rect 15 1781 73 1793
rect -73 1551 -15 1563
rect -73 1375 -61 1551
rect -27 1375 -15 1551
rect -73 1363 -15 1375
rect 15 1551 73 1563
rect 15 1375 27 1551
rect 61 1375 73 1551
rect 15 1363 73 1375
rect -73 1133 -15 1145
rect -73 957 -61 1133
rect -27 957 -15 1133
rect -73 945 -15 957
rect 15 1133 73 1145
rect 15 957 27 1133
rect 61 957 73 1133
rect 15 945 73 957
rect -73 715 -15 727
rect -73 539 -61 715
rect -27 539 -15 715
rect -73 527 -15 539
rect 15 715 73 727
rect 15 539 27 715
rect 61 539 73 715
rect 15 527 73 539
rect -73 297 -15 309
rect -73 121 -61 297
rect -27 121 -15 297
rect -73 109 -15 121
rect 15 297 73 309
rect 15 121 27 297
rect 61 121 73 297
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -297 -61 -121
rect -27 -297 -15 -121
rect -73 -309 -15 -297
rect 15 -121 73 -109
rect 15 -297 27 -121
rect 61 -297 73 -121
rect 15 -309 73 -297
rect -73 -539 -15 -527
rect -73 -715 -61 -539
rect -27 -715 -15 -539
rect -73 -727 -15 -715
rect 15 -539 73 -527
rect 15 -715 27 -539
rect 61 -715 73 -539
rect 15 -727 73 -715
rect -73 -957 -15 -945
rect -73 -1133 -61 -957
rect -27 -1133 -15 -957
rect -73 -1145 -15 -1133
rect 15 -957 73 -945
rect 15 -1133 27 -957
rect 61 -1133 73 -957
rect 15 -1145 73 -1133
rect -73 -1375 -15 -1363
rect -73 -1551 -61 -1375
rect -27 -1551 -15 -1375
rect -73 -1563 -15 -1551
rect 15 -1375 73 -1363
rect 15 -1551 27 -1375
rect 61 -1551 73 -1375
rect 15 -1563 73 -1551
rect -73 -1793 -15 -1781
rect -73 -1969 -61 -1793
rect -27 -1969 -15 -1793
rect -73 -1981 -15 -1969
rect 15 -1793 73 -1781
rect 15 -1969 27 -1793
rect 61 -1969 73 -1793
rect 15 -1981 73 -1969
rect -73 -2211 -15 -2199
rect -73 -2387 -61 -2211
rect -27 -2387 -15 -2211
rect -73 -2399 -15 -2387
rect 15 -2211 73 -2199
rect 15 -2387 27 -2211
rect 61 -2387 73 -2211
rect 15 -2399 73 -2387
rect -73 -2629 -15 -2617
rect -73 -2805 -61 -2629
rect -27 -2805 -15 -2629
rect -73 -2817 -15 -2805
rect 15 -2629 73 -2617
rect 15 -2805 27 -2629
rect 61 -2805 73 -2629
rect 15 -2817 73 -2805
rect -73 -3047 -15 -3035
rect -73 -3223 -61 -3047
rect -27 -3223 -15 -3047
rect -73 -3235 -15 -3223
rect 15 -3047 73 -3035
rect 15 -3223 27 -3047
rect 61 -3223 73 -3047
rect 15 -3235 73 -3223
rect -73 -3465 -15 -3453
rect -73 -3641 -61 -3465
rect -27 -3641 -15 -3465
rect -73 -3653 -15 -3641
rect 15 -3465 73 -3453
rect 15 -3641 27 -3465
rect 61 -3641 73 -3465
rect 15 -3653 73 -3641
rect -73 -3883 -15 -3871
rect -73 -4059 -61 -3883
rect -27 -4059 -15 -3883
rect -73 -4071 -15 -4059
rect 15 -3883 73 -3871
rect 15 -4059 27 -3883
rect 61 -4059 73 -3883
rect 15 -4071 73 -4059
rect -73 -4301 -15 -4289
rect -73 -4477 -61 -4301
rect -27 -4477 -15 -4301
rect -73 -4489 -15 -4477
rect 15 -4301 73 -4289
rect 15 -4477 27 -4301
rect 61 -4477 73 -4301
rect 15 -4489 73 -4477
rect -73 -4719 -15 -4707
rect -73 -4895 -61 -4719
rect -27 -4895 -15 -4719
rect -73 -4907 -15 -4895
rect 15 -4719 73 -4707
rect 15 -4895 27 -4719
rect 61 -4895 73 -4719
rect 15 -4907 73 -4895
rect -73 -5137 -15 -5125
rect -73 -5313 -61 -5137
rect -27 -5313 -15 -5137
rect -73 -5325 -15 -5313
rect 15 -5137 73 -5125
rect 15 -5313 27 -5137
rect 61 -5313 73 -5137
rect 15 -5325 73 -5313
rect -73 -5555 -15 -5543
rect -73 -5731 -61 -5555
rect -27 -5731 -15 -5555
rect -73 -5743 -15 -5731
rect 15 -5555 73 -5543
rect 15 -5731 27 -5555
rect 61 -5731 73 -5555
rect 15 -5743 73 -5731
rect -73 -5973 -15 -5961
rect -73 -6149 -61 -5973
rect -27 -6149 -15 -5973
rect -73 -6161 -15 -6149
rect 15 -5973 73 -5961
rect 15 -6149 27 -5973
rect 61 -6149 73 -5973
rect 15 -6161 73 -6149
rect -73 -6391 -15 -6379
rect -73 -6567 -61 -6391
rect -27 -6567 -15 -6391
rect -73 -6579 -15 -6567
rect 15 -6391 73 -6379
rect 15 -6567 27 -6391
rect 61 -6567 73 -6391
rect 15 -6579 73 -6567
rect -73 -6809 -15 -6797
rect -73 -6985 -61 -6809
rect -27 -6985 -15 -6809
rect -73 -6997 -15 -6985
rect 15 -6809 73 -6797
rect 15 -6985 27 -6809
rect 61 -6985 73 -6809
rect 15 -6997 73 -6985
rect -73 -7227 -15 -7215
rect -73 -7403 -61 -7227
rect -27 -7403 -15 -7227
rect -73 -7415 -15 -7403
rect 15 -7227 73 -7215
rect 15 -7403 27 -7227
rect 61 -7403 73 -7227
rect 15 -7415 73 -7403
rect -73 -7645 -15 -7633
rect -73 -7821 -61 -7645
rect -27 -7821 -15 -7645
rect -73 -7833 -15 -7821
rect 15 -7645 73 -7633
rect 15 -7821 27 -7645
rect 61 -7821 73 -7645
rect 15 -7833 73 -7821
rect -73 -8063 -15 -8051
rect -73 -8239 -61 -8063
rect -27 -8239 -15 -8063
rect -73 -8251 -15 -8239
rect 15 -8063 73 -8051
rect 15 -8239 27 -8063
rect 61 -8239 73 -8063
rect 15 -8251 73 -8239
rect -73 -8481 -15 -8469
rect -73 -8657 -61 -8481
rect -27 -8657 -15 -8481
rect -73 -8669 -15 -8657
rect 15 -8481 73 -8469
rect 15 -8657 27 -8481
rect 61 -8657 73 -8481
rect 15 -8669 73 -8657
rect -73 -8899 -15 -8887
rect -73 -9075 -61 -8899
rect -27 -9075 -15 -8899
rect -73 -9087 -15 -9075
rect 15 -8899 73 -8887
rect 15 -9075 27 -8899
rect 61 -9075 73 -8899
rect 15 -9087 73 -9075
rect -73 -9317 -15 -9305
rect -73 -9493 -61 -9317
rect -27 -9493 -15 -9317
rect -73 -9505 -15 -9493
rect 15 -9317 73 -9305
rect 15 -9493 27 -9317
rect 61 -9493 73 -9317
rect 15 -9505 73 -9493
rect -73 -9735 -15 -9723
rect -73 -9911 -61 -9735
rect -27 -9911 -15 -9735
rect -73 -9923 -15 -9911
rect 15 -9735 73 -9723
rect 15 -9911 27 -9735
rect 61 -9911 73 -9735
rect 15 -9923 73 -9911
rect -73 -10153 -15 -10141
rect -73 -10329 -61 -10153
rect -27 -10329 -15 -10153
rect -73 -10341 -15 -10329
rect 15 -10153 73 -10141
rect 15 -10329 27 -10153
rect 61 -10329 73 -10153
rect 15 -10341 73 -10329
rect -73 -10571 -15 -10559
rect -73 -10747 -61 -10571
rect -27 -10747 -15 -10571
rect -73 -10759 -15 -10747
rect 15 -10571 73 -10559
rect 15 -10747 27 -10571
rect 61 -10747 73 -10571
rect 15 -10759 73 -10747
rect -73 -10989 -15 -10977
rect -73 -11165 -61 -10989
rect -27 -11165 -15 -10989
rect -73 -11177 -15 -11165
rect 15 -10989 73 -10977
rect 15 -11165 27 -10989
rect 61 -11165 73 -10989
rect 15 -11177 73 -11165
rect -73 -11407 -15 -11395
rect -73 -11583 -61 -11407
rect -27 -11583 -15 -11407
rect -73 -11595 -15 -11583
rect 15 -11407 73 -11395
rect 15 -11583 27 -11407
rect 61 -11583 73 -11407
rect 15 -11595 73 -11583
rect -73 -11825 -15 -11813
rect -73 -12001 -61 -11825
rect -27 -12001 -15 -11825
rect -73 -12013 -15 -12001
rect 15 -11825 73 -11813
rect 15 -12001 27 -11825
rect 61 -12001 73 -11825
rect 15 -12013 73 -12001
rect -73 -12243 -15 -12231
rect -73 -12419 -61 -12243
rect -27 -12419 -15 -12243
rect -73 -12431 -15 -12419
rect 15 -12243 73 -12231
rect 15 -12419 27 -12243
rect 61 -12419 73 -12243
rect 15 -12431 73 -12419
rect -73 -12661 -15 -12649
rect -73 -12837 -61 -12661
rect -27 -12837 -15 -12661
rect -73 -12849 -15 -12837
rect 15 -12661 73 -12649
rect 15 -12837 27 -12661
rect 61 -12837 73 -12661
rect 15 -12849 73 -12837
rect -73 -13079 -15 -13067
rect -73 -13255 -61 -13079
rect -27 -13255 -15 -13079
rect -73 -13267 -15 -13255
rect 15 -13079 73 -13067
rect 15 -13255 27 -13079
rect 61 -13255 73 -13079
rect 15 -13267 73 -13255
<< ndiffc >>
rect -61 13079 -27 13255
rect 27 13079 61 13255
rect -61 12661 -27 12837
rect 27 12661 61 12837
rect -61 12243 -27 12419
rect 27 12243 61 12419
rect -61 11825 -27 12001
rect 27 11825 61 12001
rect -61 11407 -27 11583
rect 27 11407 61 11583
rect -61 10989 -27 11165
rect 27 10989 61 11165
rect -61 10571 -27 10747
rect 27 10571 61 10747
rect -61 10153 -27 10329
rect 27 10153 61 10329
rect -61 9735 -27 9911
rect 27 9735 61 9911
rect -61 9317 -27 9493
rect 27 9317 61 9493
rect -61 8899 -27 9075
rect 27 8899 61 9075
rect -61 8481 -27 8657
rect 27 8481 61 8657
rect -61 8063 -27 8239
rect 27 8063 61 8239
rect -61 7645 -27 7821
rect 27 7645 61 7821
rect -61 7227 -27 7403
rect 27 7227 61 7403
rect -61 6809 -27 6985
rect 27 6809 61 6985
rect -61 6391 -27 6567
rect 27 6391 61 6567
rect -61 5973 -27 6149
rect 27 5973 61 6149
rect -61 5555 -27 5731
rect 27 5555 61 5731
rect -61 5137 -27 5313
rect 27 5137 61 5313
rect -61 4719 -27 4895
rect 27 4719 61 4895
rect -61 4301 -27 4477
rect 27 4301 61 4477
rect -61 3883 -27 4059
rect 27 3883 61 4059
rect -61 3465 -27 3641
rect 27 3465 61 3641
rect -61 3047 -27 3223
rect 27 3047 61 3223
rect -61 2629 -27 2805
rect 27 2629 61 2805
rect -61 2211 -27 2387
rect 27 2211 61 2387
rect -61 1793 -27 1969
rect 27 1793 61 1969
rect -61 1375 -27 1551
rect 27 1375 61 1551
rect -61 957 -27 1133
rect 27 957 61 1133
rect -61 539 -27 715
rect 27 539 61 715
rect -61 121 -27 297
rect 27 121 61 297
rect -61 -297 -27 -121
rect 27 -297 61 -121
rect -61 -715 -27 -539
rect 27 -715 61 -539
rect -61 -1133 -27 -957
rect 27 -1133 61 -957
rect -61 -1551 -27 -1375
rect 27 -1551 61 -1375
rect -61 -1969 -27 -1793
rect 27 -1969 61 -1793
rect -61 -2387 -27 -2211
rect 27 -2387 61 -2211
rect -61 -2805 -27 -2629
rect 27 -2805 61 -2629
rect -61 -3223 -27 -3047
rect 27 -3223 61 -3047
rect -61 -3641 -27 -3465
rect 27 -3641 61 -3465
rect -61 -4059 -27 -3883
rect 27 -4059 61 -3883
rect -61 -4477 -27 -4301
rect 27 -4477 61 -4301
rect -61 -4895 -27 -4719
rect 27 -4895 61 -4719
rect -61 -5313 -27 -5137
rect 27 -5313 61 -5137
rect -61 -5731 -27 -5555
rect 27 -5731 61 -5555
rect -61 -6149 -27 -5973
rect 27 -6149 61 -5973
rect -61 -6567 -27 -6391
rect 27 -6567 61 -6391
rect -61 -6985 -27 -6809
rect 27 -6985 61 -6809
rect -61 -7403 -27 -7227
rect 27 -7403 61 -7227
rect -61 -7821 -27 -7645
rect 27 -7821 61 -7645
rect -61 -8239 -27 -8063
rect 27 -8239 61 -8063
rect -61 -8657 -27 -8481
rect 27 -8657 61 -8481
rect -61 -9075 -27 -8899
rect 27 -9075 61 -8899
rect -61 -9493 -27 -9317
rect 27 -9493 61 -9317
rect -61 -9911 -27 -9735
rect 27 -9911 61 -9735
rect -61 -10329 -27 -10153
rect 27 -10329 61 -10153
rect -61 -10747 -27 -10571
rect 27 -10747 61 -10571
rect -61 -11165 -27 -10989
rect 27 -11165 61 -10989
rect -61 -11583 -27 -11407
rect 27 -11583 61 -11407
rect -61 -12001 -27 -11825
rect 27 -12001 61 -11825
rect -61 -12419 -27 -12243
rect 27 -12419 61 -12243
rect -61 -12837 -27 -12661
rect 27 -12837 61 -12661
rect -61 -13255 -27 -13079
rect 27 -13255 61 -13079
<< psubdiff >>
rect -175 13407 -79 13441
rect 79 13407 175 13441
rect -175 13345 -141 13407
rect 141 13345 175 13407
rect -175 -13407 -141 -13345
rect 141 -13407 175 -13345
rect -175 -13441 -79 -13407
rect 79 -13441 175 -13407
<< psubdiffcont >>
rect -79 13407 79 13441
rect -175 -13345 -141 13345
rect 141 -13345 175 13345
rect -79 -13441 79 -13407
<< poly >>
rect -33 13339 33 13355
rect -33 13305 -17 13339
rect 17 13305 33 13339
rect -33 13289 33 13305
rect -15 13267 15 13289
rect -15 13045 15 13067
rect -33 13029 33 13045
rect -33 12995 -17 13029
rect 17 12995 33 13029
rect -33 12979 33 12995
rect -33 12921 33 12937
rect -33 12887 -17 12921
rect 17 12887 33 12921
rect -33 12871 33 12887
rect -15 12849 15 12871
rect -15 12627 15 12649
rect -33 12611 33 12627
rect -33 12577 -17 12611
rect 17 12577 33 12611
rect -33 12561 33 12577
rect -33 12503 33 12519
rect -33 12469 -17 12503
rect 17 12469 33 12503
rect -33 12453 33 12469
rect -15 12431 15 12453
rect -15 12209 15 12231
rect -33 12193 33 12209
rect -33 12159 -17 12193
rect 17 12159 33 12193
rect -33 12143 33 12159
rect -33 12085 33 12101
rect -33 12051 -17 12085
rect 17 12051 33 12085
rect -33 12035 33 12051
rect -15 12013 15 12035
rect -15 11791 15 11813
rect -33 11775 33 11791
rect -33 11741 -17 11775
rect 17 11741 33 11775
rect -33 11725 33 11741
rect -33 11667 33 11683
rect -33 11633 -17 11667
rect 17 11633 33 11667
rect -33 11617 33 11633
rect -15 11595 15 11617
rect -15 11373 15 11395
rect -33 11357 33 11373
rect -33 11323 -17 11357
rect 17 11323 33 11357
rect -33 11307 33 11323
rect -33 11249 33 11265
rect -33 11215 -17 11249
rect 17 11215 33 11249
rect -33 11199 33 11215
rect -15 11177 15 11199
rect -15 10955 15 10977
rect -33 10939 33 10955
rect -33 10905 -17 10939
rect 17 10905 33 10939
rect -33 10889 33 10905
rect -33 10831 33 10847
rect -33 10797 -17 10831
rect 17 10797 33 10831
rect -33 10781 33 10797
rect -15 10759 15 10781
rect -15 10537 15 10559
rect -33 10521 33 10537
rect -33 10487 -17 10521
rect 17 10487 33 10521
rect -33 10471 33 10487
rect -33 10413 33 10429
rect -33 10379 -17 10413
rect 17 10379 33 10413
rect -33 10363 33 10379
rect -15 10341 15 10363
rect -15 10119 15 10141
rect -33 10103 33 10119
rect -33 10069 -17 10103
rect 17 10069 33 10103
rect -33 10053 33 10069
rect -33 9995 33 10011
rect -33 9961 -17 9995
rect 17 9961 33 9995
rect -33 9945 33 9961
rect -15 9923 15 9945
rect -15 9701 15 9723
rect -33 9685 33 9701
rect -33 9651 -17 9685
rect 17 9651 33 9685
rect -33 9635 33 9651
rect -33 9577 33 9593
rect -33 9543 -17 9577
rect 17 9543 33 9577
rect -33 9527 33 9543
rect -15 9505 15 9527
rect -15 9283 15 9305
rect -33 9267 33 9283
rect -33 9233 -17 9267
rect 17 9233 33 9267
rect -33 9217 33 9233
rect -33 9159 33 9175
rect -33 9125 -17 9159
rect 17 9125 33 9159
rect -33 9109 33 9125
rect -15 9087 15 9109
rect -15 8865 15 8887
rect -33 8849 33 8865
rect -33 8815 -17 8849
rect 17 8815 33 8849
rect -33 8799 33 8815
rect -33 8741 33 8757
rect -33 8707 -17 8741
rect 17 8707 33 8741
rect -33 8691 33 8707
rect -15 8669 15 8691
rect -15 8447 15 8469
rect -33 8431 33 8447
rect -33 8397 -17 8431
rect 17 8397 33 8431
rect -33 8381 33 8397
rect -33 8323 33 8339
rect -33 8289 -17 8323
rect 17 8289 33 8323
rect -33 8273 33 8289
rect -15 8251 15 8273
rect -15 8029 15 8051
rect -33 8013 33 8029
rect -33 7979 -17 8013
rect 17 7979 33 8013
rect -33 7963 33 7979
rect -33 7905 33 7921
rect -33 7871 -17 7905
rect 17 7871 33 7905
rect -33 7855 33 7871
rect -15 7833 15 7855
rect -15 7611 15 7633
rect -33 7595 33 7611
rect -33 7561 -17 7595
rect 17 7561 33 7595
rect -33 7545 33 7561
rect -33 7487 33 7503
rect -33 7453 -17 7487
rect 17 7453 33 7487
rect -33 7437 33 7453
rect -15 7415 15 7437
rect -15 7193 15 7215
rect -33 7177 33 7193
rect -33 7143 -17 7177
rect 17 7143 33 7177
rect -33 7127 33 7143
rect -33 7069 33 7085
rect -33 7035 -17 7069
rect 17 7035 33 7069
rect -33 7019 33 7035
rect -15 6997 15 7019
rect -15 6775 15 6797
rect -33 6759 33 6775
rect -33 6725 -17 6759
rect 17 6725 33 6759
rect -33 6709 33 6725
rect -33 6651 33 6667
rect -33 6617 -17 6651
rect 17 6617 33 6651
rect -33 6601 33 6617
rect -15 6579 15 6601
rect -15 6357 15 6379
rect -33 6341 33 6357
rect -33 6307 -17 6341
rect 17 6307 33 6341
rect -33 6291 33 6307
rect -33 6233 33 6249
rect -33 6199 -17 6233
rect 17 6199 33 6233
rect -33 6183 33 6199
rect -15 6161 15 6183
rect -15 5939 15 5961
rect -33 5923 33 5939
rect -33 5889 -17 5923
rect 17 5889 33 5923
rect -33 5873 33 5889
rect -33 5815 33 5831
rect -33 5781 -17 5815
rect 17 5781 33 5815
rect -33 5765 33 5781
rect -15 5743 15 5765
rect -15 5521 15 5543
rect -33 5505 33 5521
rect -33 5471 -17 5505
rect 17 5471 33 5505
rect -33 5455 33 5471
rect -33 5397 33 5413
rect -33 5363 -17 5397
rect 17 5363 33 5397
rect -33 5347 33 5363
rect -15 5325 15 5347
rect -15 5103 15 5125
rect -33 5087 33 5103
rect -33 5053 -17 5087
rect 17 5053 33 5087
rect -33 5037 33 5053
rect -33 4979 33 4995
rect -33 4945 -17 4979
rect 17 4945 33 4979
rect -33 4929 33 4945
rect -15 4907 15 4929
rect -15 4685 15 4707
rect -33 4669 33 4685
rect -33 4635 -17 4669
rect 17 4635 33 4669
rect -33 4619 33 4635
rect -33 4561 33 4577
rect -33 4527 -17 4561
rect 17 4527 33 4561
rect -33 4511 33 4527
rect -15 4489 15 4511
rect -15 4267 15 4289
rect -33 4251 33 4267
rect -33 4217 -17 4251
rect 17 4217 33 4251
rect -33 4201 33 4217
rect -33 4143 33 4159
rect -33 4109 -17 4143
rect 17 4109 33 4143
rect -33 4093 33 4109
rect -15 4071 15 4093
rect -15 3849 15 3871
rect -33 3833 33 3849
rect -33 3799 -17 3833
rect 17 3799 33 3833
rect -33 3783 33 3799
rect -33 3725 33 3741
rect -33 3691 -17 3725
rect 17 3691 33 3725
rect -33 3675 33 3691
rect -15 3653 15 3675
rect -15 3431 15 3453
rect -33 3415 33 3431
rect -33 3381 -17 3415
rect 17 3381 33 3415
rect -33 3365 33 3381
rect -33 3307 33 3323
rect -33 3273 -17 3307
rect 17 3273 33 3307
rect -33 3257 33 3273
rect -15 3235 15 3257
rect -15 3013 15 3035
rect -33 2997 33 3013
rect -33 2963 -17 2997
rect 17 2963 33 2997
rect -33 2947 33 2963
rect -33 2889 33 2905
rect -33 2855 -17 2889
rect 17 2855 33 2889
rect -33 2839 33 2855
rect -15 2817 15 2839
rect -15 2595 15 2617
rect -33 2579 33 2595
rect -33 2545 -17 2579
rect 17 2545 33 2579
rect -33 2529 33 2545
rect -33 2471 33 2487
rect -33 2437 -17 2471
rect 17 2437 33 2471
rect -33 2421 33 2437
rect -15 2399 15 2421
rect -15 2177 15 2199
rect -33 2161 33 2177
rect -33 2127 -17 2161
rect 17 2127 33 2161
rect -33 2111 33 2127
rect -33 2053 33 2069
rect -33 2019 -17 2053
rect 17 2019 33 2053
rect -33 2003 33 2019
rect -15 1981 15 2003
rect -15 1759 15 1781
rect -33 1743 33 1759
rect -33 1709 -17 1743
rect 17 1709 33 1743
rect -33 1693 33 1709
rect -33 1635 33 1651
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -33 1585 33 1601
rect -15 1563 15 1585
rect -15 1341 15 1363
rect -33 1325 33 1341
rect -33 1291 -17 1325
rect 17 1291 33 1325
rect -33 1275 33 1291
rect -33 1217 33 1233
rect -33 1183 -17 1217
rect 17 1183 33 1217
rect -33 1167 33 1183
rect -15 1145 15 1167
rect -15 923 15 945
rect -33 907 33 923
rect -33 873 -17 907
rect 17 873 33 907
rect -33 857 33 873
rect -33 799 33 815
rect -33 765 -17 799
rect 17 765 33 799
rect -33 749 33 765
rect -15 727 15 749
rect -15 505 15 527
rect -33 489 33 505
rect -33 455 -17 489
rect 17 455 33 489
rect -33 439 33 455
rect -33 381 33 397
rect -33 347 -17 381
rect 17 347 33 381
rect -33 331 33 347
rect -15 309 15 331
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -331 15 -309
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
rect -33 -455 33 -439
rect -33 -489 -17 -455
rect 17 -489 33 -455
rect -33 -505 33 -489
rect -15 -527 15 -505
rect -15 -749 15 -727
rect -33 -765 33 -749
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -815 33 -799
rect -33 -873 33 -857
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -33 -923 33 -907
rect -15 -945 15 -923
rect -15 -1167 15 -1145
rect -33 -1183 33 -1167
rect -33 -1217 -17 -1183
rect 17 -1217 33 -1183
rect -33 -1233 33 -1217
rect -33 -1291 33 -1275
rect -33 -1325 -17 -1291
rect 17 -1325 33 -1291
rect -33 -1341 33 -1325
rect -15 -1363 15 -1341
rect -15 -1585 15 -1563
rect -33 -1601 33 -1585
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1651 33 -1635
rect -33 -1709 33 -1693
rect -33 -1743 -17 -1709
rect 17 -1743 33 -1709
rect -33 -1759 33 -1743
rect -15 -1781 15 -1759
rect -15 -2003 15 -1981
rect -33 -2019 33 -2003
rect -33 -2053 -17 -2019
rect 17 -2053 33 -2019
rect -33 -2069 33 -2053
rect -33 -2127 33 -2111
rect -33 -2161 -17 -2127
rect 17 -2161 33 -2127
rect -33 -2177 33 -2161
rect -15 -2199 15 -2177
rect -15 -2421 15 -2399
rect -33 -2437 33 -2421
rect -33 -2471 -17 -2437
rect 17 -2471 33 -2437
rect -33 -2487 33 -2471
rect -33 -2545 33 -2529
rect -33 -2579 -17 -2545
rect 17 -2579 33 -2545
rect -33 -2595 33 -2579
rect -15 -2617 15 -2595
rect -15 -2839 15 -2817
rect -33 -2855 33 -2839
rect -33 -2889 -17 -2855
rect 17 -2889 33 -2855
rect -33 -2905 33 -2889
rect -33 -2963 33 -2947
rect -33 -2997 -17 -2963
rect 17 -2997 33 -2963
rect -33 -3013 33 -2997
rect -15 -3035 15 -3013
rect -15 -3257 15 -3235
rect -33 -3273 33 -3257
rect -33 -3307 -17 -3273
rect 17 -3307 33 -3273
rect -33 -3323 33 -3307
rect -33 -3381 33 -3365
rect -33 -3415 -17 -3381
rect 17 -3415 33 -3381
rect -33 -3431 33 -3415
rect -15 -3453 15 -3431
rect -15 -3675 15 -3653
rect -33 -3691 33 -3675
rect -33 -3725 -17 -3691
rect 17 -3725 33 -3691
rect -33 -3741 33 -3725
rect -33 -3799 33 -3783
rect -33 -3833 -17 -3799
rect 17 -3833 33 -3799
rect -33 -3849 33 -3833
rect -15 -3871 15 -3849
rect -15 -4093 15 -4071
rect -33 -4109 33 -4093
rect -33 -4143 -17 -4109
rect 17 -4143 33 -4109
rect -33 -4159 33 -4143
rect -33 -4217 33 -4201
rect -33 -4251 -17 -4217
rect 17 -4251 33 -4217
rect -33 -4267 33 -4251
rect -15 -4289 15 -4267
rect -15 -4511 15 -4489
rect -33 -4527 33 -4511
rect -33 -4561 -17 -4527
rect 17 -4561 33 -4527
rect -33 -4577 33 -4561
rect -33 -4635 33 -4619
rect -33 -4669 -17 -4635
rect 17 -4669 33 -4635
rect -33 -4685 33 -4669
rect -15 -4707 15 -4685
rect -15 -4929 15 -4907
rect -33 -4945 33 -4929
rect -33 -4979 -17 -4945
rect 17 -4979 33 -4945
rect -33 -4995 33 -4979
rect -33 -5053 33 -5037
rect -33 -5087 -17 -5053
rect 17 -5087 33 -5053
rect -33 -5103 33 -5087
rect -15 -5125 15 -5103
rect -15 -5347 15 -5325
rect -33 -5363 33 -5347
rect -33 -5397 -17 -5363
rect 17 -5397 33 -5363
rect -33 -5413 33 -5397
rect -33 -5471 33 -5455
rect -33 -5505 -17 -5471
rect 17 -5505 33 -5471
rect -33 -5521 33 -5505
rect -15 -5543 15 -5521
rect -15 -5765 15 -5743
rect -33 -5781 33 -5765
rect -33 -5815 -17 -5781
rect 17 -5815 33 -5781
rect -33 -5831 33 -5815
rect -33 -5889 33 -5873
rect -33 -5923 -17 -5889
rect 17 -5923 33 -5889
rect -33 -5939 33 -5923
rect -15 -5961 15 -5939
rect -15 -6183 15 -6161
rect -33 -6199 33 -6183
rect -33 -6233 -17 -6199
rect 17 -6233 33 -6199
rect -33 -6249 33 -6233
rect -33 -6307 33 -6291
rect -33 -6341 -17 -6307
rect 17 -6341 33 -6307
rect -33 -6357 33 -6341
rect -15 -6379 15 -6357
rect -15 -6601 15 -6579
rect -33 -6617 33 -6601
rect -33 -6651 -17 -6617
rect 17 -6651 33 -6617
rect -33 -6667 33 -6651
rect -33 -6725 33 -6709
rect -33 -6759 -17 -6725
rect 17 -6759 33 -6725
rect -33 -6775 33 -6759
rect -15 -6797 15 -6775
rect -15 -7019 15 -6997
rect -33 -7035 33 -7019
rect -33 -7069 -17 -7035
rect 17 -7069 33 -7035
rect -33 -7085 33 -7069
rect -33 -7143 33 -7127
rect -33 -7177 -17 -7143
rect 17 -7177 33 -7143
rect -33 -7193 33 -7177
rect -15 -7215 15 -7193
rect -15 -7437 15 -7415
rect -33 -7453 33 -7437
rect -33 -7487 -17 -7453
rect 17 -7487 33 -7453
rect -33 -7503 33 -7487
rect -33 -7561 33 -7545
rect -33 -7595 -17 -7561
rect 17 -7595 33 -7561
rect -33 -7611 33 -7595
rect -15 -7633 15 -7611
rect -15 -7855 15 -7833
rect -33 -7871 33 -7855
rect -33 -7905 -17 -7871
rect 17 -7905 33 -7871
rect -33 -7921 33 -7905
rect -33 -7979 33 -7963
rect -33 -8013 -17 -7979
rect 17 -8013 33 -7979
rect -33 -8029 33 -8013
rect -15 -8051 15 -8029
rect -15 -8273 15 -8251
rect -33 -8289 33 -8273
rect -33 -8323 -17 -8289
rect 17 -8323 33 -8289
rect -33 -8339 33 -8323
rect -33 -8397 33 -8381
rect -33 -8431 -17 -8397
rect 17 -8431 33 -8397
rect -33 -8447 33 -8431
rect -15 -8469 15 -8447
rect -15 -8691 15 -8669
rect -33 -8707 33 -8691
rect -33 -8741 -17 -8707
rect 17 -8741 33 -8707
rect -33 -8757 33 -8741
rect -33 -8815 33 -8799
rect -33 -8849 -17 -8815
rect 17 -8849 33 -8815
rect -33 -8865 33 -8849
rect -15 -8887 15 -8865
rect -15 -9109 15 -9087
rect -33 -9125 33 -9109
rect -33 -9159 -17 -9125
rect 17 -9159 33 -9125
rect -33 -9175 33 -9159
rect -33 -9233 33 -9217
rect -33 -9267 -17 -9233
rect 17 -9267 33 -9233
rect -33 -9283 33 -9267
rect -15 -9305 15 -9283
rect -15 -9527 15 -9505
rect -33 -9543 33 -9527
rect -33 -9577 -17 -9543
rect 17 -9577 33 -9543
rect -33 -9593 33 -9577
rect -33 -9651 33 -9635
rect -33 -9685 -17 -9651
rect 17 -9685 33 -9651
rect -33 -9701 33 -9685
rect -15 -9723 15 -9701
rect -15 -9945 15 -9923
rect -33 -9961 33 -9945
rect -33 -9995 -17 -9961
rect 17 -9995 33 -9961
rect -33 -10011 33 -9995
rect -33 -10069 33 -10053
rect -33 -10103 -17 -10069
rect 17 -10103 33 -10069
rect -33 -10119 33 -10103
rect -15 -10141 15 -10119
rect -15 -10363 15 -10341
rect -33 -10379 33 -10363
rect -33 -10413 -17 -10379
rect 17 -10413 33 -10379
rect -33 -10429 33 -10413
rect -33 -10487 33 -10471
rect -33 -10521 -17 -10487
rect 17 -10521 33 -10487
rect -33 -10537 33 -10521
rect -15 -10559 15 -10537
rect -15 -10781 15 -10759
rect -33 -10797 33 -10781
rect -33 -10831 -17 -10797
rect 17 -10831 33 -10797
rect -33 -10847 33 -10831
rect -33 -10905 33 -10889
rect -33 -10939 -17 -10905
rect 17 -10939 33 -10905
rect -33 -10955 33 -10939
rect -15 -10977 15 -10955
rect -15 -11199 15 -11177
rect -33 -11215 33 -11199
rect -33 -11249 -17 -11215
rect 17 -11249 33 -11215
rect -33 -11265 33 -11249
rect -33 -11323 33 -11307
rect -33 -11357 -17 -11323
rect 17 -11357 33 -11323
rect -33 -11373 33 -11357
rect -15 -11395 15 -11373
rect -15 -11617 15 -11595
rect -33 -11633 33 -11617
rect -33 -11667 -17 -11633
rect 17 -11667 33 -11633
rect -33 -11683 33 -11667
rect -33 -11741 33 -11725
rect -33 -11775 -17 -11741
rect 17 -11775 33 -11741
rect -33 -11791 33 -11775
rect -15 -11813 15 -11791
rect -15 -12035 15 -12013
rect -33 -12051 33 -12035
rect -33 -12085 -17 -12051
rect 17 -12085 33 -12051
rect -33 -12101 33 -12085
rect -33 -12159 33 -12143
rect -33 -12193 -17 -12159
rect 17 -12193 33 -12159
rect -33 -12209 33 -12193
rect -15 -12231 15 -12209
rect -15 -12453 15 -12431
rect -33 -12469 33 -12453
rect -33 -12503 -17 -12469
rect 17 -12503 33 -12469
rect -33 -12519 33 -12503
rect -33 -12577 33 -12561
rect -33 -12611 -17 -12577
rect 17 -12611 33 -12577
rect -33 -12627 33 -12611
rect -15 -12649 15 -12627
rect -15 -12871 15 -12849
rect -33 -12887 33 -12871
rect -33 -12921 -17 -12887
rect 17 -12921 33 -12887
rect -33 -12937 33 -12921
rect -33 -12995 33 -12979
rect -33 -13029 -17 -12995
rect 17 -13029 33 -12995
rect -33 -13045 33 -13029
rect -15 -13067 15 -13045
rect -15 -13289 15 -13267
rect -33 -13305 33 -13289
rect -33 -13339 -17 -13305
rect 17 -13339 33 -13305
rect -33 -13355 33 -13339
<< polycont >>
rect -17 13305 17 13339
rect -17 12995 17 13029
rect -17 12887 17 12921
rect -17 12577 17 12611
rect -17 12469 17 12503
rect -17 12159 17 12193
rect -17 12051 17 12085
rect -17 11741 17 11775
rect -17 11633 17 11667
rect -17 11323 17 11357
rect -17 11215 17 11249
rect -17 10905 17 10939
rect -17 10797 17 10831
rect -17 10487 17 10521
rect -17 10379 17 10413
rect -17 10069 17 10103
rect -17 9961 17 9995
rect -17 9651 17 9685
rect -17 9543 17 9577
rect -17 9233 17 9267
rect -17 9125 17 9159
rect -17 8815 17 8849
rect -17 8707 17 8741
rect -17 8397 17 8431
rect -17 8289 17 8323
rect -17 7979 17 8013
rect -17 7871 17 7905
rect -17 7561 17 7595
rect -17 7453 17 7487
rect -17 7143 17 7177
rect -17 7035 17 7069
rect -17 6725 17 6759
rect -17 6617 17 6651
rect -17 6307 17 6341
rect -17 6199 17 6233
rect -17 5889 17 5923
rect -17 5781 17 5815
rect -17 5471 17 5505
rect -17 5363 17 5397
rect -17 5053 17 5087
rect -17 4945 17 4979
rect -17 4635 17 4669
rect -17 4527 17 4561
rect -17 4217 17 4251
rect -17 4109 17 4143
rect -17 3799 17 3833
rect -17 3691 17 3725
rect -17 3381 17 3415
rect -17 3273 17 3307
rect -17 2963 17 2997
rect -17 2855 17 2889
rect -17 2545 17 2579
rect -17 2437 17 2471
rect -17 2127 17 2161
rect -17 2019 17 2053
rect -17 1709 17 1743
rect -17 1601 17 1635
rect -17 1291 17 1325
rect -17 1183 17 1217
rect -17 873 17 907
rect -17 765 17 799
rect -17 455 17 489
rect -17 347 17 381
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -381 17 -347
rect -17 -489 17 -455
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -17 -1217 17 -1183
rect -17 -1325 17 -1291
rect -17 -1635 17 -1601
rect -17 -1743 17 -1709
rect -17 -2053 17 -2019
rect -17 -2161 17 -2127
rect -17 -2471 17 -2437
rect -17 -2579 17 -2545
rect -17 -2889 17 -2855
rect -17 -2997 17 -2963
rect -17 -3307 17 -3273
rect -17 -3415 17 -3381
rect -17 -3725 17 -3691
rect -17 -3833 17 -3799
rect -17 -4143 17 -4109
rect -17 -4251 17 -4217
rect -17 -4561 17 -4527
rect -17 -4669 17 -4635
rect -17 -4979 17 -4945
rect -17 -5087 17 -5053
rect -17 -5397 17 -5363
rect -17 -5505 17 -5471
rect -17 -5815 17 -5781
rect -17 -5923 17 -5889
rect -17 -6233 17 -6199
rect -17 -6341 17 -6307
rect -17 -6651 17 -6617
rect -17 -6759 17 -6725
rect -17 -7069 17 -7035
rect -17 -7177 17 -7143
rect -17 -7487 17 -7453
rect -17 -7595 17 -7561
rect -17 -7905 17 -7871
rect -17 -8013 17 -7979
rect -17 -8323 17 -8289
rect -17 -8431 17 -8397
rect -17 -8741 17 -8707
rect -17 -8849 17 -8815
rect -17 -9159 17 -9125
rect -17 -9267 17 -9233
rect -17 -9577 17 -9543
rect -17 -9685 17 -9651
rect -17 -9995 17 -9961
rect -17 -10103 17 -10069
rect -17 -10413 17 -10379
rect -17 -10521 17 -10487
rect -17 -10831 17 -10797
rect -17 -10939 17 -10905
rect -17 -11249 17 -11215
rect -17 -11357 17 -11323
rect -17 -11667 17 -11633
rect -17 -11775 17 -11741
rect -17 -12085 17 -12051
rect -17 -12193 17 -12159
rect -17 -12503 17 -12469
rect -17 -12611 17 -12577
rect -17 -12921 17 -12887
rect -17 -13029 17 -12995
rect -17 -13339 17 -13305
<< locali >>
rect -175 13407 -79 13441
rect 79 13407 175 13441
rect -175 13345 -141 13407
rect 141 13345 175 13407
rect -33 13305 -17 13339
rect 17 13305 33 13339
rect -61 13255 -27 13271
rect -61 13063 -27 13079
rect 27 13255 61 13271
rect 27 13063 61 13079
rect -33 12995 -17 13029
rect 17 12995 33 13029
rect -33 12887 -17 12921
rect 17 12887 33 12921
rect -61 12837 -27 12853
rect -61 12645 -27 12661
rect 27 12837 61 12853
rect 27 12645 61 12661
rect -33 12577 -17 12611
rect 17 12577 33 12611
rect -33 12469 -17 12503
rect 17 12469 33 12503
rect -61 12419 -27 12435
rect -61 12227 -27 12243
rect 27 12419 61 12435
rect 27 12227 61 12243
rect -33 12159 -17 12193
rect 17 12159 33 12193
rect -33 12051 -17 12085
rect 17 12051 33 12085
rect -61 12001 -27 12017
rect -61 11809 -27 11825
rect 27 12001 61 12017
rect 27 11809 61 11825
rect -33 11741 -17 11775
rect 17 11741 33 11775
rect -33 11633 -17 11667
rect 17 11633 33 11667
rect -61 11583 -27 11599
rect -61 11391 -27 11407
rect 27 11583 61 11599
rect 27 11391 61 11407
rect -33 11323 -17 11357
rect 17 11323 33 11357
rect -33 11215 -17 11249
rect 17 11215 33 11249
rect -61 11165 -27 11181
rect -61 10973 -27 10989
rect 27 11165 61 11181
rect 27 10973 61 10989
rect -33 10905 -17 10939
rect 17 10905 33 10939
rect -33 10797 -17 10831
rect 17 10797 33 10831
rect -61 10747 -27 10763
rect -61 10555 -27 10571
rect 27 10747 61 10763
rect 27 10555 61 10571
rect -33 10487 -17 10521
rect 17 10487 33 10521
rect -33 10379 -17 10413
rect 17 10379 33 10413
rect -61 10329 -27 10345
rect -61 10137 -27 10153
rect 27 10329 61 10345
rect 27 10137 61 10153
rect -33 10069 -17 10103
rect 17 10069 33 10103
rect -33 9961 -17 9995
rect 17 9961 33 9995
rect -61 9911 -27 9927
rect -61 9719 -27 9735
rect 27 9911 61 9927
rect 27 9719 61 9735
rect -33 9651 -17 9685
rect 17 9651 33 9685
rect -33 9543 -17 9577
rect 17 9543 33 9577
rect -61 9493 -27 9509
rect -61 9301 -27 9317
rect 27 9493 61 9509
rect 27 9301 61 9317
rect -33 9233 -17 9267
rect 17 9233 33 9267
rect -33 9125 -17 9159
rect 17 9125 33 9159
rect -61 9075 -27 9091
rect -61 8883 -27 8899
rect 27 9075 61 9091
rect 27 8883 61 8899
rect -33 8815 -17 8849
rect 17 8815 33 8849
rect -33 8707 -17 8741
rect 17 8707 33 8741
rect -61 8657 -27 8673
rect -61 8465 -27 8481
rect 27 8657 61 8673
rect 27 8465 61 8481
rect -33 8397 -17 8431
rect 17 8397 33 8431
rect -33 8289 -17 8323
rect 17 8289 33 8323
rect -61 8239 -27 8255
rect -61 8047 -27 8063
rect 27 8239 61 8255
rect 27 8047 61 8063
rect -33 7979 -17 8013
rect 17 7979 33 8013
rect -33 7871 -17 7905
rect 17 7871 33 7905
rect -61 7821 -27 7837
rect -61 7629 -27 7645
rect 27 7821 61 7837
rect 27 7629 61 7645
rect -33 7561 -17 7595
rect 17 7561 33 7595
rect -33 7453 -17 7487
rect 17 7453 33 7487
rect -61 7403 -27 7419
rect -61 7211 -27 7227
rect 27 7403 61 7419
rect 27 7211 61 7227
rect -33 7143 -17 7177
rect 17 7143 33 7177
rect -33 7035 -17 7069
rect 17 7035 33 7069
rect -61 6985 -27 7001
rect -61 6793 -27 6809
rect 27 6985 61 7001
rect 27 6793 61 6809
rect -33 6725 -17 6759
rect 17 6725 33 6759
rect -33 6617 -17 6651
rect 17 6617 33 6651
rect -61 6567 -27 6583
rect -61 6375 -27 6391
rect 27 6567 61 6583
rect 27 6375 61 6391
rect -33 6307 -17 6341
rect 17 6307 33 6341
rect -33 6199 -17 6233
rect 17 6199 33 6233
rect -61 6149 -27 6165
rect -61 5957 -27 5973
rect 27 6149 61 6165
rect 27 5957 61 5973
rect -33 5889 -17 5923
rect 17 5889 33 5923
rect -33 5781 -17 5815
rect 17 5781 33 5815
rect -61 5731 -27 5747
rect -61 5539 -27 5555
rect 27 5731 61 5747
rect 27 5539 61 5555
rect -33 5471 -17 5505
rect 17 5471 33 5505
rect -33 5363 -17 5397
rect 17 5363 33 5397
rect -61 5313 -27 5329
rect -61 5121 -27 5137
rect 27 5313 61 5329
rect 27 5121 61 5137
rect -33 5053 -17 5087
rect 17 5053 33 5087
rect -33 4945 -17 4979
rect 17 4945 33 4979
rect -61 4895 -27 4911
rect -61 4703 -27 4719
rect 27 4895 61 4911
rect 27 4703 61 4719
rect -33 4635 -17 4669
rect 17 4635 33 4669
rect -33 4527 -17 4561
rect 17 4527 33 4561
rect -61 4477 -27 4493
rect -61 4285 -27 4301
rect 27 4477 61 4493
rect 27 4285 61 4301
rect -33 4217 -17 4251
rect 17 4217 33 4251
rect -33 4109 -17 4143
rect 17 4109 33 4143
rect -61 4059 -27 4075
rect -61 3867 -27 3883
rect 27 4059 61 4075
rect 27 3867 61 3883
rect -33 3799 -17 3833
rect 17 3799 33 3833
rect -33 3691 -17 3725
rect 17 3691 33 3725
rect -61 3641 -27 3657
rect -61 3449 -27 3465
rect 27 3641 61 3657
rect 27 3449 61 3465
rect -33 3381 -17 3415
rect 17 3381 33 3415
rect -33 3273 -17 3307
rect 17 3273 33 3307
rect -61 3223 -27 3239
rect -61 3031 -27 3047
rect 27 3223 61 3239
rect 27 3031 61 3047
rect -33 2963 -17 2997
rect 17 2963 33 2997
rect -33 2855 -17 2889
rect 17 2855 33 2889
rect -61 2805 -27 2821
rect -61 2613 -27 2629
rect 27 2805 61 2821
rect 27 2613 61 2629
rect -33 2545 -17 2579
rect 17 2545 33 2579
rect -33 2437 -17 2471
rect 17 2437 33 2471
rect -61 2387 -27 2403
rect -61 2195 -27 2211
rect 27 2387 61 2403
rect 27 2195 61 2211
rect -33 2127 -17 2161
rect 17 2127 33 2161
rect -33 2019 -17 2053
rect 17 2019 33 2053
rect -61 1969 -27 1985
rect -61 1777 -27 1793
rect 27 1969 61 1985
rect 27 1777 61 1793
rect -33 1709 -17 1743
rect 17 1709 33 1743
rect -33 1601 -17 1635
rect 17 1601 33 1635
rect -61 1551 -27 1567
rect -61 1359 -27 1375
rect 27 1551 61 1567
rect 27 1359 61 1375
rect -33 1291 -17 1325
rect 17 1291 33 1325
rect -33 1183 -17 1217
rect 17 1183 33 1217
rect -61 1133 -27 1149
rect -61 941 -27 957
rect 27 1133 61 1149
rect 27 941 61 957
rect -33 873 -17 907
rect 17 873 33 907
rect -33 765 -17 799
rect 17 765 33 799
rect -61 715 -27 731
rect -61 523 -27 539
rect 27 715 61 731
rect 27 523 61 539
rect -33 455 -17 489
rect 17 455 33 489
rect -33 347 -17 381
rect 17 347 33 381
rect -61 297 -27 313
rect -61 105 -27 121
rect 27 297 61 313
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -313 -27 -297
rect 27 -121 61 -105
rect 27 -313 61 -297
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -489 -17 -455
rect 17 -489 33 -455
rect -61 -539 -27 -523
rect -61 -731 -27 -715
rect 27 -539 61 -523
rect 27 -731 61 -715
rect -33 -799 -17 -765
rect 17 -799 33 -765
rect -33 -907 -17 -873
rect 17 -907 33 -873
rect -61 -957 -27 -941
rect -61 -1149 -27 -1133
rect 27 -957 61 -941
rect 27 -1149 61 -1133
rect -33 -1217 -17 -1183
rect 17 -1217 33 -1183
rect -33 -1325 -17 -1291
rect 17 -1325 33 -1291
rect -61 -1375 -27 -1359
rect -61 -1567 -27 -1551
rect 27 -1375 61 -1359
rect 27 -1567 61 -1551
rect -33 -1635 -17 -1601
rect 17 -1635 33 -1601
rect -33 -1743 -17 -1709
rect 17 -1743 33 -1709
rect -61 -1793 -27 -1777
rect -61 -1985 -27 -1969
rect 27 -1793 61 -1777
rect 27 -1985 61 -1969
rect -33 -2053 -17 -2019
rect 17 -2053 33 -2019
rect -33 -2161 -17 -2127
rect 17 -2161 33 -2127
rect -61 -2211 -27 -2195
rect -61 -2403 -27 -2387
rect 27 -2211 61 -2195
rect 27 -2403 61 -2387
rect -33 -2471 -17 -2437
rect 17 -2471 33 -2437
rect -33 -2579 -17 -2545
rect 17 -2579 33 -2545
rect -61 -2629 -27 -2613
rect -61 -2821 -27 -2805
rect 27 -2629 61 -2613
rect 27 -2821 61 -2805
rect -33 -2889 -17 -2855
rect 17 -2889 33 -2855
rect -33 -2997 -17 -2963
rect 17 -2997 33 -2963
rect -61 -3047 -27 -3031
rect -61 -3239 -27 -3223
rect 27 -3047 61 -3031
rect 27 -3239 61 -3223
rect -33 -3307 -17 -3273
rect 17 -3307 33 -3273
rect -33 -3415 -17 -3381
rect 17 -3415 33 -3381
rect -61 -3465 -27 -3449
rect -61 -3657 -27 -3641
rect 27 -3465 61 -3449
rect 27 -3657 61 -3641
rect -33 -3725 -17 -3691
rect 17 -3725 33 -3691
rect -33 -3833 -17 -3799
rect 17 -3833 33 -3799
rect -61 -3883 -27 -3867
rect -61 -4075 -27 -4059
rect 27 -3883 61 -3867
rect 27 -4075 61 -4059
rect -33 -4143 -17 -4109
rect 17 -4143 33 -4109
rect -33 -4251 -17 -4217
rect 17 -4251 33 -4217
rect -61 -4301 -27 -4285
rect -61 -4493 -27 -4477
rect 27 -4301 61 -4285
rect 27 -4493 61 -4477
rect -33 -4561 -17 -4527
rect 17 -4561 33 -4527
rect -33 -4669 -17 -4635
rect 17 -4669 33 -4635
rect -61 -4719 -27 -4703
rect -61 -4911 -27 -4895
rect 27 -4719 61 -4703
rect 27 -4911 61 -4895
rect -33 -4979 -17 -4945
rect 17 -4979 33 -4945
rect -33 -5087 -17 -5053
rect 17 -5087 33 -5053
rect -61 -5137 -27 -5121
rect -61 -5329 -27 -5313
rect 27 -5137 61 -5121
rect 27 -5329 61 -5313
rect -33 -5397 -17 -5363
rect 17 -5397 33 -5363
rect -33 -5505 -17 -5471
rect 17 -5505 33 -5471
rect -61 -5555 -27 -5539
rect -61 -5747 -27 -5731
rect 27 -5555 61 -5539
rect 27 -5747 61 -5731
rect -33 -5815 -17 -5781
rect 17 -5815 33 -5781
rect -33 -5923 -17 -5889
rect 17 -5923 33 -5889
rect -61 -5973 -27 -5957
rect -61 -6165 -27 -6149
rect 27 -5973 61 -5957
rect 27 -6165 61 -6149
rect -33 -6233 -17 -6199
rect 17 -6233 33 -6199
rect -33 -6341 -17 -6307
rect 17 -6341 33 -6307
rect -61 -6391 -27 -6375
rect -61 -6583 -27 -6567
rect 27 -6391 61 -6375
rect 27 -6583 61 -6567
rect -33 -6651 -17 -6617
rect 17 -6651 33 -6617
rect -33 -6759 -17 -6725
rect 17 -6759 33 -6725
rect -61 -6809 -27 -6793
rect -61 -7001 -27 -6985
rect 27 -6809 61 -6793
rect 27 -7001 61 -6985
rect -33 -7069 -17 -7035
rect 17 -7069 33 -7035
rect -33 -7177 -17 -7143
rect 17 -7177 33 -7143
rect -61 -7227 -27 -7211
rect -61 -7419 -27 -7403
rect 27 -7227 61 -7211
rect 27 -7419 61 -7403
rect -33 -7487 -17 -7453
rect 17 -7487 33 -7453
rect -33 -7595 -17 -7561
rect 17 -7595 33 -7561
rect -61 -7645 -27 -7629
rect -61 -7837 -27 -7821
rect 27 -7645 61 -7629
rect 27 -7837 61 -7821
rect -33 -7905 -17 -7871
rect 17 -7905 33 -7871
rect -33 -8013 -17 -7979
rect 17 -8013 33 -7979
rect -61 -8063 -27 -8047
rect -61 -8255 -27 -8239
rect 27 -8063 61 -8047
rect 27 -8255 61 -8239
rect -33 -8323 -17 -8289
rect 17 -8323 33 -8289
rect -33 -8431 -17 -8397
rect 17 -8431 33 -8397
rect -61 -8481 -27 -8465
rect -61 -8673 -27 -8657
rect 27 -8481 61 -8465
rect 27 -8673 61 -8657
rect -33 -8741 -17 -8707
rect 17 -8741 33 -8707
rect -33 -8849 -17 -8815
rect 17 -8849 33 -8815
rect -61 -8899 -27 -8883
rect -61 -9091 -27 -9075
rect 27 -8899 61 -8883
rect 27 -9091 61 -9075
rect -33 -9159 -17 -9125
rect 17 -9159 33 -9125
rect -33 -9267 -17 -9233
rect 17 -9267 33 -9233
rect -61 -9317 -27 -9301
rect -61 -9509 -27 -9493
rect 27 -9317 61 -9301
rect 27 -9509 61 -9493
rect -33 -9577 -17 -9543
rect 17 -9577 33 -9543
rect -33 -9685 -17 -9651
rect 17 -9685 33 -9651
rect -61 -9735 -27 -9719
rect -61 -9927 -27 -9911
rect 27 -9735 61 -9719
rect 27 -9927 61 -9911
rect -33 -9995 -17 -9961
rect 17 -9995 33 -9961
rect -33 -10103 -17 -10069
rect 17 -10103 33 -10069
rect -61 -10153 -27 -10137
rect -61 -10345 -27 -10329
rect 27 -10153 61 -10137
rect 27 -10345 61 -10329
rect -33 -10413 -17 -10379
rect 17 -10413 33 -10379
rect -33 -10521 -17 -10487
rect 17 -10521 33 -10487
rect -61 -10571 -27 -10555
rect -61 -10763 -27 -10747
rect 27 -10571 61 -10555
rect 27 -10763 61 -10747
rect -33 -10831 -17 -10797
rect 17 -10831 33 -10797
rect -33 -10939 -17 -10905
rect 17 -10939 33 -10905
rect -61 -10989 -27 -10973
rect -61 -11181 -27 -11165
rect 27 -10989 61 -10973
rect 27 -11181 61 -11165
rect -33 -11249 -17 -11215
rect 17 -11249 33 -11215
rect -33 -11357 -17 -11323
rect 17 -11357 33 -11323
rect -61 -11407 -27 -11391
rect -61 -11599 -27 -11583
rect 27 -11407 61 -11391
rect 27 -11599 61 -11583
rect -33 -11667 -17 -11633
rect 17 -11667 33 -11633
rect -33 -11775 -17 -11741
rect 17 -11775 33 -11741
rect -61 -11825 -27 -11809
rect -61 -12017 -27 -12001
rect 27 -11825 61 -11809
rect 27 -12017 61 -12001
rect -33 -12085 -17 -12051
rect 17 -12085 33 -12051
rect -33 -12193 -17 -12159
rect 17 -12193 33 -12159
rect -61 -12243 -27 -12227
rect -61 -12435 -27 -12419
rect 27 -12243 61 -12227
rect 27 -12435 61 -12419
rect -33 -12503 -17 -12469
rect 17 -12503 33 -12469
rect -33 -12611 -17 -12577
rect 17 -12611 33 -12577
rect -61 -12661 -27 -12645
rect -61 -12853 -27 -12837
rect 27 -12661 61 -12645
rect 27 -12853 61 -12837
rect -33 -12921 -17 -12887
rect 17 -12921 33 -12887
rect -33 -13029 -17 -12995
rect 17 -13029 33 -12995
rect -61 -13079 -27 -13063
rect -61 -13271 -27 -13255
rect 27 -13079 61 -13063
rect 27 -13271 61 -13255
rect -33 -13339 -17 -13305
rect 17 -13339 33 -13305
rect -175 -13407 -141 -13345
rect 141 -13407 175 -13345
rect -175 -13441 -79 -13407
rect 79 -13441 175 -13407
<< viali >>
rect -17 13305 17 13339
rect -61 13079 -27 13255
rect 27 13079 61 13255
rect -17 12995 17 13029
rect -17 12887 17 12921
rect -61 12661 -27 12837
rect 27 12661 61 12837
rect -17 12577 17 12611
rect -17 12469 17 12503
rect -61 12243 -27 12419
rect 27 12243 61 12419
rect -17 12159 17 12193
rect -17 12051 17 12085
rect -61 11825 -27 12001
rect 27 11825 61 12001
rect -17 11741 17 11775
rect -17 11633 17 11667
rect -61 11407 -27 11583
rect 27 11407 61 11583
rect -17 11323 17 11357
rect -17 11215 17 11249
rect -61 10989 -27 11165
rect 27 10989 61 11165
rect -17 10905 17 10939
rect -17 10797 17 10831
rect -61 10571 -27 10747
rect 27 10571 61 10747
rect -17 10487 17 10521
rect -17 10379 17 10413
rect -61 10153 -27 10329
rect 27 10153 61 10329
rect -17 10069 17 10103
rect -17 9961 17 9995
rect -61 9735 -27 9911
rect 27 9735 61 9911
rect -17 9651 17 9685
rect -17 9543 17 9577
rect -61 9317 -27 9493
rect 27 9317 61 9493
rect -17 9233 17 9267
rect -17 9125 17 9159
rect -61 8899 -27 9075
rect 27 8899 61 9075
rect -17 8815 17 8849
rect -17 8707 17 8741
rect -61 8481 -27 8657
rect 27 8481 61 8657
rect -17 8397 17 8431
rect -17 8289 17 8323
rect -61 8063 -27 8239
rect 27 8063 61 8239
rect -17 7979 17 8013
rect -17 7871 17 7905
rect -61 7645 -27 7821
rect 27 7645 61 7821
rect -17 7561 17 7595
rect -17 7453 17 7487
rect -61 7227 -27 7403
rect 27 7227 61 7403
rect -17 7143 17 7177
rect -17 7035 17 7069
rect -61 6809 -27 6985
rect 27 6809 61 6985
rect -17 6725 17 6759
rect -17 6617 17 6651
rect -61 6391 -27 6567
rect 27 6391 61 6567
rect -17 6307 17 6341
rect -17 6199 17 6233
rect -61 5973 -27 6149
rect 27 5973 61 6149
rect -17 5889 17 5923
rect -17 5781 17 5815
rect -61 5555 -27 5731
rect 27 5555 61 5731
rect -17 5471 17 5505
rect -17 5363 17 5397
rect -61 5137 -27 5313
rect 27 5137 61 5313
rect -17 5053 17 5087
rect -17 4945 17 4979
rect -61 4719 -27 4895
rect 27 4719 61 4895
rect -17 4635 17 4669
rect -17 4527 17 4561
rect -61 4301 -27 4477
rect 27 4301 61 4477
rect -17 4217 17 4251
rect -17 4109 17 4143
rect -61 3883 -27 4059
rect 27 3883 61 4059
rect -17 3799 17 3833
rect -17 3691 17 3725
rect -61 3465 -27 3641
rect 27 3465 61 3641
rect -17 3381 17 3415
rect -17 3273 17 3307
rect -61 3047 -27 3223
rect 27 3047 61 3223
rect -17 2963 17 2997
rect -17 2855 17 2889
rect -61 2629 -27 2805
rect 27 2629 61 2805
rect -17 2545 17 2579
rect -17 2437 17 2471
rect -61 2211 -27 2387
rect 27 2211 61 2387
rect -17 2127 17 2161
rect -17 2019 17 2053
rect -61 1793 -27 1969
rect 27 1793 61 1969
rect -17 1709 17 1743
rect -17 1601 17 1635
rect -61 1375 -27 1551
rect 27 1375 61 1551
rect -17 1291 17 1325
rect -17 1183 17 1217
rect -61 957 -27 1133
rect 27 957 61 1133
rect -17 873 17 907
rect -17 765 17 799
rect -61 539 -27 715
rect 27 539 61 715
rect -17 455 17 489
rect -17 347 17 381
rect -61 121 -27 297
rect 27 121 61 297
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -297 -27 -121
rect 27 -297 61 -121
rect -17 -381 17 -347
rect -17 -489 17 -455
rect -61 -715 -27 -539
rect 27 -715 61 -539
rect -17 -799 17 -765
rect -17 -907 17 -873
rect -61 -1133 -27 -957
rect 27 -1133 61 -957
rect -17 -1217 17 -1183
rect -17 -1325 17 -1291
rect -61 -1551 -27 -1375
rect 27 -1551 61 -1375
rect -17 -1635 17 -1601
rect -17 -1743 17 -1709
rect -61 -1969 -27 -1793
rect 27 -1969 61 -1793
rect -17 -2053 17 -2019
rect -17 -2161 17 -2127
rect -61 -2387 -27 -2211
rect 27 -2387 61 -2211
rect -17 -2471 17 -2437
rect -17 -2579 17 -2545
rect -61 -2805 -27 -2629
rect 27 -2805 61 -2629
rect -17 -2889 17 -2855
rect -17 -2997 17 -2963
rect -61 -3223 -27 -3047
rect 27 -3223 61 -3047
rect -17 -3307 17 -3273
rect -17 -3415 17 -3381
rect -61 -3641 -27 -3465
rect 27 -3641 61 -3465
rect -17 -3725 17 -3691
rect -17 -3833 17 -3799
rect -61 -4059 -27 -3883
rect 27 -4059 61 -3883
rect -17 -4143 17 -4109
rect -17 -4251 17 -4217
rect -61 -4477 -27 -4301
rect 27 -4477 61 -4301
rect -17 -4561 17 -4527
rect -17 -4669 17 -4635
rect -61 -4895 -27 -4719
rect 27 -4895 61 -4719
rect -17 -4979 17 -4945
rect -17 -5087 17 -5053
rect -61 -5313 -27 -5137
rect 27 -5313 61 -5137
rect -17 -5397 17 -5363
rect -17 -5505 17 -5471
rect -61 -5731 -27 -5555
rect 27 -5731 61 -5555
rect -17 -5815 17 -5781
rect -17 -5923 17 -5889
rect -61 -6149 -27 -5973
rect 27 -6149 61 -5973
rect -17 -6233 17 -6199
rect -17 -6341 17 -6307
rect -61 -6567 -27 -6391
rect 27 -6567 61 -6391
rect -17 -6651 17 -6617
rect -17 -6759 17 -6725
rect -61 -6985 -27 -6809
rect 27 -6985 61 -6809
rect -17 -7069 17 -7035
rect -17 -7177 17 -7143
rect -61 -7403 -27 -7227
rect 27 -7403 61 -7227
rect -17 -7487 17 -7453
rect -17 -7595 17 -7561
rect -61 -7821 -27 -7645
rect 27 -7821 61 -7645
rect -17 -7905 17 -7871
rect -17 -8013 17 -7979
rect -61 -8239 -27 -8063
rect 27 -8239 61 -8063
rect -17 -8323 17 -8289
rect -17 -8431 17 -8397
rect -61 -8657 -27 -8481
rect 27 -8657 61 -8481
rect -17 -8741 17 -8707
rect -17 -8849 17 -8815
rect -61 -9075 -27 -8899
rect 27 -9075 61 -8899
rect -17 -9159 17 -9125
rect -17 -9267 17 -9233
rect -61 -9493 -27 -9317
rect 27 -9493 61 -9317
rect -17 -9577 17 -9543
rect -17 -9685 17 -9651
rect -61 -9911 -27 -9735
rect 27 -9911 61 -9735
rect -17 -9995 17 -9961
rect -17 -10103 17 -10069
rect -61 -10329 -27 -10153
rect 27 -10329 61 -10153
rect -17 -10413 17 -10379
rect -17 -10521 17 -10487
rect -61 -10747 -27 -10571
rect 27 -10747 61 -10571
rect -17 -10831 17 -10797
rect -17 -10939 17 -10905
rect -61 -11165 -27 -10989
rect 27 -11165 61 -10989
rect -17 -11249 17 -11215
rect -17 -11357 17 -11323
rect -61 -11583 -27 -11407
rect 27 -11583 61 -11407
rect -17 -11667 17 -11633
rect -17 -11775 17 -11741
rect -61 -12001 -27 -11825
rect 27 -12001 61 -11825
rect -17 -12085 17 -12051
rect -17 -12193 17 -12159
rect -61 -12419 -27 -12243
rect 27 -12419 61 -12243
rect -17 -12503 17 -12469
rect -17 -12611 17 -12577
rect -61 -12837 -27 -12661
rect 27 -12837 61 -12661
rect -17 -12921 17 -12887
rect -17 -13029 17 -12995
rect -61 -13255 -27 -13079
rect 27 -13255 61 -13079
rect -17 -13339 17 -13305
<< metal1 >>
rect -29 13339 29 13345
rect -29 13305 -17 13339
rect 17 13305 29 13339
rect -29 13299 29 13305
rect -67 13255 -21 13267
rect -67 13079 -61 13255
rect -27 13079 -21 13255
rect -67 13067 -21 13079
rect 21 13255 67 13267
rect 21 13079 27 13255
rect 61 13079 67 13255
rect 21 13067 67 13079
rect -29 13029 29 13035
rect -29 12995 -17 13029
rect 17 12995 29 13029
rect -29 12989 29 12995
rect -29 12921 29 12927
rect -29 12887 -17 12921
rect 17 12887 29 12921
rect -29 12881 29 12887
rect -67 12837 -21 12849
rect -67 12661 -61 12837
rect -27 12661 -21 12837
rect -67 12649 -21 12661
rect 21 12837 67 12849
rect 21 12661 27 12837
rect 61 12661 67 12837
rect 21 12649 67 12661
rect -29 12611 29 12617
rect -29 12577 -17 12611
rect 17 12577 29 12611
rect -29 12571 29 12577
rect -29 12503 29 12509
rect -29 12469 -17 12503
rect 17 12469 29 12503
rect -29 12463 29 12469
rect -67 12419 -21 12431
rect -67 12243 -61 12419
rect -27 12243 -21 12419
rect -67 12231 -21 12243
rect 21 12419 67 12431
rect 21 12243 27 12419
rect 61 12243 67 12419
rect 21 12231 67 12243
rect -29 12193 29 12199
rect -29 12159 -17 12193
rect 17 12159 29 12193
rect -29 12153 29 12159
rect -29 12085 29 12091
rect -29 12051 -17 12085
rect 17 12051 29 12085
rect -29 12045 29 12051
rect -67 12001 -21 12013
rect -67 11825 -61 12001
rect -27 11825 -21 12001
rect -67 11813 -21 11825
rect 21 12001 67 12013
rect 21 11825 27 12001
rect 61 11825 67 12001
rect 21 11813 67 11825
rect -29 11775 29 11781
rect -29 11741 -17 11775
rect 17 11741 29 11775
rect -29 11735 29 11741
rect -29 11667 29 11673
rect -29 11633 -17 11667
rect 17 11633 29 11667
rect -29 11627 29 11633
rect -67 11583 -21 11595
rect -67 11407 -61 11583
rect -27 11407 -21 11583
rect -67 11395 -21 11407
rect 21 11583 67 11595
rect 21 11407 27 11583
rect 61 11407 67 11583
rect 21 11395 67 11407
rect -29 11357 29 11363
rect -29 11323 -17 11357
rect 17 11323 29 11357
rect -29 11317 29 11323
rect -29 11249 29 11255
rect -29 11215 -17 11249
rect 17 11215 29 11249
rect -29 11209 29 11215
rect -67 11165 -21 11177
rect -67 10989 -61 11165
rect -27 10989 -21 11165
rect -67 10977 -21 10989
rect 21 11165 67 11177
rect 21 10989 27 11165
rect 61 10989 67 11165
rect 21 10977 67 10989
rect -29 10939 29 10945
rect -29 10905 -17 10939
rect 17 10905 29 10939
rect -29 10899 29 10905
rect -29 10831 29 10837
rect -29 10797 -17 10831
rect 17 10797 29 10831
rect -29 10791 29 10797
rect -67 10747 -21 10759
rect -67 10571 -61 10747
rect -27 10571 -21 10747
rect -67 10559 -21 10571
rect 21 10747 67 10759
rect 21 10571 27 10747
rect 61 10571 67 10747
rect 21 10559 67 10571
rect -29 10521 29 10527
rect -29 10487 -17 10521
rect 17 10487 29 10521
rect -29 10481 29 10487
rect -29 10413 29 10419
rect -29 10379 -17 10413
rect 17 10379 29 10413
rect -29 10373 29 10379
rect -67 10329 -21 10341
rect -67 10153 -61 10329
rect -27 10153 -21 10329
rect -67 10141 -21 10153
rect 21 10329 67 10341
rect 21 10153 27 10329
rect 61 10153 67 10329
rect 21 10141 67 10153
rect -29 10103 29 10109
rect -29 10069 -17 10103
rect 17 10069 29 10103
rect -29 10063 29 10069
rect -29 9995 29 10001
rect -29 9961 -17 9995
rect 17 9961 29 9995
rect -29 9955 29 9961
rect -67 9911 -21 9923
rect -67 9735 -61 9911
rect -27 9735 -21 9911
rect -67 9723 -21 9735
rect 21 9911 67 9923
rect 21 9735 27 9911
rect 61 9735 67 9911
rect 21 9723 67 9735
rect -29 9685 29 9691
rect -29 9651 -17 9685
rect 17 9651 29 9685
rect -29 9645 29 9651
rect -29 9577 29 9583
rect -29 9543 -17 9577
rect 17 9543 29 9577
rect -29 9537 29 9543
rect -67 9493 -21 9505
rect -67 9317 -61 9493
rect -27 9317 -21 9493
rect -67 9305 -21 9317
rect 21 9493 67 9505
rect 21 9317 27 9493
rect 61 9317 67 9493
rect 21 9305 67 9317
rect -29 9267 29 9273
rect -29 9233 -17 9267
rect 17 9233 29 9267
rect -29 9227 29 9233
rect -29 9159 29 9165
rect -29 9125 -17 9159
rect 17 9125 29 9159
rect -29 9119 29 9125
rect -67 9075 -21 9087
rect -67 8899 -61 9075
rect -27 8899 -21 9075
rect -67 8887 -21 8899
rect 21 9075 67 9087
rect 21 8899 27 9075
rect 61 8899 67 9075
rect 21 8887 67 8899
rect -29 8849 29 8855
rect -29 8815 -17 8849
rect 17 8815 29 8849
rect -29 8809 29 8815
rect -29 8741 29 8747
rect -29 8707 -17 8741
rect 17 8707 29 8741
rect -29 8701 29 8707
rect -67 8657 -21 8669
rect -67 8481 -61 8657
rect -27 8481 -21 8657
rect -67 8469 -21 8481
rect 21 8657 67 8669
rect 21 8481 27 8657
rect 61 8481 67 8657
rect 21 8469 67 8481
rect -29 8431 29 8437
rect -29 8397 -17 8431
rect 17 8397 29 8431
rect -29 8391 29 8397
rect -29 8323 29 8329
rect -29 8289 -17 8323
rect 17 8289 29 8323
rect -29 8283 29 8289
rect -67 8239 -21 8251
rect -67 8063 -61 8239
rect -27 8063 -21 8239
rect -67 8051 -21 8063
rect 21 8239 67 8251
rect 21 8063 27 8239
rect 61 8063 67 8239
rect 21 8051 67 8063
rect -29 8013 29 8019
rect -29 7979 -17 8013
rect 17 7979 29 8013
rect -29 7973 29 7979
rect -29 7905 29 7911
rect -29 7871 -17 7905
rect 17 7871 29 7905
rect -29 7865 29 7871
rect -67 7821 -21 7833
rect -67 7645 -61 7821
rect -27 7645 -21 7821
rect -67 7633 -21 7645
rect 21 7821 67 7833
rect 21 7645 27 7821
rect 61 7645 67 7821
rect 21 7633 67 7645
rect -29 7595 29 7601
rect -29 7561 -17 7595
rect 17 7561 29 7595
rect -29 7555 29 7561
rect -29 7487 29 7493
rect -29 7453 -17 7487
rect 17 7453 29 7487
rect -29 7447 29 7453
rect -67 7403 -21 7415
rect -67 7227 -61 7403
rect -27 7227 -21 7403
rect -67 7215 -21 7227
rect 21 7403 67 7415
rect 21 7227 27 7403
rect 61 7227 67 7403
rect 21 7215 67 7227
rect -29 7177 29 7183
rect -29 7143 -17 7177
rect 17 7143 29 7177
rect -29 7137 29 7143
rect -29 7069 29 7075
rect -29 7035 -17 7069
rect 17 7035 29 7069
rect -29 7029 29 7035
rect -67 6985 -21 6997
rect -67 6809 -61 6985
rect -27 6809 -21 6985
rect -67 6797 -21 6809
rect 21 6985 67 6997
rect 21 6809 27 6985
rect 61 6809 67 6985
rect 21 6797 67 6809
rect -29 6759 29 6765
rect -29 6725 -17 6759
rect 17 6725 29 6759
rect -29 6719 29 6725
rect -29 6651 29 6657
rect -29 6617 -17 6651
rect 17 6617 29 6651
rect -29 6611 29 6617
rect -67 6567 -21 6579
rect -67 6391 -61 6567
rect -27 6391 -21 6567
rect -67 6379 -21 6391
rect 21 6567 67 6579
rect 21 6391 27 6567
rect 61 6391 67 6567
rect 21 6379 67 6391
rect -29 6341 29 6347
rect -29 6307 -17 6341
rect 17 6307 29 6341
rect -29 6301 29 6307
rect -29 6233 29 6239
rect -29 6199 -17 6233
rect 17 6199 29 6233
rect -29 6193 29 6199
rect -67 6149 -21 6161
rect -67 5973 -61 6149
rect -27 5973 -21 6149
rect -67 5961 -21 5973
rect 21 6149 67 6161
rect 21 5973 27 6149
rect 61 5973 67 6149
rect 21 5961 67 5973
rect -29 5923 29 5929
rect -29 5889 -17 5923
rect 17 5889 29 5923
rect -29 5883 29 5889
rect -29 5815 29 5821
rect -29 5781 -17 5815
rect 17 5781 29 5815
rect -29 5775 29 5781
rect -67 5731 -21 5743
rect -67 5555 -61 5731
rect -27 5555 -21 5731
rect -67 5543 -21 5555
rect 21 5731 67 5743
rect 21 5555 27 5731
rect 61 5555 67 5731
rect 21 5543 67 5555
rect -29 5505 29 5511
rect -29 5471 -17 5505
rect 17 5471 29 5505
rect -29 5465 29 5471
rect -29 5397 29 5403
rect -29 5363 -17 5397
rect 17 5363 29 5397
rect -29 5357 29 5363
rect -67 5313 -21 5325
rect -67 5137 -61 5313
rect -27 5137 -21 5313
rect -67 5125 -21 5137
rect 21 5313 67 5325
rect 21 5137 27 5313
rect 61 5137 67 5313
rect 21 5125 67 5137
rect -29 5087 29 5093
rect -29 5053 -17 5087
rect 17 5053 29 5087
rect -29 5047 29 5053
rect -29 4979 29 4985
rect -29 4945 -17 4979
rect 17 4945 29 4979
rect -29 4939 29 4945
rect -67 4895 -21 4907
rect -67 4719 -61 4895
rect -27 4719 -21 4895
rect -67 4707 -21 4719
rect 21 4895 67 4907
rect 21 4719 27 4895
rect 61 4719 67 4895
rect 21 4707 67 4719
rect -29 4669 29 4675
rect -29 4635 -17 4669
rect 17 4635 29 4669
rect -29 4629 29 4635
rect -29 4561 29 4567
rect -29 4527 -17 4561
rect 17 4527 29 4561
rect -29 4521 29 4527
rect -67 4477 -21 4489
rect -67 4301 -61 4477
rect -27 4301 -21 4477
rect -67 4289 -21 4301
rect 21 4477 67 4489
rect 21 4301 27 4477
rect 61 4301 67 4477
rect 21 4289 67 4301
rect -29 4251 29 4257
rect -29 4217 -17 4251
rect 17 4217 29 4251
rect -29 4211 29 4217
rect -29 4143 29 4149
rect -29 4109 -17 4143
rect 17 4109 29 4143
rect -29 4103 29 4109
rect -67 4059 -21 4071
rect -67 3883 -61 4059
rect -27 3883 -21 4059
rect -67 3871 -21 3883
rect 21 4059 67 4071
rect 21 3883 27 4059
rect 61 3883 67 4059
rect 21 3871 67 3883
rect -29 3833 29 3839
rect -29 3799 -17 3833
rect 17 3799 29 3833
rect -29 3793 29 3799
rect -29 3725 29 3731
rect -29 3691 -17 3725
rect 17 3691 29 3725
rect -29 3685 29 3691
rect -67 3641 -21 3653
rect -67 3465 -61 3641
rect -27 3465 -21 3641
rect -67 3453 -21 3465
rect 21 3641 67 3653
rect 21 3465 27 3641
rect 61 3465 67 3641
rect 21 3453 67 3465
rect -29 3415 29 3421
rect -29 3381 -17 3415
rect 17 3381 29 3415
rect -29 3375 29 3381
rect -29 3307 29 3313
rect -29 3273 -17 3307
rect 17 3273 29 3307
rect -29 3267 29 3273
rect -67 3223 -21 3235
rect -67 3047 -61 3223
rect -27 3047 -21 3223
rect -67 3035 -21 3047
rect 21 3223 67 3235
rect 21 3047 27 3223
rect 61 3047 67 3223
rect 21 3035 67 3047
rect -29 2997 29 3003
rect -29 2963 -17 2997
rect 17 2963 29 2997
rect -29 2957 29 2963
rect -29 2889 29 2895
rect -29 2855 -17 2889
rect 17 2855 29 2889
rect -29 2849 29 2855
rect -67 2805 -21 2817
rect -67 2629 -61 2805
rect -27 2629 -21 2805
rect -67 2617 -21 2629
rect 21 2805 67 2817
rect 21 2629 27 2805
rect 61 2629 67 2805
rect 21 2617 67 2629
rect -29 2579 29 2585
rect -29 2545 -17 2579
rect 17 2545 29 2579
rect -29 2539 29 2545
rect -29 2471 29 2477
rect -29 2437 -17 2471
rect 17 2437 29 2471
rect -29 2431 29 2437
rect -67 2387 -21 2399
rect -67 2211 -61 2387
rect -27 2211 -21 2387
rect -67 2199 -21 2211
rect 21 2387 67 2399
rect 21 2211 27 2387
rect 61 2211 67 2387
rect 21 2199 67 2211
rect -29 2161 29 2167
rect -29 2127 -17 2161
rect 17 2127 29 2161
rect -29 2121 29 2127
rect -29 2053 29 2059
rect -29 2019 -17 2053
rect 17 2019 29 2053
rect -29 2013 29 2019
rect -67 1969 -21 1981
rect -67 1793 -61 1969
rect -27 1793 -21 1969
rect -67 1781 -21 1793
rect 21 1969 67 1981
rect 21 1793 27 1969
rect 61 1793 67 1969
rect 21 1781 67 1793
rect -29 1743 29 1749
rect -29 1709 -17 1743
rect 17 1709 29 1743
rect -29 1703 29 1709
rect -29 1635 29 1641
rect -29 1601 -17 1635
rect 17 1601 29 1635
rect -29 1595 29 1601
rect -67 1551 -21 1563
rect -67 1375 -61 1551
rect -27 1375 -21 1551
rect -67 1363 -21 1375
rect 21 1551 67 1563
rect 21 1375 27 1551
rect 61 1375 67 1551
rect 21 1363 67 1375
rect -29 1325 29 1331
rect -29 1291 -17 1325
rect 17 1291 29 1325
rect -29 1285 29 1291
rect -29 1217 29 1223
rect -29 1183 -17 1217
rect 17 1183 29 1217
rect -29 1177 29 1183
rect -67 1133 -21 1145
rect -67 957 -61 1133
rect -27 957 -21 1133
rect -67 945 -21 957
rect 21 1133 67 1145
rect 21 957 27 1133
rect 61 957 67 1133
rect 21 945 67 957
rect -29 907 29 913
rect -29 873 -17 907
rect 17 873 29 907
rect -29 867 29 873
rect -29 799 29 805
rect -29 765 -17 799
rect 17 765 29 799
rect -29 759 29 765
rect -67 715 -21 727
rect -67 539 -61 715
rect -27 539 -21 715
rect -67 527 -21 539
rect 21 715 67 727
rect 21 539 27 715
rect 61 539 67 715
rect 21 527 67 539
rect -29 489 29 495
rect -29 455 -17 489
rect 17 455 29 489
rect -29 449 29 455
rect -29 381 29 387
rect -29 347 -17 381
rect 17 347 29 381
rect -29 341 29 347
rect -67 297 -21 309
rect -67 121 -61 297
rect -27 121 -21 297
rect -67 109 -21 121
rect 21 297 67 309
rect 21 121 27 297
rect 61 121 67 297
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -297 -61 -121
rect -27 -297 -21 -121
rect -67 -309 -21 -297
rect 21 -121 67 -109
rect 21 -297 27 -121
rect 61 -297 67 -121
rect 21 -309 67 -297
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
rect -29 -455 29 -449
rect -29 -489 -17 -455
rect 17 -489 29 -455
rect -29 -495 29 -489
rect -67 -539 -21 -527
rect -67 -715 -61 -539
rect -27 -715 -21 -539
rect -67 -727 -21 -715
rect 21 -539 67 -527
rect 21 -715 27 -539
rect 61 -715 67 -539
rect 21 -727 67 -715
rect -29 -765 29 -759
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -805 29 -799
rect -29 -873 29 -867
rect -29 -907 -17 -873
rect 17 -907 29 -873
rect -29 -913 29 -907
rect -67 -957 -21 -945
rect -67 -1133 -61 -957
rect -27 -1133 -21 -957
rect -67 -1145 -21 -1133
rect 21 -957 67 -945
rect 21 -1133 27 -957
rect 61 -1133 67 -957
rect 21 -1145 67 -1133
rect -29 -1183 29 -1177
rect -29 -1217 -17 -1183
rect 17 -1217 29 -1183
rect -29 -1223 29 -1217
rect -29 -1291 29 -1285
rect -29 -1325 -17 -1291
rect 17 -1325 29 -1291
rect -29 -1331 29 -1325
rect -67 -1375 -21 -1363
rect -67 -1551 -61 -1375
rect -27 -1551 -21 -1375
rect -67 -1563 -21 -1551
rect 21 -1375 67 -1363
rect 21 -1551 27 -1375
rect 61 -1551 67 -1375
rect 21 -1563 67 -1551
rect -29 -1601 29 -1595
rect -29 -1635 -17 -1601
rect 17 -1635 29 -1601
rect -29 -1641 29 -1635
rect -29 -1709 29 -1703
rect -29 -1743 -17 -1709
rect 17 -1743 29 -1709
rect -29 -1749 29 -1743
rect -67 -1793 -21 -1781
rect -67 -1969 -61 -1793
rect -27 -1969 -21 -1793
rect -67 -1981 -21 -1969
rect 21 -1793 67 -1781
rect 21 -1969 27 -1793
rect 61 -1969 67 -1793
rect 21 -1981 67 -1969
rect -29 -2019 29 -2013
rect -29 -2053 -17 -2019
rect 17 -2053 29 -2019
rect -29 -2059 29 -2053
rect -29 -2127 29 -2121
rect -29 -2161 -17 -2127
rect 17 -2161 29 -2127
rect -29 -2167 29 -2161
rect -67 -2211 -21 -2199
rect -67 -2387 -61 -2211
rect -27 -2387 -21 -2211
rect -67 -2399 -21 -2387
rect 21 -2211 67 -2199
rect 21 -2387 27 -2211
rect 61 -2387 67 -2211
rect 21 -2399 67 -2387
rect -29 -2437 29 -2431
rect -29 -2471 -17 -2437
rect 17 -2471 29 -2437
rect -29 -2477 29 -2471
rect -29 -2545 29 -2539
rect -29 -2579 -17 -2545
rect 17 -2579 29 -2545
rect -29 -2585 29 -2579
rect -67 -2629 -21 -2617
rect -67 -2805 -61 -2629
rect -27 -2805 -21 -2629
rect -67 -2817 -21 -2805
rect 21 -2629 67 -2617
rect 21 -2805 27 -2629
rect 61 -2805 67 -2629
rect 21 -2817 67 -2805
rect -29 -2855 29 -2849
rect -29 -2889 -17 -2855
rect 17 -2889 29 -2855
rect -29 -2895 29 -2889
rect -29 -2963 29 -2957
rect -29 -2997 -17 -2963
rect 17 -2997 29 -2963
rect -29 -3003 29 -2997
rect -67 -3047 -21 -3035
rect -67 -3223 -61 -3047
rect -27 -3223 -21 -3047
rect -67 -3235 -21 -3223
rect 21 -3047 67 -3035
rect 21 -3223 27 -3047
rect 61 -3223 67 -3047
rect 21 -3235 67 -3223
rect -29 -3273 29 -3267
rect -29 -3307 -17 -3273
rect 17 -3307 29 -3273
rect -29 -3313 29 -3307
rect -29 -3381 29 -3375
rect -29 -3415 -17 -3381
rect 17 -3415 29 -3381
rect -29 -3421 29 -3415
rect -67 -3465 -21 -3453
rect -67 -3641 -61 -3465
rect -27 -3641 -21 -3465
rect -67 -3653 -21 -3641
rect 21 -3465 67 -3453
rect 21 -3641 27 -3465
rect 61 -3641 67 -3465
rect 21 -3653 67 -3641
rect -29 -3691 29 -3685
rect -29 -3725 -17 -3691
rect 17 -3725 29 -3691
rect -29 -3731 29 -3725
rect -29 -3799 29 -3793
rect -29 -3833 -17 -3799
rect 17 -3833 29 -3799
rect -29 -3839 29 -3833
rect -67 -3883 -21 -3871
rect -67 -4059 -61 -3883
rect -27 -4059 -21 -3883
rect -67 -4071 -21 -4059
rect 21 -3883 67 -3871
rect 21 -4059 27 -3883
rect 61 -4059 67 -3883
rect 21 -4071 67 -4059
rect -29 -4109 29 -4103
rect -29 -4143 -17 -4109
rect 17 -4143 29 -4109
rect -29 -4149 29 -4143
rect -29 -4217 29 -4211
rect -29 -4251 -17 -4217
rect 17 -4251 29 -4217
rect -29 -4257 29 -4251
rect -67 -4301 -21 -4289
rect -67 -4477 -61 -4301
rect -27 -4477 -21 -4301
rect -67 -4489 -21 -4477
rect 21 -4301 67 -4289
rect 21 -4477 27 -4301
rect 61 -4477 67 -4301
rect 21 -4489 67 -4477
rect -29 -4527 29 -4521
rect -29 -4561 -17 -4527
rect 17 -4561 29 -4527
rect -29 -4567 29 -4561
rect -29 -4635 29 -4629
rect -29 -4669 -17 -4635
rect 17 -4669 29 -4635
rect -29 -4675 29 -4669
rect -67 -4719 -21 -4707
rect -67 -4895 -61 -4719
rect -27 -4895 -21 -4719
rect -67 -4907 -21 -4895
rect 21 -4719 67 -4707
rect 21 -4895 27 -4719
rect 61 -4895 67 -4719
rect 21 -4907 67 -4895
rect -29 -4945 29 -4939
rect -29 -4979 -17 -4945
rect 17 -4979 29 -4945
rect -29 -4985 29 -4979
rect -29 -5053 29 -5047
rect -29 -5087 -17 -5053
rect 17 -5087 29 -5053
rect -29 -5093 29 -5087
rect -67 -5137 -21 -5125
rect -67 -5313 -61 -5137
rect -27 -5313 -21 -5137
rect -67 -5325 -21 -5313
rect 21 -5137 67 -5125
rect 21 -5313 27 -5137
rect 61 -5313 67 -5137
rect 21 -5325 67 -5313
rect -29 -5363 29 -5357
rect -29 -5397 -17 -5363
rect 17 -5397 29 -5363
rect -29 -5403 29 -5397
rect -29 -5471 29 -5465
rect -29 -5505 -17 -5471
rect 17 -5505 29 -5471
rect -29 -5511 29 -5505
rect -67 -5555 -21 -5543
rect -67 -5731 -61 -5555
rect -27 -5731 -21 -5555
rect -67 -5743 -21 -5731
rect 21 -5555 67 -5543
rect 21 -5731 27 -5555
rect 61 -5731 67 -5555
rect 21 -5743 67 -5731
rect -29 -5781 29 -5775
rect -29 -5815 -17 -5781
rect 17 -5815 29 -5781
rect -29 -5821 29 -5815
rect -29 -5889 29 -5883
rect -29 -5923 -17 -5889
rect 17 -5923 29 -5889
rect -29 -5929 29 -5923
rect -67 -5973 -21 -5961
rect -67 -6149 -61 -5973
rect -27 -6149 -21 -5973
rect -67 -6161 -21 -6149
rect 21 -5973 67 -5961
rect 21 -6149 27 -5973
rect 61 -6149 67 -5973
rect 21 -6161 67 -6149
rect -29 -6199 29 -6193
rect -29 -6233 -17 -6199
rect 17 -6233 29 -6199
rect -29 -6239 29 -6233
rect -29 -6307 29 -6301
rect -29 -6341 -17 -6307
rect 17 -6341 29 -6307
rect -29 -6347 29 -6341
rect -67 -6391 -21 -6379
rect -67 -6567 -61 -6391
rect -27 -6567 -21 -6391
rect -67 -6579 -21 -6567
rect 21 -6391 67 -6379
rect 21 -6567 27 -6391
rect 61 -6567 67 -6391
rect 21 -6579 67 -6567
rect -29 -6617 29 -6611
rect -29 -6651 -17 -6617
rect 17 -6651 29 -6617
rect -29 -6657 29 -6651
rect -29 -6725 29 -6719
rect -29 -6759 -17 -6725
rect 17 -6759 29 -6725
rect -29 -6765 29 -6759
rect -67 -6809 -21 -6797
rect -67 -6985 -61 -6809
rect -27 -6985 -21 -6809
rect -67 -6997 -21 -6985
rect 21 -6809 67 -6797
rect 21 -6985 27 -6809
rect 61 -6985 67 -6809
rect 21 -6997 67 -6985
rect -29 -7035 29 -7029
rect -29 -7069 -17 -7035
rect 17 -7069 29 -7035
rect -29 -7075 29 -7069
rect -29 -7143 29 -7137
rect -29 -7177 -17 -7143
rect 17 -7177 29 -7143
rect -29 -7183 29 -7177
rect -67 -7227 -21 -7215
rect -67 -7403 -61 -7227
rect -27 -7403 -21 -7227
rect -67 -7415 -21 -7403
rect 21 -7227 67 -7215
rect 21 -7403 27 -7227
rect 61 -7403 67 -7227
rect 21 -7415 67 -7403
rect -29 -7453 29 -7447
rect -29 -7487 -17 -7453
rect 17 -7487 29 -7453
rect -29 -7493 29 -7487
rect -29 -7561 29 -7555
rect -29 -7595 -17 -7561
rect 17 -7595 29 -7561
rect -29 -7601 29 -7595
rect -67 -7645 -21 -7633
rect -67 -7821 -61 -7645
rect -27 -7821 -21 -7645
rect -67 -7833 -21 -7821
rect 21 -7645 67 -7633
rect 21 -7821 27 -7645
rect 61 -7821 67 -7645
rect 21 -7833 67 -7821
rect -29 -7871 29 -7865
rect -29 -7905 -17 -7871
rect 17 -7905 29 -7871
rect -29 -7911 29 -7905
rect -29 -7979 29 -7973
rect -29 -8013 -17 -7979
rect 17 -8013 29 -7979
rect -29 -8019 29 -8013
rect -67 -8063 -21 -8051
rect -67 -8239 -61 -8063
rect -27 -8239 -21 -8063
rect -67 -8251 -21 -8239
rect 21 -8063 67 -8051
rect 21 -8239 27 -8063
rect 61 -8239 67 -8063
rect 21 -8251 67 -8239
rect -29 -8289 29 -8283
rect -29 -8323 -17 -8289
rect 17 -8323 29 -8289
rect -29 -8329 29 -8323
rect -29 -8397 29 -8391
rect -29 -8431 -17 -8397
rect 17 -8431 29 -8397
rect -29 -8437 29 -8431
rect -67 -8481 -21 -8469
rect -67 -8657 -61 -8481
rect -27 -8657 -21 -8481
rect -67 -8669 -21 -8657
rect 21 -8481 67 -8469
rect 21 -8657 27 -8481
rect 61 -8657 67 -8481
rect 21 -8669 67 -8657
rect -29 -8707 29 -8701
rect -29 -8741 -17 -8707
rect 17 -8741 29 -8707
rect -29 -8747 29 -8741
rect -29 -8815 29 -8809
rect -29 -8849 -17 -8815
rect 17 -8849 29 -8815
rect -29 -8855 29 -8849
rect -67 -8899 -21 -8887
rect -67 -9075 -61 -8899
rect -27 -9075 -21 -8899
rect -67 -9087 -21 -9075
rect 21 -8899 67 -8887
rect 21 -9075 27 -8899
rect 61 -9075 67 -8899
rect 21 -9087 67 -9075
rect -29 -9125 29 -9119
rect -29 -9159 -17 -9125
rect 17 -9159 29 -9125
rect -29 -9165 29 -9159
rect -29 -9233 29 -9227
rect -29 -9267 -17 -9233
rect 17 -9267 29 -9233
rect -29 -9273 29 -9267
rect -67 -9317 -21 -9305
rect -67 -9493 -61 -9317
rect -27 -9493 -21 -9317
rect -67 -9505 -21 -9493
rect 21 -9317 67 -9305
rect 21 -9493 27 -9317
rect 61 -9493 67 -9317
rect 21 -9505 67 -9493
rect -29 -9543 29 -9537
rect -29 -9577 -17 -9543
rect 17 -9577 29 -9543
rect -29 -9583 29 -9577
rect -29 -9651 29 -9645
rect -29 -9685 -17 -9651
rect 17 -9685 29 -9651
rect -29 -9691 29 -9685
rect -67 -9735 -21 -9723
rect -67 -9911 -61 -9735
rect -27 -9911 -21 -9735
rect -67 -9923 -21 -9911
rect 21 -9735 67 -9723
rect 21 -9911 27 -9735
rect 61 -9911 67 -9735
rect 21 -9923 67 -9911
rect -29 -9961 29 -9955
rect -29 -9995 -17 -9961
rect 17 -9995 29 -9961
rect -29 -10001 29 -9995
rect -29 -10069 29 -10063
rect -29 -10103 -17 -10069
rect 17 -10103 29 -10069
rect -29 -10109 29 -10103
rect -67 -10153 -21 -10141
rect -67 -10329 -61 -10153
rect -27 -10329 -21 -10153
rect -67 -10341 -21 -10329
rect 21 -10153 67 -10141
rect 21 -10329 27 -10153
rect 61 -10329 67 -10153
rect 21 -10341 67 -10329
rect -29 -10379 29 -10373
rect -29 -10413 -17 -10379
rect 17 -10413 29 -10379
rect -29 -10419 29 -10413
rect -29 -10487 29 -10481
rect -29 -10521 -17 -10487
rect 17 -10521 29 -10487
rect -29 -10527 29 -10521
rect -67 -10571 -21 -10559
rect -67 -10747 -61 -10571
rect -27 -10747 -21 -10571
rect -67 -10759 -21 -10747
rect 21 -10571 67 -10559
rect 21 -10747 27 -10571
rect 61 -10747 67 -10571
rect 21 -10759 67 -10747
rect -29 -10797 29 -10791
rect -29 -10831 -17 -10797
rect 17 -10831 29 -10797
rect -29 -10837 29 -10831
rect -29 -10905 29 -10899
rect -29 -10939 -17 -10905
rect 17 -10939 29 -10905
rect -29 -10945 29 -10939
rect -67 -10989 -21 -10977
rect -67 -11165 -61 -10989
rect -27 -11165 -21 -10989
rect -67 -11177 -21 -11165
rect 21 -10989 67 -10977
rect 21 -11165 27 -10989
rect 61 -11165 67 -10989
rect 21 -11177 67 -11165
rect -29 -11215 29 -11209
rect -29 -11249 -17 -11215
rect 17 -11249 29 -11215
rect -29 -11255 29 -11249
rect -29 -11323 29 -11317
rect -29 -11357 -17 -11323
rect 17 -11357 29 -11323
rect -29 -11363 29 -11357
rect -67 -11407 -21 -11395
rect -67 -11583 -61 -11407
rect -27 -11583 -21 -11407
rect -67 -11595 -21 -11583
rect 21 -11407 67 -11395
rect 21 -11583 27 -11407
rect 61 -11583 67 -11407
rect 21 -11595 67 -11583
rect -29 -11633 29 -11627
rect -29 -11667 -17 -11633
rect 17 -11667 29 -11633
rect -29 -11673 29 -11667
rect -29 -11741 29 -11735
rect -29 -11775 -17 -11741
rect 17 -11775 29 -11741
rect -29 -11781 29 -11775
rect -67 -11825 -21 -11813
rect -67 -12001 -61 -11825
rect -27 -12001 -21 -11825
rect -67 -12013 -21 -12001
rect 21 -11825 67 -11813
rect 21 -12001 27 -11825
rect 61 -12001 67 -11825
rect 21 -12013 67 -12001
rect -29 -12051 29 -12045
rect -29 -12085 -17 -12051
rect 17 -12085 29 -12051
rect -29 -12091 29 -12085
rect -29 -12159 29 -12153
rect -29 -12193 -17 -12159
rect 17 -12193 29 -12159
rect -29 -12199 29 -12193
rect -67 -12243 -21 -12231
rect -67 -12419 -61 -12243
rect -27 -12419 -21 -12243
rect -67 -12431 -21 -12419
rect 21 -12243 67 -12231
rect 21 -12419 27 -12243
rect 61 -12419 67 -12243
rect 21 -12431 67 -12419
rect -29 -12469 29 -12463
rect -29 -12503 -17 -12469
rect 17 -12503 29 -12469
rect -29 -12509 29 -12503
rect -29 -12577 29 -12571
rect -29 -12611 -17 -12577
rect 17 -12611 29 -12577
rect -29 -12617 29 -12611
rect -67 -12661 -21 -12649
rect -67 -12837 -61 -12661
rect -27 -12837 -21 -12661
rect -67 -12849 -21 -12837
rect 21 -12661 67 -12649
rect 21 -12837 27 -12661
rect 61 -12837 67 -12661
rect 21 -12849 67 -12837
rect -29 -12887 29 -12881
rect -29 -12921 -17 -12887
rect 17 -12921 29 -12887
rect -29 -12927 29 -12921
rect -29 -12995 29 -12989
rect -29 -13029 -17 -12995
rect 17 -13029 29 -12995
rect -29 -13035 29 -13029
rect -67 -13079 -21 -13067
rect -67 -13255 -61 -13079
rect -27 -13255 -21 -13079
rect -67 -13267 -21 -13255
rect 21 -13079 67 -13067
rect 21 -13255 27 -13079
rect 61 -13255 67 -13079
rect 21 -13267 67 -13255
rect -29 -13305 29 -13299
rect -29 -13339 -17 -13305
rect 17 -13339 29 -13305
rect -29 -13345 29 -13339
<< properties >>
string FIXED_BBOX -158 -13424 158 13424
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 64 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
