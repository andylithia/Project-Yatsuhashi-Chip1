magic
tech sky130B
magscale 1 2
timestamp 1659585137
<< error_p >>
rect -653 472 -595 478
rect -461 472 -403 478
rect -269 472 -211 478
rect -77 472 -19 478
rect 115 472 173 478
rect 307 472 365 478
rect 499 472 557 478
rect 691 472 749 478
rect -653 438 -641 472
rect -461 438 -449 472
rect -269 438 -257 472
rect -77 438 -65 472
rect 115 438 127 472
rect 307 438 319 472
rect 499 438 511 472
rect 691 438 703 472
rect -653 432 -595 438
rect -461 432 -403 438
rect -269 432 -211 438
rect -77 432 -19 438
rect 115 432 173 438
rect 307 432 365 438
rect 499 432 557 438
rect 691 432 749 438
rect -749 -438 -691 -432
rect -557 -438 -499 -432
rect -365 -438 -307 -432
rect -173 -438 -115 -432
rect 19 -438 77 -432
rect 211 -438 269 -432
rect 403 -438 461 -432
rect 595 -438 653 -432
rect -749 -472 -737 -438
rect -557 -472 -545 -438
rect -365 -472 -353 -438
rect -173 -472 -161 -438
rect 19 -472 31 -438
rect 211 -472 223 -438
rect 403 -472 415 -438
rect 595 -472 607 -438
rect -749 -478 -691 -472
rect -557 -478 -499 -472
rect -365 -478 -307 -472
rect -173 -478 -115 -472
rect 19 -478 77 -472
rect 211 -478 269 -472
rect 403 -478 461 -472
rect 595 -478 653 -472
<< pwell >>
rect -935 -610 935 610
<< nmos >>
rect -735 -400 -705 400
rect -639 -400 -609 400
rect -543 -400 -513 400
rect -447 -400 -417 400
rect -351 -400 -321 400
rect -255 -400 -225 400
rect -159 -400 -129 400
rect -63 -400 -33 400
rect 33 -400 63 400
rect 129 -400 159 400
rect 225 -400 255 400
rect 321 -400 351 400
rect 417 -400 447 400
rect 513 -400 543 400
rect 609 -400 639 400
rect 705 -400 735 400
<< ndiff >>
rect -797 388 -735 400
rect -797 -388 -785 388
rect -751 -388 -735 388
rect -797 -400 -735 -388
rect -705 388 -639 400
rect -705 -388 -689 388
rect -655 -388 -639 388
rect -705 -400 -639 -388
rect -609 388 -543 400
rect -609 -388 -593 388
rect -559 -388 -543 388
rect -609 -400 -543 -388
rect -513 388 -447 400
rect -513 -388 -497 388
rect -463 -388 -447 388
rect -513 -400 -447 -388
rect -417 388 -351 400
rect -417 -388 -401 388
rect -367 -388 -351 388
rect -417 -400 -351 -388
rect -321 388 -255 400
rect -321 -388 -305 388
rect -271 -388 -255 388
rect -321 -400 -255 -388
rect -225 388 -159 400
rect -225 -388 -209 388
rect -175 -388 -159 388
rect -225 -400 -159 -388
rect -129 388 -63 400
rect -129 -388 -113 388
rect -79 -388 -63 388
rect -129 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 129 400
rect 63 -388 79 388
rect 113 -388 129 388
rect 63 -400 129 -388
rect 159 388 225 400
rect 159 -388 175 388
rect 209 -388 225 388
rect 159 -400 225 -388
rect 255 388 321 400
rect 255 -388 271 388
rect 305 -388 321 388
rect 255 -400 321 -388
rect 351 388 417 400
rect 351 -388 367 388
rect 401 -388 417 388
rect 351 -400 417 -388
rect 447 388 513 400
rect 447 -388 463 388
rect 497 -388 513 388
rect 447 -400 513 -388
rect 543 388 609 400
rect 543 -388 559 388
rect 593 -388 609 388
rect 543 -400 609 -388
rect 639 388 705 400
rect 639 -388 655 388
rect 689 -388 705 388
rect 639 -400 705 -388
rect 735 388 797 400
rect 735 -388 751 388
rect 785 -388 797 388
rect 735 -400 797 -388
<< ndiffc >>
rect -785 -388 -751 388
rect -689 -388 -655 388
rect -593 -388 -559 388
rect -497 -388 -463 388
rect -401 -388 -367 388
rect -305 -388 -271 388
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect 271 -388 305 388
rect 367 -388 401 388
rect 463 -388 497 388
rect 559 -388 593 388
rect 655 -388 689 388
rect 751 -388 785 388
<< psubdiff >>
rect -899 540 899 574
rect -899 478 -865 540
rect 865 478 899 540
rect -899 -540 -865 -478
rect 865 -540 899 -478
rect -899 -574 -803 -540
rect 803 -574 899 -540
<< psubdiffcont >>
rect -899 -478 -865 478
rect 865 -478 899 478
rect -803 -574 803 -540
<< poly >>
rect -657 472 -591 488
rect -657 438 -641 472
rect -607 438 -591 472
rect -735 400 -705 426
rect -657 422 -591 438
rect -465 472 -399 488
rect -465 438 -449 472
rect -415 438 -399 472
rect -639 400 -609 422
rect -543 400 -513 426
rect -465 422 -399 438
rect -273 472 -207 488
rect -273 438 -257 472
rect -223 438 -207 472
rect -447 400 -417 422
rect -351 400 -321 426
rect -273 422 -207 438
rect -81 472 -15 488
rect -81 438 -65 472
rect -31 438 -15 472
rect -255 400 -225 422
rect -159 400 -129 426
rect -81 422 -15 438
rect 111 472 177 488
rect 111 438 127 472
rect 161 438 177 472
rect -63 400 -33 422
rect 33 400 63 426
rect 111 422 177 438
rect 303 472 369 488
rect 303 438 319 472
rect 353 438 369 472
rect 129 400 159 422
rect 225 400 255 426
rect 303 422 369 438
rect 495 472 561 488
rect 495 438 511 472
rect 545 438 561 472
rect 321 400 351 422
rect 417 400 447 426
rect 495 422 561 438
rect 687 472 753 488
rect 687 438 703 472
rect 737 438 753 472
rect 513 400 543 422
rect 609 400 639 426
rect 687 422 753 438
rect 705 400 735 422
rect -735 -422 -705 -400
rect -753 -438 -687 -422
rect -639 -426 -609 -400
rect -543 -422 -513 -400
rect -753 -472 -737 -438
rect -703 -472 -687 -438
rect -753 -488 -687 -472
rect -561 -438 -495 -422
rect -447 -426 -417 -400
rect -351 -422 -321 -400
rect -561 -472 -545 -438
rect -511 -472 -495 -438
rect -561 -488 -495 -472
rect -369 -438 -303 -422
rect -255 -426 -225 -400
rect -159 -422 -129 -400
rect -369 -472 -353 -438
rect -319 -472 -303 -438
rect -369 -488 -303 -472
rect -177 -438 -111 -422
rect -63 -426 -33 -400
rect 33 -422 63 -400
rect -177 -472 -161 -438
rect -127 -472 -111 -438
rect -177 -488 -111 -472
rect 15 -438 81 -422
rect 129 -426 159 -400
rect 225 -422 255 -400
rect 15 -472 31 -438
rect 65 -472 81 -438
rect 15 -488 81 -472
rect 207 -438 273 -422
rect 321 -426 351 -400
rect 417 -422 447 -400
rect 207 -472 223 -438
rect 257 -472 273 -438
rect 207 -488 273 -472
rect 399 -438 465 -422
rect 513 -426 543 -400
rect 609 -422 639 -400
rect 399 -472 415 -438
rect 449 -472 465 -438
rect 399 -488 465 -472
rect 591 -438 657 -422
rect 705 -426 735 -400
rect 591 -472 607 -438
rect 641 -472 657 -438
rect 591 -488 657 -472
<< polycont >>
rect -641 438 -607 472
rect -449 438 -415 472
rect -257 438 -223 472
rect -65 438 -31 472
rect 127 438 161 472
rect 319 438 353 472
rect 511 438 545 472
rect 703 438 737 472
rect -737 -472 -703 -438
rect -545 -472 -511 -438
rect -353 -472 -319 -438
rect -161 -472 -127 -438
rect 31 -472 65 -438
rect 223 -472 257 -438
rect 415 -472 449 -438
rect 607 -472 641 -438
<< locali >>
rect -899 540 899 574
rect -899 478 -865 540
rect 865 478 899 540
rect -657 438 -641 472
rect -607 438 -591 472
rect -465 438 -449 472
rect -415 438 -399 472
rect -273 438 -257 472
rect -223 438 -207 472
rect -81 438 -65 472
rect -31 438 -15 472
rect 111 438 127 472
rect 161 438 177 472
rect 303 438 319 472
rect 353 438 369 472
rect 495 438 511 472
rect 545 438 561 472
rect 687 438 703 472
rect 737 438 753 472
rect -785 388 -751 404
rect -785 -404 -751 -388
rect -689 388 -655 404
rect -689 -404 -655 -388
rect -593 388 -559 404
rect -593 -404 -559 -388
rect -497 388 -463 404
rect -497 -404 -463 -388
rect -401 388 -367 404
rect -401 -404 -367 -388
rect -305 388 -271 404
rect -305 -404 -271 -388
rect -209 388 -175 404
rect -209 -404 -175 -388
rect -113 388 -79 404
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 79 388 113 404
rect 79 -404 113 -388
rect 175 388 209 404
rect 175 -404 209 -388
rect 271 388 305 404
rect 271 -404 305 -388
rect 367 388 401 404
rect 367 -404 401 -388
rect 463 388 497 404
rect 463 -404 497 -388
rect 559 388 593 404
rect 559 -404 593 -388
rect 655 388 689 404
rect 655 -404 689 -388
rect 751 388 785 404
rect 751 -404 785 -388
rect -753 -472 -737 -438
rect -703 -472 -687 -438
rect -561 -472 -545 -438
rect -511 -472 -495 -438
rect -369 -472 -353 -438
rect -319 -472 -303 -438
rect -177 -472 -161 -438
rect -127 -472 -111 -438
rect 15 -472 31 -438
rect 65 -472 81 -438
rect 207 -472 223 -438
rect 257 -472 273 -438
rect 399 -472 415 -438
rect 449 -472 465 -438
rect 591 -472 607 -438
rect 641 -472 657 -438
rect -899 -540 -865 -478
rect 865 -540 899 -478
rect -899 -574 -803 -540
rect 803 -574 899 -540
<< viali >>
rect -641 438 -607 472
rect -449 438 -415 472
rect -257 438 -223 472
rect -65 438 -31 472
rect 127 438 161 472
rect 319 438 353 472
rect 511 438 545 472
rect 703 438 737 472
rect -785 -388 -751 388
rect -689 -388 -655 388
rect -593 -388 -559 388
rect -497 -388 -463 388
rect -401 -388 -367 388
rect -305 -388 -271 388
rect -209 -388 -175 388
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect 175 -388 209 388
rect 271 -388 305 388
rect 367 -388 401 388
rect 463 -388 497 388
rect 559 -388 593 388
rect 655 -388 689 388
rect 751 -388 785 388
rect -737 -472 -703 -438
rect -545 -472 -511 -438
rect -353 -472 -319 -438
rect -161 -472 -127 -438
rect 31 -472 65 -438
rect 223 -472 257 -438
rect 415 -472 449 -438
rect 607 -472 641 -438
<< metal1 >>
rect -653 472 -595 478
rect -653 438 -641 472
rect -607 438 -595 472
rect -653 432 -595 438
rect -461 472 -403 478
rect -461 438 -449 472
rect -415 438 -403 472
rect -461 432 -403 438
rect -269 472 -211 478
rect -269 438 -257 472
rect -223 438 -211 472
rect -269 432 -211 438
rect -77 472 -19 478
rect -77 438 -65 472
rect -31 438 -19 472
rect -77 432 -19 438
rect 115 472 173 478
rect 115 438 127 472
rect 161 438 173 472
rect 115 432 173 438
rect 307 472 365 478
rect 307 438 319 472
rect 353 438 365 472
rect 307 432 365 438
rect 499 472 557 478
rect 499 438 511 472
rect 545 438 557 472
rect 499 432 557 438
rect 691 472 749 478
rect 691 438 703 472
rect 737 438 749 472
rect 691 432 749 438
rect -791 388 -745 400
rect -791 -388 -785 388
rect -751 -388 -745 388
rect -791 -400 -745 -388
rect -695 388 -649 400
rect -695 -388 -689 388
rect -655 -388 -649 388
rect -695 -400 -649 -388
rect -599 388 -553 400
rect -599 -388 -593 388
rect -559 -388 -553 388
rect -599 -400 -553 -388
rect -503 388 -457 400
rect -503 -388 -497 388
rect -463 -388 -457 388
rect -503 -400 -457 -388
rect -407 388 -361 400
rect -407 -388 -401 388
rect -367 -388 -361 388
rect -407 -400 -361 -388
rect -311 388 -265 400
rect -311 -388 -305 388
rect -271 -388 -265 388
rect -311 -400 -265 -388
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect -119 388 -73 400
rect -119 -388 -113 388
rect -79 -388 -73 388
rect -119 -400 -73 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 73 388 119 400
rect 73 -388 79 388
rect 113 -388 119 388
rect 73 -400 119 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
rect 265 388 311 400
rect 265 -388 271 388
rect 305 -388 311 388
rect 265 -400 311 -388
rect 361 388 407 400
rect 361 -388 367 388
rect 401 -388 407 388
rect 361 -400 407 -388
rect 457 388 503 400
rect 457 -388 463 388
rect 497 -388 503 388
rect 457 -400 503 -388
rect 553 388 599 400
rect 553 -388 559 388
rect 593 -388 599 388
rect 553 -400 599 -388
rect 649 388 695 400
rect 649 -388 655 388
rect 689 -388 695 388
rect 649 -400 695 -388
rect 745 388 791 400
rect 745 -388 751 388
rect 785 -388 791 388
rect 745 -400 791 -388
rect -749 -438 -691 -432
rect -749 -472 -737 -438
rect -703 -472 -691 -438
rect -749 -478 -691 -472
rect -557 -438 -499 -432
rect -557 -472 -545 -438
rect -511 -472 -499 -438
rect -557 -478 -499 -472
rect -365 -438 -307 -432
rect -365 -472 -353 -438
rect -319 -472 -307 -438
rect -365 -478 -307 -472
rect -173 -438 -115 -432
rect -173 -472 -161 -438
rect -127 -472 -115 -438
rect -173 -478 -115 -472
rect 19 -438 77 -432
rect 19 -472 31 -438
rect 65 -472 77 -438
rect 19 -478 77 -472
rect 211 -438 269 -432
rect 211 -472 223 -438
rect 257 -472 269 -438
rect 211 -478 269 -472
rect 403 -438 461 -432
rect 403 -472 415 -438
rect 449 -472 461 -438
rect 403 -478 461 -472
rect 595 -438 653 -432
rect 595 -472 607 -438
rect 641 -472 653 -438
rect 595 -478 653 -472
<< properties >>
string FIXED_BBOX -882 -557 882 557
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 0.150 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
