magic
tech sky130A
magscale 1 2
timestamp 1665275929
<< metal4 >>
rect -6000 -18137 21000 -18025
rect -6000 -23913 -5888 -18137
rect -112 -23913 15112 -18137
rect 20888 -23913 21000 -18137
rect -6000 -24025 21000 -23913
<< via4 >>
rect -5888 -23913 -112 -18137
rect 15112 -23913 20888 -18137
<< metal5 >>
tri -51477 -3000 -45477 3000 se
rect -45477 -3000 -1523 3000
tri -1523 -3000 4477 3000 sw
tri -55000 -6523 -51477 -3000 se
rect -51477 -4000 -43991 -3000
tri -43991 -4000 -42991 -3000 nw
tri -4009 -4000 -3009 -3000 ne
rect -3009 -4000 4477 -3000
rect -51477 -5414 -45405 -4000
tri -45405 -5414 -43991 -4000 nw
tri -43991 -5414 -42577 -4000 se
rect -42577 -5414 -4423 -4000
tri -4423 -5414 -3009 -4000 sw
tri -3009 -5414 -1595 -4000 ne
rect -1595 -5414 4477 -4000
rect -51477 -6523 -46586 -5414
tri -56486 -8009 -55000 -6523 se
rect -55000 -6595 -46586 -6523
tri -46586 -6595 -45405 -5414 nw
tri -45172 -6595 -43991 -5414 se
rect -43991 -6595 -3009 -5414
rect -55000 -8009 -48000 -6595
tri -48000 -8009 -46586 -6595 nw
tri -46586 -8009 -45172 -6595 se
rect -45172 -6828 -3009 -6595
tri -3009 -6828 -1595 -5414 sw
tri -1595 -6828 -181 -5414 ne
rect -181 -6828 4477 -5414
rect -45172 -7172 -1595 -6828
tri -1595 -7172 -1251 -6828 sw
tri -181 -7172 163 -6828 ne
rect 163 -7172 4477 -6828
rect -45172 -8009 -1251 -7172
tri -59385 -10908 -56486 -8009 se
rect -56486 -9423 -49414 -8009
tri -49414 -9423 -48000 -8009 nw
tri -48000 -9423 -46586 -8009 se
rect -46586 -8586 -1251 -8009
tri -1251 -8586 163 -7172 sw
tri 163 -8586 1577 -7172 ne
rect 1577 -8586 4477 -7172
rect -46586 -9423 163 -8586
rect -56486 -10000 -49991 -9423
tri -49991 -10000 -49414 -9423 nw
tri -48577 -10000 -48000 -9423 se
rect -48000 -10000 163 -9423
tri 163 -10000 1577 -8586 sw
tri 1577 -10000 2991 -8586 ne
rect 2991 -10000 4477 -8586
tri 4477 -10000 11477 -3000 sw
rect -56486 -10908 -50899 -10000
tri -50899 -10908 -49991 -10000 nw
tri -49485 -10908 -48577 -10000 se
rect -48577 -10908 -41092 -10000
tri -61000 -12523 -59385 -10908 se
rect -59385 -12322 -52313 -10908
tri -52313 -12322 -50899 -10908 nw
tri -50899 -12322 -49485 -10908 se
rect -49485 -11000 -41092 -10908
tri -41092 -11000 -40092 -10000 nw
tri -6908 -11000 -5908 -10000 ne
rect -5908 -11000 1577 -10000
rect -49485 -12322 -42414 -11000
tri -42414 -12322 -41092 -11000 nw
tri -41000 -12322 -39678 -11000 se
rect -39678 -11414 -7322 -11000
tri -7322 -11414 -6908 -11000 sw
tri -5908 -11414 -5494 -11000 ne
rect -5494 -11414 1577 -11000
tri 1577 -11414 2991 -10000 sw
tri 2991 -11414 4405 -10000 ne
rect 4405 -11414 11477 -10000
rect -39678 -12322 -6908 -11414
rect -59385 -12523 -52586 -12322
rect -61000 -12595 -52586 -12523
tri -52586 -12595 -52313 -12322 nw
tri -51172 -12595 -50899 -12322 se
rect -50899 -12595 -43828 -12322
rect -61000 -14009 -54000 -12595
tri -54000 -14009 -52586 -12595 nw
tri -52586 -14009 -51172 -12595 se
rect -51172 -13736 -43828 -12595
tri -43828 -13736 -42414 -12322 nw
tri -42414 -13736 -41000 -12322 se
rect -41000 -12414 -6908 -12322
tri -6908 -12414 -5908 -11414 sw
tri -5494 -12414 -4494 -11414 ne
rect -4494 -12414 2991 -11414
rect -41000 -13736 -5908 -12414
rect -51172 -14009 -45242 -13736
rect -61000 -15000 -55000 -14009
rect -56600 -15200 -55000 -15000
tri -55000 -15009 -54000 -14009 nw
tri -53586 -15009 -52586 -14009 se
rect -52586 -15009 -45242 -14009
tri -54000 -15423 -53586 -15009 se
rect -53586 -15150 -45242 -15009
tri -45242 -15150 -43828 -13736 nw
tri -43828 -15150 -42414 -13736 se
rect -42414 -13828 -5908 -13736
tri -5908 -13828 -4494 -12414 sw
tri -4494 -13828 -3080 -12414 ne
rect -3080 -12595 2991 -12414
tri 2991 -12595 4172 -11414 sw
tri 4405 -12595 5586 -11414 ne
rect 5586 -12523 11477 -11414
tri 11477 -12523 14000 -10000 sw
rect 5586 -12595 14000 -12523
rect -3080 -13828 4172 -12595
rect -42414 -14172 -4494 -13828
tri -4494 -14172 -4150 -13828 sw
tri -3080 -14172 -2736 -13828 ne
rect -2736 -14009 4172 -13828
tri 4172 -14009 5586 -12595 sw
tri 5586 -14009 7000 -12595 ne
rect 7000 -14009 14000 -12595
rect -2736 -14172 5586 -14009
rect -42414 -15150 -4150 -14172
rect -53586 -15423 -45586 -15150
rect -54000 -15494 -45586 -15423
tri -45586 -15494 -45242 -15150 nw
tri -44172 -15494 -43828 -15150 se
rect -43828 -15494 -4150 -15150
rect -54000 -16908 -47000 -15494
tri -47000 -16908 -45586 -15494 nw
tri -45586 -16908 -44172 -15494 se
rect -44172 -15586 -4150 -15494
tri -4150 -15586 -2736 -14172 sw
tri -2736 -15586 -1322 -14172 ne
rect -1322 -15423 5586 -14172
tri 5586 -15423 7000 -14009 sw
tri 7000 -15009 8000 -14009 ne
rect -1322 -15586 7000 -15423
rect -44172 -16908 -2736 -15586
rect -54000 -28042 -48000 -16908
tri -48000 -17908 -47000 -16908 nw
tri -47000 -18322 -45586 -16908 se
rect -45586 -17000 -2736 -16908
tri -2736 -17000 -1322 -15586 sw
tri -1322 -17000 92 -15586 ne
rect 92 -17000 7000 -15586
rect -45586 -18322 -41000 -17000
rect -47000 -26627 -41000 -18322
tri -41000 -20808 -37192 -17000 nw
tri -9808 -18137 -8671 -17000 ne
rect -8671 -18025 -1322 -17000
tri -1322 -18025 -297 -17000 sw
tri 92 -17908 1000 -17000 ne
rect -8671 -18137 0 -18025
tri -8671 -20808 -6000 -18137 ne
rect -6000 -23913 -5888 -18137
rect -112 -23913 0 -18137
rect -6000 -24025 0 -23913
tri -48000 -28042 -47000 -27042 sw
tri -47000 -28042 -45585 -26627 ne
rect -45585 -28042 -41000 -26627
rect -54000 -28585 -47000 -28042
tri -47000 -28585 -46457 -28042 sw
tri -45585 -28585 -45042 -28042 ne
rect -45042 -28585 -41000 -28042
rect -54000 -29527 -46457 -28585
tri -54000 -30000 -53527 -29527 ne
rect -53527 -30000 -46457 -29527
tri -46457 -30000 -45042 -28585 sw
tri -45042 -30000 -43627 -28585 ne
rect -43627 -30000 -41000 -28585
tri -41000 -30000 -35142 -24142 sw
tri -4858 -30000 1000 -24142 se
rect 1000 -26627 7000 -17000
rect 1000 -28042 5585 -26627
tri 5585 -28042 7000 -26627 nw
tri 7000 -28042 8000 -27042 se
rect 8000 -28042 14000 -14009
rect 15000 -18137 21000 -18025
rect 15000 -23913 15112 -18137
rect 20888 -23913 21000 -18137
rect 15000 -24025 21000 -23913
rect 1000 -28585 5042 -28042
tri 5042 -28585 5585 -28042 nw
tri 6457 -28585 7000 -28042 se
rect 7000 -28585 14000 -28042
rect 1000 -30000 3627 -28585
tri 3627 -30000 5042 -28585 nw
tri 5042 -30000 6457 -28585 se
rect 6457 -29527 14000 -28585
rect 6457 -30000 6527 -29527
tri -53527 -31415 -52112 -30000 ne
rect -52112 -31415 -45042 -30000
tri -45042 -31415 -43627 -30000 sw
tri -43627 -31415 -42212 -30000 ne
rect -42212 -31212 2415 -30000
tri 2415 -31212 3627 -30000 nw
tri 3830 -31212 5042 -30000 se
rect 5042 -31212 6527 -30000
rect -42212 -31415 1000 -31212
tri -52112 -32830 -50697 -31415 ne
rect -50697 -32830 -43627 -31415
tri -43627 -32830 -42212 -31415 sw
tri -42212 -32830 -40797 -31415 ne
rect -40797 -32627 1000 -31415
tri 1000 -32627 2415 -31212 nw
tri 2415 -32627 3830 -31212 se
rect 3830 -32627 6527 -31212
rect -40797 -32830 -415 -32627
tri -50697 -33464 -50063 -32830 ne
rect -50063 -33170 -42212 -32830
tri -42212 -33170 -41872 -32830 sw
tri -40797 -33170 -40457 -32830 ne
rect -40457 -33170 -415 -32830
rect -50063 -33464 -41872 -33170
tri -50063 -34585 -48942 -33464 ne
rect -48942 -34042 -41872 -33464
tri -41872 -34042 -41000 -33170 sw
tri -40457 -34042 -39585 -33170 ne
rect -39585 -34042 -415 -33170
tri -415 -34042 1000 -32627 nw
tri 1000 -34042 2415 -32627 se
rect 2415 -34042 6527 -32627
rect -48942 -34585 -41000 -34042
tri -41000 -34585 -40457 -34042 sw
tri -39585 -34585 -39042 -34042 ne
rect -39042 -34585 -958 -34042
tri -958 -34585 -415 -34042 nw
tri 457 -34585 1000 -34042 se
rect 1000 -34585 6527 -34042
tri -48942 -35527 -48000 -34585 ne
rect -48000 -35527 -40457 -34585
tri -48000 -37000 -46527 -35527 ne
rect -46527 -36000 -40457 -35527
tri -40457 -36000 -39042 -34585 sw
tri -39042 -36000 -37627 -34585 ne
rect -37627 -36000 -2373 -34585
tri -2373 -36000 -958 -34585 nw
tri -958 -36000 457 -34585 se
rect 457 -36000 6527 -34585
rect -46527 -37000 -39042 -36000
tri -39042 -37000 -38042 -36000 sw
tri -1958 -37000 -958 -36000 se
rect -958 -37000 6527 -36000
tri 6527 -37000 14000 -29527 nw
tri -46527 -43000 -40527 -37000 ne
rect -40527 -43000 527 -37000
tri 527 -43000 6527 -37000 nw
<< end >>
