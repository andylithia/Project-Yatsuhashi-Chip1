magic
tech sky130B
timestamp 1659324110
<< metal4 >>
rect 6800 3550 7900 3600
rect 2900 3400 3700 3500
rect 2900 2900 3000 3400
rect 3600 2900 3700 3400
rect 6800 2950 6850 3550
rect 7450 2950 7900 3550
rect 6800 2900 7900 2950
rect 2900 2800 3700 2900
<< via4 >>
rect 3000 2900 3600 3400
rect 6850 2950 7450 3550
<< metal5 >>
rect 0 6000 6500 6500
rect 0 -300 500 6000
rect 800 5200 5700 5700
rect 800 500 1300 5200
rect 1600 4400 4900 4900
rect 1600 1300 2100 4400
rect 2400 3400 3700 3500
rect 2400 2900 3000 3400
rect 3600 2900 3700 3400
rect 2400 2800 3700 2900
rect 2400 2100 2900 2800
rect 4400 2100 4900 4400
rect 2400 1600 4900 2100
rect 5200 1300 5700 5200
rect 1600 800 5700 1300
rect 6000 500 6500 6000
rect 800 0 6500 500
rect 6800 3550 7500 3600
rect 6800 2950 6850 3550
rect 7450 2950 7500 3550
rect 6800 2900 7500 2950
rect 6800 2850 7450 2900
rect 6800 2800 7400 2850
rect 6800 2750 7350 2800
rect 6800 -300 7300 2750
rect 0 -800 7300 -300
<< labels >>
rlabel metal5 2900 2800 3700 3500 1 B
rlabel metal4 7500 2900 7900 3600 1 A
<< end >>
