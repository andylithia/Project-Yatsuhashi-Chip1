magic
tech sky130A
timestamp 1658705077
<< metal2 >>
rect 0 1100 600 1200
rect 0 900 100 1100
rect 500 900 600 1100
rect 0 800 600 900
rect 0 -100 200 800
rect 400 -100 600 800
rect 0 -200 600 -100
rect 0 -400 100 -200
rect 500 -400 600 -200
rect 0 -500 600 -400
<< via2 >>
rect 100 900 500 1100
rect 100 -400 500 -200
<< metal3 >>
rect 0 1100 600 1200
rect 0 900 100 1100
rect 500 900 600 1100
rect 0 800 600 900
rect 0 -100 200 800
rect 400 -100 600 800
rect 0 -200 600 -100
rect 0 -400 100 -200
rect 500 -400 600 -200
rect 0 -500 600 -400
<< via3 >>
rect 100 900 500 1100
rect 100 -400 500 -200
<< metal4 >>
rect 0 1100 600 1200
rect 0 900 100 1100
rect 500 900 600 1100
rect 0 800 600 900
rect 0 -200 600 -100
rect 0 -400 100 -200
rect 500 -400 600 -200
rect 0 -500 600 -400
<< via4 >>
rect 100 900 500 1100
rect 100 -400 500 -200
<< metal5 >>
rect 0 1100 600 1200
rect 0 900 100 1100
rect 500 900 600 1100
rect 0 800 600 900
rect 0 200 600 500
rect 0 -200 600 -100
rect 0 -400 100 -200
rect 500 -400 600 -200
rect 0 -500 600 -400
<< labels >>
rlabel metal5 500 800 600 1200 1 gnd
rlabel metal5 0 200 100 500 1 l
rlabel metal5 500 200 600 500 1 r
<< end >>
