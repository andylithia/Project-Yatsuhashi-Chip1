* NGSPICE file created from ./CLASSE/cascode_complete_3_flat.ext - technology: sky130A

X0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t239 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t238 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t239 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t237 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t236 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__res_high_po_0p35 l=1.6e+06u
X18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t235 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t234 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t233 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t232 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t238 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t231 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t230 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t237 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t229 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t236 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t228 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t227 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t235 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t234 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t233 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t226 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t232 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t231 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t225 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t230 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t224 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t223 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t225 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t229 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t228 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t222 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t224 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t227 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t226 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t221 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t220 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t225 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t224 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t219 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t223 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t222 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t221 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t120 sky130_fd_pr__cap_mim_m3_2 l=2.5e+07u w=3.9e+07u
X117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t220 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t219 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t218 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t218 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t231 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t217 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t217 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t230 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 sky130_fd_pr__cap_mim_m3_2 l=2.5e+07u w=2e+07u
X142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
R0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 sky130_fd_pr__res_generic_po w=330000u l=6.5e+06u
X144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
R1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 sky130_fd_pr__res_generic_po w=330000u l=6.5e+06u
X161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t233 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
R2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 sky130_fd_pr__res_generic_po w=330000u l=6.5e+06u
X184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t232 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X217 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X218 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X219 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X220 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X221 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X222 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X223 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X224 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X225 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X226 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X227 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X228 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X229 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X230 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X231 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X232 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X233 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X234 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X235 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X236 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X237 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X238 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X239 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X240 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X241 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X242 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X243 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X244 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X245 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X246 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t0 sky130_fd_pr__cap_mim_m3_2 l=2.5e+07u w=3.9e+07u
X247 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X248 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X249 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X250 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X251 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X252 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X253 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X254 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X255 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X256 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X257 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X258 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X259 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X260 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X261 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X262 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X263 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X264 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X265 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X266 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X267 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X268 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X269 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X270 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X271 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X272 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X273 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X274 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X275 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X276 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X277 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X278 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X279 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X280 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X281 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X282 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X283 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X284 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X285 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X286 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X287 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X288 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X289 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X290 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X291 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X292 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X293 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X294 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X295 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X296 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X297 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X298 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X299 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X300 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X301 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X302 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X303 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X304 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X305 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X306 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X307 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X308 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X309 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X310 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X311 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X312 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X313 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X314 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X315 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X316 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X317 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X318 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X319 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X320 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X321 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X322 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X323 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X324 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X325 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X326 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X327 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X328 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X329 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X330 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X331 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X332 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X333 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X334 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X335 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X336 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X337 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X338 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X339 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X340 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X341 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X342 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X343 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X344 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X345 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X346 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X347 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t3 sky130_fd_pr__cap_mim_m3_2 l=5.2e+07u w=2.3e+07u
X348 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X349 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X350 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X351 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X352 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X353 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X354 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X355 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X356 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X357 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X358 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X359 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X360 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X361 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X362 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X363 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X364 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X365 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X366 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X367 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X368 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X369 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X370 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X371 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X372 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X373 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X374 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X375 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X376 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X377 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X378 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X379 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X380 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X381 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X382 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X383 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X384 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X385 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X386 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X387 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X388 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X389 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X390 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X391 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X392 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X393 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X394 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X395 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X396 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X397 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X398 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X399 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X400 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X401 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X402 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X403 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X404 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X405 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X406 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X407 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X408 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X409 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X410 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X411 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X412 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X413 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X414 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X415 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X416 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X417 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t227 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X418 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X419 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X420 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t226 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X421 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X422 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X423 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X424 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X425 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t217 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X426 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X427 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X428 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X429 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X430 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X431 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X432 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X433 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X434 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X435 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X436 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X437 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X438 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X439 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X440 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X441 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X442 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X443 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X444 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X445 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X446 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X447 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X448 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X449 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X450 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X451 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X452 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X453 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X454 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X455 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t235 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X456 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X457 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X458 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X459 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X460 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X461 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X462 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X463 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X464 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X465 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X466 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X467 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t234 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X468 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X469 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X470 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X471 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X472 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X473 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X474 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X475 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X476 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X477 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t219 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X478 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X479 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X480 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t218 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X481 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X482 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X483 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X484 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X485 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X486 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X487 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X488 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X489 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X490 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X491 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X492 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X493 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X494 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X495 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X496 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X497 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X498 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t237 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X499 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X500 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X501 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X502 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X503 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X504 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X505 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__res_high_po w=350000u l=1.6e+06u
X506 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X507 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t236 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X508 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t221 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X509 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X510 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X511 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X512 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X513 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X514 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X515 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X516 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X517 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X518 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X519 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X520 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X521 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X522 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X523 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X524 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X525 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X526 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X527 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X528 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X529 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t220 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X530 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X531 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X532 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X533 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X534 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X535 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X536 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X537 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X538 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X539 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X540 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X541 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X542 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X543 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X544 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X545 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
R3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 sky130_fd_pr__res_generic_po w=330000u l=6.5e+06u
X546 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X547 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X548 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X549 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X550 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X551 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X552 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X553 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X554 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X555 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X556 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X557 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X558 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X559 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X560 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X561 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X562 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X563 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X564 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X565 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X566 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X567 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X568 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X569 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X570 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X571 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X572 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X573 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X574 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X575 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X576 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X577 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X578 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X579 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X580 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X581 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X582 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X583 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X584 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X585 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X586 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X587 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X588 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X589 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X590 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X591 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X592 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X593 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X594 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X595 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X596 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X597 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X598 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X599 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X600 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X601 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X602 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X603 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X604 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X605 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X606 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X607 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X608 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X609 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X610 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X611 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X612 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X613 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X614 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X615 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X616 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X617 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X618 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X619 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X620 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X621 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X622 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X623 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X624 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X625 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X626 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X627 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X628 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X629 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X630 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X631 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X632 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X633 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X634 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X635 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X636 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X637 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X638 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X639 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X640 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X641 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X642 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X643 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X644 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X645 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X646 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t1 sky130_fd_pr__cap_mim_m3_2 l=5.2e+07u w=8e+06u
X647 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X648 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X649 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t229 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X650 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X651 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X652 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X653 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X654 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X655 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X656 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t228 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X657 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X658 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X659 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X660 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X661 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X662 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X663 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X664 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X665 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X666 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X667 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t223 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X668 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t222 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X669 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X670 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X671 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X672 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X673 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X674 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X675 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X676 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X677 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X678 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X679 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X680 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X681 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X682 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X683 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X684 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X685 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X686 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X687 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X688 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X689 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X690 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X691 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X692 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X693 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X694 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X695 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X696 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X697 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X698 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X699 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X700 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X701 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X702 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X703 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t123 sky130_fd_pr__cap_mim_m3_2 l=5.2e+07u w=2.3e+07u
X704 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X705 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X706 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X707 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X708 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X709 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X710 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X711 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X712 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X713 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X714 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t239 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X715 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X716 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X717 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X718 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X719 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X720 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X721 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X722 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 sky130_fd_pr__cap_mim_m3_2 l=2.5e+07u w=2e+07u
X723 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X724 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X725 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X726 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t238 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X727 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t121 sky130_fd_pr__cap_mim_m3_2 l=5.2e+07u w=8e+06u
X728 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X729 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
C0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 89.46fF
C1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G 96.34fF
C2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 837.22fF
C3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 136.24fF
C4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 831.50fF
C5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G 21.28fF
C6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 110.88fF
C7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G 33.77fF
C8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 89.53fF
C9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G 14.33fF
C10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G 100.66fF
C11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 103.99fF
C12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G 33.77fF
C13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 110.88fF
C14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 94.93fF
C15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 37.67fF
C16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G 17.28fF
C17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G 95.91fF
C18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 113.57fF
C19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 135.82fF
C20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G 16.33fF
C21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G 13.23fF
C22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G 28.21fF
C23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 56.34fF
C24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G 96.60fF
C25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 886.00fF
C26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 97.88fF
C27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 832.19fF
C28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 935.79fF
C29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 16.33fF
C30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 132.68fF
C31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 4.98fF
C32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 98.97fF
C33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 37.51fF
C34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 16.01fF
C35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 4.98fF
C36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 45.03fF
C37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G 29.89fF
C38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 882.00fF
C39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 16.70fF
C40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 103.03fF
C41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 126.91fF
R4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t122 9.377
R5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t31 1.965
R6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t62 1.965
R7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t89 1.963
R8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t39 1.96
R9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n35 1.435
R10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n64 1.435
R11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n31 1.428
R12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n32 1.428
R13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n33 1.428
R14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n34 1.428
R15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n30 1.428
R16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n29 1.428
R17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n28 1.428
R18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n27 1.428
R19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n26 1.428
R20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n25 1.428
R21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n60 1.428
R22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n61 1.428
R23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n62 1.428
R24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n63 1.428
R25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n59 1.428
R26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n58 1.428
R27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n57 1.428
R28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n56 1.428
R29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n55 1.428
R30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n54 1.428
R31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n20 1.414
R32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n19 1.414
R33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n18 1.414
R34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n17 1.414
R35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n16 1.414
R36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n15 1.414
R37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n14 1.414
R38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n13 1.414
R39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n12 1.414
R40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n11 1.414
R41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n50 1.414
R42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n49 1.414
R43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n48 1.414
R44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n47 1.414
R45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n46 1.414
R46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n45 1.414
R47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n44 1.414
R48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n43 1.414
R49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n42 1.414
R50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n41 1.414
R51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n40 1.414
R52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n72 1.413
R53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n21 1.412
R54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n22 1.412
R55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n23 1.412
R56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n51 1.41
R57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n52 1.409
R58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n53 1.409
R59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n36 1.28
R60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n37 1.28
R61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n38 1.28
R62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n39 1.28
R63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n65 1.28
R64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n66 1.28
R65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n67 1.28
R66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n68 1.28
R67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t105 0.551
R68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t108 0.551
R69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t20 0.551
R70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t69 0.551
R71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t77 0.551
R72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t32 0.551
R73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t87 0.551
R74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t36 0.551
R75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t21 0.551
R76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t24 0.551
R77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t1 0.551
R78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t3 0.551
R79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t88 0.551
R80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t13 0.551
R81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t82 0.551
R82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t19 0.551
R83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t51 0.551
R84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t107 0.551
R85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t25 0.551
R86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t70 0.551
R87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t56 0.551
R88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t94 0.551
R89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t119 0.551
R90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t111 0.551
R91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t65 0.551
R92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t79 0.551
R93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t63 0.551
R94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t2 0.551
R95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t6 0.551
R96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t33 0.551
R97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t45 0.551
R98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t113 0.551
R99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t97 0.551
R100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t93 0.551
R101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t83 0.551
R102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t106 0.551
R103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t59 0.551
R104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t112 0.551
R105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t72 0.551
R106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t14 0.551
R107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t58 0.551
R108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t92 0.551
R109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t61 0.551
R110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t26 0.551
R111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t30 0.551
R112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t46 0.551
R113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t47 0.551
R114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t60 0.551
R115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t27 0.551
R116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t76 0.551
R117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t68 0.551
R118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t23 0.551
R119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t16 0.551
R120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t49 0.551
R121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t64 0.551
R122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t85 0.551
R123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t5 0.551
R124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t17 0.551
R125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t100 0.551
R126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t71 0.551
R127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t22 0.551
R128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t86 0.551
R129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t66 0.551
R130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t67 0.551
R131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t9 0.551
R132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t43 0.551
R133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t90 0.551
R134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t41 0.551
R135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t37 0.551
R136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t81 0.551
R137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t80 0.551
R138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t117 0.551
R139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t54 0.551
R140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t99 0.551
R141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t104 0.551
R142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t44 0.551
R143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t8 0.551
R144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t91 0.551
R145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t95 0.551
R146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t4 0.551
R147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t118 0.551
R148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t12 0.551
R149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t38 0.551
R150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t96 0.551
R151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t78 0.551
R152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t53 0.551
R153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t15 0.551
R154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t98 0.551
R155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t110 0.551
R156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t73 0.551
R157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t29 0.551
R158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t42 0.551
R159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t115 0.551
R160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t40 0.551
R161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t34 0.551
R162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t101 0.551
R163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t57 0.551
R164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t50 0.551
R165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t52 0.551
R166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t18 0.551
R167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t7 0.551
R168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t74 0.551
R169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t55 0.551
R170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t84 0.551
R171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t114 0.551
R172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t109 0.551
R173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t35 0.551
R174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t75 0.551
R175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t116 0.551
R176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t11 0.551
R177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t102 0.551
R178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t48 0.551
R179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t10 0.551
R180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t28 0.551
R181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t103 0.551
R182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t0 0.551
R183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 0.349
R184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 0.306
R185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n71 0.279
R186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t121 0.231
R187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 0.18
R188 VSSH cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n70 0.154
R189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n24 0.137
R190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n69 0.091
R191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t123 0.061
R192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n6 0.043
R193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 0.042
R194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n71 VSSH 0.034
R195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD1 0.028
R196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD1 0.028
R197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n1 0.028
R198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n2 0.028
R199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 0.027
R200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t120 0.022
R201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n9 0.021
R202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n7 0.021
R203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n10 0.016
R204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n8 0.016
R205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n214 2.204
R206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n212 2.204
R207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n183 2.204
R208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t113 1.965
R209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t180 1.965
R210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t57 1.965
R211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t164 1.965
R212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t43 1.963
R213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t215 1.963
R214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t80 1.963
R215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t191 1.96
R216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n197 1.435
R217 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n95 1.435
R218 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n169 1.435
R219 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n16 1.435
R220 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n188 1.428
R221 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n189 1.428
R222 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n190 1.428
R223 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n191 1.428
R224 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n192 1.428
R225 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n193 1.428
R226 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n194 1.428
R227 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n195 1.428
R228 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n196 1.428
R229 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n91 1.428
R230 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n92 1.428
R231 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n93 1.428
R232 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n94 1.428
R233 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n84 1.428
R234 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n83 1.428
R235 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n82 1.428
R236 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n81 1.428
R237 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n80 1.428
R238 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n79 1.428
R239 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n159 1.428
R240 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n160 1.428
R241 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n161 1.428
R242 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n162 1.428
R243 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n163 1.428
R244 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n164 1.428
R245 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n165 1.428
R246 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n166 1.428
R247 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n167 1.428
R248 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n168 1.428
R249 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n12 1.428
R250 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n13 1.428
R251 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n14 1.428
R252 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n15 1.428
R253 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n5 1.428
R254 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n4 1.428
R255 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n3 1.428
R256 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n2 1.428
R257 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n1 1.428
R258 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n0 1.428
R259 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n202 1.427
R260 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n62 1.414
R261 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n61 1.414
R262 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n60 1.414
R263 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n59 1.414
R264 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n58 1.414
R265 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n57 1.414
R266 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n56 1.414
R267 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n55 1.414
R268 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n54 1.414
R269 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n53 1.414
R270 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n52 1.414
R271 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n105 1.414
R272 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n106 1.414
R273 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n107 1.414
R274 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n108 1.414
R275 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n109 1.414
R276 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n110 1.414
R277 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n111 1.414
R278 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n112 1.414
R279 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n113 1.414
R280 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n114 1.414
R281 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n115 1.414
R282 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n131 1.414
R283 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n132 1.414
R284 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n133 1.414
R285 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n134 1.414
R286 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n135 1.414
R287 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n136 1.414
R288 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n137 1.414
R289 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n138 1.414
R290 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n139 1.414
R291 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n140 1.414
R292 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n141 1.414
R293 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n26 1.414
R294 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n27 1.414
R295 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n28 1.414
R296 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n29 1.414
R297 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n30 1.414
R298 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n31 1.414
R299 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n32 1.414
R300 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n33 1.414
R301 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n34 1.414
R302 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n35 1.414
R303 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n36 1.414
R304 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n129 1.412
R305 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n128 1.412
R306 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n127 1.412
R307 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n155 1.412
R308 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n154 1.412
R309 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n153 1.412
R310 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n50 1.412
R311 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n49 1.412
R312 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n48 1.412
R313 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n74 1.41
R314 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n76 1.409
R315 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n77 1.409
R316 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n183 1.302
R317 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n212 1.302
R318 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n214 1.302
R319 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n209 1.282
R320 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n180 1.282
R321 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n100 1.28
R322 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n101 1.28
R323 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n102 1.28
R324 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n103 1.28
R325 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n21 1.28
R326 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n22 1.28
R327 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n23 1.28
R328 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n24 1.28
R329 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n187 1.278
R330 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n157 1.278
R331 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n158 1.278
R332 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t71 0.551
R333 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t103 0.551
R334 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t23 0.551
R335 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t77 0.551
R336 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t56 0.551
R337 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t116 0.551
R338 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t111 0.551
R339 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t15 0.551
R340 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t51 0.551
R341 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t81 0.551
R342 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t0 0.551
R343 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t62 0.551
R344 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t30 0.551
R345 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t90 0.551
R346 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t105 0.551
R347 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t11 0.551
R348 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t96 0.551
R349 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t73 0.551
R350 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t40 0.551
R351 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t68 0.551
R352 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t76 0.551
R353 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t110 0.551
R354 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t66 0.551
R355 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t6 0.551
R356 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t36 0.551
R357 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t33 0.551
R358 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t93 0.551
R359 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t4 0.551
R360 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t238 0.551
R361 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t220 0.551
R362 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t125 0.551
R363 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t121 0.551
R364 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t142 0.551
R365 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t147 0.551
R366 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t199 0.551
R367 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t127 0.551
R368 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t175 0.551
R369 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t139 0.551
R370 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t223 0.551
R371 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t206 0.551
R372 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t124 0.551
R373 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t140 0.551
R374 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t225 0.551
R375 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t189 0.551
R376 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t227 0.551
R377 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t126 0.551
R378 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t232 0.551
R379 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t152 0.551
R380 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t222 0.551
R381 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t149 0.551
R382 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t205 0.551
R383 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t193 0.551
R384 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t171 0.551
R385 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t187 0.551
R386 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t181 0.551
R387 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t169 0.551
R388 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t176 0.551
R389 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t184 0.551
R390 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t197 0.551
R391 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t178 0.551
R392 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t130 0.551
R393 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t165 0.551
R394 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t173 0.551
R395 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t158 0.551
R396 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t203 0.551
R397 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t237 0.551
R398 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t143 0.551
R399 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t123 0.551
R400 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t150 0.551
R401 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t137 0.551
R402 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t217 0.551
R403 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t153 0.551
R404 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t228 0.551
R405 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t207 0.551
R406 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t135 0.551
R407 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t141 0.551
R408 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t155 0.551
R409 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t168 0.551
R410 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t210 0.551
R411 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t208 0.551
R412 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t177 0.551
R413 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t182 0.551
R414 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t170 0.551
R415 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t129 0.551
R416 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t204 0.551
R417 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t172 0.551
R418 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t94 0.551
R419 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t5 0.551
R420 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t26 0.551
R421 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t49 0.551
R422 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t3 0.551
R423 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t55 0.551
R424 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t85 0.551
R425 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t114 0.551
R426 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t19 0.551
R427 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t39 0.551
R428 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t102 0.551
R429 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t44 0.551
R430 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t109 0.551
R431 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t101 0.551
R432 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t10 0.551
R433 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t59 0.551
R434 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t88 0.551
R435 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t65 0.551
R436 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t60 0.551
R437 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t2 0.551
R438 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t25 0.551
R439 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t50 0.551
R440 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t72 0.551
R441 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t104 0.551
R442 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t34 0.551
R443 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t61 0.551
R444 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t14 0.551
R445 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t32 0.551
R446 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t52 0.551
R447 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t82 0.551
R448 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t84 0.551
R449 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t21 0.551
R450 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t1 0.551
R451 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t53 0.551
R452 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t64 0.551
R453 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t91 0.551
R454 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t92 0.551
R455 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t35 0.551
R456 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t12 0.551
R457 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t31 0.551
R458 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t75 0.551
R459 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t108 0.551
R460 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t70 0.551
R461 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t45 0.551
R462 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t22 0.551
R463 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t42 0.551
R464 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t54 0.551
R465 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t115 0.551
R466 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t83 0.551
R467 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t27 0.551
R468 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t20 0.551
R469 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t41 0.551
R470 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t13 0.551
R471 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t63 0.551
R472 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t107 0.551
R473 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t98 0.551
R474 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t74 0.551
R475 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t106 0.551
R476 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t148 0.551
R477 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t211 0.551
R478 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t128 0.551
R479 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t198 0.551
R480 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t122 0.551
R481 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t195 0.551
R482 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t188 0.551
R483 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t134 0.551
R484 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t133 0.551
R485 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t186 0.551
R486 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t235 0.551
R487 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t179 0.551
R488 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t156 0.551
R489 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t219 0.551
R490 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t214 0.551
R491 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t212 0.551
R492 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t166 0.551
R493 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t190 0.551
R494 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t224 0.551
R495 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t230 0.551
R496 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t167 0.551
R497 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t183 0.551
R498 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t239 0.551
R499 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t163 0.551
R500 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t145 0.551
R501 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t157 0.551
R502 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t209 0.551
R503 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t161 0.551
R504 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t226 0.551
R505 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t231 0.551
R506 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t229 0.551
R507 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t138 0.551
R508 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t216 0.551
R509 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t196 0.551
R510 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t194 0.551
R511 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t192 0.551
R512 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t236 0.551
R513 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t120 0.551
R514 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t131 0.551
R515 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t200 0.551
R516 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t136 0.551
R517 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t159 0.551
R518 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t213 0.551
R519 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t144 0.551
R520 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t234 0.551
R521 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t233 0.551
R522 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t202 0.551
R523 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t221 0.551
R524 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t218 0.551
R525 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t162 0.551
R526 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t151 0.551
R527 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t174 0.551
R528 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t185 0.551
R529 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t132 0.551
R530 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t201 0.551
R531 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t160 0.551
R532 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t146 0.551
R533 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t154 0.551
R534 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t9 0.551
R535 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t69 0.551
R536 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t100 0.551
R537 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t8 0.551
R538 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t29 0.551
R539 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t87 0.551
R540 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t118 0.551
R541 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t58 0.551
R542 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t86 0.551
R543 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t117 0.551
R544 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t47 0.551
R545 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t79 0.551
R546 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t17 0.551
R547 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t46 0.551
R548 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t78 0.551
R549 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t16 0.551
R550 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t38 0.551
R551 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t99 0.551
R552 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t95 0.551
R553 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t28 0.551
R554 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t97 0.551
R555 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t7 0.551
R556 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t24 0.551
R557 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t48 0.551
R558 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t112 0.551
R559 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t18 0.551
R560 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t37 0.551
R561 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t67 0.551
R562 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t89 0.551
R563 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t119 0.551
R564 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n213 0.46
R565 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n211 0.46
R566 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n182 0.46
R567 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n156 0.429
R568 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n78 0.35
R569 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n130 0.347
R570 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n51 0.347
R571 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n104 0.224
R572 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n25 0.224
R573 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n185 0.091
R574 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n186 0.078
R575 cascode_1_0/SD2R cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n216 0.054
R576 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1 0.05
R577 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 0.05
R578 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n184 0.039
R579 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n215 0.039
R580 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n73 0.007
R581 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n72 0.007
R582 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n71 0.007
R583 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n70 0.007
R584 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n69 0.007
R585 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n68 0.007
R586 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n67 0.007
R587 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n66 0.007
R588 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n65 0.007
R589 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n64 0.007
R590 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n63 0.007
R591 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD2 0.007
R592 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n96 0.007
R593 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n97 0.007
R594 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n98 0.007
R595 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n89 0.007
R596 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n88 0.007
R597 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n87 0.007
R598 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n86 0.007
R599 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n85 0.007
R600 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n125 0.007
R601 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n124 0.007
R602 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n123 0.007
R603 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n122 0.007
R604 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n121 0.007
R605 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n120 0.007
R606 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n119 0.007
R607 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n118 0.007
R608 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n117 0.007
R609 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n116 0.007
R610 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD2 0.007
R611 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n170 0.007
R612 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n171 0.007
R613 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n172 0.007
R614 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n173 0.007
R615 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n174 0.007
R616 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n175 0.007
R617 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n176 0.007
R618 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n177 0.007
R619 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n178 0.007
R620 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n179 0.007
R621 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n151 0.007
R622 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n150 0.007
R623 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n149 0.007
R624 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n148 0.007
R625 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n147 0.007
R626 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n146 0.007
R627 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n145 0.007
R628 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n144 0.007
R629 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n143 0.007
R630 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n142 0.007
R631 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD2 0.007
R632 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n17 0.007
R633 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n18 0.007
R634 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n19 0.007
R635 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n10 0.007
R636 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n9 0.007
R637 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n8 0.007
R638 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n7 0.007
R639 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n6 0.007
R640 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n46 0.007
R641 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n45 0.007
R642 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n44 0.007
R643 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n43 0.007
R644 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n42 0.007
R645 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n41 0.007
R646 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n40 0.007
R647 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n39 0.007
R648 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n38 0.007
R649 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n37 0.007
R650 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD2 0.007
R651 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n198 0.007
R652 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n199 0.007
R653 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n200 0.007
R654 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n201 0.007
R655 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n203 0.007
R656 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n204 0.007
R657 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n205 0.007
R658 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n206 0.007
R659 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n207 0.007
R660 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n208 0.007
R661 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n126 0.006
R662 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n152 0.006
R663 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n47 0.006
R664 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n99 0.005
R665 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n20 0.005
R666 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n90 0.004
R667 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n11 0.004
R668 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/SD1 0.003
R669 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 0.003
R670 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n181 0.003
R671 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n210 0.003
R672 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n75 0.001
R673 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 3.41
R674 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 3.41
R675 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n11 2.204
R676 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n10 2.204
R677 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n13 2.204
R678 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n12 2.204
R679 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t104 1.972
R680 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t68 1.972
R681 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t116 1.965
R682 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t26 1.965
R683 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n38 1.435
R684 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n68 1.435
R685 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n28 1.428
R686 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n29 1.428
R687 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n30 1.428
R688 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n31 1.428
R689 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n32 1.428
R690 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n33 1.428
R691 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n34 1.428
R692 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n35 1.428
R693 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n36 1.428
R694 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n37 1.428
R695 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n58 1.428
R696 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n59 1.428
R697 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n60 1.428
R698 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n61 1.428
R699 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n62 1.428
R700 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n63 1.428
R701 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n64 1.428
R702 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n65 1.428
R703 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n66 1.428
R704 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n67 1.428
R705 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n20 1.414
R706 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n21 1.414
R707 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n22 1.414
R708 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n23 1.414
R709 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n24 1.414
R710 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n14 1.414
R711 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n15 1.414
R712 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n16 1.414
R713 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n17 1.414
R714 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n18 1.414
R715 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n47 1.414
R716 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n48 1.414
R717 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n49 1.414
R718 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n50 1.414
R719 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n51 1.414
R720 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n46 1.414
R721 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n45 1.414
R722 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n44 1.414
R723 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n43 1.414
R724 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n42 1.414
R725 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n55 1.412
R726 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n54 1.412
R727 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n53 1.412
R728 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n52 1.412
R729 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n75 1.412
R730 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n74 1.412
R731 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n25 1.412
R732 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n19 1.41
R733 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n10 1.302
R734 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n11 1.302
R735 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n12 1.302
R736 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n13 1.302
R737 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n26 1.278
R738 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n27 1.278
R739 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n56 1.278
R740 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n57 1.278
R741 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n73 0.573
R742 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t69 0.551
R743 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t62 0.551
R744 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t109 0.551
R745 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t34 0.551
R746 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t95 0.551
R747 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t61 0.551
R748 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t19 0.551
R749 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t57 0.551
R750 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t8 0.551
R751 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t87 0.551
R752 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t28 0.551
R753 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t59 0.551
R754 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t35 0.551
R755 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t24 0.551
R756 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t92 0.551
R757 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t30 0.551
R758 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t103 0.551
R759 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t23 0.551
R760 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t56 0.551
R761 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t112 0.551
R762 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t70 0.551
R763 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t119 0.551
R764 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t10 0.551
R765 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t114 0.551
R766 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t106 0.551
R767 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t101 0.551
R768 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t105 0.551
R769 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t46 0.551
R770 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t41 0.551
R771 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t52 0.551
R772 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t118 0.551
R773 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t82 0.551
R774 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t11 0.551
R775 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t115 0.551
R776 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t27 0.551
R777 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t9 0.551
R778 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t2 0.551
R779 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t89 0.551
R780 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t14 0.551
R781 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t17 0.551
R782 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t74 0.551
R783 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t72 0.551
R784 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t79 0.551
R785 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t63 0.551
R786 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t78 0.551
R787 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t96 0.551
R788 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t110 0.551
R789 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t55 0.551
R790 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t36 0.551
R791 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t88 0.551
R792 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t13 0.551
R793 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t83 0.551
R794 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t42 0.551
R795 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t53 0.551
R796 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t18 0.551
R797 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t7 0.551
R798 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t4 0.551
R799 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t12 0.551
R800 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t60 0.551
R801 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t84 0.551
R802 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t71 0.551
R803 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t29 0.551
R804 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t94 0.551
R805 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t16 0.551
R806 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t25 0.551
R807 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t44 0.551
R808 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t33 0.551
R809 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t77 0.551
R810 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t50 0.551
R811 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t39 0.551
R812 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t45 0.551
R813 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t67 0.551
R814 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t85 0.551
R815 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t37 0.551
R816 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t97 0.551
R817 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t66 0.551
R818 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t58 0.551
R819 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t98 0.551
R820 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t47 0.551
R821 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t111 0.551
R822 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t40 0.551
R823 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t108 0.551
R824 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t22 0.551
R825 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t81 0.551
R826 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t76 0.551
R827 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t90 0.551
R828 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t3 0.551
R829 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t113 0.551
R830 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t75 0.551
R831 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t73 0.551
R832 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t93 0.551
R833 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t64 0.551
R834 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t15 0.551
R835 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t99 0.551
R836 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t43 0.551
R837 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t54 0.551
R838 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t107 0.551
R839 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t102 0.551
R840 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t48 0.551
R841 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t31 0.551
R842 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t21 0.551
R843 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t49 0.551
R844 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t6 0.551
R845 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t1 0.551
R846 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t65 0.551
R847 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t80 0.551
R848 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t32 0.551
R849 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t91 0.551
R850 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t117 0.551
R851 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t51 0.551
R852 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t20 0.551
R853 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t38 0.551
R854 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t100 0.551
R855 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t86 0.551
R856 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t5 0.551
R857 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t0 0.551
R858 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n40 0.46
R859 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n39 0.46
R860 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n70 0.46
R861 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n69 0.46
R862 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 0.403
R863 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n72 cascode_1_0/SD4L 0.166
R864 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n72 0.091
R865 cascode_1_0/SD4L cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t120 0.068
R866 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n41 0.063
R867 cascode_1_0/SD4L cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n71 0.063
R868 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n5 0.041
R869 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n3 0.041
R870 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n7 0.028
R871 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD2 0.028
R872 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n4 0.028
R873 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n2 0.028
R874 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n1 0.028
R875 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n0 0.028
R876 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 0.027
R877 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 0.027
R878 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 0.017
R879 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n6 0.017
R880 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 3.41
R881 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 3.41
R882 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n212 2.204
R883 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n210 2.204
R884 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n26 2.204
R885 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n24 2.204
R886 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n78 2.204
R887 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n76 2.204
R888 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n131 2.204
R889 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n129 2.204
R890 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t116 1.972
R891 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t181 1.972
R892 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t68 1.972
R893 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t121 1.972
R894 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_6/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t189 1.965
R895 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_4/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t233 1.965
R896 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t69 1.962
R897 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t104 1.961
R898 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n198 1.435
R899 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n12 1.435
R900 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n64 1.435
R901 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n117 1.435
R902 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n188 1.428
R903 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n189 1.428
R904 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n190 1.428
R905 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n191 1.428
R906 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n192 1.428
R907 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n193 1.428
R908 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n194 1.428
R909 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n195 1.428
R910 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n196 1.428
R911 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n197 1.428
R912 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n2 1.428
R913 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n3 1.428
R914 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n4 1.428
R915 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n5 1.428
R916 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n6 1.428
R917 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n7 1.428
R918 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n8 1.428
R919 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n9 1.428
R920 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n10 1.428
R921 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n11 1.428
R922 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n54 1.428
R923 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n55 1.428
R924 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n56 1.428
R925 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n57 1.428
R926 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n58 1.428
R927 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n59 1.428
R928 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n60 1.428
R929 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n61 1.428
R930 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n62 1.428
R931 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n63 1.428
R932 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n107 1.428
R933 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n108 1.428
R934 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n109 1.428
R935 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n110 1.428
R936 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n111 1.428
R937 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n112 1.428
R938 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n113 1.428
R939 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n114 1.428
R940 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n115 1.428
R941 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n116 1.428
R942 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n163 1.414
R943 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n164 1.414
R944 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n165 1.414
R945 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n166 1.414
R946 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n167 1.414
R947 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n168 1.414
R948 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n169 1.414
R949 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n170 1.414
R950 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n171 1.414
R951 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n172 1.414
R952 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n37 1.414
R953 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n38 1.414
R954 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n39 1.414
R955 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n40 1.414
R956 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n41 1.414
R957 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n31 1.414
R958 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n30 1.414
R959 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n29 1.414
R960 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n28 1.414
R961 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n27 1.414
R962 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n81 1.414
R963 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n82 1.414
R964 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n83 1.414
R965 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n84 1.414
R966 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n85 1.414
R967 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n86 1.414
R968 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n87 1.414
R969 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n88 1.414
R970 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n89 1.414
R971 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n90 1.414
R972 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n91 1.414
R973 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n142 1.414
R974 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n143 1.414
R975 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n144 1.414
R976 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n145 1.414
R977 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n146 1.414
R978 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n136 1.414
R979 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n135 1.414
R980 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n134 1.414
R981 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n133 1.414
R982 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n132 1.414
R983 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n181 1.413
R984 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n50 1.412
R985 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n49 1.412
R986 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n48 1.412
R987 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n47 1.412
R988 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n155 1.412
R989 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n154 1.412
R990 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n153 1.412
R991 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n152 1.412
R992 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n161 1.411
R993 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n162 1.411
R994 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n185 1.411
R995 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n80 1.411
R996 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n104 1.411
R997 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n103 1.411
R998 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n210 1.302
R999 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n212 1.302
R1000 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n24 1.302
R1001 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n26 1.302
R1002 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n76 1.302
R1003 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n78 1.302
R1004 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n129 1.302
R1005 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n131 1.302
R1006 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n186 1.278
R1007 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n187 1.278
R1008 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n0 1.278
R1009 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n1 1.278
R1010 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n52 1.278
R1011 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n53 1.278
R1012 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n105 1.278
R1013 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n106 1.278
R1014 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t115 0.551
R1015 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t1 0.551
R1016 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t5 0.551
R1017 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t67 0.551
R1018 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t23 0.551
R1019 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t66 0.551
R1020 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t70 0.551
R1021 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t106 0.551
R1022 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t20 0.551
R1023 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t26 0.551
R1024 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t55 0.551
R1025 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t95 0.551
R1026 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t98 0.551
R1027 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t9 0.551
R1028 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t44 0.551
R1029 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t91 0.551
R1030 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t81 0.551
R1031 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t6 0.551
R1032 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t31 0.551
R1033 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t76 0.551
R1034 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t46 0.551
R1035 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t53 0.551
R1036 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t48 0.551
R1037 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t99 0.551
R1038 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t10 0.551
R1039 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t15 0.551
R1040 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t194 0.551
R1041 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t123 0.551
R1042 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t128 0.551
R1043 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t133 0.551
R1044 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t191 0.551
R1045 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t200 0.551
R1046 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t238 0.551
R1047 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t150 0.551
R1048 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t154 0.551
R1049 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t197 0.551
R1050 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t222 0.551
R1051 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t148 0.551
R1052 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t138 0.551
R1053 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t183 0.551
R1054 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t218 0.551
R1055 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t229 0.551
R1056 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t135 0.551
R1057 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t170 0.551
R1058 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t203 0.551
R1059 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t207 0.551
R1060 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t122 0.551
R1061 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t159 0.551
R1062 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t228 0.551
R1063 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t235 0.551
R1064 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t130 0.551
R1065 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t174 0.551
R1066 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t144 0.551
R1067 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t177 0.551
R1068 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t180 0.551
R1069 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t140 0.551
R1070 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t103 0.551
R1071 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t30 0.551
R1072 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t19 0.551
R1073 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t25 0.551
R1074 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t88 0.551
R1075 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t94 0.551
R1076 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t113 0.551
R1077 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t32 0.551
R1078 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t21 0.551
R1079 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t64 0.551
R1080 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t89 0.551
R1081 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t12 0.551
R1082 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t18 0.551
R1083 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t52 0.551
R1084 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t87 0.551
R1085 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t93 0.551
R1086 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t3 0.551
R1087 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t40 0.551
R1088 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t85 0.551
R1089 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t78 0.551
R1090 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t110 0.551
R1091 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t39 0.551
R1092 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t114 0.551
R1093 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t0 0.551
R1094 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t22 0.551
R1095 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t65 0.551
R1096 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t36 0.551
R1097 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t82 0.551
R1098 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t72 0.551
R1099 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t33 0.551
R1100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t124 0.551
R1101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t162 0.551
R1102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t165 0.551
R1103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t210 0.551
R1104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t236 0.551
R1105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t161 0.551
R1106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t151 0.551
R1107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t192 0.551
R1108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t234 0.551
R1109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t157 0.551
R1110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t156 0.551
R1111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t186 0.551
R1112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t224 0.551
R1113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t232 0.551
R1114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t141 0.551
R1115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t145 0.551
R1116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t221 0.551
R1117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t212 0.551
R1118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t215 0.551
R1119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t172 0.551
R1120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t204 0.551
R1121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t213 0.551
R1122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t142 0.551
R1123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t185 0.551
R1124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t225 0.551
R1125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t160 0.551
R1126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t164 0.551
R1127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t209 0.551
R1128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t166 0.551
R1129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t211 0.551
R1130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t201 0.551
R1131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t205 0.551
R1132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t163 0.551
R1133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t167 0.551
R1134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t198 0.551
R1135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t239 0.551
R1136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t231 0.551
R1137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t155 0.551
R1138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t187 0.551
R1139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t223 0.551
R1140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t230 0.551
R1141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t152 0.551
R1142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t171 0.551
R1143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t178 0.551
R1144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t226 0.551
R1145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t126 0.551
R1146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t168 0.551
R1147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t175 0.551
R1148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t195 0.551
R1149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t125 0.551
R1150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t188 0.551
R1151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t196 0.551
R1152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t216 0.551
R1153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t143 0.551
R1154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t219 0.551
R1155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t146 0.551
R1156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t136 0.551
R1157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t214 0.551
R1158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t83 0.551
R1159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t90 0.551
R1160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t79 0.551
R1161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t37 0.551
R1162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t42 0.551
R1163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t74 0.551
R1164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t108 0.551
R1165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t35 0.551
R1166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t27 0.551
R1167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t71 0.551
R1168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t96 0.551
R1169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t101 0.551
R1170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t24 0.551
R1171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t58 0.551
R1172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t49 0.551
R1173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t100 0.551
R1174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t118 0.551
R1175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t45 0.551
R1176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t47 0.551
R1177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t97 0.551
R1178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t117 0.551
R1179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t43 0.551
R1180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t16 0.551
R1181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t61 0.551
R1182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t13 0.551
R1183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t7 0.551
R1184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t86 0.551
R1185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t92 0.551
R1186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t4 0.551
R1187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t50 0.551
R1188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t54 0.551
R1189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t59 0.551
R1190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t2 0.551
R1191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t8 0.551
R1192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t41 0.551
R1193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t77 0.551
R1194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t80 0.551
R1195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t112 0.551
R1196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t29 0.551
R1197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t75 0.551
R1198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t62 0.551
R1199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t111 0.551
R1200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t28 0.551
R1201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t17 0.551
R1202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t60 0.551
R1203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t102 0.551
R1204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t11 0.551
R1205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t14 0.551
R1206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t51 0.551
R1207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t84 0.551
R1208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t34 0.551
R1209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t38 0.551
R1210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t56 0.551
R1211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t105 0.551
R1212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t57 0.551
R1213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t107 0.551
R1214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t109 0.551
R1215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t63 0.551
R1216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t182 0.551
R1217 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t220 0.551
R1218 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t208 0.551
R1219 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t137 0.551
R1220 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t169 0.551
R1221 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t217 0.551
R1222 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t206 0.551
R1223 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t134 0.551
R1224 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t158 0.551
R1225 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t202 0.551
R1226 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t176 0.551
R1227 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t227 0.551
R1228 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t139 0.551
R1229 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t131 0.551
R1230 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t173 0.551
R1231 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t179 0.551
R1232 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t120 0.551
R1233 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t129 0.551
R1234 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t132 0.551
R1235 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t193 0.551
R1236 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t147 0.551
R1237 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t153 0.551
R1238 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t184 0.551
R1239 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t237 0.551
R1240 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t149 0.551
R1241 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t190 0.551
R1242 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t199 0.551
R1243 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t127 0.551
R1244 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t73 0.551
R1245 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t119 0.551
R1246 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n211 0.46
R1247 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n209 0.46
R1248 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n25 0.46
R1249 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n23 0.46
R1250 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n77 0.46
R1251 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n75 0.46
R1252 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n130 0.46
R1253 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n128 0.46
R1254 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n156 0.455
R1255 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n51 0.416
R1256 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD2 0.281
R1257 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD2 0.281
R1258 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 0.155
R1259 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 0.155
R1260 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n157 0.13
R1261 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n160 0.13
R1262 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n158 0.091
R1263 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n79 0.076
R1264 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n214 N2 0.073
R1265 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n213 0.041
R1266 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n159 0.039
R1267 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n214 0.034
R1268 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 0.027
R1269 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 0.027
R1270 cascode_1_0/SD3L cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n215 0.015
R1271 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n199 0.007
R1272 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n200 0.007
R1273 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n201 0.007
R1274 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n202 0.007
R1275 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n203 0.007
R1276 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n204 0.007
R1277 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n205 0.007
R1278 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n206 0.007
R1279 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n207 0.007
R1280 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n13 0.007
R1281 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n14 0.007
R1282 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n15 0.007
R1283 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n16 0.007
R1284 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n17 0.007
R1285 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n18 0.007
R1286 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n19 0.007
R1287 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n20 0.007
R1288 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n21 0.007
R1289 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n42 0.007
R1290 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n43 0.007
R1291 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n44 0.007
R1292 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n45 0.007
R1293 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n35 0.007
R1294 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n34 0.007
R1295 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n33 0.007
R1296 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n32 0.007
R1297 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_6/SD2 0.007
R1298 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n65 0.007
R1299 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n66 0.007
R1300 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n67 0.007
R1301 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n68 0.007
R1302 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n69 0.007
R1303 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n70 0.007
R1304 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n71 0.007
R1305 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n72 0.007
R1306 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n73 0.007
R1307 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n92 0.007
R1308 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n93 0.007
R1309 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n94 0.007
R1310 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n95 0.007
R1311 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n96 0.007
R1312 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n97 0.007
R1313 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n98 0.007
R1314 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n99 0.007
R1315 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n100 0.007
R1316 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n101 0.007
R1317 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n118 0.007
R1318 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n119 0.007
R1319 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n120 0.007
R1320 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n121 0.007
R1321 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n122 0.007
R1322 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n123 0.007
R1323 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n124 0.007
R1324 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n125 0.007
R1325 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n126 0.007
R1326 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n147 0.007
R1327 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n148 0.007
R1328 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n149 0.007
R1329 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n150 0.007
R1330 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n140 0.007
R1331 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n139 0.007
R1332 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n138 0.007
R1333 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n137 0.007
R1334 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_4/SD2 0.007
R1335 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n173 0.007
R1336 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n174 0.007
R1337 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n175 0.007
R1338 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n176 0.007
R1339 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n177 0.007
R1340 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n178 0.007
R1341 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n179 0.007
R1342 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n180 0.007
R1343 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n182 0.007
R1344 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n183 0.007
R1345 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n208 0.006
R1346 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n22 0.006
R1347 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n36 0.006
R1348 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n74 0.006
R1349 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n127 0.006
R1350 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n141 0.006
R1351 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n46 0.004
R1352 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n102 0.004
R1353 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n151 0.004
R1354 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n184 0.004
R1355 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n177 2.204
R1356 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n207 2.204
R1357 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t231 1.965
R1358 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_3/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t69 1.965
R1359 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t146 1.965
R1360 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t25 1.965
R1361 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t229 1.963
R1362 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t77 1.963
R1363 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t156 1.963
R1364 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t17 1.96
R1365 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n88 1.435
R1366 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n163 1.435
R1367 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n193 1.435
R1368 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n14 1.434
R1369 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n10 1.428
R1370 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n11 1.428
R1371 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n12 1.428
R1372 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n13 1.428
R1373 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n0 1.428
R1374 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n1 1.428
R1375 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n2 1.428
R1376 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n3 1.428
R1377 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n4 1.428
R1378 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n5 1.428
R1379 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n84 1.428
R1380 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n85 1.428
R1381 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n86 1.428
R1382 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n87 1.428
R1383 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n77 1.428
R1384 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n76 1.428
R1385 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n75 1.428
R1386 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n74 1.428
R1387 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n73 1.428
R1388 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n72 1.428
R1389 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n153 1.428
R1390 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n154 1.428
R1391 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n155 1.428
R1392 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n156 1.428
R1393 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n157 1.428
R1394 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n158 1.428
R1395 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n159 1.428
R1396 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n160 1.428
R1397 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n161 1.428
R1398 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n162 1.428
R1399 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n183 1.428
R1400 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n184 1.428
R1401 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n185 1.428
R1402 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n186 1.428
R1403 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n187 1.428
R1404 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n188 1.428
R1405 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n189 1.428
R1406 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n190 1.428
R1407 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n191 1.428
R1408 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n192 1.428
R1409 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n55 1.414
R1410 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n54 1.414
R1411 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n53 1.414
R1412 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n52 1.414
R1413 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n51 1.414
R1414 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n50 1.414
R1415 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n49 1.414
R1416 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n48 1.414
R1417 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n47 1.414
R1418 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n46 1.414
R1419 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n45 1.414
R1420 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n98 1.414
R1421 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n99 1.414
R1422 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n100 1.414
R1423 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n101 1.414
R1424 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n102 1.414
R1425 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n103 1.414
R1426 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n104 1.414
R1427 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n105 1.414
R1428 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n106 1.414
R1429 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n107 1.414
R1430 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n108 1.414
R1431 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n124 1.414
R1432 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n125 1.414
R1433 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n126 1.414
R1434 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n127 1.414
R1435 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n128 1.414
R1436 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n129 1.414
R1437 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n130 1.414
R1438 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n131 1.414
R1439 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n132 1.414
R1440 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n133 1.414
R1441 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n134 1.414
R1442 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n19 1.414
R1443 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n20 1.414
R1444 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n21 1.414
R1445 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n22 1.414
R1446 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n23 1.414
R1447 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n24 1.414
R1448 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n25 1.414
R1449 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n26 1.414
R1450 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n27 1.414
R1451 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n28 1.414
R1452 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n29 1.414
R1453 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n122 1.412
R1454 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n121 1.412
R1455 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n120 1.412
R1456 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n148 1.412
R1457 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n147 1.412
R1458 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n146 1.412
R1459 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n43 1.412
R1460 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n42 1.412
R1461 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n41 1.412
R1462 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n67 1.41
R1463 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n69 1.409
R1464 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n70 1.409
R1465 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n177 1.302
R1466 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n207 1.302
R1467 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n174 1.282
R1468 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n204 1.282
R1469 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n93 1.28
R1470 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n94 1.28
R1471 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n95 1.28
R1472 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n96 1.28
R1473 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n9 1.28
R1474 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n8 1.28
R1475 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n7 1.28
R1476 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n6 1.28
R1477 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n151 1.278
R1478 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n152 1.278
R1479 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n181 1.278
R1480 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n182 1.278
R1481 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t98 0.551
R1482 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t23 0.551
R1483 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t59 0.551
R1484 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t67 0.551
R1485 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t96 0.551
R1486 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t9 0.551
R1487 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t41 0.551
R1488 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t49 0.551
R1489 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t66 0.551
R1490 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t74 0.551
R1491 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t104 0.551
R1492 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t15 0.551
R1493 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t21 0.551
R1494 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t99 0.551
R1495 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t89 0.551
R1496 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t12 0.551
R1497 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t32 0.551
R1498 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t81 0.551
R1499 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t87 0.551
R1500 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t92 0.551
R1501 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t62 0.551
R1502 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t107 0.551
R1503 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t114 0.551
R1504 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t36 0.551
R1505 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t75 0.551
R1506 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t109 0.551
R1507 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t30 0.551
R1508 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t38 0.551
R1509 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t110 0.551
R1510 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t22 0.551
R1511 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t58 0.551
R1512 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t64 0.551
R1513 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t95 0.551
R1514 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t100 0.551
R1515 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t55 0.551
R1516 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t48 0.551
R1517 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t51 0.551
R1518 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t6 0.551
R1519 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t1 0.551
R1520 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t45 0.551
R1521 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t57 0.551
R1522 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t117 0.551
R1523 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t94 0.551
R1524 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t20 0.551
R1525 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t40 0.551
R1526 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t47 0.551
R1527 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t79 0.551
R1528 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t118 0.551
R1529 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t0 0.551
R1530 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t44 0.551
R1531 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t72 0.551
R1532 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t116 0.551
R1533 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t105 0.551
R1534 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t27 0.551
R1535 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t70 0.551
R1536 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t113 0.551
R1537 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t68 0.551
R1538 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t111 0.551
R1539 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t10 0.551
R1540 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t16 0.551
R1541 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t65 0.551
R1542 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t85 0.551
R1543 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t7 0.551
R1544 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t13 0.551
R1545 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t33 0.551
R1546 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t83 0.551
R1547 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t28 0.551
R1548 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t34 0.551
R1549 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t60 0.551
R1550 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t106 0.551
R1551 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t97 0.551
R1552 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t52 0.551
R1553 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t56 0.551
R1554 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t102 0.551
R1555 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t3 0.551
R1556 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t50 0.551
R1557 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t39 0.551
R1558 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t46 0.551
R1559 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t24 0.551
R1560 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t63 0.551
R1561 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t71 0.551
R1562 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t115 0.551
R1563 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t37 0.551
R1564 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t76 0.551
R1565 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t2 0.551
R1566 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t5 0.551
R1567 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t212 0.551
R1568 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t142 0.551
R1569 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t188 0.551
R1570 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t220 0.551
R1571 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t136 0.551
R1572 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t143 0.551
R1573 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t192 0.551
R1574 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t234 0.551
R1575 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t151 0.551
R1576 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t198 0.551
R1577 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t202 0.551
R1578 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t237 0.551
R1579 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t122 0.551
R1580 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t201 0.551
R1581 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t127 0.551
R1582 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t132 0.551
R1583 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t177 0.551
R1584 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t169 0.551
R1585 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t129 0.551
R1586 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t134 0.551
R1587 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t181 0.551
R1588 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t225 0.551
R1589 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t157 0.551
R1590 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t203 0.551
R1591 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t210 0.551
R1592 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t138 0.551
R1593 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t159 0.551
R1594 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t205 0.551
R1595 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t163 0.551
R1596 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t206 0.551
R1597 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t213 0.551
R1598 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t218 0.551
R1599 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t160 0.551
R1600 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t165 0.551
R1601 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t200 0.551
R1602 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t233 0.551
R1603 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t239 0.551
R1604 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t152 0.551
R1605 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t186 0.551
R1606 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t230 0.551
R1607 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t221 0.551
R1608 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t150 0.551
R1609 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t185 0.551
R1610 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t174 0.551
R1611 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t219 0.551
R1612 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t137 0.551
R1613 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t167 0.551
R1614 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t173 0.551
R1615 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t207 0.551
R1616 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t121 0.551
R1617 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t214 0.551
R1618 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t144 0.551
R1619 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t193 0.551
R1620 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t196 0.551
R1621 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t148 0.551
R1622 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t222 0.551
R1623 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t216 0.551
R1624 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t145 0.551
R1625 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t43 0.551
R1626 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t91 0.551
R1627 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t18 0.551
R1628 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t54 0.551
R1629 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t101 0.551
R1630 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t108 0.551
R1631 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t19 0.551
R1632 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t73 0.551
R1633 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t103 0.551
R1634 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t26 0.551
R1635 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t31 0.551
R1636 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t80 0.551
R1637 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t88 0.551
R1638 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t29 0.551
R1639 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t78 0.551
R1640 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t84 0.551
R1641 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t8 0.551
R1642 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t14 0.551
R1643 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t93 0.551
R1644 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t86 0.551
R1645 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t11 0.551
R1646 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t61 0.551
R1647 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t112 0.551
R1648 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t35 0.551
R1649 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t42 0.551
R1650 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t90 0.551
R1651 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t4 0.551
R1652 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t53 0.551
R1653 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t140 0.551
R1654 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t170 0.551
R1655 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t217 0.551
R1656 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t135 0.551
R1657 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t182 0.551
R1658 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t189 0.551
R1659 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t232 0.551
R1660 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t147 0.551
R1661 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t184 0.551
R1662 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t226 0.551
R1663 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t236 0.551
R1664 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t162 0.551
R1665 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t166 0.551
R1666 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t228 0.551
R1667 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t155 0.551
R1668 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t164 0.551
R1669 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t209 0.551
R1670 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t215 0.551
R1671 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t172 0.551
R1672 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t180 0.551
R1673 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t211 0.551
R1674 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t139 0.551
R1675 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t194 0.551
R1676 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t238 0.551
R1677 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t124 0.551
R1678 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t168 0.551
R1679 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t204 0.551
R1680 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t133 0.551
R1681 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t141 0.551
R1682 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t187 0.551
R1683 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t176 0.551
R1684 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t183 0.551
R1685 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t126 0.551
R1686 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t131 0.551
R1687 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t153 0.551
R1688 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t190 0.551
R1689 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t178 0.551
R1690 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t223 0.551
R1691 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t128 0.551
R1692 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t171 0.551
R1693 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t175 0.551
R1694 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t208 0.551
R1695 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t125 0.551
R1696 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t130 0.551
R1697 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t161 0.551
R1698 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t199 0.551
R1699 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t123 0.551
R1700 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t235 0.551
R1701 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t149 0.551
R1702 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t197 0.551
R1703 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t179 0.551
R1704 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t224 0.551
R1705 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t154 0.551
R1706 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t158 0.551
R1707 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t227 0.551
R1708 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t191 0.551
R1709 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t195 0.551
R1710 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t120 0.551
R1711 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t82 0.551
R1712 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t119 0.551
R1713 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n176 0.46
R1714 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n206 0.46
R1715 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n71 0.35
R1716 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n123 0.347
R1717 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n44 0.347
R1718 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n149 0.315
R1719 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n97 0.224
R1720 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n209 0.224
R1721 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n150 0.113
R1722 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n179 0.091
R1723 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n180 0.079
R1724 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n209 cascode_1_0/SD3R 0.054
R1725 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1 0.05
R1726 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 0.05
R1727 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n150 P2 0.049
R1728 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n178 0.039
R1729 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n208 0.039
R1730 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n66 0.007
R1731 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n65 0.007
R1732 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n64 0.007
R1733 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n63 0.007
R1734 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n62 0.007
R1735 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n61 0.007
R1736 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n60 0.007
R1737 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n59 0.007
R1738 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n58 0.007
R1739 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n57 0.007
R1740 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n56 0.007
R1741 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/SD2 0.007
R1742 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n89 0.007
R1743 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n90 0.007
R1744 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n91 0.007
R1745 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n82 0.007
R1746 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n81 0.007
R1747 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n80 0.007
R1748 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n79 0.007
R1749 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n78 0.007
R1750 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n118 0.007
R1751 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n117 0.007
R1752 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n116 0.007
R1753 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n115 0.007
R1754 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n114 0.007
R1755 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n113 0.007
R1756 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n112 0.007
R1757 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n111 0.007
R1758 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n110 0.007
R1759 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n109 0.007
R1760 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/SD2 0.007
R1761 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n164 0.007
R1762 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n165 0.007
R1763 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n166 0.007
R1764 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n167 0.007
R1765 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n168 0.007
R1766 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n169 0.007
R1767 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n170 0.007
R1768 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n171 0.007
R1769 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n172 0.007
R1770 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n173 0.007
R1771 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n144 0.007
R1772 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n143 0.007
R1773 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n142 0.007
R1774 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n141 0.007
R1775 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n140 0.007
R1776 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n139 0.007
R1777 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n138 0.007
R1778 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n137 0.007
R1779 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n136 0.007
R1780 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n135 0.007
R1781 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_3/SD2 0.007
R1782 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n39 0.007
R1783 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n38 0.007
R1784 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n37 0.007
R1785 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n36 0.007
R1786 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n35 0.007
R1787 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n34 0.007
R1788 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n33 0.007
R1789 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n32 0.007
R1790 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n31 0.007
R1791 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n30 0.007
R1792 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD2 0.007
R1793 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n194 0.007
R1794 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n195 0.007
R1795 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n196 0.007
R1796 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n197 0.007
R1797 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n198 0.007
R1798 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n199 0.007
R1799 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n200 0.007
R1800 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n201 0.007
R1801 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n202 0.007
R1802 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n203 0.007
R1803 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n15 0.007
R1804 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n16 0.007
R1805 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n17 0.007
R1806 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n211 0.007
R1807 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n212 0.007
R1808 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n213 0.007
R1809 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n214 0.007
R1810 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n215 0.007
R1811 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n119 0.006
R1812 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n145 0.006
R1813 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n40 0.006
R1814 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n92 0.005
R1815 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n18 0.005
R1816 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n83 0.004
R1817 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n210 0.004
R1818 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_5/SD1 0.003
R1819 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n216 0.003
R1820 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n175 0.003
R1821 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n205 0.003
R1822 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n68 0.001
R1823 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t2 9.759
R1824 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n52 2.204
R1825 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n50 2.204
R1826 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n104 2.204
R1827 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n102 2.204
R1828 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t87 1.972
R1829 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t117 1.972
R1830 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t26 1.962
R1831 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t102 1.962
R1832 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n38 1.435
R1833 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n90 1.435
R1834 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n28 1.428
R1835 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n29 1.428
R1836 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n30 1.428
R1837 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n31 1.428
R1838 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n32 1.428
R1839 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n33 1.428
R1840 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n34 1.428
R1841 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n35 1.428
R1842 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n36 1.428
R1843 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n37 1.428
R1844 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n80 1.428
R1845 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n81 1.428
R1846 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n82 1.428
R1847 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n83 1.428
R1848 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n84 1.428
R1849 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n85 1.428
R1850 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n86 1.428
R1851 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n87 1.428
R1852 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n88 1.428
R1853 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n89 1.428
R1854 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n54 1.414
R1855 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n55 1.414
R1856 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n56 1.414
R1857 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n57 1.414
R1858 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n58 1.414
R1859 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n59 1.414
R1860 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n60 1.414
R1861 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n61 1.414
R1862 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n62 1.414
R1863 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n63 1.414
R1864 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n64 1.414
R1865 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n1 1.414
R1866 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n2 1.414
R1867 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n3 1.414
R1868 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n4 1.414
R1869 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n5 1.414
R1870 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n6 1.414
R1871 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n7 1.414
R1872 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n8 1.414
R1873 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n9 1.414
R1874 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n10 1.414
R1875 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n11 1.414
R1876 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n53 1.411
R1877 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n77 1.411
R1878 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n76 1.411
R1879 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n0 1.411
R1880 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n108 1.411
R1881 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n23 1.411
R1882 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n50 1.302
R1883 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n52 1.302
R1884 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n102 1.302
R1885 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n104 1.302
R1886 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n26 1.278
R1887 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n27 1.278
R1888 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n78 1.278
R1889 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n79 1.278
R1890 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t50 0.551
R1891 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t78 0.551
R1892 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t122 0.551
R1893 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t58 0.551
R1894 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t35 0.551
R1895 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t96 0.551
R1896 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t89 0.551
R1897 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t114 0.551
R1898 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t29 0.551
R1899 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t60 0.551
R1900 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t67 0.551
R1901 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t98 0.551
R1902 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t99 0.551
R1903 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t40 0.551
R1904 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t10 0.551
R1905 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t69 0.551
R1906 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t81 0.551
R1907 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t109 0.551
R1908 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t76 0.551
R1909 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t52 0.551
R1910 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t22 0.551
R1911 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t48 0.551
R1912 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t46 0.551
R1913 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t107 0.551
R1914 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t59 0.551
R1915 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t86 0.551
R1916 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t73 0.551
R1917 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t101 0.551
R1918 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t20 0.551
R1919 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t12 0.551
R1920 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t43 0.551
R1921 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t105 0.551
R1922 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t21 0.551
R1923 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t16 0.551
R1924 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t17 0.551
R1925 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t88 0.551
R1926 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t55 0.551
R1927 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t82 0.551
R1928 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t123 0.551
R1929 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t28 0.551
R1930 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t37 0.551
R1931 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t97 0.551
R1932 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t66 0.551
R1933 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t94 0.551
R1934 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t8 0.551
R1935 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t38 0.551
R1936 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t47 0.551
R1937 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t74 0.551
R1938 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t75 0.551
R1939 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t106 0.551
R1940 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t115 0.551
R1941 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t18 0.551
R1942 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t65 0.551
R1943 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t93 0.551
R1944 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t6 0.551
R1945 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t108 0.551
R1946 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t104 0.551
R1947 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t36 0.551
R1948 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t33 0.551
R1949 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t61 0.551
R1950 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t63 0.551
R1951 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t120 0.551
R1952 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t100 0.551
R1953 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t32 0.551
R1954 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t45 0.551
R1955 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t71 0.551
R1956 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t72 0.551
R1957 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t19 0.551
R1958 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t111 0.551
R1959 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t11 0.551
R1960 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t57 0.551
R1961 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t85 0.551
R1962 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t49 0.551
R1963 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t27 0.551
R1964 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t121 0.551
R1965 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t23 0.551
R1966 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t34 0.551
R1967 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t95 0.551
R1968 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t62 0.551
R1969 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t7 0.551
R1970 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t112 0.551
R1971 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t44 0.551
R1972 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t119 0.551
R1973 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t24 0.551
R1974 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t56 0.551
R1975 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t83 0.551
R1976 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t84 0.551
R1977 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t77 0.551
R1978 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t116 0.551
R1979 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t51 0.551
R1980 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t53 0.551
R1981 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t90 0.551
R1982 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t91 0.551
R1983 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t118 0.551
R1984 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t4 0.551
R1985 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t30 0.551
R1986 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t31 0.551
R1987 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t103 0.551
R1988 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t70 0.551
R1989 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t5 0.551
R1990 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t15 0.551
R1991 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t39 0.551
R1992 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t42 0.551
R1993 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t113 0.551
R1994 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t80 0.551
R1995 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t110 0.551
R1996 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t25 0.551
R1997 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t54 0.551
R1998 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t64 0.551
R1999 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t92 0.551
R2000 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t13 0.551
R2001 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t41 0.551
R2002 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t79 0.551
R2003 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t14 0.551
R2004 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t9 0.551
R2005 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t68 0.551
R2006 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n51 0.46
R2007 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n49 0.46
R2008 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n103 0.46
R2009 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n101 0.46
R2010 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 0.254
R2011 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD2 0.249
R2012 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n107 0.243
R2013 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t1 0.231
R2014 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n24 0.137
R2015 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n105 0.13
R2016 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 0.124
R2017 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n106 0.114
R2018 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t3 0.061
R2019 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n25 cascode_1_0/SD1L 0.039
R2020 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t0 0.031
R2021 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n39 0.007
R2022 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n40 0.007
R2023 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n41 0.007
R2024 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n42 0.007
R2025 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n43 0.007
R2026 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n44 0.007
R2027 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n45 0.007
R2028 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n46 0.007
R2029 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n47 0.007
R2030 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n65 0.007
R2031 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n66 0.007
R2032 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n67 0.007
R2033 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n68 0.007
R2034 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n69 0.007
R2035 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n70 0.007
R2036 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n71 0.007
R2037 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n72 0.007
R2038 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n73 0.007
R2039 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n74 0.007
R2040 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n91 0.007
R2041 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n92 0.007
R2042 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n93 0.007
R2043 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n94 0.007
R2044 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n95 0.007
R2045 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n96 0.007
R2046 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n97 0.007
R2047 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n98 0.007
R2048 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n99 0.007
R2049 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n12 0.007
R2050 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n13 0.007
R2051 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n14 0.007
R2052 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n15 0.007
R2053 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n16 0.007
R2054 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n17 0.007
R2055 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n18 0.007
R2056 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n19 0.007
R2057 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n20 0.007
R2058 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n21 0.007
R2059 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n25 0.006
R2060 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n48 0.006
R2061 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n100 0.006
R2062 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n75 0.004
R2063 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n22 0.004
C42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 139.46fF
C43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 106.66fF $ **FLOATING
C44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 107.53fF $ **FLOATING
C45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 154.39fF
C46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 170.60fF
C47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 226.65fF $ **FLOATING
C48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 240.38fF $ **FLOATING
C49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 178.26fF $ **FLOATING
C50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 112.16fF $ **FLOATING
C51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 139.45fF $ **FLOATING
C52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 114.40fF $ **FLOATING
C53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 104.54fF $ **FLOATING
C54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.06fF
C55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.78fF $ **FLOATING
C67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 8.35fF
C68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.12fF
C78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.06fF
C79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 74.34fF $ **FLOATING
C80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 157.91fF $ **FLOATING
C81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 110.09fF
C82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 203.45fF $ **FLOATING
C83 cascode_1_0/SD1L cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 14.76fF
C84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 82.29fF
C85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.05fF
C86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.05fF
C87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.09fF
C98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 8.57fF
C99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.61fF
C108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.96fF
C109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.96fF
C110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 32.97fF
C111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.06fF
C112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.78fF $ **FLOATING
C124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 8.35fF
C125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.12fF
C135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.06fF
C136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.76fF $ **FLOATING
C137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.06fF
C138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 44.47fF
C139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.05fF
C140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.05fF
C141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.07fF
C151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.09fF
C152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 8.57fF
C153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.65fF
C161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.61fF
C162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.96fF
C163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.96fF
C164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 51.09fF
C165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 76.40fF
C166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 45.97fF
C167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 52.07fF
C168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.t102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.76fF $ **FLOATING
C169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.06fF
C170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.63fF
C186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.03fF
C189 cascode_1_0/SD3R cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 10.20fF
C190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.08fF $ **FLOATING
C202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 6.90fF
C203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.34fF
C214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.07fF $ **FLOATING
C215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C217 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C218 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 79.37fF
C219 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C220 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C221 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C222 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C223 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C224 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C225 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C226 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C227 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C228 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C229 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C230 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.08fF $ **FLOATING
C231 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 6.90fF
C232 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C233 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C234 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C235 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C236 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C237 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C238 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C239 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C240 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C241 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C242 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.56fF
C243 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C244 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.36fF
C245 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C246 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C247 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.07fF $ **FLOATING
C248 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 75.27fF
C249 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C250 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C251 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C252 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C253 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C254 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C255 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_5/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.84fF
C256 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.40fF
C257 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C258 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C259 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C260 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C261 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.60fF
C262 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C263 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C264 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C265 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C266 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C267 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.63fF
C268 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C269 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C270 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.03fF
C271 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C272 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C273 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C274 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C275 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 60.87fF
C276 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C277 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C278 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C279 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C280 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C281 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C282 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C283 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C284 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C285 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C286 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C287 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t231 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.08fF $ **FLOATING
C288 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 6.90fF
C289 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C290 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C291 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C292 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C293 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C294 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C295 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C296 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C297 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C298 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C299 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.34fF
C300 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t229 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.07fF $ **FLOATING
C301 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C302 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C303 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C304 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 79.37fF
C305 P2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 38.08fF
C306 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C307 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C308 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C309 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C310 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C311 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C312 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C313 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C314 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C315 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C316 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C317 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.08fF $ **FLOATING
C318 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_3/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 6.90fF
C319 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C320 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C321 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C322 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C323 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C324 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C325 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C326 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C327 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C328 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C329 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.34fF
C330 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.t77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.07fF $ **FLOATING
C331 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C332 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C333 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C334 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 75.30fF
C335 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 72.99fF
C336 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C337 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C338 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C339 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C340 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C341 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C342 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C343 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C344 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C345 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C346 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C347 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C348 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C349 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.63fF
C350 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C351 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C352 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C353 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C354 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C355 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C356 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C357 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C358 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.31fF
C359 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C360 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.72fF
C361 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.36fF
C362 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 75.65fF
C363 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 68.25fF
C364 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 59.62fF
C365 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 83.75fF
C366 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C367 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C368 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C369 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C370 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C371 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C372 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C373 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C374 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C375 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C376 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C377 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.52fF
C378 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C379 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.63fF
C380 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C381 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C382 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C383 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C384 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C385 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C386 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C387 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C388 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.31fF
C389 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.50fF
C390 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.72fF
C391 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.36fF
C392 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 68.25fF
C393 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 52.88fF
C394 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 60.87fF
C395 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.60fF
C396 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n212 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C397 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C398 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C399 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.39fF
C400 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1.n216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.40fF
C401 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.84fF
C402 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C403 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C404 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C405 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C406 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C407 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C408 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C409 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C410 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C411 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C412 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C413 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C414 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.63fF
C415 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.82fF
C416 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C417 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C418 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C419 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C420 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C421 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C422 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C423 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C424 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C425 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.43fF
C426 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.43fF
C427 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 53.54fF
C428 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C429 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C430 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C431 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C432 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C433 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.14fF $ **FLOATING
C434 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_6/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 7.01fF
C435 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C436 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C437 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C438 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C439 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C440 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C441 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C442 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C443 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C444 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C445 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.16fF $ **FLOATING
C446 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.50fF
C447 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C448 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C449 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C450 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.66fF
C451 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C452 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C453 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C454 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C455 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 86.89fF
C456 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C457 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C458 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C459 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C460 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C461 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C462 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C463 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C464 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C465 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C466 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C467 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C468 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.63fF
C469 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.82fF
C470 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C471 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C472 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C473 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C474 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C475 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C476 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C477 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C478 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C479 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.43fF
C480 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.43fF
C481 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 36.14fF
C482 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 13.82fF
C483 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C484 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C485 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C486 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C487 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C488 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C489 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C490 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C491 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C492 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C493 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C494 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C495 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.16fF $ **FLOATING
C496 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.50fF
C497 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C498 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C499 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C500 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C501 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C502 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C503 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C504 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C505 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C506 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.67fF
C507 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C508 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C509 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C510 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 70.75fF
C511 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C512 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C513 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C514 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C515 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C516 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C517 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C518 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C519 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C520 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C521 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C522 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C523 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.63fF
C524 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.82fF
C525 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C526 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C527 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C528 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C529 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C530 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C531 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C532 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C533 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C534 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.43fF
C535 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.43fF
C536 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 53.54fF
C537 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C538 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C539 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C540 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C541 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C542 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t233 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.14fF $ **FLOATING
C543 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_4/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 7.34fF
C544 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C545 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C546 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C547 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C548 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C549 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C550 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C551 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C552 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C553 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C554 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.17fF $ **FLOATING
C555 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 14.61fF
C556 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C557 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C558 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C559 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.66fF
C560 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C561 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C562 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C563 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C564 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 94.58fF
C565 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 140.66fF
C566 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 89.55fF
C567 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 86.10fF
C568 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 58.72fF
C569 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C570 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C571 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C572 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C573 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C574 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C575 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C576 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C577 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C578 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C579 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C580 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C581 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.16fF $ **FLOATING
C582 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.50fF
C583 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C584 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C585 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C586 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C587 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C588 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C589 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C590 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C591 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C592 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n183 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C593 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.67fF
C594 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.t104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C595 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C596 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 70.74fF
C597 N2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 37.76fF
C598 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C599 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C600 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C601 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C602 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C603 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C604 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C605 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C606 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C607 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C608 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C609 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C610 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.63fF
C611 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.82fF
C612 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C613 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C614 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C615 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C616 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C617 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C618 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C619 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.47fF
C620 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C621 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.43fF
C622 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.43fF
C623 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 9.21fF
C624 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n214 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 16.31fF
C625 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 69.72fF
C626 cascode_1_0/SD3L cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.93fF
C627 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 17.40fF
C628 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 20.38fF
C629 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 18.94fF
C630 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 17.44fF
C631 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 18.94fF
C632 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 17.44fF
C633 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 9.95fF
C634 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 17.40fF
C635 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 18.69fF
C636 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 41.84fF
C637 cascode_1_0/SD4L cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 59.52fF
C638 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 76.02fF
C639 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 98.95fF
C640 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 10.22fF
C641 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.30fF $ **FLOATING
C642 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C643 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C644 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C645 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C646 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C647 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C648 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C649 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C650 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C651 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C652 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C653 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.32fF $ **FLOATING
C654 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C655 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.64fF
C656 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.64fF
C657 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C658 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C659 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C660 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C661 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C662 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C663 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C664 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C665 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C666 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C667 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.69fF
C668 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.53fF
C669 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.53fF
C670 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 9.68fF
C671 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C672 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C673 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C674 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C675 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C676 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.30fF $ **FLOATING
C677 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C678 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C679 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C680 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C681 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C682 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.32fF $ **FLOATING
C683 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C684 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C685 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C686 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C687 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.64fF
C688 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.64fF
C689 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C690 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C691 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C692 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C693 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C694 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C695 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C696 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C697 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C698 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C699 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.69fF
C700 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.53fF
C701 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.53fF
C702 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 9.68fF
C703 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.t120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 186.51fF $ **FLOATING
C704 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 86.50fF
C705 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 105.67fF
C706 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C707 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.66fF
C708 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C709 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C710 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C711 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C712 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C713 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C714 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.88fF
C715 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.46fF
C716 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C717 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C718 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C719 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C720 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.66fF
C721 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C722 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C723 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C724 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C725 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.62fF
C726 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.80fF
C727 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C728 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C729 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.09fF
C730 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C731 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C732 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C733 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C734 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 61.69fF
C735 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C736 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C737 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C738 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C739 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C740 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C741 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C742 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C743 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C744 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C745 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C746 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C747 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 7.00fF
C748 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C749 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C750 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C751 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C752 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C753 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C754 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C755 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C756 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C757 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C758 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C759 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C760 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C761 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C762 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C763 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 80.44fF
C764 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C765 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C766 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C767 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C768 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C769 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C770 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C771 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C772 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C773 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C774 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C775 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C776 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 7.00fF
C777 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C778 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C779 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C780 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C781 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C782 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C783 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C784 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C785 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C786 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C787 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n73 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.63fF
C788 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n74 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C789 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n75 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.42fF
C790 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n76 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C791 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n77 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C792 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C793 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n78 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 76.28fF
C794 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n79 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C795 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n80 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C796 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n81 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C797 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n82 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C798 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n83 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C799 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n84 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C800 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.88fF
C801 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n85 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.46fF
C802 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n86 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C803 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n87 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C804 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n88 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C805 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C806 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n90 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.66fF
C807 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n91 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C808 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n92 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C809 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n93 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C810 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n94 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C811 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n95 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.62fF
C812 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n96 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.80fF
C813 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n97 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C814 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n98 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C815 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n99 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.09fF
C816 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n100 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C817 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n101 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C818 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n102 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C819 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n103 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C820 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n104 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 61.69fF
C821 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n105 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C822 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n106 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C823 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n107 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C824 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n108 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C825 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n109 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C826 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n110 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C827 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n111 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C828 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n112 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C829 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C830 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n114 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C831 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n115 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C832 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t113 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C833 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 7.00fF
C834 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n116 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C835 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n117 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C836 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n118 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C837 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n119 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C838 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C839 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C840 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n122 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C841 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C842 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n124 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C843 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n125 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C844 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n126 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C845 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C846 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n127 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C847 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n128 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C848 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n129 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C849 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n130 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 80.44fF
C850 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n131 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C851 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n132 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C852 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n133 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C853 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n134 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C854 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n135 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C855 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n136 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C856 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n137 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C857 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n138 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C858 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n139 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C859 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n140 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C860 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n141 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C861 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C862 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 7.00fF
C863 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n142 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C864 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n143 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C865 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n144 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C866 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n145 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C867 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n146 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C868 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n147 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C869 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n148 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C870 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n149 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C871 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n150 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C872 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n151 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C873 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n152 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.41fF
C874 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.t215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.13fF $ **FLOATING
C875 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n153 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C876 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n154 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C877 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n155 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.58fF
C878 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n156 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 94.52fF
C879 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n157 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C880 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n158 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C881 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n159 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C882 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n160 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C883 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n161 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C884 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n162 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C885 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n163 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C886 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n164 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C887 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n165 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C888 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n166 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C889 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n167 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C890 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n168 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C891 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n169 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.62fF
C892 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n170 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.80fF
C893 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n171 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C894 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n172 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C895 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n173 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C896 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n174 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C897 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n175 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C898 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n176 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C899 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n177 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C900 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n178 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C901 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n179 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.38fF
C902 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n180 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C903 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n181 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.79fF
C904 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n182 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.42fF
C905 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 127.20fF
C906 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n184 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 69.17fF
C907 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n185 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 60.42fF
C908 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n186 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 84.69fF
C909 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n187 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C910 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n188 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C911 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n189 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C912 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n190 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C913 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n191 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C914 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n192 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C915 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n193 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C916 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n194 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C917 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n195 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C918 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n196 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C919 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n197 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.62fF
C920 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n198 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 12.80fF
C921 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n199 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C922 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n200 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C923 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n201 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C924 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n202 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.59fF
C925 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n203 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C926 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n204 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C927 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n205 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C928 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n206 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C929 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n207 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.46fF
C930 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n208 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 5.38fF
C931 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n209 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.56fF
C932 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n210 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.79fF
C933 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n211 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.42fF
C934 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n213 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 4.42fF
C935 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n215 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 69.17fF
C936 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1.n216 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 53.59fF
C937 cascode_1_0/SD2R cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 10.34fF
C938 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n0 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 63.48fF
C939 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 14.32fF
C940 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 14.32fF
C941 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n3 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 54.02fF
C942 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 8.38fF
C943 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n4 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 71.91fF
C944 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 8.38fF
C945 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n5 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 50.39fF
C946 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n6 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 14.32fF
C947 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n7 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 11.97fF
C948 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n8 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 6.92fF
C949 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n9 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 11.97fF
C950 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n10 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 6.92fF
C951 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD2 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 8.17fF
C952 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.71fF $ **FLOATING
C953 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n11 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C954 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n12 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C955 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n13 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C956 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n14 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C957 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n15 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C958 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n16 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C959 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n17 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C960 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n18 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C961 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n19 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C962 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n20 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C963 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n21 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C964 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n22 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C965 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n23 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C966 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t89 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.71fF $ **FLOATING
C967 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t121 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 72.80fF $ **FLOATING
C968 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t123 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 154.65fF $ **FLOATING
C969 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n24 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 107.81fF
C970 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t120 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 167.05fF $ **FLOATING
C971 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n25 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C972 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n26 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C973 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n27 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C974 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n28 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C975 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n29 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C976 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n30 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C977 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n31 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C978 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n32 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C979 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n33 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C980 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n34 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C981 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n35 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.03fF
C982 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n36 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.99fF
C983 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n37 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.99fF
C984 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n38 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.99fF
C985 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.99fF
C986 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n40 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C987 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n41 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C988 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n42 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C989 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n43 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C990 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n44 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C991 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n45 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C992 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n46 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C993 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n47 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C994 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n48 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C995 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n49 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C996 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n50 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C997 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.71fF $ **FLOATING
C998 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n51 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C999 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n52 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C1000 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n53 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
C1001 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.t39 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.70fF $ **FLOATING
C1002 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n54 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1003 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n55 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1004 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n56 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1005 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n57 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1006 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n58 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1007 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n59 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1008 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n60 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1009 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n61 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1010 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n62 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1011 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n63 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.01fF
C1012 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n64 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.03fF
C1013 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n65 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.99fF
C1014 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n66 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.99fF
C1015 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n67 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.99fF
C1016 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n68 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 2.99fF
C1017 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n69 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 85.76fF
C1018 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n70 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 49.95fF
C1019 VSSH cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 37.72fF
C1020 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n71 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 131.34fF
C1021 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2.n72 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB 3.00fF
