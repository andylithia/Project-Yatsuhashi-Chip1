magic
tech sky130A
timestamp 1664506494
<< metal4 >>
rect -6700 25850 -5950 25900
rect -6700 25250 -6650 25850
rect -6000 25250 -5950 25850
rect -6700 24250 -5950 25250
rect -2600 25850 -1850 25900
rect -2600 25250 -2550 25850
rect -1900 25250 -1850 25850
rect -4800 24950 -4050 25000
rect -4800 24350 -4750 24950
rect -4100 24350 -4050 24950
rect -4800 24200 -4050 24350
rect -3550 24950 -2800 25000
rect -3550 24350 -3500 24950
rect -2850 24350 -2800 24950
rect -3550 24200 -2800 24350
rect -2600 24300 -1850 25250
rect -400 25850 350 25900
rect -400 25250 -350 25850
rect 300 25250 350 25850
rect -400 24300 350 25250
rect 3700 25850 4450 25900
rect 3700 25250 3750 25850
rect 4400 25250 4450 25850
rect 1500 24950 2250 25000
rect 1500 24350 1550 24950
rect 2200 24350 2250 24950
rect 1500 24200 2250 24350
rect 2750 24950 3500 25000
rect 2750 24350 2800 24950
rect 3450 24350 3500 24950
rect 2750 24200 3500 24350
rect 3700 24250 4450 25250
rect -6700 18400 -5950 18450
rect -6700 17800 -6650 18400
rect -6000 17800 -5950 18400
rect -6700 17350 -5950 17800
rect -5750 17300 -5000 18500
rect -3550 18400 -2800 18900
rect -3550 17800 -3500 18400
rect -2850 17800 -2800 18400
rect -3550 17750 -2800 17800
rect -2600 18400 -1850 18450
rect -2600 17800 -2550 18400
rect -1900 17800 -1850 18400
rect -5750 16700 -5700 17300
rect -5050 16700 -5000 17300
rect -5750 16650 -5000 16700
rect -4800 17300 -4050 17350
rect -4800 16700 -4750 17300
rect -4100 16700 -4050 17300
rect -4800 16650 -4050 16700
rect -3550 17300 -2800 17350
rect -3550 16700 -3500 17300
rect -2850 16700 -2800 17300
rect -3550 16650 -2800 16700
rect -2600 16650 -1850 17800
rect -1650 17300 -900 18500
rect -1650 16700 -1600 17300
rect -950 16700 -900 17300
rect -1650 16650 -900 16700
rect -400 18400 350 18450
rect -400 17800 -350 18400
rect 300 17800 350 18400
rect 2750 18400 3500 18500
rect -400 16650 350 17800
rect 550 17300 1300 18300
rect 2750 17800 2800 18400
rect 3450 17800 3500 18400
rect 2750 17750 3500 17800
rect 3700 18400 4450 18450
rect 3700 17800 3750 18400
rect 4400 17800 4450 18400
rect 550 16700 600 17300
rect 1250 16700 1300 17300
rect 550 16650 1300 16700
rect 1500 17300 2250 17350
rect 1500 16700 1550 17300
rect 2200 16700 2250 17300
rect 1500 16600 2250 16700
rect 2750 17300 3500 17350
rect 2750 16700 2800 17300
rect 3450 16700 3500 17300
rect 2750 16600 3500 16700
rect 3700 16600 4450 17800
rect 4650 17300 5400 18450
rect 4650 16700 4700 17300
rect 5350 16700 5400 17300
rect 4650 16650 5400 16700
rect -6700 10750 -5950 10850
rect -6700 10150 -6650 10750
rect -6000 10150 -5950 10750
rect -6700 9700 -5950 10150
rect -5750 9650 -5000 10850
rect -3550 10750 -2800 11250
rect -3550 10150 -3500 10750
rect -2850 10150 -2800 10750
rect -3550 10100 -2800 10150
rect -2600 10750 -1850 10800
rect -2600 10150 -2550 10750
rect -1900 10150 -1850 10750
rect -5750 9050 -5700 9650
rect -5050 9050 -5000 9650
rect -5750 9000 -5000 9050
rect -4800 9650 -4050 9700
rect -4800 9050 -4750 9650
rect -4100 9050 -4050 9650
rect -4800 8550 -4050 9050
rect -3550 9650 -2800 9700
rect -3550 9050 -3500 9650
rect -2850 9050 -2800 9650
rect -2600 9600 -1850 10150
rect -1650 9650 -900 10850
rect -3550 8550 -2800 9050
rect -1650 9050 -1600 9650
rect -950 9050 -900 9650
rect -1650 9000 -900 9050
rect -400 10750 350 10800
rect -400 10150 -350 10750
rect 300 10150 350 10750
rect 2750 10750 3500 10850
rect -400 9000 350 10150
rect 550 9650 1300 10650
rect 2750 10150 2800 10750
rect 3450 10150 3500 10750
rect 2750 10100 3500 10150
rect 3700 10750 4450 10800
rect 3700 10150 3750 10750
rect 4400 10150 4450 10750
rect 550 9050 600 9650
rect 1250 9050 1300 9650
rect 550 9000 1300 9050
rect 1500 9650 2250 9700
rect 1500 9050 1550 9650
rect 2200 9050 2250 9650
rect 1500 9000 2250 9050
rect 2750 9650 3500 9700
rect 2750 9050 2800 9650
rect 3450 9050 3500 9650
rect 2750 9000 3500 9050
rect 3700 8950 4450 10150
rect 4650 9650 5400 10800
rect 4650 9050 4700 9650
rect 5350 9050 5400 9650
rect 4650 9000 5400 9050
rect -5750 2700 -5000 3650
rect -5750 2100 -5700 2700
rect -5050 2100 -5000 2700
rect -5750 2050 -5000 2100
rect -1650 2700 -900 3650
rect -1650 2100 -1600 2700
rect -950 2100 -900 2700
rect -1650 2050 -900 2100
rect 550 2700 1300 3650
rect 550 2100 600 2700
rect 1250 2100 1300 2700
rect 550 2050 1300 2100
rect 4650 2700 5400 3650
rect 4650 2100 4700 2700
rect 5350 2100 5400 2700
rect 4650 2050 5400 2100
<< via4 >>
rect -6650 25250 -6000 25850
rect -2550 25250 -1900 25850
rect -4750 24350 -4100 24950
rect -3500 24350 -2850 24950
rect -350 25250 300 25850
rect 3750 25250 4400 25850
rect 1550 24350 2200 24950
rect 2800 24350 3450 24950
rect -6650 17800 -6000 18400
rect -3500 17800 -2850 18400
rect -2550 17800 -1900 18400
rect -5700 16700 -5050 17300
rect -4750 16700 -4100 17300
rect -3500 16700 -2850 17300
rect -1600 16700 -950 17300
rect -350 17800 300 18400
rect 2800 17800 3450 18400
rect 3750 17800 4400 18400
rect 600 16700 1250 17300
rect 1550 16700 2200 17300
rect 2800 16700 3450 17300
rect 4700 16700 5350 17300
rect -6650 10150 -6000 10750
rect -3500 10150 -2850 10750
rect -2550 10150 -1900 10750
rect -5700 9050 -5050 9650
rect -4750 9050 -4100 9650
rect -3500 9050 -2850 9650
rect -1600 9050 -950 9650
rect -350 10150 300 10750
rect 2800 10150 3450 10750
rect 3750 10150 4400 10750
rect 600 9050 1250 9650
rect 1550 9050 2200 9650
rect 2800 9050 3450 9650
rect 4700 9050 5350 9650
rect -6650 3000 -6000 3600
rect -3500 3000 -2850 3600
rect -5700 2100 -5050 2700
rect -350 3000 300 3600
rect -1600 2100 -950 2700
rect 2800 3000 3450 3600
rect 600 2100 1250 2700
rect 4700 2100 5350 2700
<< metal5 >>
rect -6700 25900 -5950 26100
rect -6700 25850 4450 25900
rect -6700 25250 -6650 25850
rect -6000 25250 -2550 25850
rect -1900 25250 -350 25850
rect 300 25250 3750 25850
rect 4400 25250 4450 25850
rect -6700 25200 4450 25250
rect 4650 25000 5400 26100
rect -4800 24950 5400 25000
rect -4800 24350 -4750 24950
rect -4100 24350 -3500 24950
rect -2850 24350 1550 24950
rect 2200 24350 2800 24950
rect 3450 24350 5400 24950
rect -4800 24300 5400 24350
rect -6750 21700 -6700 21950
rect -6750 21250 -6700 21500
rect -6700 18400 5400 18450
rect -6700 17800 -6650 18400
rect -6000 17800 -3500 18400
rect -2850 17800 -2550 18400
rect -1900 17800 -350 18400
rect 300 17800 2800 18400
rect 3450 17800 3750 18400
rect 4400 17800 5400 18400
rect -6700 17750 5400 17800
rect -6700 17300 5400 17350
rect -6700 16700 -5700 17300
rect -5050 16700 -4750 17300
rect -4100 16700 -3500 17300
rect -2850 16700 -1600 17300
rect -950 16700 600 17300
rect 1250 16700 1550 17300
rect 2200 16700 2800 17300
rect 3450 16700 4700 17300
rect 5350 16700 5400 17300
rect -6700 16650 5400 16700
rect -6750 14050 -6700 14300
rect -6750 13600 -6700 13850
rect -6700 10750 5400 10800
rect -6700 10150 -6650 10750
rect -6000 10150 -3500 10750
rect -2850 10150 -2550 10750
rect -1900 10150 -350 10750
rect 300 10150 2800 10750
rect 3450 10150 3750 10750
rect 4400 10150 5400 10750
rect -6700 10100 5400 10150
rect -6700 9650 5400 9700
rect -6700 9050 -5700 9650
rect -5050 9050 -4750 9650
rect -4100 9050 -3500 9650
rect -2850 9050 -1600 9650
rect -950 9050 600 9650
rect 1250 9050 1550 9650
rect 2200 9050 2800 9650
rect 3450 9050 4700 9650
rect 5350 9050 5400 9650
rect -6700 9000 5400 9050
rect -6750 6400 -6700 6650
rect -6750 5950 -6700 6200
rect -6700 3600 3500 3650
rect -6700 3000 -6650 3600
rect -6000 3000 -3500 3600
rect -2850 3000 -350 3600
rect 300 3000 2800 3600
rect 3450 3000 3500 3600
rect -6700 2950 3500 3000
rect -6700 1850 -5950 2950
rect -5750 2700 5400 2750
rect -5750 2100 -5700 2700
rect -5050 2100 -1600 2700
rect -950 2100 600 2700
rect 1250 2100 4700 2700
rect 5350 2100 5400 2700
rect -5750 2050 5400 2100
rect 4650 1850 5400 2050
<< comment >>
rect -7250 24900 -7200 24950
rect -7300 24800 -7250 24900
rect -7200 24800 -7150 24850
rect -7300 24750 -7150 24800
rect -7200 24700 -7150 24750
rect -7350 17550 -7200 17600
rect -7250 17500 -7200 17550
rect -7300 17450 -7200 17500
rect -7250 17400 -7200 17450
rect -7350 17350 -7200 17400
rect -7300 9650 -7150 9700
rect -7200 9600 -7150 9650
rect -7250 9550 -7150 9600
rect -7300 9500 -7250 9550
rect -7300 9450 -7150 9500
rect -7150 2250 -7100 2300
rect -7200 2200 -7100 2250
rect -7150 2100 -7100 2200
rect -7200 2050 -7050 2100
use NMOS_30_0p5_30_diff4x_2s  NMOS_30_0p5_30_diff4x_2s_0
timestamp 1664504783
transform 1 0 -7400 0 1 6400
box 650 -3650 12800 3500
use NMOS_30_0p5_30_diff4x_2s  NMOS_30_0p5_30_diff4x_2s_1
timestamp 1664504783
transform 1 0 -7400 0 1 14050
box 650 -3650 12800 3500
use NMOS_30_0p5_30_diff4x_2s  NMOS_30_0p5_30_diff4x_2s_2
timestamp 1664504783
transform 1 0 -7400 0 1 21700
box 650 -3650 12800 3500
<< labels >>
rlabel metal5 -6700 1850 -5950 2050 1 SD1L
rlabel metal5 4650 1850 5400 2050 1 SD1R
rlabel metal5 -6700 9000 -6550 9700 1 SD2R
rlabel metal5 -6700 10100 -6550 10800 1 SD2L
rlabel metal5 -6700 16650 -6550 17350 1 SD3R
rlabel metal5 -6700 17750 -6550 18450 1 SD3L
rlabel metal5 -6700 25900 -5950 26100 1 SD4L
rlabel metal5 4650 25900 5400 26100 1 SD4R
rlabel metal5 -6750 6400 -6700 6650 1 G12L
rlabel metal5 -6750 5950 -6700 6200 1 G12R
rlabel metal5 -6750 13600 -6700 13850 1 G23R
rlabel metal5 -6750 14050 -6700 14300 1 G23L
rlabel metal5 -6750 21250 -6700 21500 1 G34R
rlabel metal5 -6750 21700 -6700 21950 1 G34L
<< end >>
