magic
tech sky130B
timestamp 1661296025
<< error_p >>
rect 5 23 28 29
rect 5 6 8 23
rect 5 0 28 6
<< locali >>
rect 0 6 8 23
rect 25 6 33 23
<< viali >>
rect 8 6 25 23
<< metal1 >>
rect 5 23 28 29
rect 5 6 8 23
rect 25 6 28 23
rect 5 0 28 6
<< properties >>
string FIXED_BBOX 0 0 33 29
<< end >>
