magic
tech sky130B
magscale 1 2
timestamp 1606074388
<< pwell >>
rect -5446 -3098 5446 3098
<< psubdiff >>
rect -5410 3028 -5314 3062
rect 5314 3028 5410 3062
rect -5410 2966 -5376 3028
rect 5376 2966 5410 3028
rect -5410 -3028 -5376 -2966
rect 5376 -3028 5410 -2966
rect -5410 -3062 -5314 -3028
rect 5314 -3062 5410 -3028
<< psubdiffcont >>
rect -5314 3028 5314 3062
rect -5410 -2966 -5376 2966
rect 5376 -2966 5410 2966
rect -5314 -3062 5314 -3028
<< xpolycontact >>
rect -5280 2500 -5142 2932
rect -5280 -2932 -5142 -2500
rect -4894 2500 -4756 2932
rect -4894 -2932 -4756 -2500
rect -4508 2500 -4370 2932
rect -4508 -2932 -4370 -2500
rect -4122 2500 -3984 2932
rect -4122 -2932 -3984 -2500
rect -3736 2500 -3598 2932
rect -3736 -2932 -3598 -2500
rect -3350 2500 -3212 2932
rect -3350 -2932 -3212 -2500
rect -2964 2500 -2826 2932
rect -2964 -2932 -2826 -2500
rect -2578 2500 -2440 2932
rect -2578 -2932 -2440 -2500
rect -2192 2500 -2054 2932
rect -2192 -2932 -2054 -2500
rect -1806 2500 -1668 2932
rect -1806 -2932 -1668 -2500
rect -1420 2500 -1282 2932
rect -1420 -2932 -1282 -2500
rect -1034 2500 -896 2932
rect -1034 -2932 -896 -2500
rect -648 2500 -510 2932
rect -648 -2932 -510 -2500
rect -262 2500 -124 2932
rect -262 -2932 -124 -2500
rect 124 2500 262 2932
rect 124 -2932 262 -2500
rect 510 2500 648 2932
rect 510 -2932 648 -2500
rect 896 2500 1034 2932
rect 896 -2932 1034 -2500
rect 1282 2500 1420 2932
rect 1282 -2932 1420 -2500
rect 1668 2500 1806 2932
rect 1668 -2932 1806 -2500
rect 2054 2500 2192 2932
rect 2054 -2932 2192 -2500
rect 2440 2500 2578 2932
rect 2440 -2932 2578 -2500
rect 2826 2500 2964 2932
rect 2826 -2932 2964 -2500
rect 3212 2500 3350 2932
rect 3212 -2932 3350 -2500
rect 3598 2500 3736 2932
rect 3598 -2932 3736 -2500
rect 3984 2500 4122 2932
rect 3984 -2932 4122 -2500
rect 4370 2500 4508 2932
rect 4370 -2932 4508 -2500
rect 4756 2500 4894 2932
rect 4756 -2932 4894 -2500
rect 5142 2500 5280 2932
rect 5142 -2932 5280 -2500
<< xpolyres >>
rect -5280 -2500 -5142 2500
rect -4894 -2500 -4756 2500
rect -4508 -2500 -4370 2500
rect -4122 -2500 -3984 2500
rect -3736 -2500 -3598 2500
rect -3350 -2500 -3212 2500
rect -2964 -2500 -2826 2500
rect -2578 -2500 -2440 2500
rect -2192 -2500 -2054 2500
rect -1806 -2500 -1668 2500
rect -1420 -2500 -1282 2500
rect -1034 -2500 -896 2500
rect -648 -2500 -510 2500
rect -262 -2500 -124 2500
rect 124 -2500 262 2500
rect 510 -2500 648 2500
rect 896 -2500 1034 2500
rect 1282 -2500 1420 2500
rect 1668 -2500 1806 2500
rect 2054 -2500 2192 2500
rect 2440 -2500 2578 2500
rect 2826 -2500 2964 2500
rect 3212 -2500 3350 2500
rect 3598 -2500 3736 2500
rect 3984 -2500 4122 2500
rect 4370 -2500 4508 2500
rect 4756 -2500 4894 2500
rect 5142 -2500 5280 2500
<< locali >>
rect -5410 3028 -5314 3062
rect 5314 3028 5410 3062
rect -5410 2966 -5376 3028
rect 5376 2966 5410 3028
rect -5410 -3028 -5376 -2966
rect 5376 -3028 5410 -2966
rect -5410 -3062 -5314 -3028
rect 5314 -3062 5410 -3028
<< viali >>
rect -5410 -2725 -5376 2725
rect 5376 -2725 5410 2725
rect -4838 -3062 4838 -3028
<< metal1 >>
rect -5416 2725 -5370 2737
rect -5416 -2725 -5410 2725
rect -5376 -2725 -5370 2725
rect -5416 -2737 -5370 -2725
rect 5370 2725 5416 2737
rect 5370 -2725 5376 2725
rect 5410 -2725 5416 2725
rect 5370 -2737 5416 -2725
rect -4850 -3028 4850 -3022
rect -4850 -3062 -4838 -3028
rect 4838 -3062 4850 -3028
rect -4850 -3068 4850 -3062
<< res0p69 >>
rect -5282 -2502 -5140 2502
rect -4896 -2502 -4754 2502
rect -4510 -2502 -4368 2502
rect -4124 -2502 -3982 2502
rect -3738 -2502 -3596 2502
rect -3352 -2502 -3210 2502
rect -2966 -2502 -2824 2502
rect -2580 -2502 -2438 2502
rect -2194 -2502 -2052 2502
rect -1808 -2502 -1666 2502
rect -1422 -2502 -1280 2502
rect -1036 -2502 -894 2502
rect -650 -2502 -508 2502
rect -264 -2502 -122 2502
rect 122 -2502 264 2502
rect 508 -2502 650 2502
rect 894 -2502 1036 2502
rect 1280 -2502 1422 2502
rect 1666 -2502 1808 2502
rect 2052 -2502 2194 2502
rect 2438 -2502 2580 2502
rect 2824 -2502 2966 2502
rect 3210 -2502 3352 2502
rect 3596 -2502 3738 2502
rect 3982 -2502 4124 2502
rect 4368 -2502 4510 2502
rect 4754 -2502 4896 2502
rect 5140 -2502 5282 2502
<< properties >>
string FIXED_BBOX -5393 -3045 5393 3045
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.69 l 25.0 m 1 nx 28 wmin 0.690 lmin 0.50 rho 2000 val 72.811k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 vias 0 viagb 90 viagt 0 viagl 90 viagr 90
<< end >>
