magic
tech sky130B
magscale 1 2
timestamp 1660188747
<< pwell >>
rect -2727 -2185 2727 2185
<< nnmos >>
rect -2499 1127 -2399 1927
rect -2341 1127 -2241 1927
rect -2183 1127 -2083 1927
rect -2025 1127 -1925 1927
rect -1867 1127 -1767 1927
rect -1709 1127 -1609 1927
rect -1551 1127 -1451 1927
rect -1393 1127 -1293 1927
rect -1235 1127 -1135 1927
rect -1077 1127 -977 1927
rect -919 1127 -819 1927
rect -761 1127 -661 1927
rect -603 1127 -503 1927
rect -445 1127 -345 1927
rect -287 1127 -187 1927
rect -129 1127 -29 1927
rect 29 1127 129 1927
rect 187 1127 287 1927
rect 345 1127 445 1927
rect 503 1127 603 1927
rect 661 1127 761 1927
rect 819 1127 919 1927
rect 977 1127 1077 1927
rect 1135 1127 1235 1927
rect 1293 1127 1393 1927
rect 1451 1127 1551 1927
rect 1609 1127 1709 1927
rect 1767 1127 1867 1927
rect 1925 1127 2025 1927
rect 2083 1127 2183 1927
rect 2241 1127 2341 1927
rect 2399 1127 2499 1927
rect -2499 109 -2399 909
rect -2341 109 -2241 909
rect -2183 109 -2083 909
rect -2025 109 -1925 909
rect -1867 109 -1767 909
rect -1709 109 -1609 909
rect -1551 109 -1451 909
rect -1393 109 -1293 909
rect -1235 109 -1135 909
rect -1077 109 -977 909
rect -919 109 -819 909
rect -761 109 -661 909
rect -603 109 -503 909
rect -445 109 -345 909
rect -287 109 -187 909
rect -129 109 -29 909
rect 29 109 129 909
rect 187 109 287 909
rect 345 109 445 909
rect 503 109 603 909
rect 661 109 761 909
rect 819 109 919 909
rect 977 109 1077 909
rect 1135 109 1235 909
rect 1293 109 1393 909
rect 1451 109 1551 909
rect 1609 109 1709 909
rect 1767 109 1867 909
rect 1925 109 2025 909
rect 2083 109 2183 909
rect 2241 109 2341 909
rect 2399 109 2499 909
rect -2499 -909 -2399 -109
rect -2341 -909 -2241 -109
rect -2183 -909 -2083 -109
rect -2025 -909 -1925 -109
rect -1867 -909 -1767 -109
rect -1709 -909 -1609 -109
rect -1551 -909 -1451 -109
rect -1393 -909 -1293 -109
rect -1235 -909 -1135 -109
rect -1077 -909 -977 -109
rect -919 -909 -819 -109
rect -761 -909 -661 -109
rect -603 -909 -503 -109
rect -445 -909 -345 -109
rect -287 -909 -187 -109
rect -129 -909 -29 -109
rect 29 -909 129 -109
rect 187 -909 287 -109
rect 345 -909 445 -109
rect 503 -909 603 -109
rect 661 -909 761 -109
rect 819 -909 919 -109
rect 977 -909 1077 -109
rect 1135 -909 1235 -109
rect 1293 -909 1393 -109
rect 1451 -909 1551 -109
rect 1609 -909 1709 -109
rect 1767 -909 1867 -109
rect 1925 -909 2025 -109
rect 2083 -909 2183 -109
rect 2241 -909 2341 -109
rect 2399 -909 2499 -109
rect -2499 -1927 -2399 -1127
rect -2341 -1927 -2241 -1127
rect -2183 -1927 -2083 -1127
rect -2025 -1927 -1925 -1127
rect -1867 -1927 -1767 -1127
rect -1709 -1927 -1609 -1127
rect -1551 -1927 -1451 -1127
rect -1393 -1927 -1293 -1127
rect -1235 -1927 -1135 -1127
rect -1077 -1927 -977 -1127
rect -919 -1927 -819 -1127
rect -761 -1927 -661 -1127
rect -603 -1927 -503 -1127
rect -445 -1927 -345 -1127
rect -287 -1927 -187 -1127
rect -129 -1927 -29 -1127
rect 29 -1927 129 -1127
rect 187 -1927 287 -1127
rect 345 -1927 445 -1127
rect 503 -1927 603 -1127
rect 661 -1927 761 -1127
rect 819 -1927 919 -1127
rect 977 -1927 1077 -1127
rect 1135 -1927 1235 -1127
rect 1293 -1927 1393 -1127
rect 1451 -1927 1551 -1127
rect 1609 -1927 1709 -1127
rect 1767 -1927 1867 -1127
rect 1925 -1927 2025 -1127
rect 2083 -1927 2183 -1127
rect 2241 -1927 2341 -1127
rect 2399 -1927 2499 -1127
<< mvndiff >>
rect -2557 1915 -2499 1927
rect -2557 1139 -2545 1915
rect -2511 1139 -2499 1915
rect -2557 1127 -2499 1139
rect -2399 1915 -2341 1927
rect -2399 1139 -2387 1915
rect -2353 1139 -2341 1915
rect -2399 1127 -2341 1139
rect -2241 1915 -2183 1927
rect -2241 1139 -2229 1915
rect -2195 1139 -2183 1915
rect -2241 1127 -2183 1139
rect -2083 1915 -2025 1927
rect -2083 1139 -2071 1915
rect -2037 1139 -2025 1915
rect -2083 1127 -2025 1139
rect -1925 1915 -1867 1927
rect -1925 1139 -1913 1915
rect -1879 1139 -1867 1915
rect -1925 1127 -1867 1139
rect -1767 1915 -1709 1927
rect -1767 1139 -1755 1915
rect -1721 1139 -1709 1915
rect -1767 1127 -1709 1139
rect -1609 1915 -1551 1927
rect -1609 1139 -1597 1915
rect -1563 1139 -1551 1915
rect -1609 1127 -1551 1139
rect -1451 1915 -1393 1927
rect -1451 1139 -1439 1915
rect -1405 1139 -1393 1915
rect -1451 1127 -1393 1139
rect -1293 1915 -1235 1927
rect -1293 1139 -1281 1915
rect -1247 1139 -1235 1915
rect -1293 1127 -1235 1139
rect -1135 1915 -1077 1927
rect -1135 1139 -1123 1915
rect -1089 1139 -1077 1915
rect -1135 1127 -1077 1139
rect -977 1915 -919 1927
rect -977 1139 -965 1915
rect -931 1139 -919 1915
rect -977 1127 -919 1139
rect -819 1915 -761 1927
rect -819 1139 -807 1915
rect -773 1139 -761 1915
rect -819 1127 -761 1139
rect -661 1915 -603 1927
rect -661 1139 -649 1915
rect -615 1139 -603 1915
rect -661 1127 -603 1139
rect -503 1915 -445 1927
rect -503 1139 -491 1915
rect -457 1139 -445 1915
rect -503 1127 -445 1139
rect -345 1915 -287 1927
rect -345 1139 -333 1915
rect -299 1139 -287 1915
rect -345 1127 -287 1139
rect -187 1915 -129 1927
rect -187 1139 -175 1915
rect -141 1139 -129 1915
rect -187 1127 -129 1139
rect -29 1915 29 1927
rect -29 1139 -17 1915
rect 17 1139 29 1915
rect -29 1127 29 1139
rect 129 1915 187 1927
rect 129 1139 141 1915
rect 175 1139 187 1915
rect 129 1127 187 1139
rect 287 1915 345 1927
rect 287 1139 299 1915
rect 333 1139 345 1915
rect 287 1127 345 1139
rect 445 1915 503 1927
rect 445 1139 457 1915
rect 491 1139 503 1915
rect 445 1127 503 1139
rect 603 1915 661 1927
rect 603 1139 615 1915
rect 649 1139 661 1915
rect 603 1127 661 1139
rect 761 1915 819 1927
rect 761 1139 773 1915
rect 807 1139 819 1915
rect 761 1127 819 1139
rect 919 1915 977 1927
rect 919 1139 931 1915
rect 965 1139 977 1915
rect 919 1127 977 1139
rect 1077 1915 1135 1927
rect 1077 1139 1089 1915
rect 1123 1139 1135 1915
rect 1077 1127 1135 1139
rect 1235 1915 1293 1927
rect 1235 1139 1247 1915
rect 1281 1139 1293 1915
rect 1235 1127 1293 1139
rect 1393 1915 1451 1927
rect 1393 1139 1405 1915
rect 1439 1139 1451 1915
rect 1393 1127 1451 1139
rect 1551 1915 1609 1927
rect 1551 1139 1563 1915
rect 1597 1139 1609 1915
rect 1551 1127 1609 1139
rect 1709 1915 1767 1927
rect 1709 1139 1721 1915
rect 1755 1139 1767 1915
rect 1709 1127 1767 1139
rect 1867 1915 1925 1927
rect 1867 1139 1879 1915
rect 1913 1139 1925 1915
rect 1867 1127 1925 1139
rect 2025 1915 2083 1927
rect 2025 1139 2037 1915
rect 2071 1139 2083 1915
rect 2025 1127 2083 1139
rect 2183 1915 2241 1927
rect 2183 1139 2195 1915
rect 2229 1139 2241 1915
rect 2183 1127 2241 1139
rect 2341 1915 2399 1927
rect 2341 1139 2353 1915
rect 2387 1139 2399 1915
rect 2341 1127 2399 1139
rect 2499 1915 2557 1927
rect 2499 1139 2511 1915
rect 2545 1139 2557 1915
rect 2499 1127 2557 1139
rect -2557 897 -2499 909
rect -2557 121 -2545 897
rect -2511 121 -2499 897
rect -2557 109 -2499 121
rect -2399 897 -2341 909
rect -2399 121 -2387 897
rect -2353 121 -2341 897
rect -2399 109 -2341 121
rect -2241 897 -2183 909
rect -2241 121 -2229 897
rect -2195 121 -2183 897
rect -2241 109 -2183 121
rect -2083 897 -2025 909
rect -2083 121 -2071 897
rect -2037 121 -2025 897
rect -2083 109 -2025 121
rect -1925 897 -1867 909
rect -1925 121 -1913 897
rect -1879 121 -1867 897
rect -1925 109 -1867 121
rect -1767 897 -1709 909
rect -1767 121 -1755 897
rect -1721 121 -1709 897
rect -1767 109 -1709 121
rect -1609 897 -1551 909
rect -1609 121 -1597 897
rect -1563 121 -1551 897
rect -1609 109 -1551 121
rect -1451 897 -1393 909
rect -1451 121 -1439 897
rect -1405 121 -1393 897
rect -1451 109 -1393 121
rect -1293 897 -1235 909
rect -1293 121 -1281 897
rect -1247 121 -1235 897
rect -1293 109 -1235 121
rect -1135 897 -1077 909
rect -1135 121 -1123 897
rect -1089 121 -1077 897
rect -1135 109 -1077 121
rect -977 897 -919 909
rect -977 121 -965 897
rect -931 121 -919 897
rect -977 109 -919 121
rect -819 897 -761 909
rect -819 121 -807 897
rect -773 121 -761 897
rect -819 109 -761 121
rect -661 897 -603 909
rect -661 121 -649 897
rect -615 121 -603 897
rect -661 109 -603 121
rect -503 897 -445 909
rect -503 121 -491 897
rect -457 121 -445 897
rect -503 109 -445 121
rect -345 897 -287 909
rect -345 121 -333 897
rect -299 121 -287 897
rect -345 109 -287 121
rect -187 897 -129 909
rect -187 121 -175 897
rect -141 121 -129 897
rect -187 109 -129 121
rect -29 897 29 909
rect -29 121 -17 897
rect 17 121 29 897
rect -29 109 29 121
rect 129 897 187 909
rect 129 121 141 897
rect 175 121 187 897
rect 129 109 187 121
rect 287 897 345 909
rect 287 121 299 897
rect 333 121 345 897
rect 287 109 345 121
rect 445 897 503 909
rect 445 121 457 897
rect 491 121 503 897
rect 445 109 503 121
rect 603 897 661 909
rect 603 121 615 897
rect 649 121 661 897
rect 603 109 661 121
rect 761 897 819 909
rect 761 121 773 897
rect 807 121 819 897
rect 761 109 819 121
rect 919 897 977 909
rect 919 121 931 897
rect 965 121 977 897
rect 919 109 977 121
rect 1077 897 1135 909
rect 1077 121 1089 897
rect 1123 121 1135 897
rect 1077 109 1135 121
rect 1235 897 1293 909
rect 1235 121 1247 897
rect 1281 121 1293 897
rect 1235 109 1293 121
rect 1393 897 1451 909
rect 1393 121 1405 897
rect 1439 121 1451 897
rect 1393 109 1451 121
rect 1551 897 1609 909
rect 1551 121 1563 897
rect 1597 121 1609 897
rect 1551 109 1609 121
rect 1709 897 1767 909
rect 1709 121 1721 897
rect 1755 121 1767 897
rect 1709 109 1767 121
rect 1867 897 1925 909
rect 1867 121 1879 897
rect 1913 121 1925 897
rect 1867 109 1925 121
rect 2025 897 2083 909
rect 2025 121 2037 897
rect 2071 121 2083 897
rect 2025 109 2083 121
rect 2183 897 2241 909
rect 2183 121 2195 897
rect 2229 121 2241 897
rect 2183 109 2241 121
rect 2341 897 2399 909
rect 2341 121 2353 897
rect 2387 121 2399 897
rect 2341 109 2399 121
rect 2499 897 2557 909
rect 2499 121 2511 897
rect 2545 121 2557 897
rect 2499 109 2557 121
rect -2557 -121 -2499 -109
rect -2557 -897 -2545 -121
rect -2511 -897 -2499 -121
rect -2557 -909 -2499 -897
rect -2399 -121 -2341 -109
rect -2399 -897 -2387 -121
rect -2353 -897 -2341 -121
rect -2399 -909 -2341 -897
rect -2241 -121 -2183 -109
rect -2241 -897 -2229 -121
rect -2195 -897 -2183 -121
rect -2241 -909 -2183 -897
rect -2083 -121 -2025 -109
rect -2083 -897 -2071 -121
rect -2037 -897 -2025 -121
rect -2083 -909 -2025 -897
rect -1925 -121 -1867 -109
rect -1925 -897 -1913 -121
rect -1879 -897 -1867 -121
rect -1925 -909 -1867 -897
rect -1767 -121 -1709 -109
rect -1767 -897 -1755 -121
rect -1721 -897 -1709 -121
rect -1767 -909 -1709 -897
rect -1609 -121 -1551 -109
rect -1609 -897 -1597 -121
rect -1563 -897 -1551 -121
rect -1609 -909 -1551 -897
rect -1451 -121 -1393 -109
rect -1451 -897 -1439 -121
rect -1405 -897 -1393 -121
rect -1451 -909 -1393 -897
rect -1293 -121 -1235 -109
rect -1293 -897 -1281 -121
rect -1247 -897 -1235 -121
rect -1293 -909 -1235 -897
rect -1135 -121 -1077 -109
rect -1135 -897 -1123 -121
rect -1089 -897 -1077 -121
rect -1135 -909 -1077 -897
rect -977 -121 -919 -109
rect -977 -897 -965 -121
rect -931 -897 -919 -121
rect -977 -909 -919 -897
rect -819 -121 -761 -109
rect -819 -897 -807 -121
rect -773 -897 -761 -121
rect -819 -909 -761 -897
rect -661 -121 -603 -109
rect -661 -897 -649 -121
rect -615 -897 -603 -121
rect -661 -909 -603 -897
rect -503 -121 -445 -109
rect -503 -897 -491 -121
rect -457 -897 -445 -121
rect -503 -909 -445 -897
rect -345 -121 -287 -109
rect -345 -897 -333 -121
rect -299 -897 -287 -121
rect -345 -909 -287 -897
rect -187 -121 -129 -109
rect -187 -897 -175 -121
rect -141 -897 -129 -121
rect -187 -909 -129 -897
rect -29 -121 29 -109
rect -29 -897 -17 -121
rect 17 -897 29 -121
rect -29 -909 29 -897
rect 129 -121 187 -109
rect 129 -897 141 -121
rect 175 -897 187 -121
rect 129 -909 187 -897
rect 287 -121 345 -109
rect 287 -897 299 -121
rect 333 -897 345 -121
rect 287 -909 345 -897
rect 445 -121 503 -109
rect 445 -897 457 -121
rect 491 -897 503 -121
rect 445 -909 503 -897
rect 603 -121 661 -109
rect 603 -897 615 -121
rect 649 -897 661 -121
rect 603 -909 661 -897
rect 761 -121 819 -109
rect 761 -897 773 -121
rect 807 -897 819 -121
rect 761 -909 819 -897
rect 919 -121 977 -109
rect 919 -897 931 -121
rect 965 -897 977 -121
rect 919 -909 977 -897
rect 1077 -121 1135 -109
rect 1077 -897 1089 -121
rect 1123 -897 1135 -121
rect 1077 -909 1135 -897
rect 1235 -121 1293 -109
rect 1235 -897 1247 -121
rect 1281 -897 1293 -121
rect 1235 -909 1293 -897
rect 1393 -121 1451 -109
rect 1393 -897 1405 -121
rect 1439 -897 1451 -121
rect 1393 -909 1451 -897
rect 1551 -121 1609 -109
rect 1551 -897 1563 -121
rect 1597 -897 1609 -121
rect 1551 -909 1609 -897
rect 1709 -121 1767 -109
rect 1709 -897 1721 -121
rect 1755 -897 1767 -121
rect 1709 -909 1767 -897
rect 1867 -121 1925 -109
rect 1867 -897 1879 -121
rect 1913 -897 1925 -121
rect 1867 -909 1925 -897
rect 2025 -121 2083 -109
rect 2025 -897 2037 -121
rect 2071 -897 2083 -121
rect 2025 -909 2083 -897
rect 2183 -121 2241 -109
rect 2183 -897 2195 -121
rect 2229 -897 2241 -121
rect 2183 -909 2241 -897
rect 2341 -121 2399 -109
rect 2341 -897 2353 -121
rect 2387 -897 2399 -121
rect 2341 -909 2399 -897
rect 2499 -121 2557 -109
rect 2499 -897 2511 -121
rect 2545 -897 2557 -121
rect 2499 -909 2557 -897
rect -2557 -1139 -2499 -1127
rect -2557 -1915 -2545 -1139
rect -2511 -1915 -2499 -1139
rect -2557 -1927 -2499 -1915
rect -2399 -1139 -2341 -1127
rect -2399 -1915 -2387 -1139
rect -2353 -1915 -2341 -1139
rect -2399 -1927 -2341 -1915
rect -2241 -1139 -2183 -1127
rect -2241 -1915 -2229 -1139
rect -2195 -1915 -2183 -1139
rect -2241 -1927 -2183 -1915
rect -2083 -1139 -2025 -1127
rect -2083 -1915 -2071 -1139
rect -2037 -1915 -2025 -1139
rect -2083 -1927 -2025 -1915
rect -1925 -1139 -1867 -1127
rect -1925 -1915 -1913 -1139
rect -1879 -1915 -1867 -1139
rect -1925 -1927 -1867 -1915
rect -1767 -1139 -1709 -1127
rect -1767 -1915 -1755 -1139
rect -1721 -1915 -1709 -1139
rect -1767 -1927 -1709 -1915
rect -1609 -1139 -1551 -1127
rect -1609 -1915 -1597 -1139
rect -1563 -1915 -1551 -1139
rect -1609 -1927 -1551 -1915
rect -1451 -1139 -1393 -1127
rect -1451 -1915 -1439 -1139
rect -1405 -1915 -1393 -1139
rect -1451 -1927 -1393 -1915
rect -1293 -1139 -1235 -1127
rect -1293 -1915 -1281 -1139
rect -1247 -1915 -1235 -1139
rect -1293 -1927 -1235 -1915
rect -1135 -1139 -1077 -1127
rect -1135 -1915 -1123 -1139
rect -1089 -1915 -1077 -1139
rect -1135 -1927 -1077 -1915
rect -977 -1139 -919 -1127
rect -977 -1915 -965 -1139
rect -931 -1915 -919 -1139
rect -977 -1927 -919 -1915
rect -819 -1139 -761 -1127
rect -819 -1915 -807 -1139
rect -773 -1915 -761 -1139
rect -819 -1927 -761 -1915
rect -661 -1139 -603 -1127
rect -661 -1915 -649 -1139
rect -615 -1915 -603 -1139
rect -661 -1927 -603 -1915
rect -503 -1139 -445 -1127
rect -503 -1915 -491 -1139
rect -457 -1915 -445 -1139
rect -503 -1927 -445 -1915
rect -345 -1139 -287 -1127
rect -345 -1915 -333 -1139
rect -299 -1915 -287 -1139
rect -345 -1927 -287 -1915
rect -187 -1139 -129 -1127
rect -187 -1915 -175 -1139
rect -141 -1915 -129 -1139
rect -187 -1927 -129 -1915
rect -29 -1139 29 -1127
rect -29 -1915 -17 -1139
rect 17 -1915 29 -1139
rect -29 -1927 29 -1915
rect 129 -1139 187 -1127
rect 129 -1915 141 -1139
rect 175 -1915 187 -1139
rect 129 -1927 187 -1915
rect 287 -1139 345 -1127
rect 287 -1915 299 -1139
rect 333 -1915 345 -1139
rect 287 -1927 345 -1915
rect 445 -1139 503 -1127
rect 445 -1915 457 -1139
rect 491 -1915 503 -1139
rect 445 -1927 503 -1915
rect 603 -1139 661 -1127
rect 603 -1915 615 -1139
rect 649 -1915 661 -1139
rect 603 -1927 661 -1915
rect 761 -1139 819 -1127
rect 761 -1915 773 -1139
rect 807 -1915 819 -1139
rect 761 -1927 819 -1915
rect 919 -1139 977 -1127
rect 919 -1915 931 -1139
rect 965 -1915 977 -1139
rect 919 -1927 977 -1915
rect 1077 -1139 1135 -1127
rect 1077 -1915 1089 -1139
rect 1123 -1915 1135 -1139
rect 1077 -1927 1135 -1915
rect 1235 -1139 1293 -1127
rect 1235 -1915 1247 -1139
rect 1281 -1915 1293 -1139
rect 1235 -1927 1293 -1915
rect 1393 -1139 1451 -1127
rect 1393 -1915 1405 -1139
rect 1439 -1915 1451 -1139
rect 1393 -1927 1451 -1915
rect 1551 -1139 1609 -1127
rect 1551 -1915 1563 -1139
rect 1597 -1915 1609 -1139
rect 1551 -1927 1609 -1915
rect 1709 -1139 1767 -1127
rect 1709 -1915 1721 -1139
rect 1755 -1915 1767 -1139
rect 1709 -1927 1767 -1915
rect 1867 -1139 1925 -1127
rect 1867 -1915 1879 -1139
rect 1913 -1915 1925 -1139
rect 1867 -1927 1925 -1915
rect 2025 -1139 2083 -1127
rect 2025 -1915 2037 -1139
rect 2071 -1915 2083 -1139
rect 2025 -1927 2083 -1915
rect 2183 -1139 2241 -1127
rect 2183 -1915 2195 -1139
rect 2229 -1915 2241 -1139
rect 2183 -1927 2241 -1915
rect 2341 -1139 2399 -1127
rect 2341 -1915 2353 -1139
rect 2387 -1915 2399 -1139
rect 2341 -1927 2399 -1915
rect 2499 -1139 2557 -1127
rect 2499 -1915 2511 -1139
rect 2545 -1915 2557 -1139
rect 2499 -1927 2557 -1915
<< mvndiffc >>
rect -2545 1139 -2511 1915
rect -2387 1139 -2353 1915
rect -2229 1139 -2195 1915
rect -2071 1139 -2037 1915
rect -1913 1139 -1879 1915
rect -1755 1139 -1721 1915
rect -1597 1139 -1563 1915
rect -1439 1139 -1405 1915
rect -1281 1139 -1247 1915
rect -1123 1139 -1089 1915
rect -965 1139 -931 1915
rect -807 1139 -773 1915
rect -649 1139 -615 1915
rect -491 1139 -457 1915
rect -333 1139 -299 1915
rect -175 1139 -141 1915
rect -17 1139 17 1915
rect 141 1139 175 1915
rect 299 1139 333 1915
rect 457 1139 491 1915
rect 615 1139 649 1915
rect 773 1139 807 1915
rect 931 1139 965 1915
rect 1089 1139 1123 1915
rect 1247 1139 1281 1915
rect 1405 1139 1439 1915
rect 1563 1139 1597 1915
rect 1721 1139 1755 1915
rect 1879 1139 1913 1915
rect 2037 1139 2071 1915
rect 2195 1139 2229 1915
rect 2353 1139 2387 1915
rect 2511 1139 2545 1915
rect -2545 121 -2511 897
rect -2387 121 -2353 897
rect -2229 121 -2195 897
rect -2071 121 -2037 897
rect -1913 121 -1879 897
rect -1755 121 -1721 897
rect -1597 121 -1563 897
rect -1439 121 -1405 897
rect -1281 121 -1247 897
rect -1123 121 -1089 897
rect -965 121 -931 897
rect -807 121 -773 897
rect -649 121 -615 897
rect -491 121 -457 897
rect -333 121 -299 897
rect -175 121 -141 897
rect -17 121 17 897
rect 141 121 175 897
rect 299 121 333 897
rect 457 121 491 897
rect 615 121 649 897
rect 773 121 807 897
rect 931 121 965 897
rect 1089 121 1123 897
rect 1247 121 1281 897
rect 1405 121 1439 897
rect 1563 121 1597 897
rect 1721 121 1755 897
rect 1879 121 1913 897
rect 2037 121 2071 897
rect 2195 121 2229 897
rect 2353 121 2387 897
rect 2511 121 2545 897
rect -2545 -897 -2511 -121
rect -2387 -897 -2353 -121
rect -2229 -897 -2195 -121
rect -2071 -897 -2037 -121
rect -1913 -897 -1879 -121
rect -1755 -897 -1721 -121
rect -1597 -897 -1563 -121
rect -1439 -897 -1405 -121
rect -1281 -897 -1247 -121
rect -1123 -897 -1089 -121
rect -965 -897 -931 -121
rect -807 -897 -773 -121
rect -649 -897 -615 -121
rect -491 -897 -457 -121
rect -333 -897 -299 -121
rect -175 -897 -141 -121
rect -17 -897 17 -121
rect 141 -897 175 -121
rect 299 -897 333 -121
rect 457 -897 491 -121
rect 615 -897 649 -121
rect 773 -897 807 -121
rect 931 -897 965 -121
rect 1089 -897 1123 -121
rect 1247 -897 1281 -121
rect 1405 -897 1439 -121
rect 1563 -897 1597 -121
rect 1721 -897 1755 -121
rect 1879 -897 1913 -121
rect 2037 -897 2071 -121
rect 2195 -897 2229 -121
rect 2353 -897 2387 -121
rect 2511 -897 2545 -121
rect -2545 -1915 -2511 -1139
rect -2387 -1915 -2353 -1139
rect -2229 -1915 -2195 -1139
rect -2071 -1915 -2037 -1139
rect -1913 -1915 -1879 -1139
rect -1755 -1915 -1721 -1139
rect -1597 -1915 -1563 -1139
rect -1439 -1915 -1405 -1139
rect -1281 -1915 -1247 -1139
rect -1123 -1915 -1089 -1139
rect -965 -1915 -931 -1139
rect -807 -1915 -773 -1139
rect -649 -1915 -615 -1139
rect -491 -1915 -457 -1139
rect -333 -1915 -299 -1139
rect -175 -1915 -141 -1139
rect -17 -1915 17 -1139
rect 141 -1915 175 -1139
rect 299 -1915 333 -1139
rect 457 -1915 491 -1139
rect 615 -1915 649 -1139
rect 773 -1915 807 -1139
rect 931 -1915 965 -1139
rect 1089 -1915 1123 -1139
rect 1247 -1915 1281 -1139
rect 1405 -1915 1439 -1139
rect 1563 -1915 1597 -1139
rect 1721 -1915 1755 -1139
rect 1879 -1915 1913 -1139
rect 2037 -1915 2071 -1139
rect 2195 -1915 2229 -1139
rect 2353 -1915 2387 -1139
rect 2511 -1915 2545 -1139
<< mvpsubdiff >>
rect -2691 2137 2691 2149
rect -2691 2103 -2583 2137
rect 2583 2103 2691 2137
rect -2691 2091 2691 2103
rect -2691 2041 -2633 2091
rect -2691 -2041 -2679 2041
rect -2645 -2041 -2633 2041
rect 2633 2041 2691 2091
rect -2691 -2091 -2633 -2041
rect 2633 -2041 2645 2041
rect 2679 -2041 2691 2041
rect 2633 -2091 2691 -2041
rect -2691 -2103 2691 -2091
rect -2691 -2137 -2583 -2103
rect 2583 -2137 2691 -2103
rect -2691 -2149 2691 -2137
<< mvpsubdiffcont >>
rect -2583 2103 2583 2137
rect -2679 -2041 -2645 2041
rect 2645 -2041 2679 2041
rect -2583 -2137 2583 -2103
<< poly >>
rect -2499 1999 -2399 2015
rect -2499 1965 -2483 1999
rect -2415 1965 -2399 1999
rect -2499 1927 -2399 1965
rect -2341 1999 -2241 2015
rect -2341 1965 -2325 1999
rect -2257 1965 -2241 1999
rect -2341 1927 -2241 1965
rect -2183 1999 -2083 2015
rect -2183 1965 -2167 1999
rect -2099 1965 -2083 1999
rect -2183 1927 -2083 1965
rect -2025 1999 -1925 2015
rect -2025 1965 -2009 1999
rect -1941 1965 -1925 1999
rect -2025 1927 -1925 1965
rect -1867 1999 -1767 2015
rect -1867 1965 -1851 1999
rect -1783 1965 -1767 1999
rect -1867 1927 -1767 1965
rect -1709 1999 -1609 2015
rect -1709 1965 -1693 1999
rect -1625 1965 -1609 1999
rect -1709 1927 -1609 1965
rect -1551 1999 -1451 2015
rect -1551 1965 -1535 1999
rect -1467 1965 -1451 1999
rect -1551 1927 -1451 1965
rect -1393 1999 -1293 2015
rect -1393 1965 -1377 1999
rect -1309 1965 -1293 1999
rect -1393 1927 -1293 1965
rect -1235 1999 -1135 2015
rect -1235 1965 -1219 1999
rect -1151 1965 -1135 1999
rect -1235 1927 -1135 1965
rect -1077 1999 -977 2015
rect -1077 1965 -1061 1999
rect -993 1965 -977 1999
rect -1077 1927 -977 1965
rect -919 1999 -819 2015
rect -919 1965 -903 1999
rect -835 1965 -819 1999
rect -919 1927 -819 1965
rect -761 1999 -661 2015
rect -761 1965 -745 1999
rect -677 1965 -661 1999
rect -761 1927 -661 1965
rect -603 1999 -503 2015
rect -603 1965 -587 1999
rect -519 1965 -503 1999
rect -603 1927 -503 1965
rect -445 1999 -345 2015
rect -445 1965 -429 1999
rect -361 1965 -345 1999
rect -445 1927 -345 1965
rect -287 1999 -187 2015
rect -287 1965 -271 1999
rect -203 1965 -187 1999
rect -287 1927 -187 1965
rect -129 1999 -29 2015
rect -129 1965 -113 1999
rect -45 1965 -29 1999
rect -129 1927 -29 1965
rect 29 1999 129 2015
rect 29 1965 45 1999
rect 113 1965 129 1999
rect 29 1927 129 1965
rect 187 1999 287 2015
rect 187 1965 203 1999
rect 271 1965 287 1999
rect 187 1927 287 1965
rect 345 1999 445 2015
rect 345 1965 361 1999
rect 429 1965 445 1999
rect 345 1927 445 1965
rect 503 1999 603 2015
rect 503 1965 519 1999
rect 587 1965 603 1999
rect 503 1927 603 1965
rect 661 1999 761 2015
rect 661 1965 677 1999
rect 745 1965 761 1999
rect 661 1927 761 1965
rect 819 1999 919 2015
rect 819 1965 835 1999
rect 903 1965 919 1999
rect 819 1927 919 1965
rect 977 1999 1077 2015
rect 977 1965 993 1999
rect 1061 1965 1077 1999
rect 977 1927 1077 1965
rect 1135 1999 1235 2015
rect 1135 1965 1151 1999
rect 1219 1965 1235 1999
rect 1135 1927 1235 1965
rect 1293 1999 1393 2015
rect 1293 1965 1309 1999
rect 1377 1965 1393 1999
rect 1293 1927 1393 1965
rect 1451 1999 1551 2015
rect 1451 1965 1467 1999
rect 1535 1965 1551 1999
rect 1451 1927 1551 1965
rect 1609 1999 1709 2015
rect 1609 1965 1625 1999
rect 1693 1965 1709 1999
rect 1609 1927 1709 1965
rect 1767 1999 1867 2015
rect 1767 1965 1783 1999
rect 1851 1965 1867 1999
rect 1767 1927 1867 1965
rect 1925 1999 2025 2015
rect 1925 1965 1941 1999
rect 2009 1965 2025 1999
rect 1925 1927 2025 1965
rect 2083 1999 2183 2015
rect 2083 1965 2099 1999
rect 2167 1965 2183 1999
rect 2083 1927 2183 1965
rect 2241 1999 2341 2015
rect 2241 1965 2257 1999
rect 2325 1965 2341 1999
rect 2241 1927 2341 1965
rect 2399 1999 2499 2015
rect 2399 1965 2415 1999
rect 2483 1965 2499 1999
rect 2399 1927 2499 1965
rect -2499 1089 -2399 1127
rect -2499 1055 -2483 1089
rect -2415 1055 -2399 1089
rect -2499 1039 -2399 1055
rect -2341 1089 -2241 1127
rect -2341 1055 -2325 1089
rect -2257 1055 -2241 1089
rect -2341 1039 -2241 1055
rect -2183 1089 -2083 1127
rect -2183 1055 -2167 1089
rect -2099 1055 -2083 1089
rect -2183 1039 -2083 1055
rect -2025 1089 -1925 1127
rect -2025 1055 -2009 1089
rect -1941 1055 -1925 1089
rect -2025 1039 -1925 1055
rect -1867 1089 -1767 1127
rect -1867 1055 -1851 1089
rect -1783 1055 -1767 1089
rect -1867 1039 -1767 1055
rect -1709 1089 -1609 1127
rect -1709 1055 -1693 1089
rect -1625 1055 -1609 1089
rect -1709 1039 -1609 1055
rect -1551 1089 -1451 1127
rect -1551 1055 -1535 1089
rect -1467 1055 -1451 1089
rect -1551 1039 -1451 1055
rect -1393 1089 -1293 1127
rect -1393 1055 -1377 1089
rect -1309 1055 -1293 1089
rect -1393 1039 -1293 1055
rect -1235 1089 -1135 1127
rect -1235 1055 -1219 1089
rect -1151 1055 -1135 1089
rect -1235 1039 -1135 1055
rect -1077 1089 -977 1127
rect -1077 1055 -1061 1089
rect -993 1055 -977 1089
rect -1077 1039 -977 1055
rect -919 1089 -819 1127
rect -919 1055 -903 1089
rect -835 1055 -819 1089
rect -919 1039 -819 1055
rect -761 1089 -661 1127
rect -761 1055 -745 1089
rect -677 1055 -661 1089
rect -761 1039 -661 1055
rect -603 1089 -503 1127
rect -603 1055 -587 1089
rect -519 1055 -503 1089
rect -603 1039 -503 1055
rect -445 1089 -345 1127
rect -445 1055 -429 1089
rect -361 1055 -345 1089
rect -445 1039 -345 1055
rect -287 1089 -187 1127
rect -287 1055 -271 1089
rect -203 1055 -187 1089
rect -287 1039 -187 1055
rect -129 1089 -29 1127
rect -129 1055 -113 1089
rect -45 1055 -29 1089
rect -129 1039 -29 1055
rect 29 1089 129 1127
rect 29 1055 45 1089
rect 113 1055 129 1089
rect 29 1039 129 1055
rect 187 1089 287 1127
rect 187 1055 203 1089
rect 271 1055 287 1089
rect 187 1039 287 1055
rect 345 1089 445 1127
rect 345 1055 361 1089
rect 429 1055 445 1089
rect 345 1039 445 1055
rect 503 1089 603 1127
rect 503 1055 519 1089
rect 587 1055 603 1089
rect 503 1039 603 1055
rect 661 1089 761 1127
rect 661 1055 677 1089
rect 745 1055 761 1089
rect 661 1039 761 1055
rect 819 1089 919 1127
rect 819 1055 835 1089
rect 903 1055 919 1089
rect 819 1039 919 1055
rect 977 1089 1077 1127
rect 977 1055 993 1089
rect 1061 1055 1077 1089
rect 977 1039 1077 1055
rect 1135 1089 1235 1127
rect 1135 1055 1151 1089
rect 1219 1055 1235 1089
rect 1135 1039 1235 1055
rect 1293 1089 1393 1127
rect 1293 1055 1309 1089
rect 1377 1055 1393 1089
rect 1293 1039 1393 1055
rect 1451 1089 1551 1127
rect 1451 1055 1467 1089
rect 1535 1055 1551 1089
rect 1451 1039 1551 1055
rect 1609 1089 1709 1127
rect 1609 1055 1625 1089
rect 1693 1055 1709 1089
rect 1609 1039 1709 1055
rect 1767 1089 1867 1127
rect 1767 1055 1783 1089
rect 1851 1055 1867 1089
rect 1767 1039 1867 1055
rect 1925 1089 2025 1127
rect 1925 1055 1941 1089
rect 2009 1055 2025 1089
rect 1925 1039 2025 1055
rect 2083 1089 2183 1127
rect 2083 1055 2099 1089
rect 2167 1055 2183 1089
rect 2083 1039 2183 1055
rect 2241 1089 2341 1127
rect 2241 1055 2257 1089
rect 2325 1055 2341 1089
rect 2241 1039 2341 1055
rect 2399 1089 2499 1127
rect 2399 1055 2415 1089
rect 2483 1055 2499 1089
rect 2399 1039 2499 1055
rect -2499 981 -2399 997
rect -2499 947 -2483 981
rect -2415 947 -2399 981
rect -2499 909 -2399 947
rect -2341 981 -2241 997
rect -2341 947 -2325 981
rect -2257 947 -2241 981
rect -2341 909 -2241 947
rect -2183 981 -2083 997
rect -2183 947 -2167 981
rect -2099 947 -2083 981
rect -2183 909 -2083 947
rect -2025 981 -1925 997
rect -2025 947 -2009 981
rect -1941 947 -1925 981
rect -2025 909 -1925 947
rect -1867 981 -1767 997
rect -1867 947 -1851 981
rect -1783 947 -1767 981
rect -1867 909 -1767 947
rect -1709 981 -1609 997
rect -1709 947 -1693 981
rect -1625 947 -1609 981
rect -1709 909 -1609 947
rect -1551 981 -1451 997
rect -1551 947 -1535 981
rect -1467 947 -1451 981
rect -1551 909 -1451 947
rect -1393 981 -1293 997
rect -1393 947 -1377 981
rect -1309 947 -1293 981
rect -1393 909 -1293 947
rect -1235 981 -1135 997
rect -1235 947 -1219 981
rect -1151 947 -1135 981
rect -1235 909 -1135 947
rect -1077 981 -977 997
rect -1077 947 -1061 981
rect -993 947 -977 981
rect -1077 909 -977 947
rect -919 981 -819 997
rect -919 947 -903 981
rect -835 947 -819 981
rect -919 909 -819 947
rect -761 981 -661 997
rect -761 947 -745 981
rect -677 947 -661 981
rect -761 909 -661 947
rect -603 981 -503 997
rect -603 947 -587 981
rect -519 947 -503 981
rect -603 909 -503 947
rect -445 981 -345 997
rect -445 947 -429 981
rect -361 947 -345 981
rect -445 909 -345 947
rect -287 981 -187 997
rect -287 947 -271 981
rect -203 947 -187 981
rect -287 909 -187 947
rect -129 981 -29 997
rect -129 947 -113 981
rect -45 947 -29 981
rect -129 909 -29 947
rect 29 981 129 997
rect 29 947 45 981
rect 113 947 129 981
rect 29 909 129 947
rect 187 981 287 997
rect 187 947 203 981
rect 271 947 287 981
rect 187 909 287 947
rect 345 981 445 997
rect 345 947 361 981
rect 429 947 445 981
rect 345 909 445 947
rect 503 981 603 997
rect 503 947 519 981
rect 587 947 603 981
rect 503 909 603 947
rect 661 981 761 997
rect 661 947 677 981
rect 745 947 761 981
rect 661 909 761 947
rect 819 981 919 997
rect 819 947 835 981
rect 903 947 919 981
rect 819 909 919 947
rect 977 981 1077 997
rect 977 947 993 981
rect 1061 947 1077 981
rect 977 909 1077 947
rect 1135 981 1235 997
rect 1135 947 1151 981
rect 1219 947 1235 981
rect 1135 909 1235 947
rect 1293 981 1393 997
rect 1293 947 1309 981
rect 1377 947 1393 981
rect 1293 909 1393 947
rect 1451 981 1551 997
rect 1451 947 1467 981
rect 1535 947 1551 981
rect 1451 909 1551 947
rect 1609 981 1709 997
rect 1609 947 1625 981
rect 1693 947 1709 981
rect 1609 909 1709 947
rect 1767 981 1867 997
rect 1767 947 1783 981
rect 1851 947 1867 981
rect 1767 909 1867 947
rect 1925 981 2025 997
rect 1925 947 1941 981
rect 2009 947 2025 981
rect 1925 909 2025 947
rect 2083 981 2183 997
rect 2083 947 2099 981
rect 2167 947 2183 981
rect 2083 909 2183 947
rect 2241 981 2341 997
rect 2241 947 2257 981
rect 2325 947 2341 981
rect 2241 909 2341 947
rect 2399 981 2499 997
rect 2399 947 2415 981
rect 2483 947 2499 981
rect 2399 909 2499 947
rect -2499 71 -2399 109
rect -2499 37 -2483 71
rect -2415 37 -2399 71
rect -2499 21 -2399 37
rect -2341 71 -2241 109
rect -2341 37 -2325 71
rect -2257 37 -2241 71
rect -2341 21 -2241 37
rect -2183 71 -2083 109
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2183 21 -2083 37
rect -2025 71 -1925 109
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -2025 21 -1925 37
rect -1867 71 -1767 109
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1867 21 -1767 37
rect -1709 71 -1609 109
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1709 21 -1609 37
rect -1551 71 -1451 109
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1551 21 -1451 37
rect -1393 71 -1293 109
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1393 21 -1293 37
rect -1235 71 -1135 109
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1235 21 -1135 37
rect -1077 71 -977 109
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 109
rect -919 37 -903 71
rect -835 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 109
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 109
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 109
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 109
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 109
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 109
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 109
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 109
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 109
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 109
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect 819 71 919 109
rect 819 37 835 71
rect 903 37 919 71
rect 819 21 919 37
rect 977 71 1077 109
rect 977 37 993 71
rect 1061 37 1077 71
rect 977 21 1077 37
rect 1135 71 1235 109
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1135 21 1235 37
rect 1293 71 1393 109
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1293 21 1393 37
rect 1451 71 1551 109
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1451 21 1551 37
rect 1609 71 1709 109
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1609 21 1709 37
rect 1767 71 1867 109
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1767 21 1867 37
rect 1925 71 2025 109
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 1925 21 2025 37
rect 2083 71 2183 109
rect 2083 37 2099 71
rect 2167 37 2183 71
rect 2083 21 2183 37
rect 2241 71 2341 109
rect 2241 37 2257 71
rect 2325 37 2341 71
rect 2241 21 2341 37
rect 2399 71 2499 109
rect 2399 37 2415 71
rect 2483 37 2499 71
rect 2399 21 2499 37
rect -2499 -37 -2399 -21
rect -2499 -71 -2483 -37
rect -2415 -71 -2399 -37
rect -2499 -109 -2399 -71
rect -2341 -37 -2241 -21
rect -2341 -71 -2325 -37
rect -2257 -71 -2241 -37
rect -2341 -109 -2241 -71
rect -2183 -37 -2083 -21
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2183 -109 -2083 -71
rect -2025 -37 -1925 -21
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -2025 -109 -1925 -71
rect -1867 -37 -1767 -21
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1867 -109 -1767 -71
rect -1709 -37 -1609 -21
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1709 -109 -1609 -71
rect -1551 -37 -1451 -21
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1551 -109 -1451 -71
rect -1393 -37 -1293 -21
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1393 -109 -1293 -71
rect -1235 -37 -1135 -21
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1235 -109 -1135 -71
rect -1077 -37 -977 -21
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -1077 -109 -977 -71
rect -919 -37 -819 -21
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -919 -109 -819 -71
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -109 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -109 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -109 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -109 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -109 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -109 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -109 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -109 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -109 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -109 761 -71
rect 819 -37 919 -21
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 819 -109 919 -71
rect 977 -37 1077 -21
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 977 -109 1077 -71
rect 1135 -37 1235 -21
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1135 -109 1235 -71
rect 1293 -37 1393 -21
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1293 -109 1393 -71
rect 1451 -37 1551 -21
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1451 -109 1551 -71
rect 1609 -37 1709 -21
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1609 -109 1709 -71
rect 1767 -37 1867 -21
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1767 -109 1867 -71
rect 1925 -37 2025 -21
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 1925 -109 2025 -71
rect 2083 -37 2183 -21
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect 2083 -109 2183 -71
rect 2241 -37 2341 -21
rect 2241 -71 2257 -37
rect 2325 -71 2341 -37
rect 2241 -109 2341 -71
rect 2399 -37 2499 -21
rect 2399 -71 2415 -37
rect 2483 -71 2499 -37
rect 2399 -109 2499 -71
rect -2499 -947 -2399 -909
rect -2499 -981 -2483 -947
rect -2415 -981 -2399 -947
rect -2499 -997 -2399 -981
rect -2341 -947 -2241 -909
rect -2341 -981 -2325 -947
rect -2257 -981 -2241 -947
rect -2341 -997 -2241 -981
rect -2183 -947 -2083 -909
rect -2183 -981 -2167 -947
rect -2099 -981 -2083 -947
rect -2183 -997 -2083 -981
rect -2025 -947 -1925 -909
rect -2025 -981 -2009 -947
rect -1941 -981 -1925 -947
rect -2025 -997 -1925 -981
rect -1867 -947 -1767 -909
rect -1867 -981 -1851 -947
rect -1783 -981 -1767 -947
rect -1867 -997 -1767 -981
rect -1709 -947 -1609 -909
rect -1709 -981 -1693 -947
rect -1625 -981 -1609 -947
rect -1709 -997 -1609 -981
rect -1551 -947 -1451 -909
rect -1551 -981 -1535 -947
rect -1467 -981 -1451 -947
rect -1551 -997 -1451 -981
rect -1393 -947 -1293 -909
rect -1393 -981 -1377 -947
rect -1309 -981 -1293 -947
rect -1393 -997 -1293 -981
rect -1235 -947 -1135 -909
rect -1235 -981 -1219 -947
rect -1151 -981 -1135 -947
rect -1235 -997 -1135 -981
rect -1077 -947 -977 -909
rect -1077 -981 -1061 -947
rect -993 -981 -977 -947
rect -1077 -997 -977 -981
rect -919 -947 -819 -909
rect -919 -981 -903 -947
rect -835 -981 -819 -947
rect -919 -997 -819 -981
rect -761 -947 -661 -909
rect -761 -981 -745 -947
rect -677 -981 -661 -947
rect -761 -997 -661 -981
rect -603 -947 -503 -909
rect -603 -981 -587 -947
rect -519 -981 -503 -947
rect -603 -997 -503 -981
rect -445 -947 -345 -909
rect -445 -981 -429 -947
rect -361 -981 -345 -947
rect -445 -997 -345 -981
rect -287 -947 -187 -909
rect -287 -981 -271 -947
rect -203 -981 -187 -947
rect -287 -997 -187 -981
rect -129 -947 -29 -909
rect -129 -981 -113 -947
rect -45 -981 -29 -947
rect -129 -997 -29 -981
rect 29 -947 129 -909
rect 29 -981 45 -947
rect 113 -981 129 -947
rect 29 -997 129 -981
rect 187 -947 287 -909
rect 187 -981 203 -947
rect 271 -981 287 -947
rect 187 -997 287 -981
rect 345 -947 445 -909
rect 345 -981 361 -947
rect 429 -981 445 -947
rect 345 -997 445 -981
rect 503 -947 603 -909
rect 503 -981 519 -947
rect 587 -981 603 -947
rect 503 -997 603 -981
rect 661 -947 761 -909
rect 661 -981 677 -947
rect 745 -981 761 -947
rect 661 -997 761 -981
rect 819 -947 919 -909
rect 819 -981 835 -947
rect 903 -981 919 -947
rect 819 -997 919 -981
rect 977 -947 1077 -909
rect 977 -981 993 -947
rect 1061 -981 1077 -947
rect 977 -997 1077 -981
rect 1135 -947 1235 -909
rect 1135 -981 1151 -947
rect 1219 -981 1235 -947
rect 1135 -997 1235 -981
rect 1293 -947 1393 -909
rect 1293 -981 1309 -947
rect 1377 -981 1393 -947
rect 1293 -997 1393 -981
rect 1451 -947 1551 -909
rect 1451 -981 1467 -947
rect 1535 -981 1551 -947
rect 1451 -997 1551 -981
rect 1609 -947 1709 -909
rect 1609 -981 1625 -947
rect 1693 -981 1709 -947
rect 1609 -997 1709 -981
rect 1767 -947 1867 -909
rect 1767 -981 1783 -947
rect 1851 -981 1867 -947
rect 1767 -997 1867 -981
rect 1925 -947 2025 -909
rect 1925 -981 1941 -947
rect 2009 -981 2025 -947
rect 1925 -997 2025 -981
rect 2083 -947 2183 -909
rect 2083 -981 2099 -947
rect 2167 -981 2183 -947
rect 2083 -997 2183 -981
rect 2241 -947 2341 -909
rect 2241 -981 2257 -947
rect 2325 -981 2341 -947
rect 2241 -997 2341 -981
rect 2399 -947 2499 -909
rect 2399 -981 2415 -947
rect 2483 -981 2499 -947
rect 2399 -997 2499 -981
rect -2499 -1055 -2399 -1039
rect -2499 -1089 -2483 -1055
rect -2415 -1089 -2399 -1055
rect -2499 -1127 -2399 -1089
rect -2341 -1055 -2241 -1039
rect -2341 -1089 -2325 -1055
rect -2257 -1089 -2241 -1055
rect -2341 -1127 -2241 -1089
rect -2183 -1055 -2083 -1039
rect -2183 -1089 -2167 -1055
rect -2099 -1089 -2083 -1055
rect -2183 -1127 -2083 -1089
rect -2025 -1055 -1925 -1039
rect -2025 -1089 -2009 -1055
rect -1941 -1089 -1925 -1055
rect -2025 -1127 -1925 -1089
rect -1867 -1055 -1767 -1039
rect -1867 -1089 -1851 -1055
rect -1783 -1089 -1767 -1055
rect -1867 -1127 -1767 -1089
rect -1709 -1055 -1609 -1039
rect -1709 -1089 -1693 -1055
rect -1625 -1089 -1609 -1055
rect -1709 -1127 -1609 -1089
rect -1551 -1055 -1451 -1039
rect -1551 -1089 -1535 -1055
rect -1467 -1089 -1451 -1055
rect -1551 -1127 -1451 -1089
rect -1393 -1055 -1293 -1039
rect -1393 -1089 -1377 -1055
rect -1309 -1089 -1293 -1055
rect -1393 -1127 -1293 -1089
rect -1235 -1055 -1135 -1039
rect -1235 -1089 -1219 -1055
rect -1151 -1089 -1135 -1055
rect -1235 -1127 -1135 -1089
rect -1077 -1055 -977 -1039
rect -1077 -1089 -1061 -1055
rect -993 -1089 -977 -1055
rect -1077 -1127 -977 -1089
rect -919 -1055 -819 -1039
rect -919 -1089 -903 -1055
rect -835 -1089 -819 -1055
rect -919 -1127 -819 -1089
rect -761 -1055 -661 -1039
rect -761 -1089 -745 -1055
rect -677 -1089 -661 -1055
rect -761 -1127 -661 -1089
rect -603 -1055 -503 -1039
rect -603 -1089 -587 -1055
rect -519 -1089 -503 -1055
rect -603 -1127 -503 -1089
rect -445 -1055 -345 -1039
rect -445 -1089 -429 -1055
rect -361 -1089 -345 -1055
rect -445 -1127 -345 -1089
rect -287 -1055 -187 -1039
rect -287 -1089 -271 -1055
rect -203 -1089 -187 -1055
rect -287 -1127 -187 -1089
rect -129 -1055 -29 -1039
rect -129 -1089 -113 -1055
rect -45 -1089 -29 -1055
rect -129 -1127 -29 -1089
rect 29 -1055 129 -1039
rect 29 -1089 45 -1055
rect 113 -1089 129 -1055
rect 29 -1127 129 -1089
rect 187 -1055 287 -1039
rect 187 -1089 203 -1055
rect 271 -1089 287 -1055
rect 187 -1127 287 -1089
rect 345 -1055 445 -1039
rect 345 -1089 361 -1055
rect 429 -1089 445 -1055
rect 345 -1127 445 -1089
rect 503 -1055 603 -1039
rect 503 -1089 519 -1055
rect 587 -1089 603 -1055
rect 503 -1127 603 -1089
rect 661 -1055 761 -1039
rect 661 -1089 677 -1055
rect 745 -1089 761 -1055
rect 661 -1127 761 -1089
rect 819 -1055 919 -1039
rect 819 -1089 835 -1055
rect 903 -1089 919 -1055
rect 819 -1127 919 -1089
rect 977 -1055 1077 -1039
rect 977 -1089 993 -1055
rect 1061 -1089 1077 -1055
rect 977 -1127 1077 -1089
rect 1135 -1055 1235 -1039
rect 1135 -1089 1151 -1055
rect 1219 -1089 1235 -1055
rect 1135 -1127 1235 -1089
rect 1293 -1055 1393 -1039
rect 1293 -1089 1309 -1055
rect 1377 -1089 1393 -1055
rect 1293 -1127 1393 -1089
rect 1451 -1055 1551 -1039
rect 1451 -1089 1467 -1055
rect 1535 -1089 1551 -1055
rect 1451 -1127 1551 -1089
rect 1609 -1055 1709 -1039
rect 1609 -1089 1625 -1055
rect 1693 -1089 1709 -1055
rect 1609 -1127 1709 -1089
rect 1767 -1055 1867 -1039
rect 1767 -1089 1783 -1055
rect 1851 -1089 1867 -1055
rect 1767 -1127 1867 -1089
rect 1925 -1055 2025 -1039
rect 1925 -1089 1941 -1055
rect 2009 -1089 2025 -1055
rect 1925 -1127 2025 -1089
rect 2083 -1055 2183 -1039
rect 2083 -1089 2099 -1055
rect 2167 -1089 2183 -1055
rect 2083 -1127 2183 -1089
rect 2241 -1055 2341 -1039
rect 2241 -1089 2257 -1055
rect 2325 -1089 2341 -1055
rect 2241 -1127 2341 -1089
rect 2399 -1055 2499 -1039
rect 2399 -1089 2415 -1055
rect 2483 -1089 2499 -1055
rect 2399 -1127 2499 -1089
rect -2499 -1965 -2399 -1927
rect -2499 -1999 -2483 -1965
rect -2415 -1999 -2399 -1965
rect -2499 -2015 -2399 -1999
rect -2341 -1965 -2241 -1927
rect -2341 -1999 -2325 -1965
rect -2257 -1999 -2241 -1965
rect -2341 -2015 -2241 -1999
rect -2183 -1965 -2083 -1927
rect -2183 -1999 -2167 -1965
rect -2099 -1999 -2083 -1965
rect -2183 -2015 -2083 -1999
rect -2025 -1965 -1925 -1927
rect -2025 -1999 -2009 -1965
rect -1941 -1999 -1925 -1965
rect -2025 -2015 -1925 -1999
rect -1867 -1965 -1767 -1927
rect -1867 -1999 -1851 -1965
rect -1783 -1999 -1767 -1965
rect -1867 -2015 -1767 -1999
rect -1709 -1965 -1609 -1927
rect -1709 -1999 -1693 -1965
rect -1625 -1999 -1609 -1965
rect -1709 -2015 -1609 -1999
rect -1551 -1965 -1451 -1927
rect -1551 -1999 -1535 -1965
rect -1467 -1999 -1451 -1965
rect -1551 -2015 -1451 -1999
rect -1393 -1965 -1293 -1927
rect -1393 -1999 -1377 -1965
rect -1309 -1999 -1293 -1965
rect -1393 -2015 -1293 -1999
rect -1235 -1965 -1135 -1927
rect -1235 -1999 -1219 -1965
rect -1151 -1999 -1135 -1965
rect -1235 -2015 -1135 -1999
rect -1077 -1965 -977 -1927
rect -1077 -1999 -1061 -1965
rect -993 -1999 -977 -1965
rect -1077 -2015 -977 -1999
rect -919 -1965 -819 -1927
rect -919 -1999 -903 -1965
rect -835 -1999 -819 -1965
rect -919 -2015 -819 -1999
rect -761 -1965 -661 -1927
rect -761 -1999 -745 -1965
rect -677 -1999 -661 -1965
rect -761 -2015 -661 -1999
rect -603 -1965 -503 -1927
rect -603 -1999 -587 -1965
rect -519 -1999 -503 -1965
rect -603 -2015 -503 -1999
rect -445 -1965 -345 -1927
rect -445 -1999 -429 -1965
rect -361 -1999 -345 -1965
rect -445 -2015 -345 -1999
rect -287 -1965 -187 -1927
rect -287 -1999 -271 -1965
rect -203 -1999 -187 -1965
rect -287 -2015 -187 -1999
rect -129 -1965 -29 -1927
rect -129 -1999 -113 -1965
rect -45 -1999 -29 -1965
rect -129 -2015 -29 -1999
rect 29 -1965 129 -1927
rect 29 -1999 45 -1965
rect 113 -1999 129 -1965
rect 29 -2015 129 -1999
rect 187 -1965 287 -1927
rect 187 -1999 203 -1965
rect 271 -1999 287 -1965
rect 187 -2015 287 -1999
rect 345 -1965 445 -1927
rect 345 -1999 361 -1965
rect 429 -1999 445 -1965
rect 345 -2015 445 -1999
rect 503 -1965 603 -1927
rect 503 -1999 519 -1965
rect 587 -1999 603 -1965
rect 503 -2015 603 -1999
rect 661 -1965 761 -1927
rect 661 -1999 677 -1965
rect 745 -1999 761 -1965
rect 661 -2015 761 -1999
rect 819 -1965 919 -1927
rect 819 -1999 835 -1965
rect 903 -1999 919 -1965
rect 819 -2015 919 -1999
rect 977 -1965 1077 -1927
rect 977 -1999 993 -1965
rect 1061 -1999 1077 -1965
rect 977 -2015 1077 -1999
rect 1135 -1965 1235 -1927
rect 1135 -1999 1151 -1965
rect 1219 -1999 1235 -1965
rect 1135 -2015 1235 -1999
rect 1293 -1965 1393 -1927
rect 1293 -1999 1309 -1965
rect 1377 -1999 1393 -1965
rect 1293 -2015 1393 -1999
rect 1451 -1965 1551 -1927
rect 1451 -1999 1467 -1965
rect 1535 -1999 1551 -1965
rect 1451 -2015 1551 -1999
rect 1609 -1965 1709 -1927
rect 1609 -1999 1625 -1965
rect 1693 -1999 1709 -1965
rect 1609 -2015 1709 -1999
rect 1767 -1965 1867 -1927
rect 1767 -1999 1783 -1965
rect 1851 -1999 1867 -1965
rect 1767 -2015 1867 -1999
rect 1925 -1965 2025 -1927
rect 1925 -1999 1941 -1965
rect 2009 -1999 2025 -1965
rect 1925 -2015 2025 -1999
rect 2083 -1965 2183 -1927
rect 2083 -1999 2099 -1965
rect 2167 -1999 2183 -1965
rect 2083 -2015 2183 -1999
rect 2241 -1965 2341 -1927
rect 2241 -1999 2257 -1965
rect 2325 -1999 2341 -1965
rect 2241 -2015 2341 -1999
rect 2399 -1965 2499 -1927
rect 2399 -1999 2415 -1965
rect 2483 -1999 2499 -1965
rect 2399 -2015 2499 -1999
<< polycont >>
rect -2483 1965 -2415 1999
rect -2325 1965 -2257 1999
rect -2167 1965 -2099 1999
rect -2009 1965 -1941 1999
rect -1851 1965 -1783 1999
rect -1693 1965 -1625 1999
rect -1535 1965 -1467 1999
rect -1377 1965 -1309 1999
rect -1219 1965 -1151 1999
rect -1061 1965 -993 1999
rect -903 1965 -835 1999
rect -745 1965 -677 1999
rect -587 1965 -519 1999
rect -429 1965 -361 1999
rect -271 1965 -203 1999
rect -113 1965 -45 1999
rect 45 1965 113 1999
rect 203 1965 271 1999
rect 361 1965 429 1999
rect 519 1965 587 1999
rect 677 1965 745 1999
rect 835 1965 903 1999
rect 993 1965 1061 1999
rect 1151 1965 1219 1999
rect 1309 1965 1377 1999
rect 1467 1965 1535 1999
rect 1625 1965 1693 1999
rect 1783 1965 1851 1999
rect 1941 1965 2009 1999
rect 2099 1965 2167 1999
rect 2257 1965 2325 1999
rect 2415 1965 2483 1999
rect -2483 1055 -2415 1089
rect -2325 1055 -2257 1089
rect -2167 1055 -2099 1089
rect -2009 1055 -1941 1089
rect -1851 1055 -1783 1089
rect -1693 1055 -1625 1089
rect -1535 1055 -1467 1089
rect -1377 1055 -1309 1089
rect -1219 1055 -1151 1089
rect -1061 1055 -993 1089
rect -903 1055 -835 1089
rect -745 1055 -677 1089
rect -587 1055 -519 1089
rect -429 1055 -361 1089
rect -271 1055 -203 1089
rect -113 1055 -45 1089
rect 45 1055 113 1089
rect 203 1055 271 1089
rect 361 1055 429 1089
rect 519 1055 587 1089
rect 677 1055 745 1089
rect 835 1055 903 1089
rect 993 1055 1061 1089
rect 1151 1055 1219 1089
rect 1309 1055 1377 1089
rect 1467 1055 1535 1089
rect 1625 1055 1693 1089
rect 1783 1055 1851 1089
rect 1941 1055 2009 1089
rect 2099 1055 2167 1089
rect 2257 1055 2325 1089
rect 2415 1055 2483 1089
rect -2483 947 -2415 981
rect -2325 947 -2257 981
rect -2167 947 -2099 981
rect -2009 947 -1941 981
rect -1851 947 -1783 981
rect -1693 947 -1625 981
rect -1535 947 -1467 981
rect -1377 947 -1309 981
rect -1219 947 -1151 981
rect -1061 947 -993 981
rect -903 947 -835 981
rect -745 947 -677 981
rect -587 947 -519 981
rect -429 947 -361 981
rect -271 947 -203 981
rect -113 947 -45 981
rect 45 947 113 981
rect 203 947 271 981
rect 361 947 429 981
rect 519 947 587 981
rect 677 947 745 981
rect 835 947 903 981
rect 993 947 1061 981
rect 1151 947 1219 981
rect 1309 947 1377 981
rect 1467 947 1535 981
rect 1625 947 1693 981
rect 1783 947 1851 981
rect 1941 947 2009 981
rect 2099 947 2167 981
rect 2257 947 2325 981
rect 2415 947 2483 981
rect -2483 37 -2415 71
rect -2325 37 -2257 71
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect 2257 37 2325 71
rect 2415 37 2483 71
rect -2483 -71 -2415 -37
rect -2325 -71 -2257 -37
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect 2257 -71 2325 -37
rect 2415 -71 2483 -37
rect -2483 -981 -2415 -947
rect -2325 -981 -2257 -947
rect -2167 -981 -2099 -947
rect -2009 -981 -1941 -947
rect -1851 -981 -1783 -947
rect -1693 -981 -1625 -947
rect -1535 -981 -1467 -947
rect -1377 -981 -1309 -947
rect -1219 -981 -1151 -947
rect -1061 -981 -993 -947
rect -903 -981 -835 -947
rect -745 -981 -677 -947
rect -587 -981 -519 -947
rect -429 -981 -361 -947
rect -271 -981 -203 -947
rect -113 -981 -45 -947
rect 45 -981 113 -947
rect 203 -981 271 -947
rect 361 -981 429 -947
rect 519 -981 587 -947
rect 677 -981 745 -947
rect 835 -981 903 -947
rect 993 -981 1061 -947
rect 1151 -981 1219 -947
rect 1309 -981 1377 -947
rect 1467 -981 1535 -947
rect 1625 -981 1693 -947
rect 1783 -981 1851 -947
rect 1941 -981 2009 -947
rect 2099 -981 2167 -947
rect 2257 -981 2325 -947
rect 2415 -981 2483 -947
rect -2483 -1089 -2415 -1055
rect -2325 -1089 -2257 -1055
rect -2167 -1089 -2099 -1055
rect -2009 -1089 -1941 -1055
rect -1851 -1089 -1783 -1055
rect -1693 -1089 -1625 -1055
rect -1535 -1089 -1467 -1055
rect -1377 -1089 -1309 -1055
rect -1219 -1089 -1151 -1055
rect -1061 -1089 -993 -1055
rect -903 -1089 -835 -1055
rect -745 -1089 -677 -1055
rect -587 -1089 -519 -1055
rect -429 -1089 -361 -1055
rect -271 -1089 -203 -1055
rect -113 -1089 -45 -1055
rect 45 -1089 113 -1055
rect 203 -1089 271 -1055
rect 361 -1089 429 -1055
rect 519 -1089 587 -1055
rect 677 -1089 745 -1055
rect 835 -1089 903 -1055
rect 993 -1089 1061 -1055
rect 1151 -1089 1219 -1055
rect 1309 -1089 1377 -1055
rect 1467 -1089 1535 -1055
rect 1625 -1089 1693 -1055
rect 1783 -1089 1851 -1055
rect 1941 -1089 2009 -1055
rect 2099 -1089 2167 -1055
rect 2257 -1089 2325 -1055
rect 2415 -1089 2483 -1055
rect -2483 -1999 -2415 -1965
rect -2325 -1999 -2257 -1965
rect -2167 -1999 -2099 -1965
rect -2009 -1999 -1941 -1965
rect -1851 -1999 -1783 -1965
rect -1693 -1999 -1625 -1965
rect -1535 -1999 -1467 -1965
rect -1377 -1999 -1309 -1965
rect -1219 -1999 -1151 -1965
rect -1061 -1999 -993 -1965
rect -903 -1999 -835 -1965
rect -745 -1999 -677 -1965
rect -587 -1999 -519 -1965
rect -429 -1999 -361 -1965
rect -271 -1999 -203 -1965
rect -113 -1999 -45 -1965
rect 45 -1999 113 -1965
rect 203 -1999 271 -1965
rect 361 -1999 429 -1965
rect 519 -1999 587 -1965
rect 677 -1999 745 -1965
rect 835 -1999 903 -1965
rect 993 -1999 1061 -1965
rect 1151 -1999 1219 -1965
rect 1309 -1999 1377 -1965
rect 1467 -1999 1535 -1965
rect 1625 -1999 1693 -1965
rect 1783 -1999 1851 -1965
rect 1941 -1999 2009 -1965
rect 2099 -1999 2167 -1965
rect 2257 -1999 2325 -1965
rect 2415 -1999 2483 -1965
<< locali >>
rect -2679 2103 -2583 2137
rect 2583 2103 2679 2137
rect -2679 2041 -2645 2103
rect 2645 2041 2679 2103
rect -2499 1965 -2483 1999
rect -2415 1965 -2399 1999
rect -2341 1965 -2325 1999
rect -2257 1965 -2241 1999
rect -2183 1965 -2167 1999
rect -2099 1965 -2083 1999
rect -2025 1965 -2009 1999
rect -1941 1965 -1925 1999
rect -1867 1965 -1851 1999
rect -1783 1965 -1767 1999
rect -1709 1965 -1693 1999
rect -1625 1965 -1609 1999
rect -1551 1965 -1535 1999
rect -1467 1965 -1451 1999
rect -1393 1965 -1377 1999
rect -1309 1965 -1293 1999
rect -1235 1965 -1219 1999
rect -1151 1965 -1135 1999
rect -1077 1965 -1061 1999
rect -993 1965 -977 1999
rect -919 1965 -903 1999
rect -835 1965 -819 1999
rect -761 1965 -745 1999
rect -677 1965 -661 1999
rect -603 1965 -587 1999
rect -519 1965 -503 1999
rect -445 1965 -429 1999
rect -361 1965 -345 1999
rect -287 1965 -271 1999
rect -203 1965 -187 1999
rect -129 1965 -113 1999
rect -45 1965 -29 1999
rect 29 1965 45 1999
rect 113 1965 129 1999
rect 187 1965 203 1999
rect 271 1965 287 1999
rect 345 1965 361 1999
rect 429 1965 445 1999
rect 503 1965 519 1999
rect 587 1965 603 1999
rect 661 1965 677 1999
rect 745 1965 761 1999
rect 819 1965 835 1999
rect 903 1965 919 1999
rect 977 1965 993 1999
rect 1061 1965 1077 1999
rect 1135 1965 1151 1999
rect 1219 1965 1235 1999
rect 1293 1965 1309 1999
rect 1377 1965 1393 1999
rect 1451 1965 1467 1999
rect 1535 1965 1551 1999
rect 1609 1965 1625 1999
rect 1693 1965 1709 1999
rect 1767 1965 1783 1999
rect 1851 1965 1867 1999
rect 1925 1965 1941 1999
rect 2009 1965 2025 1999
rect 2083 1965 2099 1999
rect 2167 1965 2183 1999
rect 2241 1965 2257 1999
rect 2325 1965 2341 1999
rect 2399 1965 2415 1999
rect 2483 1965 2499 1999
rect -2545 1915 -2511 1931
rect -2545 1123 -2511 1139
rect -2387 1915 -2353 1931
rect -2387 1123 -2353 1139
rect -2229 1915 -2195 1931
rect -2229 1123 -2195 1139
rect -2071 1915 -2037 1931
rect -2071 1123 -2037 1139
rect -1913 1915 -1879 1931
rect -1913 1123 -1879 1139
rect -1755 1915 -1721 1931
rect -1755 1123 -1721 1139
rect -1597 1915 -1563 1931
rect -1597 1123 -1563 1139
rect -1439 1915 -1405 1931
rect -1439 1123 -1405 1139
rect -1281 1915 -1247 1931
rect -1281 1123 -1247 1139
rect -1123 1915 -1089 1931
rect -1123 1123 -1089 1139
rect -965 1915 -931 1931
rect -965 1123 -931 1139
rect -807 1915 -773 1931
rect -807 1123 -773 1139
rect -649 1915 -615 1931
rect -649 1123 -615 1139
rect -491 1915 -457 1931
rect -491 1123 -457 1139
rect -333 1915 -299 1931
rect -333 1123 -299 1139
rect -175 1915 -141 1931
rect -175 1123 -141 1139
rect -17 1915 17 1931
rect -17 1123 17 1139
rect 141 1915 175 1931
rect 141 1123 175 1139
rect 299 1915 333 1931
rect 299 1123 333 1139
rect 457 1915 491 1931
rect 457 1123 491 1139
rect 615 1915 649 1931
rect 615 1123 649 1139
rect 773 1915 807 1931
rect 773 1123 807 1139
rect 931 1915 965 1931
rect 931 1123 965 1139
rect 1089 1915 1123 1931
rect 1089 1123 1123 1139
rect 1247 1915 1281 1931
rect 1247 1123 1281 1139
rect 1405 1915 1439 1931
rect 1405 1123 1439 1139
rect 1563 1915 1597 1931
rect 1563 1123 1597 1139
rect 1721 1915 1755 1931
rect 1721 1123 1755 1139
rect 1879 1915 1913 1931
rect 1879 1123 1913 1139
rect 2037 1915 2071 1931
rect 2037 1123 2071 1139
rect 2195 1915 2229 1931
rect 2195 1123 2229 1139
rect 2353 1915 2387 1931
rect 2353 1123 2387 1139
rect 2511 1915 2545 1931
rect 2511 1123 2545 1139
rect -2499 1055 -2483 1089
rect -2415 1055 -2399 1089
rect -2341 1055 -2325 1089
rect -2257 1055 -2241 1089
rect -2183 1055 -2167 1089
rect -2099 1055 -2083 1089
rect -2025 1055 -2009 1089
rect -1941 1055 -1925 1089
rect -1867 1055 -1851 1089
rect -1783 1055 -1767 1089
rect -1709 1055 -1693 1089
rect -1625 1055 -1609 1089
rect -1551 1055 -1535 1089
rect -1467 1055 -1451 1089
rect -1393 1055 -1377 1089
rect -1309 1055 -1293 1089
rect -1235 1055 -1219 1089
rect -1151 1055 -1135 1089
rect -1077 1055 -1061 1089
rect -993 1055 -977 1089
rect -919 1055 -903 1089
rect -835 1055 -819 1089
rect -761 1055 -745 1089
rect -677 1055 -661 1089
rect -603 1055 -587 1089
rect -519 1055 -503 1089
rect -445 1055 -429 1089
rect -361 1055 -345 1089
rect -287 1055 -271 1089
rect -203 1055 -187 1089
rect -129 1055 -113 1089
rect -45 1055 -29 1089
rect 29 1055 45 1089
rect 113 1055 129 1089
rect 187 1055 203 1089
rect 271 1055 287 1089
rect 345 1055 361 1089
rect 429 1055 445 1089
rect 503 1055 519 1089
rect 587 1055 603 1089
rect 661 1055 677 1089
rect 745 1055 761 1089
rect 819 1055 835 1089
rect 903 1055 919 1089
rect 977 1055 993 1089
rect 1061 1055 1077 1089
rect 1135 1055 1151 1089
rect 1219 1055 1235 1089
rect 1293 1055 1309 1089
rect 1377 1055 1393 1089
rect 1451 1055 1467 1089
rect 1535 1055 1551 1089
rect 1609 1055 1625 1089
rect 1693 1055 1709 1089
rect 1767 1055 1783 1089
rect 1851 1055 1867 1089
rect 1925 1055 1941 1089
rect 2009 1055 2025 1089
rect 2083 1055 2099 1089
rect 2167 1055 2183 1089
rect 2241 1055 2257 1089
rect 2325 1055 2341 1089
rect 2399 1055 2415 1089
rect 2483 1055 2499 1089
rect -2499 947 -2483 981
rect -2415 947 -2399 981
rect -2341 947 -2325 981
rect -2257 947 -2241 981
rect -2183 947 -2167 981
rect -2099 947 -2083 981
rect -2025 947 -2009 981
rect -1941 947 -1925 981
rect -1867 947 -1851 981
rect -1783 947 -1767 981
rect -1709 947 -1693 981
rect -1625 947 -1609 981
rect -1551 947 -1535 981
rect -1467 947 -1451 981
rect -1393 947 -1377 981
rect -1309 947 -1293 981
rect -1235 947 -1219 981
rect -1151 947 -1135 981
rect -1077 947 -1061 981
rect -993 947 -977 981
rect -919 947 -903 981
rect -835 947 -819 981
rect -761 947 -745 981
rect -677 947 -661 981
rect -603 947 -587 981
rect -519 947 -503 981
rect -445 947 -429 981
rect -361 947 -345 981
rect -287 947 -271 981
rect -203 947 -187 981
rect -129 947 -113 981
rect -45 947 -29 981
rect 29 947 45 981
rect 113 947 129 981
rect 187 947 203 981
rect 271 947 287 981
rect 345 947 361 981
rect 429 947 445 981
rect 503 947 519 981
rect 587 947 603 981
rect 661 947 677 981
rect 745 947 761 981
rect 819 947 835 981
rect 903 947 919 981
rect 977 947 993 981
rect 1061 947 1077 981
rect 1135 947 1151 981
rect 1219 947 1235 981
rect 1293 947 1309 981
rect 1377 947 1393 981
rect 1451 947 1467 981
rect 1535 947 1551 981
rect 1609 947 1625 981
rect 1693 947 1709 981
rect 1767 947 1783 981
rect 1851 947 1867 981
rect 1925 947 1941 981
rect 2009 947 2025 981
rect 2083 947 2099 981
rect 2167 947 2183 981
rect 2241 947 2257 981
rect 2325 947 2341 981
rect 2399 947 2415 981
rect 2483 947 2499 981
rect -2545 897 -2511 913
rect -2545 105 -2511 121
rect -2387 897 -2353 913
rect -2387 105 -2353 121
rect -2229 897 -2195 913
rect -2229 105 -2195 121
rect -2071 897 -2037 913
rect -2071 105 -2037 121
rect -1913 897 -1879 913
rect -1913 105 -1879 121
rect -1755 897 -1721 913
rect -1755 105 -1721 121
rect -1597 897 -1563 913
rect -1597 105 -1563 121
rect -1439 897 -1405 913
rect -1439 105 -1405 121
rect -1281 897 -1247 913
rect -1281 105 -1247 121
rect -1123 897 -1089 913
rect -1123 105 -1089 121
rect -965 897 -931 913
rect -965 105 -931 121
rect -807 897 -773 913
rect -807 105 -773 121
rect -649 897 -615 913
rect -649 105 -615 121
rect -491 897 -457 913
rect -491 105 -457 121
rect -333 897 -299 913
rect -333 105 -299 121
rect -175 897 -141 913
rect -175 105 -141 121
rect -17 897 17 913
rect -17 105 17 121
rect 141 897 175 913
rect 141 105 175 121
rect 299 897 333 913
rect 299 105 333 121
rect 457 897 491 913
rect 457 105 491 121
rect 615 897 649 913
rect 615 105 649 121
rect 773 897 807 913
rect 773 105 807 121
rect 931 897 965 913
rect 931 105 965 121
rect 1089 897 1123 913
rect 1089 105 1123 121
rect 1247 897 1281 913
rect 1247 105 1281 121
rect 1405 897 1439 913
rect 1405 105 1439 121
rect 1563 897 1597 913
rect 1563 105 1597 121
rect 1721 897 1755 913
rect 1721 105 1755 121
rect 1879 897 1913 913
rect 1879 105 1913 121
rect 2037 897 2071 913
rect 2037 105 2071 121
rect 2195 897 2229 913
rect 2195 105 2229 121
rect 2353 897 2387 913
rect 2353 105 2387 121
rect 2511 897 2545 913
rect 2511 105 2545 121
rect -2499 37 -2483 71
rect -2415 37 -2399 71
rect -2341 37 -2325 71
rect -2257 37 -2241 71
rect -2183 37 -2167 71
rect -2099 37 -2083 71
rect -2025 37 -2009 71
rect -1941 37 -1925 71
rect -1867 37 -1851 71
rect -1783 37 -1767 71
rect -1709 37 -1693 71
rect -1625 37 -1609 71
rect -1551 37 -1535 71
rect -1467 37 -1451 71
rect -1393 37 -1377 71
rect -1309 37 -1293 71
rect -1235 37 -1219 71
rect -1151 37 -1135 71
rect -1077 37 -1061 71
rect -993 37 -977 71
rect -919 37 -903 71
rect -835 37 -819 71
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect 819 37 835 71
rect 903 37 919 71
rect 977 37 993 71
rect 1061 37 1077 71
rect 1135 37 1151 71
rect 1219 37 1235 71
rect 1293 37 1309 71
rect 1377 37 1393 71
rect 1451 37 1467 71
rect 1535 37 1551 71
rect 1609 37 1625 71
rect 1693 37 1709 71
rect 1767 37 1783 71
rect 1851 37 1867 71
rect 1925 37 1941 71
rect 2009 37 2025 71
rect 2083 37 2099 71
rect 2167 37 2183 71
rect 2241 37 2257 71
rect 2325 37 2341 71
rect 2399 37 2415 71
rect 2483 37 2499 71
rect -2499 -71 -2483 -37
rect -2415 -71 -2399 -37
rect -2341 -71 -2325 -37
rect -2257 -71 -2241 -37
rect -2183 -71 -2167 -37
rect -2099 -71 -2083 -37
rect -2025 -71 -2009 -37
rect -1941 -71 -1925 -37
rect -1867 -71 -1851 -37
rect -1783 -71 -1767 -37
rect -1709 -71 -1693 -37
rect -1625 -71 -1609 -37
rect -1551 -71 -1535 -37
rect -1467 -71 -1451 -37
rect -1393 -71 -1377 -37
rect -1309 -71 -1293 -37
rect -1235 -71 -1219 -37
rect -1151 -71 -1135 -37
rect -1077 -71 -1061 -37
rect -993 -71 -977 -37
rect -919 -71 -903 -37
rect -835 -71 -819 -37
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 819 -71 835 -37
rect 903 -71 919 -37
rect 977 -71 993 -37
rect 1061 -71 1077 -37
rect 1135 -71 1151 -37
rect 1219 -71 1235 -37
rect 1293 -71 1309 -37
rect 1377 -71 1393 -37
rect 1451 -71 1467 -37
rect 1535 -71 1551 -37
rect 1609 -71 1625 -37
rect 1693 -71 1709 -37
rect 1767 -71 1783 -37
rect 1851 -71 1867 -37
rect 1925 -71 1941 -37
rect 2009 -71 2025 -37
rect 2083 -71 2099 -37
rect 2167 -71 2183 -37
rect 2241 -71 2257 -37
rect 2325 -71 2341 -37
rect 2399 -71 2415 -37
rect 2483 -71 2499 -37
rect -2545 -121 -2511 -105
rect -2545 -913 -2511 -897
rect -2387 -121 -2353 -105
rect -2387 -913 -2353 -897
rect -2229 -121 -2195 -105
rect -2229 -913 -2195 -897
rect -2071 -121 -2037 -105
rect -2071 -913 -2037 -897
rect -1913 -121 -1879 -105
rect -1913 -913 -1879 -897
rect -1755 -121 -1721 -105
rect -1755 -913 -1721 -897
rect -1597 -121 -1563 -105
rect -1597 -913 -1563 -897
rect -1439 -121 -1405 -105
rect -1439 -913 -1405 -897
rect -1281 -121 -1247 -105
rect -1281 -913 -1247 -897
rect -1123 -121 -1089 -105
rect -1123 -913 -1089 -897
rect -965 -121 -931 -105
rect -965 -913 -931 -897
rect -807 -121 -773 -105
rect -807 -913 -773 -897
rect -649 -121 -615 -105
rect -649 -913 -615 -897
rect -491 -121 -457 -105
rect -491 -913 -457 -897
rect -333 -121 -299 -105
rect -333 -913 -299 -897
rect -175 -121 -141 -105
rect -175 -913 -141 -897
rect -17 -121 17 -105
rect -17 -913 17 -897
rect 141 -121 175 -105
rect 141 -913 175 -897
rect 299 -121 333 -105
rect 299 -913 333 -897
rect 457 -121 491 -105
rect 457 -913 491 -897
rect 615 -121 649 -105
rect 615 -913 649 -897
rect 773 -121 807 -105
rect 773 -913 807 -897
rect 931 -121 965 -105
rect 931 -913 965 -897
rect 1089 -121 1123 -105
rect 1089 -913 1123 -897
rect 1247 -121 1281 -105
rect 1247 -913 1281 -897
rect 1405 -121 1439 -105
rect 1405 -913 1439 -897
rect 1563 -121 1597 -105
rect 1563 -913 1597 -897
rect 1721 -121 1755 -105
rect 1721 -913 1755 -897
rect 1879 -121 1913 -105
rect 1879 -913 1913 -897
rect 2037 -121 2071 -105
rect 2037 -913 2071 -897
rect 2195 -121 2229 -105
rect 2195 -913 2229 -897
rect 2353 -121 2387 -105
rect 2353 -913 2387 -897
rect 2511 -121 2545 -105
rect 2511 -913 2545 -897
rect -2499 -981 -2483 -947
rect -2415 -981 -2399 -947
rect -2341 -981 -2325 -947
rect -2257 -981 -2241 -947
rect -2183 -981 -2167 -947
rect -2099 -981 -2083 -947
rect -2025 -981 -2009 -947
rect -1941 -981 -1925 -947
rect -1867 -981 -1851 -947
rect -1783 -981 -1767 -947
rect -1709 -981 -1693 -947
rect -1625 -981 -1609 -947
rect -1551 -981 -1535 -947
rect -1467 -981 -1451 -947
rect -1393 -981 -1377 -947
rect -1309 -981 -1293 -947
rect -1235 -981 -1219 -947
rect -1151 -981 -1135 -947
rect -1077 -981 -1061 -947
rect -993 -981 -977 -947
rect -919 -981 -903 -947
rect -835 -981 -819 -947
rect -761 -981 -745 -947
rect -677 -981 -661 -947
rect -603 -981 -587 -947
rect -519 -981 -503 -947
rect -445 -981 -429 -947
rect -361 -981 -345 -947
rect -287 -981 -271 -947
rect -203 -981 -187 -947
rect -129 -981 -113 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 113 -981 129 -947
rect 187 -981 203 -947
rect 271 -981 287 -947
rect 345 -981 361 -947
rect 429 -981 445 -947
rect 503 -981 519 -947
rect 587 -981 603 -947
rect 661 -981 677 -947
rect 745 -981 761 -947
rect 819 -981 835 -947
rect 903 -981 919 -947
rect 977 -981 993 -947
rect 1061 -981 1077 -947
rect 1135 -981 1151 -947
rect 1219 -981 1235 -947
rect 1293 -981 1309 -947
rect 1377 -981 1393 -947
rect 1451 -981 1467 -947
rect 1535 -981 1551 -947
rect 1609 -981 1625 -947
rect 1693 -981 1709 -947
rect 1767 -981 1783 -947
rect 1851 -981 1867 -947
rect 1925 -981 1941 -947
rect 2009 -981 2025 -947
rect 2083 -981 2099 -947
rect 2167 -981 2183 -947
rect 2241 -981 2257 -947
rect 2325 -981 2341 -947
rect 2399 -981 2415 -947
rect 2483 -981 2499 -947
rect -2499 -1089 -2483 -1055
rect -2415 -1089 -2399 -1055
rect -2341 -1089 -2325 -1055
rect -2257 -1089 -2241 -1055
rect -2183 -1089 -2167 -1055
rect -2099 -1089 -2083 -1055
rect -2025 -1089 -2009 -1055
rect -1941 -1089 -1925 -1055
rect -1867 -1089 -1851 -1055
rect -1783 -1089 -1767 -1055
rect -1709 -1089 -1693 -1055
rect -1625 -1089 -1609 -1055
rect -1551 -1089 -1535 -1055
rect -1467 -1089 -1451 -1055
rect -1393 -1089 -1377 -1055
rect -1309 -1089 -1293 -1055
rect -1235 -1089 -1219 -1055
rect -1151 -1089 -1135 -1055
rect -1077 -1089 -1061 -1055
rect -993 -1089 -977 -1055
rect -919 -1089 -903 -1055
rect -835 -1089 -819 -1055
rect -761 -1089 -745 -1055
rect -677 -1089 -661 -1055
rect -603 -1089 -587 -1055
rect -519 -1089 -503 -1055
rect -445 -1089 -429 -1055
rect -361 -1089 -345 -1055
rect -287 -1089 -271 -1055
rect -203 -1089 -187 -1055
rect -129 -1089 -113 -1055
rect -45 -1089 -29 -1055
rect 29 -1089 45 -1055
rect 113 -1089 129 -1055
rect 187 -1089 203 -1055
rect 271 -1089 287 -1055
rect 345 -1089 361 -1055
rect 429 -1089 445 -1055
rect 503 -1089 519 -1055
rect 587 -1089 603 -1055
rect 661 -1089 677 -1055
rect 745 -1089 761 -1055
rect 819 -1089 835 -1055
rect 903 -1089 919 -1055
rect 977 -1089 993 -1055
rect 1061 -1089 1077 -1055
rect 1135 -1089 1151 -1055
rect 1219 -1089 1235 -1055
rect 1293 -1089 1309 -1055
rect 1377 -1089 1393 -1055
rect 1451 -1089 1467 -1055
rect 1535 -1089 1551 -1055
rect 1609 -1089 1625 -1055
rect 1693 -1089 1709 -1055
rect 1767 -1089 1783 -1055
rect 1851 -1089 1867 -1055
rect 1925 -1089 1941 -1055
rect 2009 -1089 2025 -1055
rect 2083 -1089 2099 -1055
rect 2167 -1089 2183 -1055
rect 2241 -1089 2257 -1055
rect 2325 -1089 2341 -1055
rect 2399 -1089 2415 -1055
rect 2483 -1089 2499 -1055
rect -2545 -1139 -2511 -1123
rect -2545 -1931 -2511 -1915
rect -2387 -1139 -2353 -1123
rect -2387 -1931 -2353 -1915
rect -2229 -1139 -2195 -1123
rect -2229 -1931 -2195 -1915
rect -2071 -1139 -2037 -1123
rect -2071 -1931 -2037 -1915
rect -1913 -1139 -1879 -1123
rect -1913 -1931 -1879 -1915
rect -1755 -1139 -1721 -1123
rect -1755 -1931 -1721 -1915
rect -1597 -1139 -1563 -1123
rect -1597 -1931 -1563 -1915
rect -1439 -1139 -1405 -1123
rect -1439 -1931 -1405 -1915
rect -1281 -1139 -1247 -1123
rect -1281 -1931 -1247 -1915
rect -1123 -1139 -1089 -1123
rect -1123 -1931 -1089 -1915
rect -965 -1139 -931 -1123
rect -965 -1931 -931 -1915
rect -807 -1139 -773 -1123
rect -807 -1931 -773 -1915
rect -649 -1139 -615 -1123
rect -649 -1931 -615 -1915
rect -491 -1139 -457 -1123
rect -491 -1931 -457 -1915
rect -333 -1139 -299 -1123
rect -333 -1931 -299 -1915
rect -175 -1139 -141 -1123
rect -175 -1931 -141 -1915
rect -17 -1139 17 -1123
rect -17 -1931 17 -1915
rect 141 -1139 175 -1123
rect 141 -1931 175 -1915
rect 299 -1139 333 -1123
rect 299 -1931 333 -1915
rect 457 -1139 491 -1123
rect 457 -1931 491 -1915
rect 615 -1139 649 -1123
rect 615 -1931 649 -1915
rect 773 -1139 807 -1123
rect 773 -1931 807 -1915
rect 931 -1139 965 -1123
rect 931 -1931 965 -1915
rect 1089 -1139 1123 -1123
rect 1089 -1931 1123 -1915
rect 1247 -1139 1281 -1123
rect 1247 -1931 1281 -1915
rect 1405 -1139 1439 -1123
rect 1405 -1931 1439 -1915
rect 1563 -1139 1597 -1123
rect 1563 -1931 1597 -1915
rect 1721 -1139 1755 -1123
rect 1721 -1931 1755 -1915
rect 1879 -1139 1913 -1123
rect 1879 -1931 1913 -1915
rect 2037 -1139 2071 -1123
rect 2037 -1931 2071 -1915
rect 2195 -1139 2229 -1123
rect 2195 -1931 2229 -1915
rect 2353 -1139 2387 -1123
rect 2353 -1931 2387 -1915
rect 2511 -1139 2545 -1123
rect 2511 -1931 2545 -1915
rect -2499 -1999 -2483 -1965
rect -2415 -1999 -2399 -1965
rect -2341 -1999 -2325 -1965
rect -2257 -1999 -2241 -1965
rect -2183 -1999 -2167 -1965
rect -2099 -1999 -2083 -1965
rect -2025 -1999 -2009 -1965
rect -1941 -1999 -1925 -1965
rect -1867 -1999 -1851 -1965
rect -1783 -1999 -1767 -1965
rect -1709 -1999 -1693 -1965
rect -1625 -1999 -1609 -1965
rect -1551 -1999 -1535 -1965
rect -1467 -1999 -1451 -1965
rect -1393 -1999 -1377 -1965
rect -1309 -1999 -1293 -1965
rect -1235 -1999 -1219 -1965
rect -1151 -1999 -1135 -1965
rect -1077 -1999 -1061 -1965
rect -993 -1999 -977 -1965
rect -919 -1999 -903 -1965
rect -835 -1999 -819 -1965
rect -761 -1999 -745 -1965
rect -677 -1999 -661 -1965
rect -603 -1999 -587 -1965
rect -519 -1999 -503 -1965
rect -445 -1999 -429 -1965
rect -361 -1999 -345 -1965
rect -287 -1999 -271 -1965
rect -203 -1999 -187 -1965
rect -129 -1999 -113 -1965
rect -45 -1999 -29 -1965
rect 29 -1999 45 -1965
rect 113 -1999 129 -1965
rect 187 -1999 203 -1965
rect 271 -1999 287 -1965
rect 345 -1999 361 -1965
rect 429 -1999 445 -1965
rect 503 -1999 519 -1965
rect 587 -1999 603 -1965
rect 661 -1999 677 -1965
rect 745 -1999 761 -1965
rect 819 -1999 835 -1965
rect 903 -1999 919 -1965
rect 977 -1999 993 -1965
rect 1061 -1999 1077 -1965
rect 1135 -1999 1151 -1965
rect 1219 -1999 1235 -1965
rect 1293 -1999 1309 -1965
rect 1377 -1999 1393 -1965
rect 1451 -1999 1467 -1965
rect 1535 -1999 1551 -1965
rect 1609 -1999 1625 -1965
rect 1693 -1999 1709 -1965
rect 1767 -1999 1783 -1965
rect 1851 -1999 1867 -1965
rect 1925 -1999 1941 -1965
rect 2009 -1999 2025 -1965
rect 2083 -1999 2099 -1965
rect 2167 -1999 2183 -1965
rect 2241 -1999 2257 -1965
rect 2325 -1999 2341 -1965
rect 2399 -1999 2415 -1965
rect 2483 -1999 2499 -1965
rect -2679 -2103 -2645 -2041
rect 2645 -2103 2679 -2041
rect -2679 -2137 -2583 -2103
rect 2583 -2137 2679 -2103
<< viali >>
rect -2483 1965 -2415 1999
rect -2325 1965 -2257 1999
rect -2167 1965 -2099 1999
rect -2009 1965 -1941 1999
rect -1851 1965 -1783 1999
rect -1693 1965 -1625 1999
rect -1535 1965 -1467 1999
rect -1377 1965 -1309 1999
rect -1219 1965 -1151 1999
rect -1061 1965 -993 1999
rect -903 1965 -835 1999
rect -745 1965 -677 1999
rect -587 1965 -519 1999
rect -429 1965 -361 1999
rect -271 1965 -203 1999
rect -113 1965 -45 1999
rect 45 1965 113 1999
rect 203 1965 271 1999
rect 361 1965 429 1999
rect 519 1965 587 1999
rect 677 1965 745 1999
rect 835 1965 903 1999
rect 993 1965 1061 1999
rect 1151 1965 1219 1999
rect 1309 1965 1377 1999
rect 1467 1965 1535 1999
rect 1625 1965 1693 1999
rect 1783 1965 1851 1999
rect 1941 1965 2009 1999
rect 2099 1965 2167 1999
rect 2257 1965 2325 1999
rect 2415 1965 2483 1999
rect -2545 1139 -2511 1915
rect -2387 1139 -2353 1915
rect -2229 1139 -2195 1915
rect -2071 1139 -2037 1915
rect -1913 1139 -1879 1915
rect -1755 1139 -1721 1915
rect -1597 1139 -1563 1915
rect -1439 1139 -1405 1915
rect -1281 1139 -1247 1915
rect -1123 1139 -1089 1915
rect -965 1139 -931 1915
rect -807 1139 -773 1915
rect -649 1139 -615 1915
rect -491 1139 -457 1915
rect -333 1139 -299 1915
rect -175 1139 -141 1915
rect -17 1139 17 1915
rect 141 1139 175 1915
rect 299 1139 333 1915
rect 457 1139 491 1915
rect 615 1139 649 1915
rect 773 1139 807 1915
rect 931 1139 965 1915
rect 1089 1139 1123 1915
rect 1247 1139 1281 1915
rect 1405 1139 1439 1915
rect 1563 1139 1597 1915
rect 1721 1139 1755 1915
rect 1879 1139 1913 1915
rect 2037 1139 2071 1915
rect 2195 1139 2229 1915
rect 2353 1139 2387 1915
rect 2511 1139 2545 1915
rect -2483 1055 -2415 1089
rect -2325 1055 -2257 1089
rect -2167 1055 -2099 1089
rect -2009 1055 -1941 1089
rect -1851 1055 -1783 1089
rect -1693 1055 -1625 1089
rect -1535 1055 -1467 1089
rect -1377 1055 -1309 1089
rect -1219 1055 -1151 1089
rect -1061 1055 -993 1089
rect -903 1055 -835 1089
rect -745 1055 -677 1089
rect -587 1055 -519 1089
rect -429 1055 -361 1089
rect -271 1055 -203 1089
rect -113 1055 -45 1089
rect 45 1055 113 1089
rect 203 1055 271 1089
rect 361 1055 429 1089
rect 519 1055 587 1089
rect 677 1055 745 1089
rect 835 1055 903 1089
rect 993 1055 1061 1089
rect 1151 1055 1219 1089
rect 1309 1055 1377 1089
rect 1467 1055 1535 1089
rect 1625 1055 1693 1089
rect 1783 1055 1851 1089
rect 1941 1055 2009 1089
rect 2099 1055 2167 1089
rect 2257 1055 2325 1089
rect 2415 1055 2483 1089
rect -2483 947 -2415 981
rect -2325 947 -2257 981
rect -2167 947 -2099 981
rect -2009 947 -1941 981
rect -1851 947 -1783 981
rect -1693 947 -1625 981
rect -1535 947 -1467 981
rect -1377 947 -1309 981
rect -1219 947 -1151 981
rect -1061 947 -993 981
rect -903 947 -835 981
rect -745 947 -677 981
rect -587 947 -519 981
rect -429 947 -361 981
rect -271 947 -203 981
rect -113 947 -45 981
rect 45 947 113 981
rect 203 947 271 981
rect 361 947 429 981
rect 519 947 587 981
rect 677 947 745 981
rect 835 947 903 981
rect 993 947 1061 981
rect 1151 947 1219 981
rect 1309 947 1377 981
rect 1467 947 1535 981
rect 1625 947 1693 981
rect 1783 947 1851 981
rect 1941 947 2009 981
rect 2099 947 2167 981
rect 2257 947 2325 981
rect 2415 947 2483 981
rect -2545 121 -2511 897
rect -2387 121 -2353 897
rect -2229 121 -2195 897
rect -2071 121 -2037 897
rect -1913 121 -1879 897
rect -1755 121 -1721 897
rect -1597 121 -1563 897
rect -1439 121 -1405 897
rect -1281 121 -1247 897
rect -1123 121 -1089 897
rect -965 121 -931 897
rect -807 121 -773 897
rect -649 121 -615 897
rect -491 121 -457 897
rect -333 121 -299 897
rect -175 121 -141 897
rect -17 121 17 897
rect 141 121 175 897
rect 299 121 333 897
rect 457 121 491 897
rect 615 121 649 897
rect 773 121 807 897
rect 931 121 965 897
rect 1089 121 1123 897
rect 1247 121 1281 897
rect 1405 121 1439 897
rect 1563 121 1597 897
rect 1721 121 1755 897
rect 1879 121 1913 897
rect 2037 121 2071 897
rect 2195 121 2229 897
rect 2353 121 2387 897
rect 2511 121 2545 897
rect -2483 37 -2415 71
rect -2325 37 -2257 71
rect -2167 37 -2099 71
rect -2009 37 -1941 71
rect -1851 37 -1783 71
rect -1693 37 -1625 71
rect -1535 37 -1467 71
rect -1377 37 -1309 71
rect -1219 37 -1151 71
rect -1061 37 -993 71
rect -903 37 -835 71
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect 835 37 903 71
rect 993 37 1061 71
rect 1151 37 1219 71
rect 1309 37 1377 71
rect 1467 37 1535 71
rect 1625 37 1693 71
rect 1783 37 1851 71
rect 1941 37 2009 71
rect 2099 37 2167 71
rect 2257 37 2325 71
rect 2415 37 2483 71
rect -2483 -71 -2415 -37
rect -2325 -71 -2257 -37
rect -2167 -71 -2099 -37
rect -2009 -71 -1941 -37
rect -1851 -71 -1783 -37
rect -1693 -71 -1625 -37
rect -1535 -71 -1467 -37
rect -1377 -71 -1309 -37
rect -1219 -71 -1151 -37
rect -1061 -71 -993 -37
rect -903 -71 -835 -37
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect 835 -71 903 -37
rect 993 -71 1061 -37
rect 1151 -71 1219 -37
rect 1309 -71 1377 -37
rect 1467 -71 1535 -37
rect 1625 -71 1693 -37
rect 1783 -71 1851 -37
rect 1941 -71 2009 -37
rect 2099 -71 2167 -37
rect 2257 -71 2325 -37
rect 2415 -71 2483 -37
rect -2545 -897 -2511 -121
rect -2387 -897 -2353 -121
rect -2229 -897 -2195 -121
rect -2071 -897 -2037 -121
rect -1913 -897 -1879 -121
rect -1755 -897 -1721 -121
rect -1597 -897 -1563 -121
rect -1439 -897 -1405 -121
rect -1281 -897 -1247 -121
rect -1123 -897 -1089 -121
rect -965 -897 -931 -121
rect -807 -897 -773 -121
rect -649 -897 -615 -121
rect -491 -897 -457 -121
rect -333 -897 -299 -121
rect -175 -897 -141 -121
rect -17 -897 17 -121
rect 141 -897 175 -121
rect 299 -897 333 -121
rect 457 -897 491 -121
rect 615 -897 649 -121
rect 773 -897 807 -121
rect 931 -897 965 -121
rect 1089 -897 1123 -121
rect 1247 -897 1281 -121
rect 1405 -897 1439 -121
rect 1563 -897 1597 -121
rect 1721 -897 1755 -121
rect 1879 -897 1913 -121
rect 2037 -897 2071 -121
rect 2195 -897 2229 -121
rect 2353 -897 2387 -121
rect 2511 -897 2545 -121
rect -2483 -981 -2415 -947
rect -2325 -981 -2257 -947
rect -2167 -981 -2099 -947
rect -2009 -981 -1941 -947
rect -1851 -981 -1783 -947
rect -1693 -981 -1625 -947
rect -1535 -981 -1467 -947
rect -1377 -981 -1309 -947
rect -1219 -981 -1151 -947
rect -1061 -981 -993 -947
rect -903 -981 -835 -947
rect -745 -981 -677 -947
rect -587 -981 -519 -947
rect -429 -981 -361 -947
rect -271 -981 -203 -947
rect -113 -981 -45 -947
rect 45 -981 113 -947
rect 203 -981 271 -947
rect 361 -981 429 -947
rect 519 -981 587 -947
rect 677 -981 745 -947
rect 835 -981 903 -947
rect 993 -981 1061 -947
rect 1151 -981 1219 -947
rect 1309 -981 1377 -947
rect 1467 -981 1535 -947
rect 1625 -981 1693 -947
rect 1783 -981 1851 -947
rect 1941 -981 2009 -947
rect 2099 -981 2167 -947
rect 2257 -981 2325 -947
rect 2415 -981 2483 -947
rect -2483 -1089 -2415 -1055
rect -2325 -1089 -2257 -1055
rect -2167 -1089 -2099 -1055
rect -2009 -1089 -1941 -1055
rect -1851 -1089 -1783 -1055
rect -1693 -1089 -1625 -1055
rect -1535 -1089 -1467 -1055
rect -1377 -1089 -1309 -1055
rect -1219 -1089 -1151 -1055
rect -1061 -1089 -993 -1055
rect -903 -1089 -835 -1055
rect -745 -1089 -677 -1055
rect -587 -1089 -519 -1055
rect -429 -1089 -361 -1055
rect -271 -1089 -203 -1055
rect -113 -1089 -45 -1055
rect 45 -1089 113 -1055
rect 203 -1089 271 -1055
rect 361 -1089 429 -1055
rect 519 -1089 587 -1055
rect 677 -1089 745 -1055
rect 835 -1089 903 -1055
rect 993 -1089 1061 -1055
rect 1151 -1089 1219 -1055
rect 1309 -1089 1377 -1055
rect 1467 -1089 1535 -1055
rect 1625 -1089 1693 -1055
rect 1783 -1089 1851 -1055
rect 1941 -1089 2009 -1055
rect 2099 -1089 2167 -1055
rect 2257 -1089 2325 -1055
rect 2415 -1089 2483 -1055
rect -2545 -1915 -2511 -1139
rect -2387 -1915 -2353 -1139
rect -2229 -1915 -2195 -1139
rect -2071 -1915 -2037 -1139
rect -1913 -1915 -1879 -1139
rect -1755 -1915 -1721 -1139
rect -1597 -1915 -1563 -1139
rect -1439 -1915 -1405 -1139
rect -1281 -1915 -1247 -1139
rect -1123 -1915 -1089 -1139
rect -965 -1915 -931 -1139
rect -807 -1915 -773 -1139
rect -649 -1915 -615 -1139
rect -491 -1915 -457 -1139
rect -333 -1915 -299 -1139
rect -175 -1915 -141 -1139
rect -17 -1915 17 -1139
rect 141 -1915 175 -1139
rect 299 -1915 333 -1139
rect 457 -1915 491 -1139
rect 615 -1915 649 -1139
rect 773 -1915 807 -1139
rect 931 -1915 965 -1139
rect 1089 -1915 1123 -1139
rect 1247 -1915 1281 -1139
rect 1405 -1915 1439 -1139
rect 1563 -1915 1597 -1139
rect 1721 -1915 1755 -1139
rect 1879 -1915 1913 -1139
rect 2037 -1915 2071 -1139
rect 2195 -1915 2229 -1139
rect 2353 -1915 2387 -1139
rect 2511 -1915 2545 -1139
rect -2483 -1999 -2415 -1965
rect -2325 -1999 -2257 -1965
rect -2167 -1999 -2099 -1965
rect -2009 -1999 -1941 -1965
rect -1851 -1999 -1783 -1965
rect -1693 -1999 -1625 -1965
rect -1535 -1999 -1467 -1965
rect -1377 -1999 -1309 -1965
rect -1219 -1999 -1151 -1965
rect -1061 -1999 -993 -1965
rect -903 -1999 -835 -1965
rect -745 -1999 -677 -1965
rect -587 -1999 -519 -1965
rect -429 -1999 -361 -1965
rect -271 -1999 -203 -1965
rect -113 -1999 -45 -1965
rect 45 -1999 113 -1965
rect 203 -1999 271 -1965
rect 361 -1999 429 -1965
rect 519 -1999 587 -1965
rect 677 -1999 745 -1965
rect 835 -1999 903 -1965
rect 993 -1999 1061 -1965
rect 1151 -1999 1219 -1965
rect 1309 -1999 1377 -1965
rect 1467 -1999 1535 -1965
rect 1625 -1999 1693 -1965
rect 1783 -1999 1851 -1965
rect 1941 -1999 2009 -1965
rect 2099 -1999 2167 -1965
rect 2257 -1999 2325 -1965
rect 2415 -1999 2483 -1965
<< metal1 >>
rect -2495 1999 -2403 2005
rect -2495 1965 -2483 1999
rect -2415 1965 -2403 1999
rect -2495 1959 -2403 1965
rect -2337 1999 -2245 2005
rect -2337 1965 -2325 1999
rect -2257 1965 -2245 1999
rect -2337 1959 -2245 1965
rect -2179 1999 -2087 2005
rect -2179 1965 -2167 1999
rect -2099 1965 -2087 1999
rect -2179 1959 -2087 1965
rect -2021 1999 -1929 2005
rect -2021 1965 -2009 1999
rect -1941 1965 -1929 1999
rect -2021 1959 -1929 1965
rect -1863 1999 -1771 2005
rect -1863 1965 -1851 1999
rect -1783 1965 -1771 1999
rect -1863 1959 -1771 1965
rect -1705 1999 -1613 2005
rect -1705 1965 -1693 1999
rect -1625 1965 -1613 1999
rect -1705 1959 -1613 1965
rect -1547 1999 -1455 2005
rect -1547 1965 -1535 1999
rect -1467 1965 -1455 1999
rect -1547 1959 -1455 1965
rect -1389 1999 -1297 2005
rect -1389 1965 -1377 1999
rect -1309 1965 -1297 1999
rect -1389 1959 -1297 1965
rect -1231 1999 -1139 2005
rect -1231 1965 -1219 1999
rect -1151 1965 -1139 1999
rect -1231 1959 -1139 1965
rect -1073 1999 -981 2005
rect -1073 1965 -1061 1999
rect -993 1965 -981 1999
rect -1073 1959 -981 1965
rect -915 1999 -823 2005
rect -915 1965 -903 1999
rect -835 1965 -823 1999
rect -915 1959 -823 1965
rect -757 1999 -665 2005
rect -757 1965 -745 1999
rect -677 1965 -665 1999
rect -757 1959 -665 1965
rect -599 1999 -507 2005
rect -599 1965 -587 1999
rect -519 1965 -507 1999
rect -599 1959 -507 1965
rect -441 1999 -349 2005
rect -441 1965 -429 1999
rect -361 1965 -349 1999
rect -441 1959 -349 1965
rect -283 1999 -191 2005
rect -283 1965 -271 1999
rect -203 1965 -191 1999
rect -283 1959 -191 1965
rect -125 1999 -33 2005
rect -125 1965 -113 1999
rect -45 1965 -33 1999
rect -125 1959 -33 1965
rect 33 1999 125 2005
rect 33 1965 45 1999
rect 113 1965 125 1999
rect 33 1959 125 1965
rect 191 1999 283 2005
rect 191 1965 203 1999
rect 271 1965 283 1999
rect 191 1959 283 1965
rect 349 1999 441 2005
rect 349 1965 361 1999
rect 429 1965 441 1999
rect 349 1959 441 1965
rect 507 1999 599 2005
rect 507 1965 519 1999
rect 587 1965 599 1999
rect 507 1959 599 1965
rect 665 1999 757 2005
rect 665 1965 677 1999
rect 745 1965 757 1999
rect 665 1959 757 1965
rect 823 1999 915 2005
rect 823 1965 835 1999
rect 903 1965 915 1999
rect 823 1959 915 1965
rect 981 1999 1073 2005
rect 981 1965 993 1999
rect 1061 1965 1073 1999
rect 981 1959 1073 1965
rect 1139 1999 1231 2005
rect 1139 1965 1151 1999
rect 1219 1965 1231 1999
rect 1139 1959 1231 1965
rect 1297 1999 1389 2005
rect 1297 1965 1309 1999
rect 1377 1965 1389 1999
rect 1297 1959 1389 1965
rect 1455 1999 1547 2005
rect 1455 1965 1467 1999
rect 1535 1965 1547 1999
rect 1455 1959 1547 1965
rect 1613 1999 1705 2005
rect 1613 1965 1625 1999
rect 1693 1965 1705 1999
rect 1613 1959 1705 1965
rect 1771 1999 1863 2005
rect 1771 1965 1783 1999
rect 1851 1965 1863 1999
rect 1771 1959 1863 1965
rect 1929 1999 2021 2005
rect 1929 1965 1941 1999
rect 2009 1965 2021 1999
rect 1929 1959 2021 1965
rect 2087 1999 2179 2005
rect 2087 1965 2099 1999
rect 2167 1965 2179 1999
rect 2087 1959 2179 1965
rect 2245 1999 2337 2005
rect 2245 1965 2257 1999
rect 2325 1965 2337 1999
rect 2245 1959 2337 1965
rect 2403 1999 2495 2005
rect 2403 1965 2415 1999
rect 2483 1965 2495 1999
rect 2403 1959 2495 1965
rect -2551 1915 -2505 1927
rect -2551 1139 -2545 1915
rect -2511 1139 -2505 1915
rect -2551 1127 -2505 1139
rect -2393 1915 -2347 1927
rect -2393 1139 -2387 1915
rect -2353 1139 -2347 1915
rect -2393 1127 -2347 1139
rect -2235 1915 -2189 1927
rect -2235 1139 -2229 1915
rect -2195 1139 -2189 1915
rect -2235 1127 -2189 1139
rect -2077 1915 -2031 1927
rect -2077 1139 -2071 1915
rect -2037 1139 -2031 1915
rect -2077 1127 -2031 1139
rect -1919 1915 -1873 1927
rect -1919 1139 -1913 1915
rect -1879 1139 -1873 1915
rect -1919 1127 -1873 1139
rect -1761 1915 -1715 1927
rect -1761 1139 -1755 1915
rect -1721 1139 -1715 1915
rect -1761 1127 -1715 1139
rect -1603 1915 -1557 1927
rect -1603 1139 -1597 1915
rect -1563 1139 -1557 1915
rect -1603 1127 -1557 1139
rect -1445 1915 -1399 1927
rect -1445 1139 -1439 1915
rect -1405 1139 -1399 1915
rect -1445 1127 -1399 1139
rect -1287 1915 -1241 1927
rect -1287 1139 -1281 1915
rect -1247 1139 -1241 1915
rect -1287 1127 -1241 1139
rect -1129 1915 -1083 1927
rect -1129 1139 -1123 1915
rect -1089 1139 -1083 1915
rect -1129 1127 -1083 1139
rect -971 1915 -925 1927
rect -971 1139 -965 1915
rect -931 1139 -925 1915
rect -971 1127 -925 1139
rect -813 1915 -767 1927
rect -813 1139 -807 1915
rect -773 1139 -767 1915
rect -813 1127 -767 1139
rect -655 1915 -609 1927
rect -655 1139 -649 1915
rect -615 1139 -609 1915
rect -655 1127 -609 1139
rect -497 1915 -451 1927
rect -497 1139 -491 1915
rect -457 1139 -451 1915
rect -497 1127 -451 1139
rect -339 1915 -293 1927
rect -339 1139 -333 1915
rect -299 1139 -293 1915
rect -339 1127 -293 1139
rect -181 1915 -135 1927
rect -181 1139 -175 1915
rect -141 1139 -135 1915
rect -181 1127 -135 1139
rect -23 1915 23 1927
rect -23 1139 -17 1915
rect 17 1139 23 1915
rect -23 1127 23 1139
rect 135 1915 181 1927
rect 135 1139 141 1915
rect 175 1139 181 1915
rect 135 1127 181 1139
rect 293 1915 339 1927
rect 293 1139 299 1915
rect 333 1139 339 1915
rect 293 1127 339 1139
rect 451 1915 497 1927
rect 451 1139 457 1915
rect 491 1139 497 1915
rect 451 1127 497 1139
rect 609 1915 655 1927
rect 609 1139 615 1915
rect 649 1139 655 1915
rect 609 1127 655 1139
rect 767 1915 813 1927
rect 767 1139 773 1915
rect 807 1139 813 1915
rect 767 1127 813 1139
rect 925 1915 971 1927
rect 925 1139 931 1915
rect 965 1139 971 1915
rect 925 1127 971 1139
rect 1083 1915 1129 1927
rect 1083 1139 1089 1915
rect 1123 1139 1129 1915
rect 1083 1127 1129 1139
rect 1241 1915 1287 1927
rect 1241 1139 1247 1915
rect 1281 1139 1287 1915
rect 1241 1127 1287 1139
rect 1399 1915 1445 1927
rect 1399 1139 1405 1915
rect 1439 1139 1445 1915
rect 1399 1127 1445 1139
rect 1557 1915 1603 1927
rect 1557 1139 1563 1915
rect 1597 1139 1603 1915
rect 1557 1127 1603 1139
rect 1715 1915 1761 1927
rect 1715 1139 1721 1915
rect 1755 1139 1761 1915
rect 1715 1127 1761 1139
rect 1873 1915 1919 1927
rect 1873 1139 1879 1915
rect 1913 1139 1919 1915
rect 1873 1127 1919 1139
rect 2031 1915 2077 1927
rect 2031 1139 2037 1915
rect 2071 1139 2077 1915
rect 2031 1127 2077 1139
rect 2189 1915 2235 1927
rect 2189 1139 2195 1915
rect 2229 1139 2235 1915
rect 2189 1127 2235 1139
rect 2347 1915 2393 1927
rect 2347 1139 2353 1915
rect 2387 1139 2393 1915
rect 2347 1127 2393 1139
rect 2505 1915 2551 1927
rect 2505 1139 2511 1915
rect 2545 1139 2551 1915
rect 2505 1127 2551 1139
rect -2495 1089 -2403 1095
rect -2495 1055 -2483 1089
rect -2415 1055 -2403 1089
rect -2495 1049 -2403 1055
rect -2337 1089 -2245 1095
rect -2337 1055 -2325 1089
rect -2257 1055 -2245 1089
rect -2337 1049 -2245 1055
rect -2179 1089 -2087 1095
rect -2179 1055 -2167 1089
rect -2099 1055 -2087 1089
rect -2179 1049 -2087 1055
rect -2021 1089 -1929 1095
rect -2021 1055 -2009 1089
rect -1941 1055 -1929 1089
rect -2021 1049 -1929 1055
rect -1863 1089 -1771 1095
rect -1863 1055 -1851 1089
rect -1783 1055 -1771 1089
rect -1863 1049 -1771 1055
rect -1705 1089 -1613 1095
rect -1705 1055 -1693 1089
rect -1625 1055 -1613 1089
rect -1705 1049 -1613 1055
rect -1547 1089 -1455 1095
rect -1547 1055 -1535 1089
rect -1467 1055 -1455 1089
rect -1547 1049 -1455 1055
rect -1389 1089 -1297 1095
rect -1389 1055 -1377 1089
rect -1309 1055 -1297 1089
rect -1389 1049 -1297 1055
rect -1231 1089 -1139 1095
rect -1231 1055 -1219 1089
rect -1151 1055 -1139 1089
rect -1231 1049 -1139 1055
rect -1073 1089 -981 1095
rect -1073 1055 -1061 1089
rect -993 1055 -981 1089
rect -1073 1049 -981 1055
rect -915 1089 -823 1095
rect -915 1055 -903 1089
rect -835 1055 -823 1089
rect -915 1049 -823 1055
rect -757 1089 -665 1095
rect -757 1055 -745 1089
rect -677 1055 -665 1089
rect -757 1049 -665 1055
rect -599 1089 -507 1095
rect -599 1055 -587 1089
rect -519 1055 -507 1089
rect -599 1049 -507 1055
rect -441 1089 -349 1095
rect -441 1055 -429 1089
rect -361 1055 -349 1089
rect -441 1049 -349 1055
rect -283 1089 -191 1095
rect -283 1055 -271 1089
rect -203 1055 -191 1089
rect -283 1049 -191 1055
rect -125 1089 -33 1095
rect -125 1055 -113 1089
rect -45 1055 -33 1089
rect -125 1049 -33 1055
rect 33 1089 125 1095
rect 33 1055 45 1089
rect 113 1055 125 1089
rect 33 1049 125 1055
rect 191 1089 283 1095
rect 191 1055 203 1089
rect 271 1055 283 1089
rect 191 1049 283 1055
rect 349 1089 441 1095
rect 349 1055 361 1089
rect 429 1055 441 1089
rect 349 1049 441 1055
rect 507 1089 599 1095
rect 507 1055 519 1089
rect 587 1055 599 1089
rect 507 1049 599 1055
rect 665 1089 757 1095
rect 665 1055 677 1089
rect 745 1055 757 1089
rect 665 1049 757 1055
rect 823 1089 915 1095
rect 823 1055 835 1089
rect 903 1055 915 1089
rect 823 1049 915 1055
rect 981 1089 1073 1095
rect 981 1055 993 1089
rect 1061 1055 1073 1089
rect 981 1049 1073 1055
rect 1139 1089 1231 1095
rect 1139 1055 1151 1089
rect 1219 1055 1231 1089
rect 1139 1049 1231 1055
rect 1297 1089 1389 1095
rect 1297 1055 1309 1089
rect 1377 1055 1389 1089
rect 1297 1049 1389 1055
rect 1455 1089 1547 1095
rect 1455 1055 1467 1089
rect 1535 1055 1547 1089
rect 1455 1049 1547 1055
rect 1613 1089 1705 1095
rect 1613 1055 1625 1089
rect 1693 1055 1705 1089
rect 1613 1049 1705 1055
rect 1771 1089 1863 1095
rect 1771 1055 1783 1089
rect 1851 1055 1863 1089
rect 1771 1049 1863 1055
rect 1929 1089 2021 1095
rect 1929 1055 1941 1089
rect 2009 1055 2021 1089
rect 1929 1049 2021 1055
rect 2087 1089 2179 1095
rect 2087 1055 2099 1089
rect 2167 1055 2179 1089
rect 2087 1049 2179 1055
rect 2245 1089 2337 1095
rect 2245 1055 2257 1089
rect 2325 1055 2337 1089
rect 2245 1049 2337 1055
rect 2403 1089 2495 1095
rect 2403 1055 2415 1089
rect 2483 1055 2495 1089
rect 2403 1049 2495 1055
rect -2495 981 -2403 987
rect -2495 947 -2483 981
rect -2415 947 -2403 981
rect -2495 941 -2403 947
rect -2337 981 -2245 987
rect -2337 947 -2325 981
rect -2257 947 -2245 981
rect -2337 941 -2245 947
rect -2179 981 -2087 987
rect -2179 947 -2167 981
rect -2099 947 -2087 981
rect -2179 941 -2087 947
rect -2021 981 -1929 987
rect -2021 947 -2009 981
rect -1941 947 -1929 981
rect -2021 941 -1929 947
rect -1863 981 -1771 987
rect -1863 947 -1851 981
rect -1783 947 -1771 981
rect -1863 941 -1771 947
rect -1705 981 -1613 987
rect -1705 947 -1693 981
rect -1625 947 -1613 981
rect -1705 941 -1613 947
rect -1547 981 -1455 987
rect -1547 947 -1535 981
rect -1467 947 -1455 981
rect -1547 941 -1455 947
rect -1389 981 -1297 987
rect -1389 947 -1377 981
rect -1309 947 -1297 981
rect -1389 941 -1297 947
rect -1231 981 -1139 987
rect -1231 947 -1219 981
rect -1151 947 -1139 981
rect -1231 941 -1139 947
rect -1073 981 -981 987
rect -1073 947 -1061 981
rect -993 947 -981 981
rect -1073 941 -981 947
rect -915 981 -823 987
rect -915 947 -903 981
rect -835 947 -823 981
rect -915 941 -823 947
rect -757 981 -665 987
rect -757 947 -745 981
rect -677 947 -665 981
rect -757 941 -665 947
rect -599 981 -507 987
rect -599 947 -587 981
rect -519 947 -507 981
rect -599 941 -507 947
rect -441 981 -349 987
rect -441 947 -429 981
rect -361 947 -349 981
rect -441 941 -349 947
rect -283 981 -191 987
rect -283 947 -271 981
rect -203 947 -191 981
rect -283 941 -191 947
rect -125 981 -33 987
rect -125 947 -113 981
rect -45 947 -33 981
rect -125 941 -33 947
rect 33 981 125 987
rect 33 947 45 981
rect 113 947 125 981
rect 33 941 125 947
rect 191 981 283 987
rect 191 947 203 981
rect 271 947 283 981
rect 191 941 283 947
rect 349 981 441 987
rect 349 947 361 981
rect 429 947 441 981
rect 349 941 441 947
rect 507 981 599 987
rect 507 947 519 981
rect 587 947 599 981
rect 507 941 599 947
rect 665 981 757 987
rect 665 947 677 981
rect 745 947 757 981
rect 665 941 757 947
rect 823 981 915 987
rect 823 947 835 981
rect 903 947 915 981
rect 823 941 915 947
rect 981 981 1073 987
rect 981 947 993 981
rect 1061 947 1073 981
rect 981 941 1073 947
rect 1139 981 1231 987
rect 1139 947 1151 981
rect 1219 947 1231 981
rect 1139 941 1231 947
rect 1297 981 1389 987
rect 1297 947 1309 981
rect 1377 947 1389 981
rect 1297 941 1389 947
rect 1455 981 1547 987
rect 1455 947 1467 981
rect 1535 947 1547 981
rect 1455 941 1547 947
rect 1613 981 1705 987
rect 1613 947 1625 981
rect 1693 947 1705 981
rect 1613 941 1705 947
rect 1771 981 1863 987
rect 1771 947 1783 981
rect 1851 947 1863 981
rect 1771 941 1863 947
rect 1929 981 2021 987
rect 1929 947 1941 981
rect 2009 947 2021 981
rect 1929 941 2021 947
rect 2087 981 2179 987
rect 2087 947 2099 981
rect 2167 947 2179 981
rect 2087 941 2179 947
rect 2245 981 2337 987
rect 2245 947 2257 981
rect 2325 947 2337 981
rect 2245 941 2337 947
rect 2403 981 2495 987
rect 2403 947 2415 981
rect 2483 947 2495 981
rect 2403 941 2495 947
rect -2551 897 -2505 909
rect -2551 121 -2545 897
rect -2511 121 -2505 897
rect -2551 109 -2505 121
rect -2393 897 -2347 909
rect -2393 121 -2387 897
rect -2353 121 -2347 897
rect -2393 109 -2347 121
rect -2235 897 -2189 909
rect -2235 121 -2229 897
rect -2195 121 -2189 897
rect -2235 109 -2189 121
rect -2077 897 -2031 909
rect -2077 121 -2071 897
rect -2037 121 -2031 897
rect -2077 109 -2031 121
rect -1919 897 -1873 909
rect -1919 121 -1913 897
rect -1879 121 -1873 897
rect -1919 109 -1873 121
rect -1761 897 -1715 909
rect -1761 121 -1755 897
rect -1721 121 -1715 897
rect -1761 109 -1715 121
rect -1603 897 -1557 909
rect -1603 121 -1597 897
rect -1563 121 -1557 897
rect -1603 109 -1557 121
rect -1445 897 -1399 909
rect -1445 121 -1439 897
rect -1405 121 -1399 897
rect -1445 109 -1399 121
rect -1287 897 -1241 909
rect -1287 121 -1281 897
rect -1247 121 -1241 897
rect -1287 109 -1241 121
rect -1129 897 -1083 909
rect -1129 121 -1123 897
rect -1089 121 -1083 897
rect -1129 109 -1083 121
rect -971 897 -925 909
rect -971 121 -965 897
rect -931 121 -925 897
rect -971 109 -925 121
rect -813 897 -767 909
rect -813 121 -807 897
rect -773 121 -767 897
rect -813 109 -767 121
rect -655 897 -609 909
rect -655 121 -649 897
rect -615 121 -609 897
rect -655 109 -609 121
rect -497 897 -451 909
rect -497 121 -491 897
rect -457 121 -451 897
rect -497 109 -451 121
rect -339 897 -293 909
rect -339 121 -333 897
rect -299 121 -293 897
rect -339 109 -293 121
rect -181 897 -135 909
rect -181 121 -175 897
rect -141 121 -135 897
rect -181 109 -135 121
rect -23 897 23 909
rect -23 121 -17 897
rect 17 121 23 897
rect -23 109 23 121
rect 135 897 181 909
rect 135 121 141 897
rect 175 121 181 897
rect 135 109 181 121
rect 293 897 339 909
rect 293 121 299 897
rect 333 121 339 897
rect 293 109 339 121
rect 451 897 497 909
rect 451 121 457 897
rect 491 121 497 897
rect 451 109 497 121
rect 609 897 655 909
rect 609 121 615 897
rect 649 121 655 897
rect 609 109 655 121
rect 767 897 813 909
rect 767 121 773 897
rect 807 121 813 897
rect 767 109 813 121
rect 925 897 971 909
rect 925 121 931 897
rect 965 121 971 897
rect 925 109 971 121
rect 1083 897 1129 909
rect 1083 121 1089 897
rect 1123 121 1129 897
rect 1083 109 1129 121
rect 1241 897 1287 909
rect 1241 121 1247 897
rect 1281 121 1287 897
rect 1241 109 1287 121
rect 1399 897 1445 909
rect 1399 121 1405 897
rect 1439 121 1445 897
rect 1399 109 1445 121
rect 1557 897 1603 909
rect 1557 121 1563 897
rect 1597 121 1603 897
rect 1557 109 1603 121
rect 1715 897 1761 909
rect 1715 121 1721 897
rect 1755 121 1761 897
rect 1715 109 1761 121
rect 1873 897 1919 909
rect 1873 121 1879 897
rect 1913 121 1919 897
rect 1873 109 1919 121
rect 2031 897 2077 909
rect 2031 121 2037 897
rect 2071 121 2077 897
rect 2031 109 2077 121
rect 2189 897 2235 909
rect 2189 121 2195 897
rect 2229 121 2235 897
rect 2189 109 2235 121
rect 2347 897 2393 909
rect 2347 121 2353 897
rect 2387 121 2393 897
rect 2347 109 2393 121
rect 2505 897 2551 909
rect 2505 121 2511 897
rect 2545 121 2551 897
rect 2505 109 2551 121
rect -2495 71 -2403 77
rect -2495 37 -2483 71
rect -2415 37 -2403 71
rect -2495 31 -2403 37
rect -2337 71 -2245 77
rect -2337 37 -2325 71
rect -2257 37 -2245 71
rect -2337 31 -2245 37
rect -2179 71 -2087 77
rect -2179 37 -2167 71
rect -2099 37 -2087 71
rect -2179 31 -2087 37
rect -2021 71 -1929 77
rect -2021 37 -2009 71
rect -1941 37 -1929 71
rect -2021 31 -1929 37
rect -1863 71 -1771 77
rect -1863 37 -1851 71
rect -1783 37 -1771 71
rect -1863 31 -1771 37
rect -1705 71 -1613 77
rect -1705 37 -1693 71
rect -1625 37 -1613 71
rect -1705 31 -1613 37
rect -1547 71 -1455 77
rect -1547 37 -1535 71
rect -1467 37 -1455 71
rect -1547 31 -1455 37
rect -1389 71 -1297 77
rect -1389 37 -1377 71
rect -1309 37 -1297 71
rect -1389 31 -1297 37
rect -1231 71 -1139 77
rect -1231 37 -1219 71
rect -1151 37 -1139 71
rect -1231 31 -1139 37
rect -1073 71 -981 77
rect -1073 37 -1061 71
rect -993 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -903 71
rect -835 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 835 71
rect 903 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 993 71
rect 1061 37 1073 71
rect 981 31 1073 37
rect 1139 71 1231 77
rect 1139 37 1151 71
rect 1219 37 1231 71
rect 1139 31 1231 37
rect 1297 71 1389 77
rect 1297 37 1309 71
rect 1377 37 1389 71
rect 1297 31 1389 37
rect 1455 71 1547 77
rect 1455 37 1467 71
rect 1535 37 1547 71
rect 1455 31 1547 37
rect 1613 71 1705 77
rect 1613 37 1625 71
rect 1693 37 1705 71
rect 1613 31 1705 37
rect 1771 71 1863 77
rect 1771 37 1783 71
rect 1851 37 1863 71
rect 1771 31 1863 37
rect 1929 71 2021 77
rect 1929 37 1941 71
rect 2009 37 2021 71
rect 1929 31 2021 37
rect 2087 71 2179 77
rect 2087 37 2099 71
rect 2167 37 2179 71
rect 2087 31 2179 37
rect 2245 71 2337 77
rect 2245 37 2257 71
rect 2325 37 2337 71
rect 2245 31 2337 37
rect 2403 71 2495 77
rect 2403 37 2415 71
rect 2483 37 2495 71
rect 2403 31 2495 37
rect -2495 -37 -2403 -31
rect -2495 -71 -2483 -37
rect -2415 -71 -2403 -37
rect -2495 -77 -2403 -71
rect -2337 -37 -2245 -31
rect -2337 -71 -2325 -37
rect -2257 -71 -2245 -37
rect -2337 -77 -2245 -71
rect -2179 -37 -2087 -31
rect -2179 -71 -2167 -37
rect -2099 -71 -2087 -37
rect -2179 -77 -2087 -71
rect -2021 -37 -1929 -31
rect -2021 -71 -2009 -37
rect -1941 -71 -1929 -37
rect -2021 -77 -1929 -71
rect -1863 -37 -1771 -31
rect -1863 -71 -1851 -37
rect -1783 -71 -1771 -37
rect -1863 -77 -1771 -71
rect -1705 -37 -1613 -31
rect -1705 -71 -1693 -37
rect -1625 -71 -1613 -37
rect -1705 -77 -1613 -71
rect -1547 -37 -1455 -31
rect -1547 -71 -1535 -37
rect -1467 -71 -1455 -37
rect -1547 -77 -1455 -71
rect -1389 -37 -1297 -31
rect -1389 -71 -1377 -37
rect -1309 -71 -1297 -37
rect -1389 -77 -1297 -71
rect -1231 -37 -1139 -31
rect -1231 -71 -1219 -37
rect -1151 -71 -1139 -37
rect -1231 -77 -1139 -71
rect -1073 -37 -981 -31
rect -1073 -71 -1061 -37
rect -993 -71 -981 -37
rect -1073 -77 -981 -71
rect -915 -37 -823 -31
rect -915 -71 -903 -37
rect -835 -71 -823 -37
rect -915 -77 -823 -71
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect 823 -37 915 -31
rect 823 -71 835 -37
rect 903 -71 915 -37
rect 823 -77 915 -71
rect 981 -37 1073 -31
rect 981 -71 993 -37
rect 1061 -71 1073 -37
rect 981 -77 1073 -71
rect 1139 -37 1231 -31
rect 1139 -71 1151 -37
rect 1219 -71 1231 -37
rect 1139 -77 1231 -71
rect 1297 -37 1389 -31
rect 1297 -71 1309 -37
rect 1377 -71 1389 -37
rect 1297 -77 1389 -71
rect 1455 -37 1547 -31
rect 1455 -71 1467 -37
rect 1535 -71 1547 -37
rect 1455 -77 1547 -71
rect 1613 -37 1705 -31
rect 1613 -71 1625 -37
rect 1693 -71 1705 -37
rect 1613 -77 1705 -71
rect 1771 -37 1863 -31
rect 1771 -71 1783 -37
rect 1851 -71 1863 -37
rect 1771 -77 1863 -71
rect 1929 -37 2021 -31
rect 1929 -71 1941 -37
rect 2009 -71 2021 -37
rect 1929 -77 2021 -71
rect 2087 -37 2179 -31
rect 2087 -71 2099 -37
rect 2167 -71 2179 -37
rect 2087 -77 2179 -71
rect 2245 -37 2337 -31
rect 2245 -71 2257 -37
rect 2325 -71 2337 -37
rect 2245 -77 2337 -71
rect 2403 -37 2495 -31
rect 2403 -71 2415 -37
rect 2483 -71 2495 -37
rect 2403 -77 2495 -71
rect -2551 -121 -2505 -109
rect -2551 -897 -2545 -121
rect -2511 -897 -2505 -121
rect -2551 -909 -2505 -897
rect -2393 -121 -2347 -109
rect -2393 -897 -2387 -121
rect -2353 -897 -2347 -121
rect -2393 -909 -2347 -897
rect -2235 -121 -2189 -109
rect -2235 -897 -2229 -121
rect -2195 -897 -2189 -121
rect -2235 -909 -2189 -897
rect -2077 -121 -2031 -109
rect -2077 -897 -2071 -121
rect -2037 -897 -2031 -121
rect -2077 -909 -2031 -897
rect -1919 -121 -1873 -109
rect -1919 -897 -1913 -121
rect -1879 -897 -1873 -121
rect -1919 -909 -1873 -897
rect -1761 -121 -1715 -109
rect -1761 -897 -1755 -121
rect -1721 -897 -1715 -121
rect -1761 -909 -1715 -897
rect -1603 -121 -1557 -109
rect -1603 -897 -1597 -121
rect -1563 -897 -1557 -121
rect -1603 -909 -1557 -897
rect -1445 -121 -1399 -109
rect -1445 -897 -1439 -121
rect -1405 -897 -1399 -121
rect -1445 -909 -1399 -897
rect -1287 -121 -1241 -109
rect -1287 -897 -1281 -121
rect -1247 -897 -1241 -121
rect -1287 -909 -1241 -897
rect -1129 -121 -1083 -109
rect -1129 -897 -1123 -121
rect -1089 -897 -1083 -121
rect -1129 -909 -1083 -897
rect -971 -121 -925 -109
rect -971 -897 -965 -121
rect -931 -897 -925 -121
rect -971 -909 -925 -897
rect -813 -121 -767 -109
rect -813 -897 -807 -121
rect -773 -897 -767 -121
rect -813 -909 -767 -897
rect -655 -121 -609 -109
rect -655 -897 -649 -121
rect -615 -897 -609 -121
rect -655 -909 -609 -897
rect -497 -121 -451 -109
rect -497 -897 -491 -121
rect -457 -897 -451 -121
rect -497 -909 -451 -897
rect -339 -121 -293 -109
rect -339 -897 -333 -121
rect -299 -897 -293 -121
rect -339 -909 -293 -897
rect -181 -121 -135 -109
rect -181 -897 -175 -121
rect -141 -897 -135 -121
rect -181 -909 -135 -897
rect -23 -121 23 -109
rect -23 -897 -17 -121
rect 17 -897 23 -121
rect -23 -909 23 -897
rect 135 -121 181 -109
rect 135 -897 141 -121
rect 175 -897 181 -121
rect 135 -909 181 -897
rect 293 -121 339 -109
rect 293 -897 299 -121
rect 333 -897 339 -121
rect 293 -909 339 -897
rect 451 -121 497 -109
rect 451 -897 457 -121
rect 491 -897 497 -121
rect 451 -909 497 -897
rect 609 -121 655 -109
rect 609 -897 615 -121
rect 649 -897 655 -121
rect 609 -909 655 -897
rect 767 -121 813 -109
rect 767 -897 773 -121
rect 807 -897 813 -121
rect 767 -909 813 -897
rect 925 -121 971 -109
rect 925 -897 931 -121
rect 965 -897 971 -121
rect 925 -909 971 -897
rect 1083 -121 1129 -109
rect 1083 -897 1089 -121
rect 1123 -897 1129 -121
rect 1083 -909 1129 -897
rect 1241 -121 1287 -109
rect 1241 -897 1247 -121
rect 1281 -897 1287 -121
rect 1241 -909 1287 -897
rect 1399 -121 1445 -109
rect 1399 -897 1405 -121
rect 1439 -897 1445 -121
rect 1399 -909 1445 -897
rect 1557 -121 1603 -109
rect 1557 -897 1563 -121
rect 1597 -897 1603 -121
rect 1557 -909 1603 -897
rect 1715 -121 1761 -109
rect 1715 -897 1721 -121
rect 1755 -897 1761 -121
rect 1715 -909 1761 -897
rect 1873 -121 1919 -109
rect 1873 -897 1879 -121
rect 1913 -897 1919 -121
rect 1873 -909 1919 -897
rect 2031 -121 2077 -109
rect 2031 -897 2037 -121
rect 2071 -897 2077 -121
rect 2031 -909 2077 -897
rect 2189 -121 2235 -109
rect 2189 -897 2195 -121
rect 2229 -897 2235 -121
rect 2189 -909 2235 -897
rect 2347 -121 2393 -109
rect 2347 -897 2353 -121
rect 2387 -897 2393 -121
rect 2347 -909 2393 -897
rect 2505 -121 2551 -109
rect 2505 -897 2511 -121
rect 2545 -897 2551 -121
rect 2505 -909 2551 -897
rect -2495 -947 -2403 -941
rect -2495 -981 -2483 -947
rect -2415 -981 -2403 -947
rect -2495 -987 -2403 -981
rect -2337 -947 -2245 -941
rect -2337 -981 -2325 -947
rect -2257 -981 -2245 -947
rect -2337 -987 -2245 -981
rect -2179 -947 -2087 -941
rect -2179 -981 -2167 -947
rect -2099 -981 -2087 -947
rect -2179 -987 -2087 -981
rect -2021 -947 -1929 -941
rect -2021 -981 -2009 -947
rect -1941 -981 -1929 -947
rect -2021 -987 -1929 -981
rect -1863 -947 -1771 -941
rect -1863 -981 -1851 -947
rect -1783 -981 -1771 -947
rect -1863 -987 -1771 -981
rect -1705 -947 -1613 -941
rect -1705 -981 -1693 -947
rect -1625 -981 -1613 -947
rect -1705 -987 -1613 -981
rect -1547 -947 -1455 -941
rect -1547 -981 -1535 -947
rect -1467 -981 -1455 -947
rect -1547 -987 -1455 -981
rect -1389 -947 -1297 -941
rect -1389 -981 -1377 -947
rect -1309 -981 -1297 -947
rect -1389 -987 -1297 -981
rect -1231 -947 -1139 -941
rect -1231 -981 -1219 -947
rect -1151 -981 -1139 -947
rect -1231 -987 -1139 -981
rect -1073 -947 -981 -941
rect -1073 -981 -1061 -947
rect -993 -981 -981 -947
rect -1073 -987 -981 -981
rect -915 -947 -823 -941
rect -915 -981 -903 -947
rect -835 -981 -823 -947
rect -915 -987 -823 -981
rect -757 -947 -665 -941
rect -757 -981 -745 -947
rect -677 -981 -665 -947
rect -757 -987 -665 -981
rect -599 -947 -507 -941
rect -599 -981 -587 -947
rect -519 -981 -507 -947
rect -599 -987 -507 -981
rect -441 -947 -349 -941
rect -441 -981 -429 -947
rect -361 -981 -349 -947
rect -441 -987 -349 -981
rect -283 -947 -191 -941
rect -283 -981 -271 -947
rect -203 -981 -191 -947
rect -283 -987 -191 -981
rect -125 -947 -33 -941
rect -125 -981 -113 -947
rect -45 -981 -33 -947
rect -125 -987 -33 -981
rect 33 -947 125 -941
rect 33 -981 45 -947
rect 113 -981 125 -947
rect 33 -987 125 -981
rect 191 -947 283 -941
rect 191 -981 203 -947
rect 271 -981 283 -947
rect 191 -987 283 -981
rect 349 -947 441 -941
rect 349 -981 361 -947
rect 429 -981 441 -947
rect 349 -987 441 -981
rect 507 -947 599 -941
rect 507 -981 519 -947
rect 587 -981 599 -947
rect 507 -987 599 -981
rect 665 -947 757 -941
rect 665 -981 677 -947
rect 745 -981 757 -947
rect 665 -987 757 -981
rect 823 -947 915 -941
rect 823 -981 835 -947
rect 903 -981 915 -947
rect 823 -987 915 -981
rect 981 -947 1073 -941
rect 981 -981 993 -947
rect 1061 -981 1073 -947
rect 981 -987 1073 -981
rect 1139 -947 1231 -941
rect 1139 -981 1151 -947
rect 1219 -981 1231 -947
rect 1139 -987 1231 -981
rect 1297 -947 1389 -941
rect 1297 -981 1309 -947
rect 1377 -981 1389 -947
rect 1297 -987 1389 -981
rect 1455 -947 1547 -941
rect 1455 -981 1467 -947
rect 1535 -981 1547 -947
rect 1455 -987 1547 -981
rect 1613 -947 1705 -941
rect 1613 -981 1625 -947
rect 1693 -981 1705 -947
rect 1613 -987 1705 -981
rect 1771 -947 1863 -941
rect 1771 -981 1783 -947
rect 1851 -981 1863 -947
rect 1771 -987 1863 -981
rect 1929 -947 2021 -941
rect 1929 -981 1941 -947
rect 2009 -981 2021 -947
rect 1929 -987 2021 -981
rect 2087 -947 2179 -941
rect 2087 -981 2099 -947
rect 2167 -981 2179 -947
rect 2087 -987 2179 -981
rect 2245 -947 2337 -941
rect 2245 -981 2257 -947
rect 2325 -981 2337 -947
rect 2245 -987 2337 -981
rect 2403 -947 2495 -941
rect 2403 -981 2415 -947
rect 2483 -981 2495 -947
rect 2403 -987 2495 -981
rect -2495 -1055 -2403 -1049
rect -2495 -1089 -2483 -1055
rect -2415 -1089 -2403 -1055
rect -2495 -1095 -2403 -1089
rect -2337 -1055 -2245 -1049
rect -2337 -1089 -2325 -1055
rect -2257 -1089 -2245 -1055
rect -2337 -1095 -2245 -1089
rect -2179 -1055 -2087 -1049
rect -2179 -1089 -2167 -1055
rect -2099 -1089 -2087 -1055
rect -2179 -1095 -2087 -1089
rect -2021 -1055 -1929 -1049
rect -2021 -1089 -2009 -1055
rect -1941 -1089 -1929 -1055
rect -2021 -1095 -1929 -1089
rect -1863 -1055 -1771 -1049
rect -1863 -1089 -1851 -1055
rect -1783 -1089 -1771 -1055
rect -1863 -1095 -1771 -1089
rect -1705 -1055 -1613 -1049
rect -1705 -1089 -1693 -1055
rect -1625 -1089 -1613 -1055
rect -1705 -1095 -1613 -1089
rect -1547 -1055 -1455 -1049
rect -1547 -1089 -1535 -1055
rect -1467 -1089 -1455 -1055
rect -1547 -1095 -1455 -1089
rect -1389 -1055 -1297 -1049
rect -1389 -1089 -1377 -1055
rect -1309 -1089 -1297 -1055
rect -1389 -1095 -1297 -1089
rect -1231 -1055 -1139 -1049
rect -1231 -1089 -1219 -1055
rect -1151 -1089 -1139 -1055
rect -1231 -1095 -1139 -1089
rect -1073 -1055 -981 -1049
rect -1073 -1089 -1061 -1055
rect -993 -1089 -981 -1055
rect -1073 -1095 -981 -1089
rect -915 -1055 -823 -1049
rect -915 -1089 -903 -1055
rect -835 -1089 -823 -1055
rect -915 -1095 -823 -1089
rect -757 -1055 -665 -1049
rect -757 -1089 -745 -1055
rect -677 -1089 -665 -1055
rect -757 -1095 -665 -1089
rect -599 -1055 -507 -1049
rect -599 -1089 -587 -1055
rect -519 -1089 -507 -1055
rect -599 -1095 -507 -1089
rect -441 -1055 -349 -1049
rect -441 -1089 -429 -1055
rect -361 -1089 -349 -1055
rect -441 -1095 -349 -1089
rect -283 -1055 -191 -1049
rect -283 -1089 -271 -1055
rect -203 -1089 -191 -1055
rect -283 -1095 -191 -1089
rect -125 -1055 -33 -1049
rect -125 -1089 -113 -1055
rect -45 -1089 -33 -1055
rect -125 -1095 -33 -1089
rect 33 -1055 125 -1049
rect 33 -1089 45 -1055
rect 113 -1089 125 -1055
rect 33 -1095 125 -1089
rect 191 -1055 283 -1049
rect 191 -1089 203 -1055
rect 271 -1089 283 -1055
rect 191 -1095 283 -1089
rect 349 -1055 441 -1049
rect 349 -1089 361 -1055
rect 429 -1089 441 -1055
rect 349 -1095 441 -1089
rect 507 -1055 599 -1049
rect 507 -1089 519 -1055
rect 587 -1089 599 -1055
rect 507 -1095 599 -1089
rect 665 -1055 757 -1049
rect 665 -1089 677 -1055
rect 745 -1089 757 -1055
rect 665 -1095 757 -1089
rect 823 -1055 915 -1049
rect 823 -1089 835 -1055
rect 903 -1089 915 -1055
rect 823 -1095 915 -1089
rect 981 -1055 1073 -1049
rect 981 -1089 993 -1055
rect 1061 -1089 1073 -1055
rect 981 -1095 1073 -1089
rect 1139 -1055 1231 -1049
rect 1139 -1089 1151 -1055
rect 1219 -1089 1231 -1055
rect 1139 -1095 1231 -1089
rect 1297 -1055 1389 -1049
rect 1297 -1089 1309 -1055
rect 1377 -1089 1389 -1055
rect 1297 -1095 1389 -1089
rect 1455 -1055 1547 -1049
rect 1455 -1089 1467 -1055
rect 1535 -1089 1547 -1055
rect 1455 -1095 1547 -1089
rect 1613 -1055 1705 -1049
rect 1613 -1089 1625 -1055
rect 1693 -1089 1705 -1055
rect 1613 -1095 1705 -1089
rect 1771 -1055 1863 -1049
rect 1771 -1089 1783 -1055
rect 1851 -1089 1863 -1055
rect 1771 -1095 1863 -1089
rect 1929 -1055 2021 -1049
rect 1929 -1089 1941 -1055
rect 2009 -1089 2021 -1055
rect 1929 -1095 2021 -1089
rect 2087 -1055 2179 -1049
rect 2087 -1089 2099 -1055
rect 2167 -1089 2179 -1055
rect 2087 -1095 2179 -1089
rect 2245 -1055 2337 -1049
rect 2245 -1089 2257 -1055
rect 2325 -1089 2337 -1055
rect 2245 -1095 2337 -1089
rect 2403 -1055 2495 -1049
rect 2403 -1089 2415 -1055
rect 2483 -1089 2495 -1055
rect 2403 -1095 2495 -1089
rect -2551 -1139 -2505 -1127
rect -2551 -1915 -2545 -1139
rect -2511 -1915 -2505 -1139
rect -2551 -1927 -2505 -1915
rect -2393 -1139 -2347 -1127
rect -2393 -1915 -2387 -1139
rect -2353 -1915 -2347 -1139
rect -2393 -1927 -2347 -1915
rect -2235 -1139 -2189 -1127
rect -2235 -1915 -2229 -1139
rect -2195 -1915 -2189 -1139
rect -2235 -1927 -2189 -1915
rect -2077 -1139 -2031 -1127
rect -2077 -1915 -2071 -1139
rect -2037 -1915 -2031 -1139
rect -2077 -1927 -2031 -1915
rect -1919 -1139 -1873 -1127
rect -1919 -1915 -1913 -1139
rect -1879 -1915 -1873 -1139
rect -1919 -1927 -1873 -1915
rect -1761 -1139 -1715 -1127
rect -1761 -1915 -1755 -1139
rect -1721 -1915 -1715 -1139
rect -1761 -1927 -1715 -1915
rect -1603 -1139 -1557 -1127
rect -1603 -1915 -1597 -1139
rect -1563 -1915 -1557 -1139
rect -1603 -1927 -1557 -1915
rect -1445 -1139 -1399 -1127
rect -1445 -1915 -1439 -1139
rect -1405 -1915 -1399 -1139
rect -1445 -1927 -1399 -1915
rect -1287 -1139 -1241 -1127
rect -1287 -1915 -1281 -1139
rect -1247 -1915 -1241 -1139
rect -1287 -1927 -1241 -1915
rect -1129 -1139 -1083 -1127
rect -1129 -1915 -1123 -1139
rect -1089 -1915 -1083 -1139
rect -1129 -1927 -1083 -1915
rect -971 -1139 -925 -1127
rect -971 -1915 -965 -1139
rect -931 -1915 -925 -1139
rect -971 -1927 -925 -1915
rect -813 -1139 -767 -1127
rect -813 -1915 -807 -1139
rect -773 -1915 -767 -1139
rect -813 -1927 -767 -1915
rect -655 -1139 -609 -1127
rect -655 -1915 -649 -1139
rect -615 -1915 -609 -1139
rect -655 -1927 -609 -1915
rect -497 -1139 -451 -1127
rect -497 -1915 -491 -1139
rect -457 -1915 -451 -1139
rect -497 -1927 -451 -1915
rect -339 -1139 -293 -1127
rect -339 -1915 -333 -1139
rect -299 -1915 -293 -1139
rect -339 -1927 -293 -1915
rect -181 -1139 -135 -1127
rect -181 -1915 -175 -1139
rect -141 -1915 -135 -1139
rect -181 -1927 -135 -1915
rect -23 -1139 23 -1127
rect -23 -1915 -17 -1139
rect 17 -1915 23 -1139
rect -23 -1927 23 -1915
rect 135 -1139 181 -1127
rect 135 -1915 141 -1139
rect 175 -1915 181 -1139
rect 135 -1927 181 -1915
rect 293 -1139 339 -1127
rect 293 -1915 299 -1139
rect 333 -1915 339 -1139
rect 293 -1927 339 -1915
rect 451 -1139 497 -1127
rect 451 -1915 457 -1139
rect 491 -1915 497 -1139
rect 451 -1927 497 -1915
rect 609 -1139 655 -1127
rect 609 -1915 615 -1139
rect 649 -1915 655 -1139
rect 609 -1927 655 -1915
rect 767 -1139 813 -1127
rect 767 -1915 773 -1139
rect 807 -1915 813 -1139
rect 767 -1927 813 -1915
rect 925 -1139 971 -1127
rect 925 -1915 931 -1139
rect 965 -1915 971 -1139
rect 925 -1927 971 -1915
rect 1083 -1139 1129 -1127
rect 1083 -1915 1089 -1139
rect 1123 -1915 1129 -1139
rect 1083 -1927 1129 -1915
rect 1241 -1139 1287 -1127
rect 1241 -1915 1247 -1139
rect 1281 -1915 1287 -1139
rect 1241 -1927 1287 -1915
rect 1399 -1139 1445 -1127
rect 1399 -1915 1405 -1139
rect 1439 -1915 1445 -1139
rect 1399 -1927 1445 -1915
rect 1557 -1139 1603 -1127
rect 1557 -1915 1563 -1139
rect 1597 -1915 1603 -1139
rect 1557 -1927 1603 -1915
rect 1715 -1139 1761 -1127
rect 1715 -1915 1721 -1139
rect 1755 -1915 1761 -1139
rect 1715 -1927 1761 -1915
rect 1873 -1139 1919 -1127
rect 1873 -1915 1879 -1139
rect 1913 -1915 1919 -1139
rect 1873 -1927 1919 -1915
rect 2031 -1139 2077 -1127
rect 2031 -1915 2037 -1139
rect 2071 -1915 2077 -1139
rect 2031 -1927 2077 -1915
rect 2189 -1139 2235 -1127
rect 2189 -1915 2195 -1139
rect 2229 -1915 2235 -1139
rect 2189 -1927 2235 -1915
rect 2347 -1139 2393 -1127
rect 2347 -1915 2353 -1139
rect 2387 -1915 2393 -1139
rect 2347 -1927 2393 -1915
rect 2505 -1139 2551 -1127
rect 2505 -1915 2511 -1139
rect 2545 -1915 2551 -1139
rect 2505 -1927 2551 -1915
rect -2495 -1965 -2403 -1959
rect -2495 -1999 -2483 -1965
rect -2415 -1999 -2403 -1965
rect -2495 -2005 -2403 -1999
rect -2337 -1965 -2245 -1959
rect -2337 -1999 -2325 -1965
rect -2257 -1999 -2245 -1965
rect -2337 -2005 -2245 -1999
rect -2179 -1965 -2087 -1959
rect -2179 -1999 -2167 -1965
rect -2099 -1999 -2087 -1965
rect -2179 -2005 -2087 -1999
rect -2021 -1965 -1929 -1959
rect -2021 -1999 -2009 -1965
rect -1941 -1999 -1929 -1965
rect -2021 -2005 -1929 -1999
rect -1863 -1965 -1771 -1959
rect -1863 -1999 -1851 -1965
rect -1783 -1999 -1771 -1965
rect -1863 -2005 -1771 -1999
rect -1705 -1965 -1613 -1959
rect -1705 -1999 -1693 -1965
rect -1625 -1999 -1613 -1965
rect -1705 -2005 -1613 -1999
rect -1547 -1965 -1455 -1959
rect -1547 -1999 -1535 -1965
rect -1467 -1999 -1455 -1965
rect -1547 -2005 -1455 -1999
rect -1389 -1965 -1297 -1959
rect -1389 -1999 -1377 -1965
rect -1309 -1999 -1297 -1965
rect -1389 -2005 -1297 -1999
rect -1231 -1965 -1139 -1959
rect -1231 -1999 -1219 -1965
rect -1151 -1999 -1139 -1965
rect -1231 -2005 -1139 -1999
rect -1073 -1965 -981 -1959
rect -1073 -1999 -1061 -1965
rect -993 -1999 -981 -1965
rect -1073 -2005 -981 -1999
rect -915 -1965 -823 -1959
rect -915 -1999 -903 -1965
rect -835 -1999 -823 -1965
rect -915 -2005 -823 -1999
rect -757 -1965 -665 -1959
rect -757 -1999 -745 -1965
rect -677 -1999 -665 -1965
rect -757 -2005 -665 -1999
rect -599 -1965 -507 -1959
rect -599 -1999 -587 -1965
rect -519 -1999 -507 -1965
rect -599 -2005 -507 -1999
rect -441 -1965 -349 -1959
rect -441 -1999 -429 -1965
rect -361 -1999 -349 -1965
rect -441 -2005 -349 -1999
rect -283 -1965 -191 -1959
rect -283 -1999 -271 -1965
rect -203 -1999 -191 -1965
rect -283 -2005 -191 -1999
rect -125 -1965 -33 -1959
rect -125 -1999 -113 -1965
rect -45 -1999 -33 -1965
rect -125 -2005 -33 -1999
rect 33 -1965 125 -1959
rect 33 -1999 45 -1965
rect 113 -1999 125 -1965
rect 33 -2005 125 -1999
rect 191 -1965 283 -1959
rect 191 -1999 203 -1965
rect 271 -1999 283 -1965
rect 191 -2005 283 -1999
rect 349 -1965 441 -1959
rect 349 -1999 361 -1965
rect 429 -1999 441 -1965
rect 349 -2005 441 -1999
rect 507 -1965 599 -1959
rect 507 -1999 519 -1965
rect 587 -1999 599 -1965
rect 507 -2005 599 -1999
rect 665 -1965 757 -1959
rect 665 -1999 677 -1965
rect 745 -1999 757 -1965
rect 665 -2005 757 -1999
rect 823 -1965 915 -1959
rect 823 -1999 835 -1965
rect 903 -1999 915 -1965
rect 823 -2005 915 -1999
rect 981 -1965 1073 -1959
rect 981 -1999 993 -1965
rect 1061 -1999 1073 -1965
rect 981 -2005 1073 -1999
rect 1139 -1965 1231 -1959
rect 1139 -1999 1151 -1965
rect 1219 -1999 1231 -1965
rect 1139 -2005 1231 -1999
rect 1297 -1965 1389 -1959
rect 1297 -1999 1309 -1965
rect 1377 -1999 1389 -1965
rect 1297 -2005 1389 -1999
rect 1455 -1965 1547 -1959
rect 1455 -1999 1467 -1965
rect 1535 -1999 1547 -1965
rect 1455 -2005 1547 -1999
rect 1613 -1965 1705 -1959
rect 1613 -1999 1625 -1965
rect 1693 -1999 1705 -1965
rect 1613 -2005 1705 -1999
rect 1771 -1965 1863 -1959
rect 1771 -1999 1783 -1965
rect 1851 -1999 1863 -1965
rect 1771 -2005 1863 -1999
rect 1929 -1965 2021 -1959
rect 1929 -1999 1941 -1965
rect 2009 -1999 2021 -1965
rect 1929 -2005 2021 -1999
rect 2087 -1965 2179 -1959
rect 2087 -1999 2099 -1965
rect 2167 -1999 2179 -1965
rect 2087 -2005 2179 -1999
rect 2245 -1965 2337 -1959
rect 2245 -1999 2257 -1965
rect 2325 -1999 2337 -1965
rect 2245 -2005 2337 -1999
rect 2403 -1965 2495 -1959
rect 2403 -1999 2415 -1965
rect 2483 -1999 2495 -1965
rect 2403 -2005 2495 -1999
<< properties >>
string FIXED_BBOX -2662 -2120 2662 2120
string gencell sky130_fd_pr__nfet_03v3_nvt
string library sky130
string parameters w 4 l 0.50 m 4 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
