magic
tech sky130B
magscale 1 2
timestamp 1659896076
<< nwell >>
rect 1941 2141 5343 3651
<< pmos >>
rect 2137 3232 2197 3432
rect 2255 3232 2315 3432
rect 2373 3232 2433 3432
rect 2491 3232 2551 3432
rect 2609 3232 2669 3432
rect 2727 3232 2787 3432
rect 2845 3232 2905 3432
rect 2963 3232 3023 3432
rect 3081 3232 3141 3432
rect 3199 3232 3259 3432
rect 3317 3232 3377 3432
rect 3435 3232 3495 3432
rect 3553 3232 3613 3432
rect 3671 3232 3731 3432
rect 3789 3232 3849 3432
rect 3907 3232 3967 3432
rect 4025 3232 4085 3432
rect 4143 3232 4203 3432
rect 4261 3232 4321 3432
rect 4379 3232 4439 3432
rect 4497 3232 4557 3432
rect 4615 3232 4675 3432
rect 4733 3232 4793 3432
rect 4851 3232 4911 3432
rect 4969 3232 5029 3432
rect 5087 3232 5147 3432
rect 2137 2796 2197 2996
rect 2255 2796 2315 2996
rect 2373 2796 2433 2996
rect 2491 2796 2551 2996
rect 2609 2796 2669 2996
rect 2727 2796 2787 2996
rect 2845 2796 2905 2996
rect 2963 2796 3023 2996
rect 3081 2796 3141 2996
rect 3199 2796 3259 2996
rect 3317 2796 3377 2996
rect 3435 2796 3495 2996
rect 3553 2796 3613 2996
rect 3671 2796 3731 2996
rect 3789 2796 3849 2996
rect 3907 2796 3967 2996
rect 4025 2796 4085 2996
rect 4143 2796 4203 2996
rect 4261 2796 4321 2996
rect 4379 2796 4439 2996
rect 4497 2796 4557 2996
rect 4615 2796 4675 2996
rect 4733 2796 4793 2996
rect 4851 2796 4911 2996
rect 4969 2796 5029 2996
rect 5087 2796 5147 2996
rect 2137 2360 2197 2560
rect 2255 2360 2315 2560
rect 2373 2360 2433 2560
rect 2491 2360 2551 2560
rect 2609 2360 2669 2560
rect 2727 2360 2787 2560
rect 2845 2360 2905 2560
rect 2963 2360 3023 2560
rect 3081 2360 3141 2560
rect 3199 2360 3259 2560
rect 3317 2360 3377 2560
rect 3435 2360 3495 2560
rect 3553 2360 3613 2560
rect 3671 2360 3731 2560
rect 3789 2360 3849 2560
rect 3907 2360 3967 2560
rect 4025 2360 4085 2560
rect 4143 2360 4203 2560
rect 4261 2360 4321 2560
rect 4379 2360 4439 2560
rect 4497 2360 4557 2560
rect 4615 2360 4675 2560
rect 4733 2360 4793 2560
rect 4851 2360 4911 2560
rect 4969 2360 5029 2560
rect 5087 2360 5147 2560
<< pdiff >>
rect 2079 3420 2137 3432
rect 2079 3244 2091 3420
rect 2125 3244 2137 3420
rect 2079 3232 2137 3244
rect 2197 3420 2255 3432
rect 2197 3244 2209 3420
rect 2243 3244 2255 3420
rect 2197 3232 2255 3244
rect 2315 3420 2373 3432
rect 2315 3244 2327 3420
rect 2361 3244 2373 3420
rect 2315 3232 2373 3244
rect 2433 3420 2491 3432
rect 2433 3244 2445 3420
rect 2479 3244 2491 3420
rect 2433 3232 2491 3244
rect 2551 3420 2609 3432
rect 2551 3244 2563 3420
rect 2597 3244 2609 3420
rect 2551 3232 2609 3244
rect 2669 3420 2727 3432
rect 2669 3244 2681 3420
rect 2715 3244 2727 3420
rect 2669 3232 2727 3244
rect 2787 3420 2845 3432
rect 2787 3244 2799 3420
rect 2833 3244 2845 3420
rect 2787 3232 2845 3244
rect 2905 3420 2963 3432
rect 2905 3244 2917 3420
rect 2951 3244 2963 3420
rect 2905 3232 2963 3244
rect 3023 3420 3081 3432
rect 3023 3244 3035 3420
rect 3069 3244 3081 3420
rect 3023 3232 3081 3244
rect 3141 3420 3199 3432
rect 3141 3244 3153 3420
rect 3187 3244 3199 3420
rect 3141 3232 3199 3244
rect 3259 3420 3317 3432
rect 3259 3244 3271 3420
rect 3305 3244 3317 3420
rect 3259 3232 3317 3244
rect 3377 3420 3435 3432
rect 3377 3244 3389 3420
rect 3423 3244 3435 3420
rect 3377 3232 3435 3244
rect 3495 3420 3553 3432
rect 3495 3244 3507 3420
rect 3541 3244 3553 3420
rect 3495 3232 3553 3244
rect 3613 3420 3671 3432
rect 3613 3244 3625 3420
rect 3659 3244 3671 3420
rect 3613 3232 3671 3244
rect 3731 3420 3789 3432
rect 3731 3244 3743 3420
rect 3777 3244 3789 3420
rect 3731 3232 3789 3244
rect 3849 3420 3907 3432
rect 3849 3244 3861 3420
rect 3895 3244 3907 3420
rect 3849 3232 3907 3244
rect 3967 3420 4025 3432
rect 3967 3244 3979 3420
rect 4013 3244 4025 3420
rect 3967 3232 4025 3244
rect 4085 3420 4143 3432
rect 4085 3244 4097 3420
rect 4131 3244 4143 3420
rect 4085 3232 4143 3244
rect 4203 3420 4261 3432
rect 4203 3244 4215 3420
rect 4249 3244 4261 3420
rect 4203 3232 4261 3244
rect 4321 3420 4379 3432
rect 4321 3244 4333 3420
rect 4367 3244 4379 3420
rect 4321 3232 4379 3244
rect 4439 3420 4497 3432
rect 4439 3244 4451 3420
rect 4485 3244 4497 3420
rect 4439 3232 4497 3244
rect 4557 3420 4615 3432
rect 4557 3244 4569 3420
rect 4603 3244 4615 3420
rect 4557 3232 4615 3244
rect 4675 3420 4733 3432
rect 4675 3244 4687 3420
rect 4721 3244 4733 3420
rect 4675 3232 4733 3244
rect 4793 3420 4851 3432
rect 4793 3244 4805 3420
rect 4839 3244 4851 3420
rect 4793 3232 4851 3244
rect 4911 3420 4969 3432
rect 4911 3244 4923 3420
rect 4957 3244 4969 3420
rect 4911 3232 4969 3244
rect 5029 3420 5087 3432
rect 5029 3244 5041 3420
rect 5075 3244 5087 3420
rect 5029 3232 5087 3244
rect 5147 3420 5205 3432
rect 5147 3244 5159 3420
rect 5193 3244 5205 3420
rect 5147 3232 5205 3244
rect 2079 2984 2137 2996
rect 2079 2808 2091 2984
rect 2125 2808 2137 2984
rect 2079 2796 2137 2808
rect 2197 2984 2255 2996
rect 2197 2808 2209 2984
rect 2243 2808 2255 2984
rect 2197 2796 2255 2808
rect 2315 2984 2373 2996
rect 2315 2808 2327 2984
rect 2361 2808 2373 2984
rect 2315 2796 2373 2808
rect 2433 2984 2491 2996
rect 2433 2808 2445 2984
rect 2479 2808 2491 2984
rect 2433 2796 2491 2808
rect 2551 2984 2609 2996
rect 2551 2808 2563 2984
rect 2597 2808 2609 2984
rect 2551 2796 2609 2808
rect 2669 2984 2727 2996
rect 2669 2808 2681 2984
rect 2715 2808 2727 2984
rect 2669 2796 2727 2808
rect 2787 2984 2845 2996
rect 2787 2808 2799 2984
rect 2833 2808 2845 2984
rect 2787 2796 2845 2808
rect 2905 2984 2963 2996
rect 2905 2808 2917 2984
rect 2951 2808 2963 2984
rect 2905 2796 2963 2808
rect 3023 2984 3081 2996
rect 3023 2808 3035 2984
rect 3069 2808 3081 2984
rect 3023 2796 3081 2808
rect 3141 2984 3199 2996
rect 3141 2808 3153 2984
rect 3187 2808 3199 2984
rect 3141 2796 3199 2808
rect 3259 2984 3317 2996
rect 3259 2808 3271 2984
rect 3305 2808 3317 2984
rect 3259 2796 3317 2808
rect 3377 2984 3435 2996
rect 3377 2808 3389 2984
rect 3423 2808 3435 2984
rect 3377 2796 3435 2808
rect 3495 2984 3553 2996
rect 3495 2808 3507 2984
rect 3541 2808 3553 2984
rect 3495 2796 3553 2808
rect 3613 2984 3671 2996
rect 3613 2808 3625 2984
rect 3659 2808 3671 2984
rect 3613 2796 3671 2808
rect 3731 2984 3789 2996
rect 3731 2808 3743 2984
rect 3777 2808 3789 2984
rect 3731 2796 3789 2808
rect 3849 2984 3907 2996
rect 3849 2808 3861 2984
rect 3895 2808 3907 2984
rect 3849 2796 3907 2808
rect 3967 2984 4025 2996
rect 3967 2808 3979 2984
rect 4013 2808 4025 2984
rect 3967 2796 4025 2808
rect 4085 2984 4143 2996
rect 4085 2808 4097 2984
rect 4131 2808 4143 2984
rect 4085 2796 4143 2808
rect 4203 2984 4261 2996
rect 4203 2808 4215 2984
rect 4249 2808 4261 2984
rect 4203 2796 4261 2808
rect 4321 2984 4379 2996
rect 4321 2808 4333 2984
rect 4367 2808 4379 2984
rect 4321 2796 4379 2808
rect 4439 2984 4497 2996
rect 4439 2808 4451 2984
rect 4485 2808 4497 2984
rect 4439 2796 4497 2808
rect 4557 2984 4615 2996
rect 4557 2808 4569 2984
rect 4603 2808 4615 2984
rect 4557 2796 4615 2808
rect 4675 2984 4733 2996
rect 4675 2808 4687 2984
rect 4721 2808 4733 2984
rect 4675 2796 4733 2808
rect 4793 2984 4851 2996
rect 4793 2808 4805 2984
rect 4839 2808 4851 2984
rect 4793 2796 4851 2808
rect 4911 2984 4969 2996
rect 4911 2808 4923 2984
rect 4957 2808 4969 2984
rect 4911 2796 4969 2808
rect 5029 2984 5087 2996
rect 5029 2808 5041 2984
rect 5075 2808 5087 2984
rect 5029 2796 5087 2808
rect 5147 2984 5205 2996
rect 5147 2808 5159 2984
rect 5193 2808 5205 2984
rect 5147 2796 5205 2808
rect 2079 2548 2137 2560
rect 2079 2372 2091 2548
rect 2125 2372 2137 2548
rect 2079 2360 2137 2372
rect 2197 2548 2255 2560
rect 2197 2372 2209 2548
rect 2243 2372 2255 2548
rect 2197 2360 2255 2372
rect 2315 2548 2373 2560
rect 2315 2372 2327 2548
rect 2361 2372 2373 2548
rect 2315 2360 2373 2372
rect 2433 2548 2491 2560
rect 2433 2372 2445 2548
rect 2479 2372 2491 2548
rect 2433 2360 2491 2372
rect 2551 2548 2609 2560
rect 2551 2372 2563 2548
rect 2597 2372 2609 2548
rect 2551 2360 2609 2372
rect 2669 2548 2727 2560
rect 2669 2372 2681 2548
rect 2715 2372 2727 2548
rect 2669 2360 2727 2372
rect 2787 2548 2845 2560
rect 2787 2372 2799 2548
rect 2833 2372 2845 2548
rect 2787 2360 2845 2372
rect 2905 2548 2963 2560
rect 2905 2372 2917 2548
rect 2951 2372 2963 2548
rect 2905 2360 2963 2372
rect 3023 2548 3081 2560
rect 3023 2372 3035 2548
rect 3069 2372 3081 2548
rect 3023 2360 3081 2372
rect 3141 2548 3199 2560
rect 3141 2372 3153 2548
rect 3187 2372 3199 2548
rect 3141 2360 3199 2372
rect 3259 2548 3317 2560
rect 3259 2372 3271 2548
rect 3305 2372 3317 2548
rect 3259 2360 3317 2372
rect 3377 2548 3435 2560
rect 3377 2372 3389 2548
rect 3423 2372 3435 2548
rect 3377 2360 3435 2372
rect 3495 2548 3553 2560
rect 3495 2372 3507 2548
rect 3541 2372 3553 2548
rect 3495 2360 3553 2372
rect 3613 2548 3671 2560
rect 3613 2372 3625 2548
rect 3659 2372 3671 2548
rect 3613 2360 3671 2372
rect 3731 2548 3789 2560
rect 3731 2372 3743 2548
rect 3777 2372 3789 2548
rect 3731 2360 3789 2372
rect 3849 2548 3907 2560
rect 3849 2372 3861 2548
rect 3895 2372 3907 2548
rect 3849 2360 3907 2372
rect 3967 2548 4025 2560
rect 3967 2372 3979 2548
rect 4013 2372 4025 2548
rect 3967 2360 4025 2372
rect 4085 2548 4143 2560
rect 4085 2372 4097 2548
rect 4131 2372 4143 2548
rect 4085 2360 4143 2372
rect 4203 2548 4261 2560
rect 4203 2372 4215 2548
rect 4249 2372 4261 2548
rect 4203 2360 4261 2372
rect 4321 2548 4379 2560
rect 4321 2372 4333 2548
rect 4367 2372 4379 2548
rect 4321 2360 4379 2372
rect 4439 2548 4497 2560
rect 4439 2372 4451 2548
rect 4485 2372 4497 2548
rect 4439 2360 4497 2372
rect 4557 2548 4615 2560
rect 4557 2372 4569 2548
rect 4603 2372 4615 2548
rect 4557 2360 4615 2372
rect 4675 2548 4733 2560
rect 4675 2372 4687 2548
rect 4721 2372 4733 2548
rect 4675 2360 4733 2372
rect 4793 2548 4851 2560
rect 4793 2372 4805 2548
rect 4839 2372 4851 2548
rect 4793 2360 4851 2372
rect 4911 2548 4969 2560
rect 4911 2372 4923 2548
rect 4957 2372 4969 2548
rect 4911 2360 4969 2372
rect 5029 2548 5087 2560
rect 5029 2372 5041 2548
rect 5075 2372 5087 2548
rect 5029 2360 5087 2372
rect 5147 2548 5205 2560
rect 5147 2372 5159 2548
rect 5193 2372 5205 2548
rect 5147 2360 5205 2372
<< pdiffc >>
rect 2091 3244 2125 3420
rect 2209 3244 2243 3420
rect 2327 3244 2361 3420
rect 2445 3244 2479 3420
rect 2563 3244 2597 3420
rect 2681 3244 2715 3420
rect 2799 3244 2833 3420
rect 2917 3244 2951 3420
rect 3035 3244 3069 3420
rect 3153 3244 3187 3420
rect 3271 3244 3305 3420
rect 3389 3244 3423 3420
rect 3507 3244 3541 3420
rect 3625 3244 3659 3420
rect 3743 3244 3777 3420
rect 3861 3244 3895 3420
rect 3979 3244 4013 3420
rect 4097 3244 4131 3420
rect 4215 3244 4249 3420
rect 4333 3244 4367 3420
rect 4451 3244 4485 3420
rect 4569 3244 4603 3420
rect 4687 3244 4721 3420
rect 4805 3244 4839 3420
rect 4923 3244 4957 3420
rect 5041 3244 5075 3420
rect 5159 3244 5193 3420
rect 2091 2808 2125 2984
rect 2209 2808 2243 2984
rect 2327 2808 2361 2984
rect 2445 2808 2479 2984
rect 2563 2808 2597 2984
rect 2681 2808 2715 2984
rect 2799 2808 2833 2984
rect 2917 2808 2951 2984
rect 3035 2808 3069 2984
rect 3153 2808 3187 2984
rect 3271 2808 3305 2984
rect 3389 2808 3423 2984
rect 3507 2808 3541 2984
rect 3625 2808 3659 2984
rect 3743 2808 3777 2984
rect 3861 2808 3895 2984
rect 3979 2808 4013 2984
rect 4097 2808 4131 2984
rect 4215 2808 4249 2984
rect 4333 2808 4367 2984
rect 4451 2808 4485 2984
rect 4569 2808 4603 2984
rect 4687 2808 4721 2984
rect 4805 2808 4839 2984
rect 4923 2808 4957 2984
rect 5041 2808 5075 2984
rect 5159 2808 5193 2984
rect 2091 2372 2125 2548
rect 2209 2372 2243 2548
rect 2327 2372 2361 2548
rect 2445 2372 2479 2548
rect 2563 2372 2597 2548
rect 2681 2372 2715 2548
rect 2799 2372 2833 2548
rect 2917 2372 2951 2548
rect 3035 2372 3069 2548
rect 3153 2372 3187 2548
rect 3271 2372 3305 2548
rect 3389 2372 3423 2548
rect 3507 2372 3541 2548
rect 3625 2372 3659 2548
rect 3743 2372 3777 2548
rect 3861 2372 3895 2548
rect 3979 2372 4013 2548
rect 4097 2372 4131 2548
rect 4215 2372 4249 2548
rect 4333 2372 4367 2548
rect 4451 2372 4485 2548
rect 4569 2372 4603 2548
rect 4687 2372 4721 2548
rect 4805 2372 4839 2548
rect 4923 2372 4957 2548
rect 5041 2372 5075 2548
rect 5159 2372 5193 2548
<< nsubdiff >>
rect 1977 3581 2073 3615
rect 5211 3581 5307 3615
rect 1977 3519 2011 3581
rect 5273 3519 5307 3581
rect 1977 2211 2011 2273
rect 5273 2211 5307 2273
rect 1977 2177 2073 2211
rect 5211 2177 5307 2211
<< nsubdiffcont >>
rect 2073 3581 5211 3615
rect 1977 2273 2011 3519
rect 5273 2273 5307 3519
rect 2073 2177 5211 2211
<< poly >>
rect 2134 3513 2200 3529
rect 2134 3479 2150 3513
rect 2184 3479 2200 3513
rect 2134 3463 2200 3479
rect 2252 3513 2318 3529
rect 2252 3479 2268 3513
rect 2302 3479 2318 3513
rect 2252 3463 2318 3479
rect 2370 3513 2436 3529
rect 2370 3479 2386 3513
rect 2420 3479 2436 3513
rect 2370 3463 2436 3479
rect 2488 3513 2554 3529
rect 2488 3479 2504 3513
rect 2538 3479 2554 3513
rect 2488 3463 2554 3479
rect 2606 3513 2672 3529
rect 2606 3479 2622 3513
rect 2656 3479 2672 3513
rect 2606 3463 2672 3479
rect 2724 3513 2790 3529
rect 2724 3479 2740 3513
rect 2774 3479 2790 3513
rect 2724 3463 2790 3479
rect 2842 3513 2908 3529
rect 2842 3479 2858 3513
rect 2892 3479 2908 3513
rect 2842 3463 2908 3479
rect 2960 3513 3026 3529
rect 2960 3479 2976 3513
rect 3010 3479 3026 3513
rect 2960 3463 3026 3479
rect 3078 3513 3144 3529
rect 3078 3479 3094 3513
rect 3128 3479 3144 3513
rect 3078 3463 3144 3479
rect 3196 3513 3262 3529
rect 3196 3479 3212 3513
rect 3246 3479 3262 3513
rect 3196 3463 3262 3479
rect 3314 3513 3380 3529
rect 3314 3479 3330 3513
rect 3364 3479 3380 3513
rect 3314 3463 3380 3479
rect 3432 3513 3498 3529
rect 3432 3479 3448 3513
rect 3482 3479 3498 3513
rect 3432 3463 3498 3479
rect 3550 3513 3616 3529
rect 3550 3479 3566 3513
rect 3600 3479 3616 3513
rect 3550 3463 3616 3479
rect 3668 3513 3734 3529
rect 3668 3479 3684 3513
rect 3718 3479 3734 3513
rect 3668 3463 3734 3479
rect 3786 3513 3852 3529
rect 3786 3479 3802 3513
rect 3836 3479 3852 3513
rect 3786 3463 3852 3479
rect 3904 3513 3970 3529
rect 3904 3479 3920 3513
rect 3954 3479 3970 3513
rect 3904 3463 3970 3479
rect 4022 3513 4088 3529
rect 4022 3479 4038 3513
rect 4072 3479 4088 3513
rect 4022 3463 4088 3479
rect 4140 3513 4206 3529
rect 4140 3479 4156 3513
rect 4190 3479 4206 3513
rect 4140 3463 4206 3479
rect 4258 3513 4324 3529
rect 4258 3479 4274 3513
rect 4308 3479 4324 3513
rect 4258 3463 4324 3479
rect 4376 3513 4442 3529
rect 4376 3479 4392 3513
rect 4426 3479 4442 3513
rect 4376 3463 4442 3479
rect 4494 3513 4560 3529
rect 4494 3479 4510 3513
rect 4544 3479 4560 3513
rect 4494 3463 4560 3479
rect 4612 3513 4678 3529
rect 4612 3479 4628 3513
rect 4662 3479 4678 3513
rect 4612 3463 4678 3479
rect 4730 3513 4796 3529
rect 4730 3479 4746 3513
rect 4780 3479 4796 3513
rect 4730 3463 4796 3479
rect 4848 3513 4914 3529
rect 4848 3479 4864 3513
rect 4898 3479 4914 3513
rect 4848 3463 4914 3479
rect 4966 3513 5032 3529
rect 4966 3479 4982 3513
rect 5016 3479 5032 3513
rect 4966 3463 5032 3479
rect 5084 3513 5150 3529
rect 5084 3479 5100 3513
rect 5134 3479 5150 3513
rect 5084 3463 5150 3479
rect 2137 3432 2197 3463
rect 2255 3432 2315 3463
rect 2373 3432 2433 3463
rect 2491 3432 2551 3463
rect 2609 3432 2669 3463
rect 2727 3432 2787 3463
rect 2845 3432 2905 3463
rect 2963 3432 3023 3463
rect 3081 3432 3141 3463
rect 3199 3432 3259 3463
rect 3317 3432 3377 3463
rect 3435 3432 3495 3463
rect 3553 3432 3613 3463
rect 3671 3432 3731 3463
rect 3789 3432 3849 3463
rect 3907 3432 3967 3463
rect 4025 3432 4085 3463
rect 4143 3432 4203 3463
rect 4261 3432 4321 3463
rect 4379 3432 4439 3463
rect 4497 3432 4557 3463
rect 4615 3432 4675 3463
rect 4733 3432 4793 3463
rect 4851 3432 4911 3463
rect 4969 3432 5029 3463
rect 5087 3432 5147 3463
rect 2137 3201 2197 3232
rect 2255 3201 2315 3232
rect 2373 3201 2433 3232
rect 2491 3201 2551 3232
rect 2609 3201 2669 3232
rect 2727 3201 2787 3232
rect 2845 3201 2905 3232
rect 2963 3201 3023 3232
rect 3081 3201 3141 3232
rect 3199 3201 3259 3232
rect 3317 3201 3377 3232
rect 3435 3201 3495 3232
rect 3553 3201 3613 3232
rect 3671 3201 3731 3232
rect 3789 3201 3849 3232
rect 3907 3201 3967 3232
rect 4025 3201 4085 3232
rect 4143 3201 4203 3232
rect 4261 3201 4321 3232
rect 4379 3201 4439 3232
rect 4497 3201 4557 3232
rect 4615 3201 4675 3232
rect 4733 3201 4793 3232
rect 4851 3201 4911 3232
rect 4969 3201 5029 3232
rect 5087 3201 5147 3232
rect 3786 3077 3852 3093
rect 3786 3043 3802 3077
rect 3836 3043 3852 3077
rect 3786 3027 3852 3043
rect 2137 2996 2197 3027
rect 2255 2996 2315 3027
rect 2373 2996 2433 3027
rect 2491 2996 2551 3027
rect 2609 2996 2669 3027
rect 2727 2996 2787 3027
rect 2845 2996 2905 3027
rect 2963 2996 3023 3027
rect 3081 2996 3141 3027
rect 3199 2996 3259 3027
rect 3317 2996 3377 3027
rect 3435 2996 3495 3027
rect 3553 2996 3613 3027
rect 3671 2996 3731 3027
rect 3789 2996 3849 3027
rect 3907 2996 3967 3027
rect 4025 2996 4085 3027
rect 4143 2996 4203 3027
rect 4261 2996 4321 3027
rect 4379 2996 4439 3027
rect 4497 2996 4557 3027
rect 4615 2996 4675 3027
rect 4733 2996 4793 3027
rect 4851 2996 4911 3027
rect 4969 2996 5029 3027
rect 5087 2996 5147 3027
rect 2137 2765 2197 2796
rect 2255 2765 2315 2796
rect 2373 2765 2433 2796
rect 2491 2765 2551 2796
rect 2609 2765 2669 2796
rect 2727 2765 2787 2796
rect 2845 2765 2905 2796
rect 2963 2765 3023 2796
rect 3081 2765 3141 2796
rect 3199 2765 3259 2796
rect 3317 2765 3377 2796
rect 3435 2765 3495 2796
rect 3553 2765 3613 2796
rect 3671 2765 3731 2796
rect 3789 2770 3849 2796
rect 3907 2765 3967 2796
rect 4025 2765 4085 2796
rect 4143 2765 4203 2796
rect 4261 2765 4321 2796
rect 4379 2765 4439 2796
rect 4497 2765 4557 2796
rect 4615 2765 4675 2796
rect 4733 2765 4793 2796
rect 4851 2765 4911 2796
rect 4969 2765 5029 2796
rect 5087 2765 5147 2796
rect 2134 2749 2200 2765
rect 2134 2715 2150 2749
rect 2184 2715 2200 2749
rect 2134 2699 2200 2715
rect 2252 2749 2318 2765
rect 2252 2715 2268 2749
rect 2302 2715 2318 2749
rect 2252 2699 2318 2715
rect 2370 2749 2436 2765
rect 2370 2715 2386 2749
rect 2420 2715 2436 2749
rect 2370 2699 2436 2715
rect 2488 2749 2554 2765
rect 2488 2715 2504 2749
rect 2538 2715 2554 2749
rect 2488 2699 2554 2715
rect 2606 2749 2672 2765
rect 2606 2715 2622 2749
rect 2656 2715 2672 2749
rect 2606 2699 2672 2715
rect 2724 2749 2790 2765
rect 2724 2715 2740 2749
rect 2774 2715 2790 2749
rect 2724 2699 2790 2715
rect 2842 2749 2908 2765
rect 2842 2715 2858 2749
rect 2892 2715 2908 2749
rect 2842 2699 2908 2715
rect 2960 2749 3026 2765
rect 2960 2715 2976 2749
rect 3010 2715 3026 2749
rect 2960 2699 3026 2715
rect 3078 2749 3144 2765
rect 3078 2715 3094 2749
rect 3128 2715 3144 2749
rect 3078 2699 3144 2715
rect 3196 2749 3262 2765
rect 3196 2715 3212 2749
rect 3246 2715 3262 2749
rect 3196 2699 3262 2715
rect 3314 2749 3380 2765
rect 3314 2715 3330 2749
rect 3364 2715 3380 2749
rect 3314 2699 3380 2715
rect 3432 2749 3498 2765
rect 3432 2715 3448 2749
rect 3482 2715 3498 2749
rect 3432 2699 3498 2715
rect 3550 2749 3616 2765
rect 3550 2715 3566 2749
rect 3600 2715 3616 2749
rect 3550 2699 3616 2715
rect 3668 2749 3734 2765
rect 3668 2715 3684 2749
rect 3718 2715 3734 2749
rect 3668 2699 3734 2715
rect 3904 2749 3970 2765
rect 3904 2715 3920 2749
rect 3954 2715 3970 2749
rect 3904 2699 3970 2715
rect 4022 2749 4088 2765
rect 4022 2715 4038 2749
rect 4072 2715 4088 2749
rect 4022 2699 4088 2715
rect 4140 2749 4206 2765
rect 4140 2715 4156 2749
rect 4190 2715 4206 2749
rect 4140 2699 4206 2715
rect 4258 2749 4324 2765
rect 4258 2715 4274 2749
rect 4308 2715 4324 2749
rect 4258 2699 4324 2715
rect 4376 2749 4442 2765
rect 4376 2715 4392 2749
rect 4426 2715 4442 2749
rect 4376 2699 4442 2715
rect 4494 2749 4560 2765
rect 4494 2715 4510 2749
rect 4544 2715 4560 2749
rect 4494 2699 4560 2715
rect 4612 2749 4678 2765
rect 4612 2715 4628 2749
rect 4662 2715 4678 2749
rect 4612 2699 4678 2715
rect 4730 2749 4796 2765
rect 4730 2715 4746 2749
rect 4780 2715 4796 2749
rect 4730 2699 4796 2715
rect 4848 2749 4914 2765
rect 4848 2715 4864 2749
rect 4898 2715 4914 2749
rect 4848 2699 4914 2715
rect 4966 2749 5032 2765
rect 4966 2715 4982 2749
rect 5016 2715 5032 2749
rect 4966 2699 5032 2715
rect 5084 2749 5150 2765
rect 5084 2715 5100 2749
rect 5134 2715 5150 2749
rect 5084 2699 5150 2715
rect 2137 2560 2197 2591
rect 2255 2560 2315 2591
rect 2373 2560 2433 2591
rect 2491 2560 2551 2591
rect 2609 2560 2669 2591
rect 2727 2560 2787 2591
rect 2845 2560 2905 2591
rect 2963 2560 3023 2591
rect 3081 2560 3141 2591
rect 3199 2560 3259 2591
rect 3317 2560 3377 2591
rect 3435 2560 3495 2591
rect 3553 2560 3613 2591
rect 3671 2560 3731 2591
rect 3789 2560 3849 2591
rect 3907 2560 3967 2591
rect 4025 2560 4085 2591
rect 4143 2560 4203 2591
rect 4261 2560 4321 2591
rect 4379 2560 4439 2591
rect 4497 2560 4557 2591
rect 4615 2560 4675 2591
rect 4733 2560 4793 2591
rect 4851 2560 4911 2591
rect 4969 2560 5029 2591
rect 5087 2560 5147 2591
rect 2137 2329 2197 2360
rect 2255 2329 2315 2360
rect 2373 2329 2433 2360
rect 2491 2329 2551 2360
rect 2609 2329 2669 2360
rect 2727 2329 2787 2360
rect 2845 2329 2905 2360
rect 2963 2329 3023 2360
rect 3081 2329 3141 2360
rect 3199 2329 3259 2360
rect 3317 2329 3377 2360
rect 3435 2329 3495 2360
rect 3553 2329 3613 2360
rect 3671 2329 3731 2360
rect 3789 2329 3849 2360
rect 3907 2329 3967 2360
rect 4025 2329 4085 2360
rect 4143 2329 4203 2360
rect 4261 2329 4321 2360
rect 4379 2329 4439 2360
rect 4497 2329 4557 2360
rect 4615 2329 4675 2360
rect 4733 2329 4793 2360
rect 4851 2329 4911 2360
rect 4969 2329 5029 2360
rect 5087 2329 5147 2360
rect 2134 2313 2200 2329
rect 2134 2279 2150 2313
rect 2184 2279 2200 2313
rect 2134 2263 2200 2279
rect 2252 2313 2318 2329
rect 2252 2279 2268 2313
rect 2302 2279 2318 2313
rect 2252 2263 2318 2279
rect 2370 2313 2436 2329
rect 2370 2279 2386 2313
rect 2420 2279 2436 2313
rect 2370 2263 2436 2279
rect 2488 2313 2554 2329
rect 2488 2279 2504 2313
rect 2538 2279 2554 2313
rect 2488 2263 2554 2279
rect 2606 2313 2672 2329
rect 2606 2279 2622 2313
rect 2656 2279 2672 2313
rect 2606 2263 2672 2279
rect 2724 2313 2790 2329
rect 2724 2279 2740 2313
rect 2774 2279 2790 2313
rect 2724 2263 2790 2279
rect 2842 2313 2908 2329
rect 2842 2279 2858 2313
rect 2892 2279 2908 2313
rect 2842 2263 2908 2279
rect 2960 2313 3026 2329
rect 2960 2279 2976 2313
rect 3010 2279 3026 2313
rect 2960 2263 3026 2279
rect 3078 2313 3144 2329
rect 3078 2279 3094 2313
rect 3128 2279 3144 2313
rect 3078 2263 3144 2279
rect 3196 2313 3262 2329
rect 3196 2279 3212 2313
rect 3246 2279 3262 2313
rect 3196 2263 3262 2279
rect 3314 2313 3380 2329
rect 3314 2279 3330 2313
rect 3364 2279 3380 2313
rect 3314 2263 3380 2279
rect 3432 2313 3498 2329
rect 3432 2279 3448 2313
rect 3482 2279 3498 2313
rect 3432 2263 3498 2279
rect 3550 2313 3616 2329
rect 3550 2279 3566 2313
rect 3600 2279 3616 2313
rect 3550 2263 3616 2279
rect 3668 2313 3734 2329
rect 3668 2279 3684 2313
rect 3718 2279 3734 2313
rect 3668 2263 3734 2279
rect 3786 2313 3852 2329
rect 3786 2279 3802 2313
rect 3836 2279 3852 2313
rect 3786 2263 3852 2279
rect 3904 2313 3970 2329
rect 3904 2279 3920 2313
rect 3954 2279 3970 2313
rect 3904 2263 3970 2279
rect 4022 2313 4088 2329
rect 4022 2279 4038 2313
rect 4072 2279 4088 2313
rect 4022 2263 4088 2279
rect 4140 2313 4206 2329
rect 4140 2279 4156 2313
rect 4190 2279 4206 2313
rect 4140 2263 4206 2279
rect 4258 2313 4324 2329
rect 4258 2279 4274 2313
rect 4308 2279 4324 2313
rect 4258 2263 4324 2279
rect 4376 2313 4442 2329
rect 4376 2279 4392 2313
rect 4426 2279 4442 2313
rect 4376 2263 4442 2279
rect 4494 2313 4560 2329
rect 4494 2279 4510 2313
rect 4544 2279 4560 2313
rect 4494 2263 4560 2279
rect 4612 2313 4678 2329
rect 4612 2279 4628 2313
rect 4662 2279 4678 2313
rect 4612 2263 4678 2279
rect 4730 2313 4796 2329
rect 4730 2279 4746 2313
rect 4780 2279 4796 2313
rect 4730 2263 4796 2279
rect 4848 2313 4914 2329
rect 4848 2279 4864 2313
rect 4898 2279 4914 2313
rect 4848 2263 4914 2279
rect 4966 2313 5032 2329
rect 4966 2279 4982 2313
rect 5016 2279 5032 2313
rect 4966 2263 5032 2279
rect 5084 2313 5150 2329
rect 5084 2279 5100 2313
rect 5134 2279 5150 2313
rect 5084 2263 5150 2279
<< polycont >>
rect 2150 3479 2184 3513
rect 2268 3479 2302 3513
rect 2386 3479 2420 3513
rect 2504 3479 2538 3513
rect 2622 3479 2656 3513
rect 2740 3479 2774 3513
rect 2858 3479 2892 3513
rect 2976 3479 3010 3513
rect 3094 3479 3128 3513
rect 3212 3479 3246 3513
rect 3330 3479 3364 3513
rect 3448 3479 3482 3513
rect 3566 3479 3600 3513
rect 3684 3479 3718 3513
rect 3802 3479 3836 3513
rect 3920 3479 3954 3513
rect 4038 3479 4072 3513
rect 4156 3479 4190 3513
rect 4274 3479 4308 3513
rect 4392 3479 4426 3513
rect 4510 3479 4544 3513
rect 4628 3479 4662 3513
rect 4746 3479 4780 3513
rect 4864 3479 4898 3513
rect 4982 3479 5016 3513
rect 5100 3479 5134 3513
rect 3802 3043 3836 3077
rect 2150 2715 2184 2749
rect 2268 2715 2302 2749
rect 2386 2715 2420 2749
rect 2504 2715 2538 2749
rect 2622 2715 2656 2749
rect 2740 2715 2774 2749
rect 2858 2715 2892 2749
rect 2976 2715 3010 2749
rect 3094 2715 3128 2749
rect 3212 2715 3246 2749
rect 3330 2715 3364 2749
rect 3448 2715 3482 2749
rect 3566 2715 3600 2749
rect 3684 2715 3718 2749
rect 3920 2715 3954 2749
rect 4038 2715 4072 2749
rect 4156 2715 4190 2749
rect 4274 2715 4308 2749
rect 4392 2715 4426 2749
rect 4510 2715 4544 2749
rect 4628 2715 4662 2749
rect 4746 2715 4780 2749
rect 4864 2715 4898 2749
rect 4982 2715 5016 2749
rect 5100 2715 5134 2749
rect 2150 2279 2184 2313
rect 2268 2279 2302 2313
rect 2386 2279 2420 2313
rect 2504 2279 2538 2313
rect 2622 2279 2656 2313
rect 2740 2279 2774 2313
rect 2858 2279 2892 2313
rect 2976 2279 3010 2313
rect 3094 2279 3128 2313
rect 3212 2279 3246 2313
rect 3330 2279 3364 2313
rect 3448 2279 3482 2313
rect 3566 2279 3600 2313
rect 3684 2279 3718 2313
rect 3802 2279 3836 2313
rect 3920 2279 3954 2313
rect 4038 2279 4072 2313
rect 4156 2279 4190 2313
rect 4274 2279 4308 2313
rect 4392 2279 4426 2313
rect 4510 2279 4544 2313
rect 4628 2279 4662 2313
rect 4746 2279 4780 2313
rect 4864 2279 4898 2313
rect 4982 2279 5016 2313
rect 5100 2279 5134 2313
<< locali >>
rect 1977 3610 2073 3615
rect 1977 3519 1980 3610
rect 2014 3581 2073 3610
rect 5211 3610 5307 3615
rect 5211 3581 5280 3610
rect 5273 3519 5280 3581
rect 2134 3479 2150 3513
rect 2184 3479 2200 3513
rect 2252 3479 2268 3513
rect 2302 3479 2318 3513
rect 2370 3479 2386 3513
rect 2420 3479 2436 3513
rect 2488 3479 2504 3513
rect 2538 3479 2554 3513
rect 2606 3479 2622 3513
rect 2656 3479 2672 3513
rect 2724 3479 2740 3513
rect 2774 3479 2790 3513
rect 2842 3479 2858 3513
rect 2892 3479 2908 3513
rect 2960 3479 2976 3513
rect 3010 3479 3026 3513
rect 3078 3479 3094 3513
rect 3128 3479 3144 3513
rect 3196 3479 3212 3513
rect 3246 3479 3262 3513
rect 3314 3479 3330 3513
rect 3364 3479 3380 3513
rect 3432 3479 3448 3513
rect 3482 3479 3498 3513
rect 3550 3479 3566 3513
rect 3600 3479 3616 3513
rect 3668 3479 3684 3513
rect 3718 3479 3734 3513
rect 3786 3479 3802 3513
rect 3836 3479 3852 3513
rect 3904 3479 3920 3513
rect 3954 3479 3970 3513
rect 4022 3479 4038 3513
rect 4072 3479 4088 3513
rect 4140 3479 4156 3513
rect 4190 3479 4206 3513
rect 4258 3479 4274 3513
rect 4308 3479 4324 3513
rect 4376 3479 4392 3513
rect 4426 3479 4442 3513
rect 4494 3479 4510 3513
rect 4544 3479 4560 3513
rect 4612 3479 4628 3513
rect 4662 3479 4678 3513
rect 4730 3479 4746 3513
rect 4780 3479 4796 3513
rect 4848 3479 4864 3513
rect 4898 3479 4914 3513
rect 4966 3479 4982 3513
rect 5016 3479 5032 3513
rect 5084 3479 5100 3513
rect 5134 3479 5150 3513
rect 2091 3420 2125 3436
rect 2091 3228 2125 3244
rect 2209 3420 2243 3436
rect 2209 3228 2243 3244
rect 2327 3420 2361 3436
rect 2327 3228 2361 3244
rect 2445 3420 2479 3436
rect 2445 3228 2479 3244
rect 2563 3420 2597 3436
rect 2563 3228 2597 3244
rect 2681 3420 2715 3436
rect 2681 3228 2715 3244
rect 2799 3420 2833 3436
rect 2799 3228 2833 3244
rect 2917 3420 2951 3436
rect 2917 3228 2951 3244
rect 3035 3420 3069 3436
rect 3035 3228 3069 3244
rect 3153 3420 3187 3436
rect 3153 3228 3187 3244
rect 3271 3420 3305 3436
rect 3271 3228 3305 3244
rect 3389 3420 3423 3436
rect 3389 3228 3423 3244
rect 3507 3420 3541 3436
rect 3507 3228 3541 3244
rect 3625 3420 3659 3436
rect 3625 3228 3659 3244
rect 3743 3420 3777 3436
rect 3743 3228 3777 3244
rect 3861 3420 3895 3436
rect 3861 3228 3895 3244
rect 3979 3420 4013 3436
rect 3979 3228 4013 3244
rect 4097 3420 4131 3436
rect 4097 3228 4131 3244
rect 4215 3420 4249 3436
rect 4215 3228 4249 3244
rect 4333 3420 4367 3436
rect 4333 3228 4367 3244
rect 4451 3420 4485 3436
rect 4451 3228 4485 3244
rect 4569 3420 4603 3436
rect 4569 3228 4603 3244
rect 4687 3420 4721 3436
rect 4687 3228 4721 3244
rect 4805 3420 4839 3436
rect 4805 3228 4839 3244
rect 4923 3420 4957 3436
rect 4923 3228 4957 3244
rect 5041 3420 5075 3436
rect 5041 3228 5075 3244
rect 5159 3420 5193 3436
rect 5159 3228 5193 3244
rect 3786 3043 3802 3077
rect 3836 3043 3852 3077
rect 2091 2984 2125 3000
rect 2091 2792 2125 2808
rect 2209 2984 2243 3000
rect 2209 2792 2243 2808
rect 2327 2984 2361 3000
rect 2327 2792 2361 2808
rect 2445 2984 2479 3000
rect 2445 2792 2479 2808
rect 2563 2984 2597 3000
rect 2563 2792 2597 2808
rect 2681 2984 2715 3000
rect 2681 2792 2715 2808
rect 2799 2984 2833 3000
rect 2799 2792 2833 2808
rect 2917 2984 2951 3000
rect 2917 2792 2951 2808
rect 3035 2984 3069 3000
rect 3035 2792 3069 2808
rect 3153 2984 3187 3000
rect 3153 2792 3187 2808
rect 3271 2984 3305 3000
rect 3271 2792 3305 2808
rect 3389 2984 3423 3000
rect 3389 2792 3423 2808
rect 3507 2984 3541 3000
rect 3507 2792 3541 2808
rect 3625 2984 3659 3000
rect 3625 2792 3659 2808
rect 3743 2984 3777 3000
rect 3743 2792 3777 2808
rect 3861 2984 3895 3000
rect 3861 2792 3895 2808
rect 3979 2984 4013 3000
rect 3979 2792 4013 2808
rect 4097 2984 4131 3000
rect 4097 2792 4131 2808
rect 4215 2984 4249 3000
rect 4215 2792 4249 2808
rect 4333 2984 4367 3000
rect 4333 2792 4367 2808
rect 4451 2984 4485 3000
rect 4451 2792 4485 2808
rect 4569 2984 4603 3000
rect 4569 2792 4603 2808
rect 4687 2984 4721 3000
rect 4687 2792 4721 2808
rect 4805 2984 4839 3000
rect 4805 2792 4839 2808
rect 4923 2984 4957 3000
rect 4923 2792 4957 2808
rect 5041 2984 5075 3000
rect 5041 2792 5075 2808
rect 5159 2984 5193 3000
rect 5159 2792 5193 2808
rect 2134 2715 2150 2749
rect 2184 2715 2200 2749
rect 2252 2715 2268 2749
rect 2302 2715 2318 2749
rect 2370 2715 2386 2749
rect 2420 2715 2436 2749
rect 2488 2715 2504 2749
rect 2538 2715 2554 2749
rect 2606 2715 2622 2749
rect 2656 2715 2672 2749
rect 2724 2715 2740 2749
rect 2774 2715 2790 2749
rect 2842 2715 2858 2749
rect 2892 2715 2908 2749
rect 2960 2715 2976 2749
rect 3010 2715 3026 2749
rect 3078 2715 3094 2749
rect 3128 2715 3144 2749
rect 3196 2715 3212 2749
rect 3246 2715 3262 2749
rect 3314 2715 3330 2749
rect 3364 2715 3380 2749
rect 3432 2715 3448 2749
rect 3482 2715 3498 2749
rect 3550 2715 3566 2749
rect 3600 2715 3616 2749
rect 3668 2715 3684 2749
rect 3718 2715 3734 2749
rect 3904 2715 3920 2749
rect 3954 2715 3970 2749
rect 4022 2715 4038 2749
rect 4072 2715 4088 2749
rect 4140 2715 4156 2749
rect 4190 2715 4206 2749
rect 4258 2715 4274 2749
rect 4308 2715 4324 2749
rect 4376 2715 4392 2749
rect 4426 2715 4442 2749
rect 4494 2715 4510 2749
rect 4544 2715 4560 2749
rect 4612 2715 4628 2749
rect 4662 2715 4678 2749
rect 4730 2715 4746 2749
rect 4780 2715 4796 2749
rect 4848 2715 4864 2749
rect 4898 2715 4914 2749
rect 4966 2715 4982 2749
rect 5016 2715 5032 2749
rect 5084 2715 5100 2749
rect 5134 2715 5150 2749
rect 2091 2548 2125 2564
rect 2091 2356 2125 2372
rect 2209 2548 2243 2564
rect 2209 2356 2243 2372
rect 2327 2548 2361 2564
rect 2327 2356 2361 2372
rect 2445 2548 2479 2564
rect 2445 2356 2479 2372
rect 2563 2548 2597 2564
rect 2563 2356 2597 2372
rect 2681 2548 2715 2564
rect 2681 2356 2715 2372
rect 2799 2548 2833 2564
rect 2799 2356 2833 2372
rect 2917 2548 2951 2564
rect 2917 2356 2951 2372
rect 3035 2548 3069 2564
rect 3035 2356 3069 2372
rect 3153 2548 3187 2564
rect 3153 2356 3187 2372
rect 3271 2548 3305 2564
rect 3271 2356 3305 2372
rect 3389 2548 3423 2564
rect 3389 2356 3423 2372
rect 3507 2548 3541 2564
rect 3507 2356 3541 2372
rect 3625 2548 3659 2564
rect 3625 2356 3659 2372
rect 3743 2548 3777 2564
rect 3743 2356 3777 2372
rect 3861 2548 3895 2564
rect 3861 2356 3895 2372
rect 3979 2548 4013 2564
rect 3979 2356 4013 2372
rect 4097 2548 4131 2564
rect 4097 2356 4131 2372
rect 4215 2548 4249 2564
rect 4215 2356 4249 2372
rect 4333 2548 4367 2564
rect 4333 2356 4367 2372
rect 4451 2548 4485 2564
rect 4451 2356 4485 2372
rect 4569 2548 4603 2564
rect 4569 2356 4603 2372
rect 4687 2548 4721 2564
rect 4687 2356 4721 2372
rect 4805 2548 4839 2564
rect 4805 2356 4839 2372
rect 4923 2548 4957 2564
rect 4923 2356 4957 2372
rect 5041 2548 5075 2564
rect 5041 2356 5075 2372
rect 5159 2548 5193 2564
rect 5159 2356 5193 2372
rect 2134 2279 2150 2313
rect 2184 2279 2200 2313
rect 2252 2279 2268 2313
rect 2302 2279 2318 2313
rect 2370 2279 2386 2313
rect 2420 2279 2436 2313
rect 2488 2279 2504 2313
rect 2538 2279 2554 2313
rect 2606 2279 2622 2313
rect 2656 2279 2672 2313
rect 2724 2279 2740 2313
rect 2774 2279 2790 2313
rect 2842 2279 2858 2313
rect 2892 2279 2908 2313
rect 2960 2279 2976 2313
rect 3010 2279 3026 2313
rect 3078 2279 3094 2313
rect 3128 2279 3144 2313
rect 3196 2279 3212 2313
rect 3246 2279 3262 2313
rect 3314 2279 3330 2313
rect 3364 2279 3380 2313
rect 3432 2279 3448 2313
rect 3482 2279 3498 2313
rect 3550 2279 3566 2313
rect 3600 2279 3616 2313
rect 3668 2279 3684 2313
rect 3718 2279 3734 2313
rect 3786 2279 3802 2313
rect 3836 2279 3852 2313
rect 3904 2279 3920 2313
rect 3954 2279 3970 2313
rect 4022 2279 4038 2313
rect 4072 2279 4088 2313
rect 4140 2279 4156 2313
rect 4190 2279 4206 2313
rect 4258 2279 4274 2313
rect 4308 2279 4324 2313
rect 4376 2279 4392 2313
rect 4426 2279 4442 2313
rect 4494 2279 4510 2313
rect 4544 2279 4560 2313
rect 4612 2279 4628 2313
rect 4662 2279 4678 2313
rect 4730 2279 4746 2313
rect 4780 2279 4796 2313
rect 4848 2279 4864 2313
rect 4898 2279 4914 2313
rect 4966 2279 4982 2313
rect 5016 2279 5032 2313
rect 5084 2279 5100 2313
rect 5134 2279 5150 2313
rect 1977 2180 1980 2273
rect 5273 2211 5280 2273
rect 2014 2180 2073 2211
rect 1977 2177 2073 2180
rect 5211 2180 5280 2211
rect 5211 2177 5307 2180
<< viali >>
rect 1980 3519 2014 3610
rect 1980 2273 2011 3519
rect 2011 2273 2014 3519
rect 5280 3519 5314 3610
rect 2150 3479 2184 3513
rect 2268 3479 2302 3513
rect 2386 3479 2420 3513
rect 2504 3479 2538 3513
rect 2622 3479 2656 3513
rect 2740 3479 2774 3513
rect 2858 3479 2892 3513
rect 2976 3479 3010 3513
rect 3094 3479 3128 3513
rect 3212 3479 3246 3513
rect 3330 3479 3364 3513
rect 3448 3479 3482 3513
rect 3566 3479 3600 3513
rect 3684 3479 3718 3513
rect 3802 3479 3836 3513
rect 3920 3479 3954 3513
rect 4038 3479 4072 3513
rect 4156 3479 4190 3513
rect 4274 3479 4308 3513
rect 4392 3479 4426 3513
rect 4510 3479 4544 3513
rect 4628 3479 4662 3513
rect 4746 3479 4780 3513
rect 4864 3479 4898 3513
rect 4982 3479 5016 3513
rect 5100 3479 5134 3513
rect 2091 3244 2125 3420
rect 2209 3244 2243 3420
rect 2327 3244 2361 3420
rect 2445 3244 2479 3420
rect 2563 3244 2597 3420
rect 2681 3244 2715 3420
rect 2799 3244 2833 3420
rect 2917 3244 2951 3420
rect 3035 3244 3069 3420
rect 3153 3244 3187 3420
rect 3271 3244 3305 3420
rect 3389 3244 3423 3420
rect 3507 3244 3541 3420
rect 3625 3244 3659 3420
rect 3743 3244 3777 3420
rect 3861 3244 3895 3420
rect 3979 3244 4013 3420
rect 4097 3244 4131 3420
rect 4215 3244 4249 3420
rect 4333 3244 4367 3420
rect 4451 3244 4485 3420
rect 4569 3244 4603 3420
rect 4687 3244 4721 3420
rect 4805 3244 4839 3420
rect 4923 3244 4957 3420
rect 5041 3244 5075 3420
rect 5159 3244 5193 3420
rect 3802 3043 3836 3077
rect 2091 2808 2125 2984
rect 2209 2808 2243 2984
rect 2327 2808 2361 2984
rect 2445 2808 2479 2984
rect 2563 2808 2597 2984
rect 2681 2808 2715 2984
rect 2799 2808 2833 2984
rect 2917 2808 2951 2984
rect 3035 2808 3069 2984
rect 3153 2808 3187 2984
rect 3271 2808 3305 2984
rect 3389 2808 3423 2984
rect 3507 2808 3541 2984
rect 3625 2808 3659 2984
rect 3743 2808 3777 2984
rect 3861 2808 3895 2984
rect 3979 2808 4013 2984
rect 4097 2808 4131 2984
rect 4215 2808 4249 2984
rect 4333 2808 4367 2984
rect 4451 2808 4485 2984
rect 4569 2808 4603 2984
rect 4687 2808 4721 2984
rect 4805 2808 4839 2984
rect 4923 2808 4957 2984
rect 5041 2808 5075 2984
rect 5159 2808 5193 2984
rect 2150 2715 2184 2749
rect 2268 2715 2302 2749
rect 2386 2715 2420 2749
rect 2504 2715 2538 2749
rect 2622 2715 2656 2749
rect 2740 2715 2774 2749
rect 2858 2715 2892 2749
rect 2976 2715 3010 2749
rect 3094 2715 3128 2749
rect 3212 2715 3246 2749
rect 3330 2715 3364 2749
rect 3448 2715 3482 2749
rect 3566 2715 3600 2749
rect 3684 2715 3718 2749
rect 3920 2715 3954 2749
rect 4038 2715 4072 2749
rect 4156 2715 4190 2749
rect 4274 2715 4308 2749
rect 4392 2715 4426 2749
rect 4510 2715 4544 2749
rect 4628 2715 4662 2749
rect 4746 2715 4780 2749
rect 4864 2715 4898 2749
rect 4982 2715 5016 2749
rect 5100 2715 5134 2749
rect 2091 2372 2125 2548
rect 2209 2372 2243 2548
rect 2327 2372 2361 2548
rect 2445 2372 2479 2548
rect 2563 2372 2597 2548
rect 2681 2372 2715 2548
rect 2799 2372 2833 2548
rect 2917 2372 2951 2548
rect 3035 2372 3069 2548
rect 3153 2372 3187 2548
rect 3271 2372 3305 2548
rect 3389 2372 3423 2548
rect 3507 2372 3541 2548
rect 3625 2372 3659 2548
rect 3743 2372 3777 2548
rect 3861 2372 3895 2548
rect 3979 2372 4013 2548
rect 4097 2372 4131 2548
rect 4215 2372 4249 2548
rect 4333 2372 4367 2548
rect 4451 2372 4485 2548
rect 4569 2372 4603 2548
rect 4687 2372 4721 2548
rect 4805 2372 4839 2548
rect 4923 2372 4957 2548
rect 5041 2372 5075 2548
rect 5159 2372 5193 2548
rect 2150 2279 2184 2313
rect 2268 2279 2302 2313
rect 2386 2279 2420 2313
rect 2504 2279 2538 2313
rect 2622 2279 2656 2313
rect 2740 2279 2774 2313
rect 2858 2279 2892 2313
rect 2976 2279 3010 2313
rect 3094 2279 3128 2313
rect 3212 2279 3246 2313
rect 3330 2279 3364 2313
rect 3448 2279 3482 2313
rect 3566 2279 3600 2313
rect 3684 2279 3718 2313
rect 3802 2279 3836 2313
rect 3920 2279 3954 2313
rect 4038 2279 4072 2313
rect 4156 2279 4190 2313
rect 4274 2279 4308 2313
rect 4392 2279 4426 2313
rect 4510 2279 4544 2313
rect 4628 2279 4662 2313
rect 4746 2279 4780 2313
rect 4864 2279 4898 2313
rect 4982 2279 5016 2313
rect 5100 2279 5134 2313
rect 1980 2180 2014 2273
rect 5280 2273 5307 3519
rect 5307 2273 5314 3519
rect 5280 2180 5314 2273
<< metal1 >>
rect 1970 3610 5320 3630
rect 1970 2180 1980 3610
rect 2014 3580 5280 3610
rect 2014 2220 2020 3580
rect 2120 3540 2210 3550
rect 2120 3470 2130 3540
rect 2200 3470 2210 3540
rect 5080 3540 5170 3550
rect 2120 3460 2210 3470
rect 2251 3513 3085 3529
rect 2251 3479 2268 3513
rect 2302 3479 2386 3513
rect 2420 3479 2504 3513
rect 2538 3479 2622 3513
rect 2656 3479 2740 3513
rect 2774 3479 2858 3513
rect 2892 3479 2976 3513
rect 3010 3479 3085 3513
rect 2251 3463 3085 3479
rect 3139 3463 3145 3529
rect 3196 3513 4029 3529
rect 3196 3479 3212 3513
rect 3246 3479 3330 3513
rect 3364 3479 3448 3513
rect 3482 3479 3566 3513
rect 3600 3479 3684 3513
rect 3718 3479 3802 3513
rect 3836 3479 3920 3513
rect 3954 3479 4029 3513
rect 3196 3463 4029 3479
rect 4083 3463 4089 3529
rect 4140 3513 4973 3529
rect 4140 3479 4156 3513
rect 4190 3479 4274 3513
rect 4308 3479 4392 3513
rect 4426 3479 4510 3513
rect 4544 3479 4628 3513
rect 4662 3479 4746 3513
rect 4780 3479 4864 3513
rect 4898 3479 4973 3513
rect 4140 3463 4973 3479
rect 5027 3463 5033 3529
rect 3078 3462 3145 3463
rect 4022 3462 4089 3463
rect 4966 3462 5033 3463
rect 5080 3470 5090 3540
rect 5160 3470 5170 3540
rect 5080 3460 5170 3470
rect 2081 3426 2135 3432
rect 2081 3232 2135 3238
rect 2199 3426 2253 3432
rect 2199 3232 2253 3238
rect 2317 3426 2371 3432
rect 2317 3232 2371 3238
rect 2435 3426 2489 3432
rect 2435 3232 2489 3238
rect 2553 3426 2607 3432
rect 2553 3232 2607 3238
rect 2671 3426 2725 3432
rect 2671 3232 2725 3238
rect 2789 3426 2843 3432
rect 2789 3232 2843 3238
rect 2907 3426 2961 3432
rect 2907 3232 2961 3238
rect 3025 3426 3079 3432
rect 3025 3232 3079 3238
rect 3143 3426 3197 3432
rect 3143 3232 3197 3238
rect 3261 3426 3315 3432
rect 3261 3232 3315 3238
rect 3379 3426 3433 3432
rect 3379 3232 3433 3238
rect 3497 3426 3551 3432
rect 3497 3232 3551 3238
rect 3615 3426 3669 3432
rect 3615 3232 3669 3238
rect 3733 3426 3787 3432
rect 3733 3232 3787 3238
rect 3851 3426 3905 3432
rect 3851 3232 3905 3238
rect 3969 3426 4023 3432
rect 3969 3232 4023 3238
rect 4087 3426 4141 3432
rect 4087 3232 4141 3238
rect 4205 3426 4259 3432
rect 4205 3232 4259 3238
rect 4323 3426 4377 3432
rect 4323 3232 4377 3238
rect 4441 3426 4495 3432
rect 4441 3232 4495 3238
rect 4559 3426 4613 3432
rect 4559 3232 4613 3238
rect 4677 3426 4731 3432
rect 4677 3232 4731 3238
rect 4795 3426 4849 3432
rect 4795 3232 4849 3238
rect 4913 3426 4967 3432
rect 4913 3232 4967 3238
rect 5031 3426 5085 3432
rect 5031 3232 5085 3238
rect 5149 3426 5203 3432
rect 5149 3232 5203 3238
rect 3786 3027 3793 3093
rect 3847 3027 3853 3093
rect 3786 3026 3853 3027
rect 2081 2990 2135 2996
rect 2081 2796 2135 2802
rect 2199 2990 2253 2996
rect 2199 2796 2253 2802
rect 2317 2990 2371 2996
rect 2317 2796 2371 2802
rect 2435 2990 2489 2996
rect 2435 2796 2489 2802
rect 2553 2990 2607 2996
rect 2553 2796 2607 2802
rect 2671 2990 2725 2996
rect 2671 2796 2725 2802
rect 2789 2990 2843 2996
rect 2789 2796 2843 2802
rect 2907 2990 2961 2996
rect 2907 2796 2961 2802
rect 3025 2990 3079 2996
rect 3025 2796 3079 2802
rect 3143 2990 3197 2996
rect 3143 2796 3197 2802
rect 3261 2990 3315 2996
rect 3261 2796 3315 2802
rect 3379 2990 3433 2996
rect 3379 2796 3433 2802
rect 3497 2990 3551 2996
rect 3497 2796 3551 2802
rect 3615 2990 3669 2996
rect 3733 2990 3787 2996
rect 3669 2802 3733 2830
rect 3615 2796 3787 2802
rect 3851 2990 3905 2996
rect 3851 2796 3905 2802
rect 3969 2990 4023 2996
rect 3969 2796 4023 2802
rect 4087 2990 4141 2996
rect 4087 2796 4141 2802
rect 4205 2990 4259 2996
rect 4205 2796 4259 2802
rect 4323 2990 4377 2996
rect 4323 2796 4377 2802
rect 4441 2990 4495 2996
rect 4441 2796 4495 2802
rect 4559 2990 4613 2996
rect 4559 2796 4613 2802
rect 4677 2990 4731 2996
rect 4677 2796 4731 2802
rect 4795 2990 4849 2996
rect 4795 2796 4849 2802
rect 4913 2990 4967 2996
rect 4913 2796 4967 2802
rect 5031 2990 5085 2996
rect 5031 2796 5085 2802
rect 5149 2990 5203 2996
rect 5149 2796 5203 2802
rect 3078 2765 3145 2766
rect 3550 2765 3617 2766
rect 2134 2760 2672 2765
rect 2120 2690 2130 2760
rect 2200 2749 2672 2760
rect 2200 2715 2268 2749
rect 2302 2715 2386 2749
rect 2420 2715 2504 2749
rect 2538 2715 2622 2749
rect 2656 2715 2672 2749
rect 2200 2699 2672 2715
rect 2723 2749 3085 2765
rect 2723 2715 2740 2749
rect 2774 2715 2858 2749
rect 2892 2715 2976 2749
rect 3010 2715 3085 2749
rect 2723 2699 3085 2715
rect 3139 2699 3145 2765
rect 3196 2749 3557 2765
rect 3196 2715 3212 2749
rect 3246 2715 3330 2749
rect 3364 2715 3448 2749
rect 3482 2715 3557 2749
rect 3196 2699 3557 2715
rect 3611 2699 3617 2765
rect 3668 2749 3734 2796
rect 4022 2765 4089 2766
rect 4494 2765 4561 2766
rect 3668 2715 3684 2749
rect 3718 2715 3734 2749
rect 3668 2699 3734 2715
rect 3904 2749 4029 2765
rect 3904 2715 3920 2749
rect 3954 2715 4029 2749
rect 3904 2699 4029 2715
rect 4083 2699 4089 2765
rect 4138 2749 4501 2765
rect 4138 2715 4156 2749
rect 4190 2715 4274 2749
rect 4308 2715 4392 2749
rect 4426 2715 4501 2749
rect 4138 2699 4501 2715
rect 4555 2699 4561 2765
rect 4611 2749 5149 2765
rect 4611 2715 4628 2749
rect 4662 2715 4746 2749
rect 4780 2715 4864 2749
rect 4898 2715 4982 2749
rect 5016 2715 5100 2749
rect 5134 2715 5149 2749
rect 4610 2699 5149 2715
rect 2200 2690 2210 2699
rect 2630 2670 2670 2699
rect 4610 2670 4650 2699
rect 2630 2600 2730 2670
rect 2660 2560 2730 2600
rect 4550 2600 4650 2670
rect 4550 2560 4620 2600
rect 2081 2554 2135 2560
rect 2081 2360 2135 2366
rect 2199 2554 2253 2560
rect 2199 2360 2253 2366
rect 2317 2554 2371 2560
rect 2317 2360 2371 2366
rect 2435 2554 2489 2560
rect 2435 2360 2489 2366
rect 2553 2554 2607 2560
rect 2553 2360 2607 2366
rect 2671 2554 2725 2560
rect 2671 2360 2725 2366
rect 2789 2554 2843 2560
rect 2789 2360 2843 2366
rect 2907 2554 2961 2560
rect 2907 2360 2961 2366
rect 3025 2554 3079 2560
rect 3025 2360 3079 2366
rect 3143 2554 3197 2560
rect 3143 2360 3197 2366
rect 3261 2554 3315 2560
rect 3261 2360 3315 2366
rect 3379 2554 3433 2560
rect 3379 2360 3433 2366
rect 3497 2554 3551 2560
rect 3497 2360 3551 2366
rect 3615 2554 3669 2560
rect 3615 2360 3669 2366
rect 3733 2554 3787 2560
rect 3733 2360 3787 2366
rect 3851 2554 3905 2560
rect 3851 2360 3905 2366
rect 3969 2554 4023 2560
rect 3969 2360 4023 2366
rect 4087 2554 4141 2560
rect 4087 2360 4141 2366
rect 4205 2554 4259 2560
rect 4205 2360 4259 2366
rect 4323 2554 4377 2560
rect 4323 2360 4377 2366
rect 4441 2554 4495 2560
rect 4441 2360 4495 2366
rect 4559 2554 4613 2560
rect 4559 2360 4613 2366
rect 4677 2554 4731 2560
rect 4677 2360 4731 2366
rect 4795 2554 4849 2560
rect 4795 2360 4849 2366
rect 4913 2554 4967 2560
rect 4913 2360 4967 2366
rect 5031 2554 5085 2560
rect 5031 2360 5085 2366
rect 5149 2554 5203 2560
rect 5149 2360 5203 2366
rect 2120 2260 2130 2330
rect 2200 2260 2210 2330
rect 3078 2329 3145 2330
rect 4022 2329 4089 2330
rect 4966 2329 5033 2330
rect 2252 2313 3085 2329
rect 2252 2279 2268 2313
rect 2302 2279 2386 2313
rect 2420 2279 2504 2313
rect 2538 2279 2622 2313
rect 2656 2279 2740 2313
rect 2774 2279 2858 2313
rect 2892 2279 2976 2313
rect 3010 2279 3085 2313
rect 2252 2263 3085 2279
rect 3139 2263 3145 2329
rect 3196 2313 4029 2329
rect 3196 2279 3212 2313
rect 3246 2279 3330 2313
rect 3364 2279 3448 2313
rect 3482 2279 3566 2313
rect 3600 2279 3684 2313
rect 3718 2279 3802 2313
rect 3836 2279 3920 2313
rect 3954 2279 4029 2313
rect 3196 2263 4029 2279
rect 4083 2263 4089 2329
rect 4140 2313 4973 2329
rect 4140 2279 4156 2313
rect 4190 2279 4274 2313
rect 4308 2279 4392 2313
rect 4426 2279 4510 2313
rect 4544 2279 4628 2313
rect 4662 2279 4746 2313
rect 4780 2279 4864 2313
rect 4898 2279 4973 2313
rect 4140 2263 4973 2279
rect 5027 2263 5033 2329
rect 5084 2313 5150 2329
rect 5084 2279 5100 2313
rect 5134 2279 5150 2313
rect 5084 2263 5150 2279
rect 5270 2220 5280 3580
rect 2014 2212 5280 2220
rect 2014 2180 2070 2212
rect 1970 2160 2070 2180
rect 5210 2180 5280 2212
rect 5314 2180 5320 3610
rect 5210 2160 5320 2180
<< via1 >>
rect 2130 3513 2200 3540
rect 2130 3479 2150 3513
rect 2150 3479 2184 3513
rect 2184 3479 2200 3513
rect 2130 3470 2200 3479
rect 3085 3513 3139 3529
rect 3085 3479 3094 3513
rect 3094 3479 3128 3513
rect 3128 3479 3139 3513
rect 3085 3463 3139 3479
rect 4029 3513 4083 3529
rect 4029 3479 4038 3513
rect 4038 3479 4072 3513
rect 4072 3479 4083 3513
rect 4029 3463 4083 3479
rect 4973 3513 5027 3529
rect 4973 3479 4982 3513
rect 4982 3479 5016 3513
rect 5016 3479 5027 3513
rect 4973 3463 5027 3479
rect 5090 3513 5160 3540
rect 5090 3479 5100 3513
rect 5100 3479 5134 3513
rect 5134 3479 5160 3513
rect 5090 3470 5160 3479
rect 2081 3420 2135 3426
rect 2081 3244 2091 3420
rect 2091 3244 2125 3420
rect 2125 3244 2135 3420
rect 2081 3238 2135 3244
rect 2199 3420 2253 3426
rect 2199 3244 2209 3420
rect 2209 3244 2243 3420
rect 2243 3244 2253 3420
rect 2199 3238 2253 3244
rect 2317 3420 2371 3426
rect 2317 3244 2327 3420
rect 2327 3244 2361 3420
rect 2361 3244 2371 3420
rect 2317 3238 2371 3244
rect 2435 3420 2489 3426
rect 2435 3244 2445 3420
rect 2445 3244 2479 3420
rect 2479 3244 2489 3420
rect 2435 3238 2489 3244
rect 2553 3420 2607 3426
rect 2553 3244 2563 3420
rect 2563 3244 2597 3420
rect 2597 3244 2607 3420
rect 2553 3238 2607 3244
rect 2671 3420 2725 3426
rect 2671 3244 2681 3420
rect 2681 3244 2715 3420
rect 2715 3244 2725 3420
rect 2671 3238 2725 3244
rect 2789 3420 2843 3426
rect 2789 3244 2799 3420
rect 2799 3244 2833 3420
rect 2833 3244 2843 3420
rect 2789 3238 2843 3244
rect 2907 3420 2961 3426
rect 2907 3244 2917 3420
rect 2917 3244 2951 3420
rect 2951 3244 2961 3420
rect 2907 3238 2961 3244
rect 3025 3420 3079 3426
rect 3025 3244 3035 3420
rect 3035 3244 3069 3420
rect 3069 3244 3079 3420
rect 3025 3238 3079 3244
rect 3143 3420 3197 3426
rect 3143 3244 3153 3420
rect 3153 3244 3187 3420
rect 3187 3244 3197 3420
rect 3143 3238 3197 3244
rect 3261 3420 3315 3426
rect 3261 3244 3271 3420
rect 3271 3244 3305 3420
rect 3305 3244 3315 3420
rect 3261 3238 3315 3244
rect 3379 3420 3433 3426
rect 3379 3244 3389 3420
rect 3389 3244 3423 3420
rect 3423 3244 3433 3420
rect 3379 3238 3433 3244
rect 3497 3420 3551 3426
rect 3497 3244 3507 3420
rect 3507 3244 3541 3420
rect 3541 3244 3551 3420
rect 3497 3238 3551 3244
rect 3615 3420 3669 3426
rect 3615 3244 3625 3420
rect 3625 3244 3659 3420
rect 3659 3244 3669 3420
rect 3615 3238 3669 3244
rect 3733 3420 3787 3426
rect 3733 3244 3743 3420
rect 3743 3244 3777 3420
rect 3777 3244 3787 3420
rect 3733 3238 3787 3244
rect 3851 3420 3905 3426
rect 3851 3244 3861 3420
rect 3861 3244 3895 3420
rect 3895 3244 3905 3420
rect 3851 3238 3905 3244
rect 3969 3420 4023 3426
rect 3969 3244 3979 3420
rect 3979 3244 4013 3420
rect 4013 3244 4023 3420
rect 3969 3238 4023 3244
rect 4087 3420 4141 3426
rect 4087 3244 4097 3420
rect 4097 3244 4131 3420
rect 4131 3244 4141 3420
rect 4087 3238 4141 3244
rect 4205 3420 4259 3426
rect 4205 3244 4215 3420
rect 4215 3244 4249 3420
rect 4249 3244 4259 3420
rect 4205 3238 4259 3244
rect 4323 3420 4377 3426
rect 4323 3244 4333 3420
rect 4333 3244 4367 3420
rect 4367 3244 4377 3420
rect 4323 3238 4377 3244
rect 4441 3420 4495 3426
rect 4441 3244 4451 3420
rect 4451 3244 4485 3420
rect 4485 3244 4495 3420
rect 4441 3238 4495 3244
rect 4559 3420 4613 3426
rect 4559 3244 4569 3420
rect 4569 3244 4603 3420
rect 4603 3244 4613 3420
rect 4559 3238 4613 3244
rect 4677 3420 4731 3426
rect 4677 3244 4687 3420
rect 4687 3244 4721 3420
rect 4721 3244 4731 3420
rect 4677 3238 4731 3244
rect 4795 3420 4849 3426
rect 4795 3244 4805 3420
rect 4805 3244 4839 3420
rect 4839 3244 4849 3420
rect 4795 3238 4849 3244
rect 4913 3420 4967 3426
rect 4913 3244 4923 3420
rect 4923 3244 4957 3420
rect 4957 3244 4967 3420
rect 4913 3238 4967 3244
rect 5031 3420 5085 3426
rect 5031 3244 5041 3420
rect 5041 3244 5075 3420
rect 5075 3244 5085 3420
rect 5031 3238 5085 3244
rect 5149 3420 5203 3426
rect 5149 3244 5159 3420
rect 5159 3244 5193 3420
rect 5193 3244 5203 3420
rect 5149 3238 5203 3244
rect 3793 3077 3847 3093
rect 3793 3043 3802 3077
rect 3802 3043 3836 3077
rect 3836 3043 3847 3077
rect 3793 3027 3847 3043
rect 2081 2984 2135 2990
rect 2081 2808 2091 2984
rect 2091 2808 2125 2984
rect 2125 2808 2135 2984
rect 2081 2802 2135 2808
rect 2199 2984 2253 2990
rect 2199 2808 2209 2984
rect 2209 2808 2243 2984
rect 2243 2808 2253 2984
rect 2199 2802 2253 2808
rect 2317 2984 2371 2990
rect 2317 2808 2327 2984
rect 2327 2808 2361 2984
rect 2361 2808 2371 2984
rect 2317 2802 2371 2808
rect 2435 2984 2489 2990
rect 2435 2808 2445 2984
rect 2445 2808 2479 2984
rect 2479 2808 2489 2984
rect 2435 2802 2489 2808
rect 2553 2984 2607 2990
rect 2553 2808 2563 2984
rect 2563 2808 2597 2984
rect 2597 2808 2607 2984
rect 2553 2802 2607 2808
rect 2671 2984 2725 2990
rect 2671 2808 2681 2984
rect 2681 2808 2715 2984
rect 2715 2808 2725 2984
rect 2671 2802 2725 2808
rect 2789 2984 2843 2990
rect 2789 2808 2799 2984
rect 2799 2808 2833 2984
rect 2833 2808 2843 2984
rect 2789 2802 2843 2808
rect 2907 2984 2961 2990
rect 2907 2808 2917 2984
rect 2917 2808 2951 2984
rect 2951 2808 2961 2984
rect 2907 2802 2961 2808
rect 3025 2984 3079 2990
rect 3025 2808 3035 2984
rect 3035 2808 3069 2984
rect 3069 2808 3079 2984
rect 3025 2802 3079 2808
rect 3143 2984 3197 2990
rect 3143 2808 3153 2984
rect 3153 2808 3187 2984
rect 3187 2808 3197 2984
rect 3143 2802 3197 2808
rect 3261 2984 3315 2990
rect 3261 2808 3271 2984
rect 3271 2808 3305 2984
rect 3305 2808 3315 2984
rect 3261 2802 3315 2808
rect 3379 2984 3433 2990
rect 3379 2808 3389 2984
rect 3389 2808 3423 2984
rect 3423 2808 3433 2984
rect 3379 2802 3433 2808
rect 3497 2984 3551 2990
rect 3497 2808 3507 2984
rect 3507 2808 3541 2984
rect 3541 2808 3551 2984
rect 3497 2802 3551 2808
rect 3615 2984 3669 2990
rect 3615 2808 3625 2984
rect 3625 2808 3659 2984
rect 3659 2808 3669 2984
rect 3733 2984 3787 2990
rect 3615 2802 3669 2808
rect 3733 2808 3743 2984
rect 3743 2808 3777 2984
rect 3777 2808 3787 2984
rect 3733 2802 3787 2808
rect 3851 2984 3905 2990
rect 3851 2808 3861 2984
rect 3861 2808 3895 2984
rect 3895 2808 3905 2984
rect 3851 2802 3905 2808
rect 3969 2984 4023 2990
rect 3969 2808 3979 2984
rect 3979 2808 4013 2984
rect 4013 2808 4023 2984
rect 3969 2802 4023 2808
rect 4087 2984 4141 2990
rect 4087 2808 4097 2984
rect 4097 2808 4131 2984
rect 4131 2808 4141 2984
rect 4087 2802 4141 2808
rect 4205 2984 4259 2990
rect 4205 2808 4215 2984
rect 4215 2808 4249 2984
rect 4249 2808 4259 2984
rect 4205 2802 4259 2808
rect 4323 2984 4377 2990
rect 4323 2808 4333 2984
rect 4333 2808 4367 2984
rect 4367 2808 4377 2984
rect 4323 2802 4377 2808
rect 4441 2984 4495 2990
rect 4441 2808 4451 2984
rect 4451 2808 4485 2984
rect 4485 2808 4495 2984
rect 4441 2802 4495 2808
rect 4559 2984 4613 2990
rect 4559 2808 4569 2984
rect 4569 2808 4603 2984
rect 4603 2808 4613 2984
rect 4559 2802 4613 2808
rect 4677 2984 4731 2990
rect 4677 2808 4687 2984
rect 4687 2808 4721 2984
rect 4721 2808 4731 2984
rect 4677 2802 4731 2808
rect 4795 2984 4849 2990
rect 4795 2808 4805 2984
rect 4805 2808 4839 2984
rect 4839 2808 4849 2984
rect 4795 2802 4849 2808
rect 4913 2984 4967 2990
rect 4913 2808 4923 2984
rect 4923 2808 4957 2984
rect 4957 2808 4967 2984
rect 4913 2802 4967 2808
rect 5031 2984 5085 2990
rect 5031 2808 5041 2984
rect 5041 2808 5075 2984
rect 5075 2808 5085 2984
rect 5031 2802 5085 2808
rect 5149 2984 5203 2990
rect 5149 2808 5159 2984
rect 5159 2808 5193 2984
rect 5193 2808 5203 2984
rect 5149 2802 5203 2808
rect 2130 2749 2200 2760
rect 2130 2715 2150 2749
rect 2150 2715 2184 2749
rect 2184 2715 2200 2749
rect 2130 2690 2200 2715
rect 3085 2749 3139 2765
rect 3085 2715 3094 2749
rect 3094 2715 3128 2749
rect 3128 2715 3139 2749
rect 3085 2699 3139 2715
rect 3557 2749 3611 2765
rect 3557 2715 3566 2749
rect 3566 2715 3600 2749
rect 3600 2715 3611 2749
rect 3557 2699 3611 2715
rect 4029 2749 4083 2765
rect 4029 2715 4038 2749
rect 4038 2715 4072 2749
rect 4072 2715 4083 2749
rect 4029 2699 4083 2715
rect 4501 2749 4555 2765
rect 4501 2715 4510 2749
rect 4510 2715 4544 2749
rect 4544 2715 4555 2749
rect 4501 2699 4555 2715
rect 2081 2548 2135 2554
rect 2081 2372 2091 2548
rect 2091 2372 2125 2548
rect 2125 2372 2135 2548
rect 2081 2366 2135 2372
rect 2199 2548 2253 2554
rect 2199 2372 2209 2548
rect 2209 2372 2243 2548
rect 2243 2372 2253 2548
rect 2199 2366 2253 2372
rect 2317 2548 2371 2554
rect 2317 2372 2327 2548
rect 2327 2372 2361 2548
rect 2361 2372 2371 2548
rect 2317 2366 2371 2372
rect 2435 2548 2489 2554
rect 2435 2372 2445 2548
rect 2445 2372 2479 2548
rect 2479 2372 2489 2548
rect 2435 2366 2489 2372
rect 2553 2548 2607 2554
rect 2553 2372 2563 2548
rect 2563 2372 2597 2548
rect 2597 2372 2607 2548
rect 2553 2366 2607 2372
rect 2671 2548 2725 2554
rect 2671 2372 2681 2548
rect 2681 2372 2715 2548
rect 2715 2372 2725 2548
rect 2671 2366 2725 2372
rect 2789 2548 2843 2554
rect 2789 2372 2799 2548
rect 2799 2372 2833 2548
rect 2833 2372 2843 2548
rect 2789 2366 2843 2372
rect 2907 2548 2961 2554
rect 2907 2372 2917 2548
rect 2917 2372 2951 2548
rect 2951 2372 2961 2548
rect 2907 2366 2961 2372
rect 3025 2548 3079 2554
rect 3025 2372 3035 2548
rect 3035 2372 3069 2548
rect 3069 2372 3079 2548
rect 3025 2366 3079 2372
rect 3143 2548 3197 2554
rect 3143 2372 3153 2548
rect 3153 2372 3187 2548
rect 3187 2372 3197 2548
rect 3143 2366 3197 2372
rect 3261 2548 3315 2554
rect 3261 2372 3271 2548
rect 3271 2372 3305 2548
rect 3305 2372 3315 2548
rect 3261 2366 3315 2372
rect 3379 2548 3433 2554
rect 3379 2372 3389 2548
rect 3389 2372 3423 2548
rect 3423 2372 3433 2548
rect 3379 2366 3433 2372
rect 3497 2548 3551 2554
rect 3497 2372 3507 2548
rect 3507 2372 3541 2548
rect 3541 2372 3551 2548
rect 3497 2366 3551 2372
rect 3615 2548 3669 2554
rect 3615 2372 3625 2548
rect 3625 2372 3659 2548
rect 3659 2372 3669 2548
rect 3615 2366 3669 2372
rect 3733 2548 3787 2554
rect 3733 2372 3743 2548
rect 3743 2372 3777 2548
rect 3777 2372 3787 2548
rect 3733 2366 3787 2372
rect 3851 2548 3905 2554
rect 3851 2372 3861 2548
rect 3861 2372 3895 2548
rect 3895 2372 3905 2548
rect 3851 2366 3905 2372
rect 3969 2548 4023 2554
rect 3969 2372 3979 2548
rect 3979 2372 4013 2548
rect 4013 2372 4023 2548
rect 3969 2366 4023 2372
rect 4087 2548 4141 2554
rect 4087 2372 4097 2548
rect 4097 2372 4131 2548
rect 4131 2372 4141 2548
rect 4087 2366 4141 2372
rect 4205 2548 4259 2554
rect 4205 2372 4215 2548
rect 4215 2372 4249 2548
rect 4249 2372 4259 2548
rect 4205 2366 4259 2372
rect 4323 2548 4377 2554
rect 4323 2372 4333 2548
rect 4333 2372 4367 2548
rect 4367 2372 4377 2548
rect 4323 2366 4377 2372
rect 4441 2548 4495 2554
rect 4441 2372 4451 2548
rect 4451 2372 4485 2548
rect 4485 2372 4495 2548
rect 4441 2366 4495 2372
rect 4559 2548 4613 2554
rect 4559 2372 4569 2548
rect 4569 2372 4603 2548
rect 4603 2372 4613 2548
rect 4559 2366 4613 2372
rect 4677 2548 4731 2554
rect 4677 2372 4687 2548
rect 4687 2372 4721 2548
rect 4721 2372 4731 2548
rect 4677 2366 4731 2372
rect 4795 2548 4849 2554
rect 4795 2372 4805 2548
rect 4805 2372 4839 2548
rect 4839 2372 4849 2548
rect 4795 2366 4849 2372
rect 4913 2548 4967 2554
rect 4913 2372 4923 2548
rect 4923 2372 4957 2548
rect 4957 2372 4967 2548
rect 4913 2366 4967 2372
rect 5031 2548 5085 2554
rect 5031 2372 5041 2548
rect 5041 2372 5075 2548
rect 5075 2372 5085 2548
rect 5031 2366 5085 2372
rect 5149 2548 5203 2554
rect 5149 2372 5159 2548
rect 5159 2372 5193 2548
rect 5193 2372 5203 2548
rect 5149 2366 5203 2372
rect 2130 2313 2200 2330
rect 2130 2279 2150 2313
rect 2150 2279 2184 2313
rect 2184 2279 2200 2313
rect 2130 2260 2200 2279
rect 3085 2313 3139 2329
rect 3085 2279 3094 2313
rect 3094 2279 3128 2313
rect 3128 2279 3139 2313
rect 3085 2263 3139 2279
rect 4029 2313 4083 2329
rect 4029 2279 4038 2313
rect 4038 2279 4072 2313
rect 4072 2279 4083 2313
rect 4029 2263 4083 2279
rect 4973 2313 5027 2329
rect 4973 2279 4982 2313
rect 4982 2279 5016 2313
rect 5016 2279 5027 2313
rect 4973 2263 5027 2279
rect 2070 2160 5210 2212
<< metal2 >>
rect 2310 3580 4930 3760
rect 2081 3540 2253 3550
rect 2081 3470 2130 3540
rect 2200 3470 2253 3540
rect 2310 3480 2380 3580
rect 2540 3480 2610 3580
rect 2780 3480 2850 3580
rect 2081 3460 2253 3470
rect 2081 3426 2135 3460
rect 2081 2990 2135 3238
rect 2081 2760 2135 2802
rect 2199 3426 2253 3460
rect 2199 2990 2253 3238
rect 2199 2760 2253 2802
rect 2081 2690 2130 2760
rect 2200 2690 2253 2760
rect 2081 2554 2135 2690
rect 2081 2360 2135 2366
rect 2199 2554 2253 2690
rect 2199 2360 2253 2366
rect 2317 3426 2371 3480
rect 2317 2990 2371 3238
rect 2317 2554 2371 2802
rect 2317 2360 2371 2366
rect 2435 3426 2489 3432
rect 2435 2990 2489 3238
rect 2435 2554 2489 2802
rect 2435 2360 2489 2366
rect 2553 3426 2607 3480
rect 2553 2990 2607 3238
rect 2553 2554 2607 2802
rect 2553 2360 2607 2366
rect 2671 3426 2725 3432
rect 2671 2990 2725 3238
rect 2671 2554 2725 2802
rect 2671 2360 2725 2366
rect 2789 3426 2843 3480
rect 2970 3460 3040 3580
rect 3070 3530 3150 3540
rect 3070 3470 3080 3530
rect 3140 3470 3150 3530
rect 3250 3480 3320 3580
rect 3490 3480 3560 3580
rect 3720 3480 3790 3580
rect 3070 3463 3085 3470
rect 3139 3463 3150 3470
rect 3070 3460 3150 3463
rect 3000 3432 3040 3460
rect 2789 2990 2843 3238
rect 2789 2554 2843 2802
rect 2789 2360 2843 2366
rect 2907 3426 2961 3432
rect 3000 3426 3079 3432
rect 3000 3390 3025 3426
rect 2907 2990 2961 3238
rect 3025 2990 3079 3238
rect 2907 2554 2961 2802
rect 3000 2802 3025 2830
rect 3000 2796 3079 2802
rect 3143 3426 3197 3432
rect 3143 2990 3197 3238
rect 3261 3426 3315 3480
rect 3261 2990 3315 3238
rect 3197 2802 3220 2830
rect 3143 2796 3220 2802
rect 3000 2660 3040 2796
rect 3070 2765 3150 2768
rect 3070 2758 3085 2765
rect 3139 2758 3150 2765
rect 3070 2698 3080 2758
rect 3140 2698 3150 2758
rect 3070 2688 3150 2698
rect 3180 2660 3220 2796
rect 3000 2630 3079 2660
rect 2907 2360 2961 2366
rect 3025 2554 3079 2630
rect 3025 2360 3079 2366
rect 3143 2630 3220 2660
rect 3143 2554 3197 2630
rect 3261 2554 3315 2802
rect 3197 2366 3220 2400
rect 3143 2360 3220 2366
rect 3261 2360 3315 2366
rect 3379 3426 3433 3432
rect 3379 2990 3433 3238
rect 3497 3426 3551 3480
rect 3497 2990 3551 3238
rect 3379 2554 3433 2802
rect 3478 2802 3497 2830
rect 3478 2796 3551 2802
rect 3615 3426 3669 3432
rect 3615 2990 3669 3238
rect 3733 3426 3787 3480
rect 3914 3460 3984 3580
rect 4014 3530 4094 3540
rect 4014 3470 4024 3530
rect 4084 3470 4094 3530
rect 4200 3480 4270 3580
rect 4430 3480 4500 3580
rect 4670 3480 4740 3580
rect 4014 3463 4029 3470
rect 4083 3463 4094 3470
rect 4014 3460 4094 3463
rect 3944 3432 3984 3460
rect 3733 3160 3787 3238
rect 3714 3132 3787 3160
rect 3851 3426 3905 3432
rect 3944 3426 4023 3432
rect 3944 3390 3969 3426
rect 3851 3160 3905 3238
rect 3851 3132 3930 3160
rect 3714 2996 3754 3132
rect 3787 3094 3853 3104
rect 3787 3034 3788 3094
rect 3848 3034 3853 3094
rect 3787 3027 3793 3034
rect 3847 3027 3853 3034
rect 3787 3024 3853 3027
rect 3890 2996 3930 3132
rect 3714 2990 3787 2996
rect 3714 2960 3733 2990
rect 3669 2802 3690 2830
rect 3615 2796 3690 2802
rect 3478 2660 3518 2796
rect 3551 2765 3617 2768
rect 3551 2758 3557 2765
rect 3611 2758 3617 2765
rect 3551 2698 3552 2758
rect 3612 2698 3617 2758
rect 3551 2688 3617 2698
rect 3650 2660 3690 2796
rect 3478 2630 3551 2660
rect 3379 2360 3433 2366
rect 3497 2554 3551 2630
rect 3497 2360 3551 2366
rect 3615 2630 3690 2660
rect 3615 2554 3669 2630
rect 3615 2360 3669 2366
rect 3733 2554 3787 2802
rect 3733 2360 3787 2366
rect 3851 2990 3930 2996
rect 3905 2960 3930 2990
rect 3969 2990 4023 3238
rect 3851 2554 3905 2802
rect 3950 2802 3969 2830
rect 3950 2796 4023 2802
rect 4087 3426 4141 3432
rect 4087 2990 4141 3238
rect 4205 3426 4259 3480
rect 4205 2990 4259 3238
rect 4141 2802 4160 2830
rect 4087 2796 4160 2802
rect 3950 2660 3990 2796
rect 4023 2765 4090 2768
rect 4023 2758 4029 2765
rect 4083 2758 4090 2765
rect 4023 2698 4024 2758
rect 4084 2698 4090 2758
rect 4023 2688 4090 2698
rect 4120 2660 4160 2796
rect 3950 2630 4023 2660
rect 3851 2360 3905 2366
rect 3969 2554 4023 2630
rect 3969 2360 4023 2366
rect 4087 2630 4160 2660
rect 4087 2554 4141 2630
rect 4205 2554 4259 2802
rect 4141 2366 4170 2390
rect 4087 2360 4170 2366
rect 4205 2360 4259 2366
rect 4323 3426 4377 3432
rect 4323 2990 4377 3238
rect 4441 3426 4495 3480
rect 4441 2990 4495 3238
rect 4323 2554 4377 2802
rect 4420 2802 4441 2830
rect 4420 2796 4495 2802
rect 4559 3426 4613 3432
rect 4559 2990 4613 3238
rect 4677 3426 4731 3480
rect 4858 3460 4930 3580
rect 5080 3540 5203 3550
rect 4958 3530 5038 3540
rect 4958 3470 4968 3530
rect 5028 3470 5038 3530
rect 4958 3463 4973 3470
rect 5027 3463 5038 3470
rect 4958 3460 5038 3463
rect 5080 3470 5090 3540
rect 5160 3470 5203 3540
rect 4888 3432 4928 3460
rect 5080 3432 5203 3470
rect 4677 2990 4731 3238
rect 4613 2802 4636 2830
rect 4559 2796 4636 2802
rect 4420 2660 4462 2796
rect 4495 2765 4561 2768
rect 4495 2758 4501 2765
rect 4555 2758 4561 2765
rect 4495 2698 4496 2758
rect 4556 2698 4561 2758
rect 4495 2688 4561 2698
rect 4593 2660 4636 2796
rect 4420 2630 4495 2660
rect 4323 2360 4377 2366
rect 4441 2554 4495 2630
rect 4441 2360 4495 2366
rect 4559 2630 4636 2660
rect 4559 2554 4613 2630
rect 4559 2360 4613 2366
rect 4677 2554 4731 2802
rect 4677 2360 4731 2366
rect 4795 3426 4849 3432
rect 4888 3426 4967 3432
rect 4888 3390 4913 3426
rect 4795 2990 4849 3238
rect 4795 2554 4849 2802
rect 4795 2360 4849 2366
rect 4913 2990 4967 3238
rect 4913 2554 4967 2802
rect 4913 2360 4967 2366
rect 5031 3426 5203 3432
rect 5085 3390 5149 3426
rect 5031 2990 5085 3238
rect 5031 2554 5085 2802
rect 5149 2990 5203 3238
rect 5149 2554 5203 2802
rect 5085 2366 5100 2400
rect 5031 2360 5100 2366
rect 5149 2360 5203 2366
rect 2070 2330 2140 2360
rect 2190 2330 2260 2360
rect 2070 2260 2130 2330
rect 2200 2260 2260 2330
rect 2070 2212 2140 2260
rect 2190 2212 2260 2260
rect 2430 2212 2500 2360
rect 2660 2212 2730 2360
rect 2900 2212 2970 2360
rect 3070 2329 3150 2332
rect 3070 2322 3085 2329
rect 3139 2322 3150 2329
rect 3070 2262 3080 2322
rect 3140 2262 3150 2322
rect 3070 2252 3150 2262
rect 3180 2330 3220 2360
rect 3180 2212 3250 2330
rect 3370 2212 3440 2360
rect 3610 2212 3680 2360
rect 3840 2212 3910 2360
rect 4014 2329 4094 2332
rect 4014 2322 4029 2329
rect 4083 2322 4094 2329
rect 4014 2262 4024 2322
rect 4084 2262 4094 2322
rect 4014 2252 4094 2262
rect 4130 2320 4170 2360
rect 4130 2212 4200 2320
rect 4310 2212 4380 2360
rect 4550 2212 4620 2360
rect 4790 2212 4860 2360
rect 4958 2329 5038 2332
rect 4958 2322 4973 2329
rect 5027 2322 5038 2329
rect 4958 2262 4968 2322
rect 5028 2262 5038 2322
rect 4958 2252 5038 2262
rect 5070 2212 5210 2360
rect 2070 1870 2090 2160
rect 3570 2040 5210 2160
rect 5190 1870 5210 2040
rect 2070 1850 5210 1870
<< via2 >>
rect 3080 3529 3140 3530
rect 3080 3470 3085 3529
rect 3085 3470 3139 3529
rect 3139 3470 3140 3529
rect 3080 2699 3085 2758
rect 3085 2699 3139 2758
rect 3139 2699 3140 2758
rect 3080 2698 3140 2699
rect 4024 3529 4084 3530
rect 4024 3470 4029 3529
rect 4029 3470 4083 3529
rect 4083 3470 4084 3529
rect 3788 3093 3848 3094
rect 3788 3034 3793 3093
rect 3793 3034 3847 3093
rect 3847 3034 3848 3093
rect 3552 2699 3557 2758
rect 3557 2699 3611 2758
rect 3611 2699 3612 2758
rect 3552 2698 3612 2699
rect 4024 2699 4029 2758
rect 4029 2699 4083 2758
rect 4083 2699 4084 2758
rect 4024 2698 4084 2699
rect 4968 3529 5028 3530
rect 4968 3470 4973 3529
rect 4973 3470 5027 3529
rect 5027 3470 5028 3529
rect 4496 2699 4501 2758
rect 4501 2699 4555 2758
rect 4555 2699 4556 2758
rect 4496 2698 4556 2699
rect 3080 2263 3085 2322
rect 3085 2263 3139 2322
rect 3139 2263 3140 2322
rect 3080 2262 3140 2263
rect 4024 2263 4029 2322
rect 4029 2263 4083 2322
rect 4083 2263 4084 2322
rect 4024 2262 4084 2263
rect 4968 2263 4973 2322
rect 4973 2263 5027 2322
rect 5027 2263 5028 2322
rect 4968 2262 5028 2263
rect 2090 2160 3570 2170
rect 2090 2040 3570 2160
rect 2090 1870 5190 2040
<< metal3 >>
rect 3660 3600 5050 3670
rect 3660 3570 3950 3600
rect 4160 3570 5050 3600
rect 3660 3540 3780 3570
rect 3070 3530 3780 3540
rect 3070 3470 3080 3530
rect 3140 3470 3780 3530
rect 3070 3390 3780 3470
rect 4010 3530 4100 3540
rect 4010 3470 4024 3530
rect 4084 3470 4100 3530
rect 4950 3530 5050 3570
rect 4720 3470 4860 3480
rect 4010 3370 4730 3470
rect 4850 3370 4860 3470
rect 4720 3360 4860 3370
rect 4950 3470 4968 3530
rect 5028 3480 5050 3530
rect 5028 3470 5090 3480
rect 4950 3370 4960 3470
rect 5080 3370 5090 3470
rect 4950 3360 5090 3370
rect 3540 3200 5270 3300
rect 3070 2758 3150 2768
rect 3070 2698 3080 2758
rect 3140 2698 3150 2758
rect 3070 2610 3150 2698
rect 3540 2758 3630 3200
rect 3780 3104 5270 3120
rect 3774 3094 5270 3104
rect 3774 3034 3788 3094
rect 3848 3034 5270 3094
rect 3774 3020 5270 3034
rect 3774 3010 3880 3020
rect 3540 2698 3552 2758
rect 3612 2698 3630 2758
rect 3540 2680 3630 2698
rect 4010 2840 5270 2940
rect 4010 2758 4100 2840
rect 4010 2698 4024 2758
rect 4084 2698 4100 2758
rect 4010 2680 4100 2698
rect 4480 2758 5270 2770
rect 4480 2698 4496 2758
rect 4556 2698 5270 2758
rect 4480 2670 5270 2698
rect 4480 2610 4580 2670
rect 3070 2510 4580 2610
rect 4710 2430 5270 2530
rect 4710 2420 4860 2430
rect 3070 2322 3780 2400
rect 3070 2262 3080 2322
rect 3140 2262 3780 2322
rect 3070 2250 3780 2262
rect 4010 2322 4730 2420
rect 4010 2262 4024 2322
rect 4084 2320 4730 2322
rect 4850 2320 4860 2420
rect 4084 2262 4100 2320
rect 4710 2310 4860 2320
rect 4950 2330 5270 2340
rect 4010 2250 4100 2262
rect 3660 2220 3780 2250
rect 4950 2230 4960 2330
rect 5080 2240 5270 2330
rect 5080 2230 5090 2240
rect 4950 2220 5090 2230
rect 2070 2180 3010 2200
rect 3660 2190 3950 2220
rect 4160 2190 5050 2220
rect 2070 2170 3590 2180
rect 2070 1870 2090 2170
rect 3570 2060 3590 2170
rect 3660 2120 5050 2190
rect 3570 2040 5210 2060
rect 5190 1870 5210 2040
rect 2070 1850 5210 1870
<< via3 >>
rect 4730 3370 4850 3470
rect 4960 3370 5080 3470
rect 4730 2320 4850 2420
rect 4960 2322 5080 2330
rect 4960 2262 4968 2322
rect 4968 2262 5028 2322
rect 5028 2262 5080 2322
rect 4960 2230 5080 2262
rect 2090 1870 5190 2040
<< metal4 >>
rect 4720 3470 4860 3480
rect 4720 3370 4730 3470
rect 4850 3370 4860 3470
rect 4720 2420 4860 3370
rect 4720 2320 4730 2420
rect 4850 2320 4860 2420
rect 4720 2310 4860 2320
rect 4950 3470 5090 3480
rect 4950 3370 4960 3470
rect 5080 3370 5090 3470
rect 4950 2330 5090 3370
rect 4950 2230 4960 2330
rect 5080 2230 5090 2330
rect 4950 2220 5090 2230
rect 2070 2040 5210 2060
rect 2070 1870 2090 2040
rect 5190 1870 5210 2040
rect 2070 1850 5210 1870
<< labels >>
rlabel metal4 2070 1850 5210 2060 1 VHI
rlabel metal2 2310 3690 4930 3760 1 IOUT
rlabel metal3 5240 3200 5270 3300 1 G2
rlabel metal3 5240 3020 5270 3120 1 VREF
rlabel metal3 5240 2840 5270 2940 1 G4
rlabel metal3 5240 2670 5270 2770 1 G8
rlabel metal3 5240 2430 5270 2530 1 G16
rlabel metal3 5240 2240 5270 2340 1 G32
<< end >>
