magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< nwell >>
rect -36 679 512 1471
<< poly >>
rect 114 714 144 1055
rect 81 648 144 714
rect 114 255 144 648
<< locali >>
rect 0 1397 476 1431
rect 62 1204 96 1397
rect 64 648 98 714
rect 166 698 200 1270
rect 270 1204 304 1397
rect 374 1297 408 1397
rect 166 664 217 698
rect 166 92 200 664
rect 62 17 96 92
rect 270 17 304 92
rect 374 17 408 104
rect 0 -17 476 17
use sky130_sram_1r1w_24x128_8_contact_15  sky130_sram_1r1w_24x128_8_contact_15_0
timestamp 1661296025
transform 1 0 48 0 1 648
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_28  sky130_sram_1r1w_24x128_8_contact_28_0
timestamp 1661296025
transform 1 0 366 0 1 1256
box -59 -43 109 125
use sky130_sram_1r1w_24x128_8_contact_29  sky130_sram_1r1w_24x128_8_contact_29_0
timestamp 1661296025
transform 1 0 366 0 1 63
box -26 -26 76 108
use sky130_sram_1r1w_24x128_8_nmos_m2_w0_740_sli_dli_da_p  sky130_sram_1r1w_24x128_8_nmos_m2_w0_740_sli_dli_da_p_0
timestamp 1661296025
transform 1 0 54 0 1 51
box -26 -26 284 204
use sky130_sram_1r1w_24x128_8_pmos_m2_w1_260_sli_dli_da_p  sky130_sram_1r1w_24x128_8_pmos_m2_w1_260_sli_dli_da_p_0
timestamp 1661296025
transform 1 0 54 0 1 1111
box -59 -56 317 306
<< labels >>
rlabel locali s 81 681 81 681 4 A
port 1 nsew
rlabel locali s 200 681 200 681 4 Z
port 2 nsew
rlabel locali s 238 0 238 0 4 gnd
port 3 nsew
rlabel locali s 238 1414 238 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 476 1414
<< end >>
