magic
tech sky130B
timestamp 1662317594
<< metal4 >>
rect 8500 -3275 8650 -3050
rect 8250 -4325 8400 -3325
rect 8750 -3425 8900 -2975
rect 9000 -3650 9150 -3000
rect 8500 -4775 8650 -3650
rect 9250 -3850 9400 -3100
rect 0 -9775 150 -8700
rect 250 -9950 400 -8925
rect 0 -41925 150 -9975
rect 0 -47375 150 -42225
rect 250 -42625 400 -10150
rect 500 -10175 650 -9175
rect 250 -46600 400 -42850
rect 500 -42975 650 -10375
rect 750 -10425 900 -9425
rect 500 -46000 650 -43250
rect 750 -43325 900 -10650
rect 1000 -10700 1150 -9625
rect 1000 -12925 1150 -10925
rect 1250 -11025 1400 -9875
rect 1250 -12450 1400 -11250
rect 1500 -11300 1650 -10150
rect 1500 -12225 1650 -11575
rect 1750 -11650 1900 -10375
rect 1750 -11950 1900 -11800
rect 2000 -11850 2150 -10450
rect 2250 -11600 2400 -10450
rect 2500 -11325 2650 -10300
rect 2750 -11075 2900 -10075
rect 3000 -10850 3150 -9875
rect 3250 -10650 3400 -9675
rect 3500 -10450 3650 -9450
rect 3750 -10225 3900 -9250
rect 4000 -10000 4150 -9025
rect 4250 -9800 4400 -8800
rect 4500 -9600 4650 -8625
rect 4750 -9400 4900 -8425
rect 5000 -9200 5150 -8250
rect 5250 -8975 5400 -8075
rect 5500 -8800 5650 -7875
rect 5750 -8650 5900 -7625
rect 6000 -8525 6150 -7350
rect 6250 -8400 6400 -7075
rect 6500 -7775 6650 -6850
rect 6750 -7575 6900 -6600
rect 7000 -7375 7150 -6400
rect 7250 -7150 7400 -6175
rect 7500 -6975 7650 -6000
rect 7750 -6750 7900 -5825
rect 8000 -6550 8150 -5625
rect 8250 -6375 8400 -5425
rect 8500 -6175 8650 -5150
rect 8750 -6025 8900 -3975
rect 9500 -4000 9650 -3175
rect 9250 -4250 9400 -4075
rect 9750 -4100 9900 -3275
rect 10000 -4150 10150 -3325
rect 10250 -4175 10400 -3375
rect 9000 -5850 9150 -4275
rect 9500 -4500 9650 -4175
rect 10500 -4200 10650 -3400
rect 10750 -4225 10900 -3425
rect 11000 -4200 11150 -3425
rect 11250 -4150 11400 -3400
rect 11500 -4125 11650 -3375
rect 11750 -4100 11900 -3350
rect 12000 -4075 12150 -3350
rect 12250 -4025 12400 -3350
rect 12500 -4000 12650 -3325
rect 12750 -4000 12900 -3325
rect 13000 -4050 13150 -3350
rect 13250 -4075 13400 -3350
rect 13500 -4100 13650 -3350
rect 13750 -4125 13900 -3400
rect 14000 -4150 14150 -3425
rect 9250 -5700 9400 -4525
rect 9750 -4750 9900 -4250
rect 9500 -5600 9650 -4750
rect 10000 -4975 10150 -4325
rect 9750 -5500 9900 -5000
rect 10250 -5200 10400 -4375
rect 10000 -5425 10150 -5225
rect 10500 -5375 10650 -4400
rect 7000 -7850 7150 -7600
rect 7250 -7850 7400 -7400
rect 7500 -7850 7650 -7175
rect 7750 -7900 7900 -6975
rect 8000 -7975 8150 -6800
rect 6500 -8300 6650 -8125
rect 6750 -8300 6900 -8025
rect 1000 -38450 1150 -13850
rect 1250 -13975 1400 -13075
rect 1250 -35800 1400 -14250
rect 1500 -14375 1650 -12750
rect 1500 -34475 1650 -14600
rect 1750 -14650 1900 -12425
rect 2000 -14875 2150 -12150
rect 1750 -31425 1900 -14900
rect 2250 -15050 2400 -11850
rect 2000 -29900 2150 -15100
rect 2500 -15200 2650 -11600
rect 2250 -19375 2400 -15250
rect 2750 -15325 2900 -11350
rect 2500 -18125 2650 -15400
rect 3000 -15500 3150 -11100
rect 2750 -17175 2900 -15525
rect 3250 -15650 3400 -10875
rect 3000 -16650 3150 -15650
rect 3250 -16250 3400 -15800
rect 2750 -18125 2900 -17700
rect 3000 -17975 3150 -17050
rect 3250 -17675 3400 -16575
rect 3500 -17400 3650 -10675
rect 3750 -17150 3900 -10450
rect 4000 -16900 4150 -10250
rect 4250 -16700 4400 -10025
rect 4500 -16500 4650 -9825
rect 4750 -16325 4900 -9625
rect 5000 -16125 5150 -9400
rect 5250 -15950 5400 -9225
rect 5500 -15800 5650 -9025
rect 5750 -15675 5900 -8875
rect 6000 -15550 6150 -8725
rect 6250 -15450 6400 -8600
rect 6500 -15325 6650 -8500
rect 6750 -15225 6900 -8450
rect 7000 -15125 7150 -8000
rect 7250 -15050 7400 -8000
rect 7500 -15000 7650 -8000
rect 8250 -8100 8400 -6600
rect 7750 -15025 7900 -8100
rect 2500 -18775 2650 -18625
rect 2250 -21425 2400 -20225
rect 2500 -21375 2650 -19175
rect 2750 -21050 2900 -18700
rect 3000 -20800 3150 -18225
rect 3250 -20625 3400 -17975
rect 2250 -28750 2400 -21800
rect 2500 -27950 2650 -21650
rect 2750 -27125 2900 -21325
rect 3000 -26550 3150 -21025
rect 3250 -25950 3400 -22350
rect 3500 -22675 3650 -17650
rect 3500 -25400 3650 -23125
rect 3750 -23175 3900 -17425
rect 3750 -25050 3900 -23550
rect 4000 -23575 4150 -17175
rect 4250 -23900 4400 -16950
rect 4000 -24775 4150 -23900
rect 4500 -23975 4650 -16725
rect 4750 -24000 4900 -16500
rect 4250 -24500 4400 -24100
rect 4500 -24350 4650 -24125
rect 4750 -24300 4900 -24150
rect 5000 -24200 5150 -16350
rect 5250 -24025 5400 -16175
rect 5500 -23875 5650 -16000
rect 5750 -23775 5900 -15875
rect 6000 -23700 6150 -15725
rect 6250 -23750 6400 -15625
rect 6500 -23775 6650 -15500
rect 6750 -23825 6900 -15400
rect 7000 -23875 7150 -15300
rect 7250 -23925 7400 -15225
rect 7500 -23950 7650 -15175
rect 7750 -19325 7900 -15200
rect 8000 -19250 8150 -8150
rect 8500 -8225 8650 -6400
rect 8250 -19150 8400 -8250
rect 8500 -8800 8650 -8375
rect 8750 -8925 8900 -6200
rect 8500 -19025 8650 -8975
rect 9000 -9125 9150 -6050
rect 8750 -14325 8900 -9175
rect 9250 -9300 9400 -5900
rect 9000 -13900 9150 -9350
rect 9500 -9450 9650 -5800
rect 9250 -13500 9400 -9500
rect 9750 -9575 9900 -5700
rect 10000 -9650 10150 -5600
rect 10250 -9650 10400 -5550
rect 10500 -9625 10650 -5525
rect 10750 -9550 10900 -4400
rect 11000 -9500 11150 -4400
rect 11250 -9425 11400 -4350
rect 11500 -9375 11650 -4275
rect 11750 -9275 11900 -4250
rect 12000 -9200 12150 -4250
rect 12250 -9125 12400 -4200
rect 12500 -9000 12650 -4200
rect 12750 -8900 12900 -4200
rect 14250 -4225 14400 -3475
rect 13000 -8825 13150 -4250
rect 13250 -8775 13400 -4250
rect 13500 -8675 13650 -4250
rect 13750 -8675 13900 -4300
rect 14500 -4325 14650 -3550
rect 14000 -8825 14150 -4375
rect 14750 -4400 14900 -3600
rect 14250 -8500 14400 -4425
rect 15000 -4475 15150 -3675
rect 14500 -8150 14650 -4500
rect 15250 -4550 15400 -3750
rect 14750 -7850 14900 -4575
rect 15500 -4650 15650 -3850
rect 15000 -7575 15150 -4650
rect 15750 -4750 15900 -3925
rect 15250 -7325 15400 -4750
rect 15500 -7050 15650 -4825
rect 16000 -4900 16150 -4050
rect 15750 -6800 15900 -4950
rect 16250 -5025 16400 -4150
rect 16000 -6575 16150 -5075
rect 16500 -5175 16650 -4300
rect 16250 -6325 16400 -5225
rect 16750 -5400 16900 -4400
rect 16500 -6075 16650 -5400
rect 17000 -5600 17150 -4500
rect 17250 -5475 17400 -4475
rect 17500 -5300 17650 -4375
rect 17750 -5125 17900 -4225
rect 18000 -4975 18150 -4075
rect 18250 -4800 18400 -3900
rect 18500 -4650 18650 -3775
rect 18750 -4500 18900 -3625
rect 19000 -4350 19150 -3500
rect 19250 -4200 19400 -3350
rect 19500 -4075 19650 -3225
rect 19750 -3950 19900 -3100
rect 20000 -3825 20150 -3000
rect 20250 -3700 20400 -2875
rect 20500 -3600 20650 -2775
rect 20750 -3475 20900 -2650
rect 21000 -3375 21150 -2550
rect 21250 -3250 21400 -2425
rect 21500 -3125 21650 -2325
rect 21750 -3000 21900 -2250
rect 22000 -2900 22150 -2200
rect 22250 -2800 22400 -2150
rect 22500 -2700 22650 -2150
rect 22750 -2650 22900 -2225
rect 9500 -13200 9650 -9650
rect 9750 -12875 9900 -9750
rect 10000 -12600 10150 -9800
rect 10250 -12350 10400 -9800
rect 10500 -12125 10650 -9775
rect 10750 -11875 10900 -9725
rect 11000 -11675 11150 -9650
rect 11250 -11475 11400 -9600
rect 11500 -11250 11650 -9525
rect 11750 -11075 11900 -9425
rect 12000 -10875 12150 -9350
rect 12250 -10725 12400 -9275
rect 12500 -10575 12650 -9200
rect 12750 -10425 12900 -9100
rect 13000 -10225 13150 -9000
rect 13250 -9900 13400 -8925
rect 13500 -9575 13650 -8850
rect 13750 -9250 13900 -8825
rect 10750 -12325 10900 -12125
rect 11000 -12150 11150 -11900
rect 11250 -12025 11400 -11700
rect 11500 -11900 11650 -11500
rect 11750 -11775 11900 -11300
rect 12000 -11650 12150 -11100
rect 12250 -11575 12400 -10900
rect 12500 -11475 12650 -10750
rect 8750 -18850 8900 -14550
rect 9000 -18650 9150 -14200
rect 9250 -18375 9400 -13975
rect 9500 -18100 9650 -13575
rect 9750 -17850 9900 -13325
rect 10000 -17575 10150 -13050
rect 10250 -17275 10400 -12875
rect 10500 -17050 10650 -12650
rect 10750 -13350 10900 -12500
rect 11000 -13050 11150 -12350
rect 11250 -12750 11400 -12200
rect 11500 -12525 11650 -12075
rect 11750 -12325 11900 -11950
rect 12000 -12125 12150 -11825
rect 12250 -11975 12400 -11725
rect 12500 -11900 12650 -11625
rect 10750 -16800 10900 -13500
rect 11000 -16550 11150 -13250
rect 11250 -16300 11400 -12975
rect 11500 -16050 11650 -12725
rect 11750 -15775 11900 -12500
rect 12000 -15550 12150 -12300
rect 12250 -15350 12400 -12150
rect 12500 -15125 12650 -12050
rect 12750 -14950 12900 -10675
rect 13000 -14750 13150 -10625
rect 13250 -14575 13400 -10175
rect 13500 -14400 13650 -9850
rect 13750 -14250 13900 -9525
rect 14000 -14075 14150 -9150
rect 14250 -13925 14400 -8775
rect 14500 -13775 14650 -8425
rect 14750 -13575 14900 -8125
rect 15000 -13450 15150 -7850
rect 15250 -13325 15400 -7550
rect 15500 -13225 15650 -7300
rect 15750 -13125 15900 -7075
rect 16000 -13000 16150 -6825
rect 16250 -12900 16400 -6550
rect 16500 -12800 16650 -6325
rect 16750 -10600 16900 -6100
rect 17000 -10150 17150 -5900
rect 17250 -9675 17400 -5675
rect 17500 -9250 17650 -5500
rect 17750 -8850 17900 -5350
rect 18000 -8475 18150 -5175
rect 18250 -8100 18400 -5025
rect 18500 -7750 18650 -4850
rect 18750 -7400 18900 -4700
rect 19000 -7100 19150 -4550
rect 19250 -6800 19400 -4400
rect 19500 -6475 19650 -4250
rect 19750 -6200 19900 -4125
rect 20000 -5900 20150 -4000
rect 20250 -5625 20400 -3875
rect 20500 -5400 20650 -3800
rect 20750 -5175 20900 -3675
rect 21000 -5000 21150 -3575
rect 21250 -4800 21400 -3425
rect 21500 -4650 21650 -3300
rect 21750 -4475 21900 -3175
rect 17250 -10550 17400 -10025
rect 17500 -10100 17650 -9600
rect 17750 -9650 17900 -9200
rect 18000 -9325 18150 -8775
rect 18250 -9025 18400 -8400
rect 18500 -8800 18650 -8025
rect 18750 -8650 18900 -7675
rect 19000 -8650 19150 -7400
rect 17500 -10400 17650 -10250
rect 17750 -10725 17900 -9925
rect 17000 -11900 17150 -11100
rect 16750 -12725 16900 -12125
rect 17250 -12225 17400 -10775
rect 17000 -12625 17150 -12225
rect 17500 -12325 17650 -10800
rect 17750 -12350 17900 -10975
rect 18000 -12350 18150 -9550
rect 18250 -12350 18400 -9275
rect 18500 -12400 18650 -9000
rect 18750 -9875 18900 -8850
rect 19000 -9975 19150 -9350
rect 19250 -9875 19400 -7075
rect 19500 -9775 19650 -6775
rect 19750 -9675 19900 -6350
rect 20000 -9600 20150 -6150
rect 20250 -9575 20400 -5900
rect 20500 -9550 20650 -5650
rect 20750 -9550 20900 -5425
rect 7750 -23900 7900 -19525
rect 8250 -19625 8400 -19325
rect 8000 -23775 8150 -19700
rect 8500 -19725 8650 -19225
rect 8750 -19800 8900 -19075
rect 8250 -23650 8400 -19825
rect 9000 -19850 9150 -18875
rect 9250 -19900 9400 -18625
rect 8500 -23500 8650 -19900
rect 9500 -19925 9650 -18375
rect 9750 -19900 9900 -18100
rect 10000 -19900 10150 -17825
rect 8750 -23325 8900 -19975
rect 9000 -23125 9150 -20025
rect 9250 -22075 9400 -20075
rect 9500 -21050 9650 -20100
rect 9750 -20325 9900 -20175
rect 9250 -22975 9400 -22825
rect 5500 -24275 5650 -24125
rect 2000 -34225 2150 -31925
rect 2250 -34050 2400 -30275
rect 2500 -33975 2650 -28825
rect 2750 -33900 2900 -28050
rect 3000 -33875 3150 -27300
rect 3250 -33875 3400 -26825
rect 3500 -33875 3650 -26400
rect 3750 -33825 3900 -25925
rect 4000 -33825 4150 -25575
rect 4250 -33850 4400 -25275
rect 4500 -33850 4650 -25025
rect 4750 -33850 4900 -24700
rect 5000 -33850 5150 -24575
rect 5250 -33900 5400 -24450
rect 5500 -33900 5650 -24425
rect 5750 -33950 5900 -24125
rect 6000 -34000 6150 -24025
rect 8250 -24050 8400 -23875
rect 2250 -34375 2400 -34200
rect 2500 -34325 2650 -34125
rect 2750 -34275 2900 -34050
rect 3000 -34250 3150 -34025
rect 3250 -34200 3400 -34025
rect 3500 -34175 3650 -34025
rect 3750 -34175 3900 -34025
rect 4000 -34200 4150 -34050
rect 4250 -34200 4400 -34050
rect 4500 -34175 4650 -34025
rect 4750 -34175 4900 -34000
rect 5000 -34175 5150 -34000
rect 5250 -34200 5400 -34050
rect 5500 -34200 5650 -34050
rect 6250 -34075 6400 -24050
rect 6500 -34200 6650 -24075
rect 1500 -35475 1650 -35325
rect 1750 -35400 1900 -35150
rect 2000 -35275 2150 -34975
rect 2250 -35225 2400 -34825
rect 2500 -35175 2650 -34675
rect 2750 -35150 2900 -34575
rect 3000 -35100 3150 -34525
rect 3250 -35075 3400 -34475
rect 3500 -35075 3650 -34425
rect 3750 -35075 3900 -34425
rect 4000 -35100 4150 -34425
rect 4250 -35150 4400 -34425
rect 4500 -35225 4650 -34450
rect 2000 -35650 2150 -35450
rect 2250 -35575 2400 -35375
rect 2500 -35500 2650 -35325
rect 2750 -35450 2900 -35300
rect 3000 -35450 3150 -35300
rect 3500 -35375 3650 -35225
rect 3750 -35375 3900 -35225
rect 4750 -35325 4900 -34475
rect 5250 -34500 5400 -34350
rect 5500 -34500 5650 -34350
rect 5750 -34525 5900 -34275
rect 6750 -34300 6900 -24075
rect 5000 -35350 5150 -34525
rect 6000 -34550 6150 -34300
rect 7000 -34350 7150 -24125
rect 6250 -34550 6400 -34350
rect 6500 -34625 6650 -34400
rect 7250 -34450 7400 -24200
rect 6750 -34650 6900 -34500
rect 7500 -34575 7650 -24250
rect 8500 -24375 8650 -23700
rect 5250 -35400 5400 -34650
rect 5500 -35400 5650 -34650
rect 5750 -35450 5900 -34675
rect 7750 -34700 7900 -24400
rect 8750 -24575 8900 -23525
rect 8000 -33875 8150 -24575
rect 8250 -32750 8400 -24750
rect 9000 -24800 9150 -23425
rect 9250 -23600 9400 -23450
rect 8500 -32200 8650 -24825
rect 9250 -24875 9400 -24225
rect 9500 -24650 9650 -21700
rect 8750 -31725 8900 -24900
rect 9000 -31100 9150 -25050
rect 9250 -30050 9400 -25275
rect 9750 -25600 9900 -20775
rect 10000 -25650 10150 -20150
rect 10250 -25600 10400 -17550
rect 9500 -26375 9650 -25650
rect 9500 -26675 9650 -26525
rect 9250 -31425 9400 -30925
rect 9500 -31250 9650 -26825
rect 9750 -28250 9900 -26025
rect 9750 -30100 9900 -28600
rect 10000 -28925 10150 -26100
rect 10250 -26200 10400 -25750
rect 10500 -26700 10650 -17300
rect 10750 -26575 10900 -17050
rect 11000 -26375 11150 -16800
rect 11250 -26175 11400 -16500
rect 11500 -26000 11650 -16275
rect 11750 -25775 11900 -16075
rect 12000 -25550 12150 -15800
rect 12250 -25350 12400 -15575
rect 12500 -25200 12650 -15375
rect 12750 -24900 12900 -15175
rect 13000 -24775 13150 -14975
rect 13250 -24525 13400 -14800
rect 13500 -24300 13650 -14625
rect 13750 -24025 13900 -14450
rect 14000 -23800 14150 -14300
rect 14250 -21050 14400 -14125
rect 14500 -20050 14650 -13975
rect 14750 -20200 14900 -13825
rect 14500 -21050 14650 -20250
rect 15000 -20425 15150 -13650
rect 15250 -20600 15400 -13525
rect 14750 -21050 14900 -20600
rect 15500 -20725 15650 -13400
rect 15750 -20875 15900 -13300
rect 15000 -21050 15150 -20900
rect 16000 -21000 16150 -13175
rect 16250 -21025 16400 -13075
rect 16500 -20775 16650 -13000
rect 16750 -20450 16900 -12925
rect 17000 -20125 17150 -12900
rect 17250 -19800 17400 -12825
rect 17500 -17275 17650 -12750
rect 17750 -16925 17900 -12675
rect 18000 -16600 18150 -12625
rect 18250 -16350 18400 -12575
rect 18500 -16100 18650 -12550
rect 18750 -15850 18900 -10400
rect 19000 -12000 19150 -10225
rect 19250 -11875 19400 -10050
rect 19500 -11775 19650 -9925
rect 19750 -11625 19900 -9825
rect 20000 -11450 20150 -9750
rect 20250 -11075 20400 -9750
rect 20500 -10475 20650 -9700
rect 19000 -15675 19150 -12150
rect 19250 -15450 19400 -12025
rect 19500 -15250 19650 -11950
rect 19750 -15050 19900 -11850
rect 20000 -12175 20150 -12025
rect 20000 -12475 20150 -12325
rect 20000 -13475 20150 -12650
rect 20250 -12700 20400 -11450
rect 20500 -12225 20650 -10975
rect 20750 -11750 20900 -10150
rect 21000 -11275 21150 -5250
rect 21250 -10600 21400 -5050
rect 21500 -9875 21650 -4850
rect 21750 -4950 21900 -4800
rect 21750 -8775 21900 -5325
rect 22000 -7150 22150 -3075
rect 22250 -4750 22400 -3000
rect 22250 -5150 22400 -5000
rect 22250 -5550 22400 -5400
rect 21000 -12000 21150 -11650
rect 20000 -14850 20150 -13750
rect 20250 -14700 20400 -13500
rect 20500 -14550 20650 -13075
rect 20750 -14450 20900 -12575
rect 18000 -17275 18150 -16875
rect 18250 -17225 18400 -16600
rect 17500 -19425 17650 -17500
rect 17750 -19025 17900 -17525
rect 18000 -18600 18150 -17475
rect 18500 -18675 18650 -16350
rect 14250 -23550 14400 -21200
rect 16750 -21250 16900 -20775
rect 14500 -23275 14650 -21250
rect 14750 -22950 14900 -21300
rect 17000 -21350 17150 -20450
rect 15000 -22650 15150 -21375
rect 17250 -21425 17400 -20100
rect 17500 -21375 17650 -19750
rect 17750 -21275 17900 -19325
rect 18000 -21225 18150 -18900
rect 18250 -21150 18400 -18700
rect 18500 -21150 18650 -19200
rect 18750 -19350 18900 -16125
rect 18750 -21150 18900 -19700
rect 19000 -19775 19150 -15900
rect 19250 -20050 19400 -15700
rect 19000 -21175 19150 -20050
rect 19500 -20325 19650 -15475
rect 19250 -21250 19400 -20325
rect 19750 -20550 19900 -15275
rect 19500 -21350 19650 -20575
rect 15250 -22275 15400 -21600
rect 15500 -22050 15650 -21625
rect 18250 -21650 18400 -21500
rect 18500 -21675 18650 -21425
rect 15750 -21825 15900 -21675
rect 15750 -22425 15900 -22025
rect 16000 -22400 16150 -21750
rect 16250 -22225 16400 -21775
rect 16500 -22000 16650 -21850
rect 13000 -25675 13150 -25025
rect 10000 -29225 10150 -29075
rect 10250 -29700 10400 -26750
rect 10500 -30425 10650 -26950
rect 9000 -32475 9150 -31725
rect 9250 -32050 9400 -31575
rect 8750 -32700 8900 -32550
rect 6000 -35450 6150 -34700
rect 6250 -35475 6400 -34725
rect 1250 -36850 1400 -36050
rect 1000 -39725 1150 -39100
rect 1250 -41875 1400 -39775
rect 1250 -42200 1400 -42025
rect 750 -45575 900 -43550
rect 1000 -43625 1150 -42825
rect 1000 -45150 1150 -43875
rect 1500 -44150 1650 -37300
rect 1750 -44050 1900 -36575
rect 2000 -42250 2150 -36200
rect 2250 -42075 2400 -36000
rect 2500 -41900 2650 -35850
rect 2750 -41750 2900 -35750
rect 3000 -41625 3150 -35675
rect 3250 -41525 3400 -35600
rect 3500 -41425 3650 -35575
rect 3750 -41350 3900 -35550
rect 4000 -41275 4150 -35500
rect 4250 -41250 4400 -35500
rect 4500 -41200 4650 -35500
rect 4750 -41125 4900 -35525
rect 6500 -35550 6650 -34800
rect 5000 -41075 5150 -35550
rect 5250 -41000 5400 -35550
rect 6750 -35600 6900 -34825
rect 5500 -40950 5650 -35600
rect 5750 -40850 5900 -35650
rect 7000 -35700 7150 -34900
rect 6000 -40800 6150 -35725
rect 7250 -35775 7400 -34950
rect 6250 -40725 6400 -35800
rect 6500 -40625 6650 -35825
rect 7500 -35875 7650 -34975
rect 6750 -40525 6900 -35875
rect 7000 -40450 7150 -35950
rect 7750 -35975 7900 -35300
rect 7250 -40300 7400 -36050
rect 7500 -40100 7650 -36175
rect 7750 -39875 7900 -36425
rect 8250 -37850 8400 -36675
rect 8250 -39000 8400 -38250
rect 8500 -39400 8650 -36225
rect 8750 -39300 8900 -35900
rect 9000 -39200 9150 -35350
rect 9250 -39125 9400 -34700
rect 9500 -38275 9650 -34075
rect 9750 -38175 9900 -33450
rect 10000 -38050 10150 -32275
rect 10250 -37975 10400 -30750
rect 10500 -37750 10650 -30950
rect 10750 -31075 10900 -26800
rect 11000 -26975 11150 -26825
rect 11250 -27100 11400 -26400
rect 10750 -31375 10900 -31225
rect 10750 -37850 10900 -31525
rect 11000 -31575 11150 -27125
rect 11500 -27350 11650 -26200
rect 11000 -37725 11150 -31875
rect 11250 -32075 11400 -27375
rect 11750 -27575 11900 -26000
rect 13250 -26050 13400 -24775
rect 11250 -37550 11400 -32300
rect 11500 -32575 11650 -27575
rect 12000 -27825 12150 -26200
rect 13500 -26325 13650 -24500
rect 11500 -37375 11650 -32850
rect 11750 -32975 11900 -27850
rect 12250 -28025 12400 -26500
rect 13750 -26575 13900 -24275
rect 14000 -24750 14150 -24050
rect 14250 -25125 14400 -23800
rect 14000 -26750 14150 -25200
rect 14500 -25425 14650 -23500
rect 11750 -37225 11900 -33250
rect 12000 -33325 12150 -28050
rect 12500 -28250 12650 -26750
rect 14250 -26925 14400 -25525
rect 14750 -25725 14900 -23250
rect 12000 -37025 12150 -33525
rect 12250 -33650 12400 -28275
rect 12750 -28425 12900 -27000
rect 14500 -27150 14650 -25800
rect 15000 -26000 15150 -22900
rect 12250 -36900 12400 -33875
rect 12500 -33925 12650 -28450
rect 13000 -28600 13150 -27225
rect 14750 -27325 14900 -26075
rect 15250 -26250 15400 -22625
rect 15000 -27450 15150 -26350
rect 15500 -26500 15650 -22650
rect 15750 -23000 15900 -22850
rect 12500 -36775 12650 -34150
rect 12750 -34200 12900 -28650
rect 13250 -28775 13400 -27450
rect 15250 -27550 15400 -26600
rect 15750 -26775 15900 -24325
rect 16000 -24350 16150 -23275
rect 16250 -24600 16400 -22775
rect 15500 -27550 15650 -26850
rect 16000 -27025 16150 -24650
rect 16500 -24725 16650 -22450
rect 16750 -24800 16900 -22225
rect 17000 -24850 17150 -22025
rect 17250 -24850 17400 -22000
rect 17500 -24825 17650 -22125
rect 17750 -24775 17900 -22200
rect 18000 -24725 18150 -22275
rect 18250 -24600 18400 -22075
rect 18500 -24500 18650 -21900
rect 18750 -24350 18900 -21425
rect 19000 -24175 19150 -21450
rect 19750 -21500 19900 -20850
rect 20000 -20900 20150 -15075
rect 20250 -21000 20400 -14900
rect 20500 -20900 20650 -14725
rect 20750 -20775 20900 -14600
rect 21000 -20650 21150 -12150
rect 21250 -20225 21400 -11100
rect 21500 -19825 21650 -10325
rect 21750 -19350 21900 -9475
rect 22000 -18850 22150 -8300
rect 22250 -18300 22400 -5775
rect 22500 -17975 22650 -4150
rect 22750 -7775 22900 -3100
rect 23000 -5900 23150 -2350
rect 23250 -4225 23400 -2650
rect 23000 -7975 23150 -6525
rect 22750 -17000 22900 -8000
rect 23250 -8200 23400 -7150
rect 23500 -8225 23650 -7375
rect 19250 -23975 19400 -21525
rect 19500 -23700 19650 -21600
rect 20000 -21775 20150 -21050
rect 19750 -23350 19900 -21775
rect 20250 -22200 20400 -21150
rect 20000 -22475 20150 -22325
rect 20000 -23775 20150 -23625
rect 20250 -23975 20400 -22950
rect 20500 -23875 20650 -21050
rect 20750 -23725 20900 -20975
rect 21000 -23600 21150 -20850
rect 21250 -21400 21400 -20475
rect 21500 -20875 21650 -20000
rect 21750 -20150 21900 -20000
rect 21500 -21800 21650 -21300
rect 21750 -21850 21900 -20600
rect 21250 -23550 21400 -21900
rect 22000 -21925 22150 -19900
rect 22250 -21925 22400 -18875
rect 22500 -21900 22650 -18125
rect 22750 -21900 22900 -17275
rect 23000 -21875 23150 -8225
rect 23750 -8400 23900 -7525
rect 23250 -21800 23400 -8425
rect 24000 -8600 24150 -7700
rect 23500 -21750 23650 -8700
rect 24250 -8825 24400 -7850
rect 24500 -8900 24650 -8025
rect 23750 -21675 23900 -8950
rect 24000 -9550 24150 -9000
rect 24250 -9675 24400 -9050
rect 24750 -9075 24900 -8200
rect 24000 -21575 24150 -9700
rect 24500 -9825 24650 -9150
rect 25000 -9225 25150 -8350
rect 24250 -21500 24400 -9925
rect 24750 -10100 24900 -9275
rect 25250 -9375 25400 -8475
rect 24500 -21425 24650 -10175
rect 24750 -21175 24900 -10425
rect 25000 -10475 25150 -9425
rect 25500 -9550 25650 -8650
rect 25000 -20850 25150 -10775
rect 25250 -10825 25400 -9575
rect 25750 -9700 25900 -8775
rect 25250 -20325 25400 -11150
rect 25500 -11250 25650 -9750
rect 26000 -9900 26150 -8950
rect 28250 -9175 28400 -5725
rect 28500 -5825 28650 -5650
rect 28750 -5800 28900 -5650
rect 29000 -5800 29150 -5650
rect 29250 -5825 29400 -5675
rect 29500 -5925 29650 -5725
rect 31000 -5800 31150 -5650
rect 31250 -5800 31400 -5650
rect 29750 -6175 29900 -5875
rect 31500 -5900 31650 -5650
rect 31750 -5850 31900 -5650
rect 32000 -5800 32150 -5650
rect 32250 -5800 32400 -5650
rect 30000 -7100 30150 -6250
rect 28500 -7725 28650 -7500
rect 28750 -7700 28900 -7525
rect 29000 -7725 29150 -7525
rect 29250 -8075 29400 -7500
rect 29500 -7650 29650 -7450
rect 29750 -7475 29900 -7200
rect 29500 -8525 29650 -8200
rect 29750 -9025 29900 -8675
rect 31600 -9000 31800 -6000
rect 33500 -6175 33650 -5850
rect 33750 -5900 33900 -5700
rect 34000 -5800 34150 -5650
rect 34250 -5800 34400 -5650
rect 34500 -5850 34650 -5675
rect 34750 -6050 34900 -5800
rect 33250 -6800 33400 -6200
rect 35000 -6425 35150 -6075
rect 33500 -7150 33650 -6825
rect 33750 -7375 33900 -7150
rect 34000 -7525 34150 -7325
rect 34250 -7650 34400 -7450
rect 34500 -7800 34650 -7575
rect 34750 -8050 34900 -7750
rect 33250 -8875 33400 -8650
rect 25500 -19575 25650 -11575
rect 25750 -19425 25900 -9900
rect 26250 -10125 26400 -9200
rect 30000 -9250 30150 -9100
rect 31000 -9375 31150 -9175
rect 31250 -9375 31400 -9175
rect 31500 -9375 31650 -9100
rect 31750 -9375 31900 -9125
rect 32000 -9375 32150 -9175
rect 32250 -9375 32400 -9175
rect 33500 -9200 33650 -8925
rect 35000 -8950 35150 -8075
rect 33750 -9350 33900 -9150
rect 34000 -9400 34150 -9200
rect 34250 -9400 34400 -9200
rect 34500 -9350 34650 -9150
rect 34750 -9200 34900 -8975
rect 36000 -9100 36150 -5725
rect 37500 -8925 37650 -5725
rect 41250 -5975 41400 -5750
rect 41500 -5800 41650 -5650
rect 41750 -5775 41900 -5625
rect 42000 -5800 42150 -5650
rect 42250 -5975 42400 -5750
rect 38500 -7725 38650 -7575
rect 38750 -7725 38900 -7575
rect 39000 -7725 39150 -7575
rect 39250 -7725 39400 -7575
rect 39500 -7725 39650 -7575
rect 39750 -7725 39900 -7575
rect 40000 -7725 40150 -7575
rect 36250 -9300 36400 -9075
rect 36500 -9375 36650 -9200
rect 36750 -9400 36900 -9200
rect 37000 -9350 37150 -9150
rect 37250 -9225 37400 -8975
rect 41000 -9050 41150 -5975
rect 42250 -7200 42400 -7000
rect 41250 -8025 41400 -7775
rect 41500 -7800 41650 -7600
rect 41750 -7625 41900 -7400
rect 42000 -7425 42150 -7200
rect 41250 -9250 41400 -9050
rect 41500 -9375 41650 -9175
rect 41750 -9400 41900 -9200
rect 42000 -9375 42150 -9175
rect 42250 -9275 42400 -9050
rect 42500 -9075 42650 -5950
rect 44250 -6250 44400 -5825
rect 47250 -5875 47400 -5725
rect 44000 -6750 44150 -6325
rect 47000 -6350 47150 -5950
rect 46750 -6825 46900 -6450
rect 43500 -8975 43650 -7400
rect 43750 -7575 43900 -6825
rect 44000 -7400 44150 -7225
rect 44250 -7350 44400 -7200
rect 44500 -7400 44650 -7225
rect 46500 -7325 46650 -6925
rect 44750 -7525 44900 -7325
rect 43750 -9250 43900 -9025
rect 44000 -9375 44150 -9175
rect 44250 -9400 44400 -9200
rect 44500 -9375 44650 -9175
rect 44750 -9275 44900 -9050
rect 45000 -9075 45150 -7500
rect 46250 -7775 46400 -7400
rect 46000 -8300 46150 -7850
rect 46250 -8300 46400 -8150
rect 46500 -8300 46650 -8150
rect 46750 -8300 46900 -8150
rect 47000 -8325 47150 -8150
rect 47250 -9225 47400 -7175
rect 47500 -8300 47650 -8150
rect 21500 -23600 21650 -21975
rect 24000 -22000 24150 -21775
rect 16250 -27275 16400 -24875
rect 16500 -27450 16650 -25000
rect 16750 -27575 16900 -25100
rect 12750 -35975 12900 -34400
rect 13000 -34450 13150 -28825
rect 13500 -28925 13650 -27600
rect 17000 -27650 17150 -25150
rect 17250 -27700 17400 -25150
rect 17500 -27650 17650 -25150
rect 17750 -27625 17900 -25100
rect 18000 -26025 18150 -25050
rect 18250 -26150 18400 -24975
rect 18500 -26175 18650 -24875
rect 18000 -27600 18150 -26175
rect 18750 -26200 18900 -24750
rect 18250 -27550 18400 -26300
rect 18500 -27500 18650 -26325
rect 18750 -27450 18900 -26400
rect 19000 -27425 19150 -24600
rect 19250 -27375 19400 -24425
rect 19500 -27350 19650 -24225
rect 19750 -27325 19900 -24050
rect 20000 -27300 20150 -24125
rect 20250 -27200 20400 -24250
rect 20500 -27175 20650 -24200
rect 20750 -25250 20900 -23950
rect 21000 -24500 21150 -23800
rect 21250 -24900 21400 -23725
rect 21000 -25400 21150 -25250
rect 21250 -25325 21400 -25175
rect 20750 -27100 20900 -25625
rect 21000 -27050 21150 -25575
rect 21250 -26950 21400 -25475
rect 21500 -26825 21650 -24000
rect 21750 -24125 21900 -22025
rect 24250 -22050 24400 -21675
rect 24500 -22025 24650 -21575
rect 24750 -22000 24900 -21425
rect 25000 -21550 25150 -21175
rect 25250 -21625 25400 -21200
rect 25500 -21500 25650 -20475
rect 25750 -21300 25900 -19575
rect 26000 -20950 26150 -10125
rect 26250 -20475 26400 -10325
rect 26500 -10375 26650 -9400
rect 26500 -19800 26650 -10625
rect 26750 -10650 26900 -9600
rect 26750 -19000 26900 -10900
rect 27000 -10950 27150 -9825
rect 27000 -18050 27150 -11225
rect 27250 -11275 27400 -10100
rect 27500 -11550 27650 -10375
rect 27250 -15400 27400 -11575
rect 27750 -11725 27900 -10675
rect 27500 -12175 27650 -11750
rect 28000 -11850 28150 -10925
rect 27750 -12400 27900 -12250
rect 28000 -12400 28150 -12100
rect 28250 -12400 28400 -11175
rect 28500 -12375 28650 -11375
rect 28750 -12400 28900 -11550
rect 27250 -16400 27400 -16150
rect 22000 -23725 22150 -22075
rect 22250 -23200 22400 -22150
rect 25250 -22200 25400 -21875
rect 25500 -22125 25650 -21700
rect 25750 -21775 25900 -21550
rect 22500 -22575 22650 -22425
rect 23000 -23900 23150 -23650
rect 22250 -24500 22400 -24325
rect 22500 -24425 22650 -24200
rect 22750 -24225 22900 -23925
rect 21750 -26675 21900 -24725
rect 22000 -24825 22150 -24600
rect 22250 -25300 22400 -24650
rect 22000 -26475 22150 -25300
rect 22500 -25425 22650 -24600
rect 22750 -25500 22900 -24500
rect 23000 -25100 23150 -24150
rect 23250 -24725 23400 -23825
rect 23500 -24400 23650 -23425
rect 23750 -23525 23900 -23025
rect 24250 -23650 24400 -23325
rect 24500 -23450 24650 -22600
rect 24750 -23200 24900 -22325
rect 25000 -22825 25150 -22325
rect 25250 -22600 25400 -22450
rect 24000 -23875 24150 -23725
rect 23750 -24100 23900 -23900
rect 24250 -24175 24400 -24025
rect 24500 -24300 24650 -23775
rect 23000 -25500 23150 -25275
rect 23250 -25450 23400 -25075
rect 23500 -25350 23650 -24825
rect 23750 -25275 23900 -24525
rect 24000 -25125 24150 -24375
rect 24750 -24500 24900 -23525
rect 25000 -24325 25150 -23225
rect 25250 -23975 25400 -22900
rect 25500 -23275 25650 -22850
rect 25750 -22900 25900 -22200
rect 24250 -25000 24400 -24525
rect 22250 -26150 22400 -25575
rect 13000 -35950 13150 -34675
rect 13250 -34700 13400 -29025
rect 13750 -29100 13900 -27850
rect 13500 -34925 13650 -29200
rect 14000 -29250 14150 -28025
rect 17000 -28100 17150 -27950
rect 17250 -28125 17400 -27900
rect 13250 -35875 13400 -34925
rect 13750 -35100 13900 -29375
rect 14250 -29400 14400 -28175
rect 17500 -28200 17650 -27875
rect 13500 -35850 13650 -35100
rect 14000 -35300 14150 -29550
rect 14500 -29600 14650 -28300
rect 14750 -29725 14900 -28375
rect 14250 -34250 14400 -29725
rect 14500 -34275 14650 -29875
rect 15000 -29900 15150 -28875
rect 17250 -29050 17400 -28375
rect 15250 -30025 15400 -29325
rect 17500 -29600 17650 -28350
rect 14750 -34450 14900 -30025
rect 15500 -30200 15650 -29600
rect 14250 -34750 14400 -34475
rect 14500 -34750 14650 -34450
rect 13750 -35800 13900 -35300
rect 14250 -35450 14400 -34950
rect 14000 -35750 14150 -35450
rect 14500 -35550 14650 -34950
rect 14750 -35450 14900 -34725
rect 15000 -35050 15150 -30225
rect 15750 -30325 15900 -29875
rect 15250 -34425 15400 -30375
rect 15500 -34050 15650 -30500
rect 15750 -33300 15900 -30650
rect 16000 -32575 16150 -30775
rect 16250 -31425 16400 -30850
rect 16500 -30950 16650 -30800
rect 16750 -31175 16900 -29975
rect 17000 -31525 17150 -30250
rect 17750 -30325 17900 -27850
rect 18000 -28250 18150 -27775
rect 18250 -28275 18400 -27700
rect 18500 -28350 18650 -27650
rect 18750 -28375 18900 -27600
rect 16750 -31875 16900 -31600
rect 15250 -34725 15400 -34575
rect 14250 -35750 14400 -35600
rect 15000 -35700 15150 -35475
rect 15250 -35700 15400 -34875
rect 15500 -35700 15650 -34200
rect 15750 -35575 15900 -33850
rect 16000 -33875 16150 -32800
rect 16250 -34000 16400 -32125
rect 16500 -33850 16650 -31950
rect 17000 -32000 17150 -31850
rect 17250 -31950 17400 -30625
rect 18000 -30975 18150 -28400
rect 16750 -33600 16900 -32050
rect 17000 -33050 17150 -32150
rect 17500 -32250 17650 -31050
rect 18250 -31450 18400 -28425
rect 19000 -28475 19150 -27575
rect 17750 -32850 17900 -31500
rect 18500 -31825 18650 -28500
rect 17000 -33825 17150 -33200
rect 17250 -33700 17400 -32850
rect 17500 -33250 17650 -32975
rect 18000 -33275 18150 -32000
rect 18250 -32250 18400 -32100
rect 18750 -32200 18900 -28525
rect 19250 -28550 19400 -27550
rect 19500 -27850 19650 -27700
rect 19500 -28375 19650 -28225
rect 19750 -28325 19900 -27475
rect 19000 -32550 19150 -28625
rect 20000 -28750 20150 -27450
rect 19500 -29025 19650 -28875
rect 19250 -32600 19400 -29075
rect 19500 -32600 19650 -29175
rect 19750 -29200 19900 -29050
rect 20250 -29125 20400 -27350
rect 19750 -32600 19900 -29350
rect 20000 -32550 20150 -29450
rect 20500 -29475 20650 -27325
rect 20250 -32525 20400 -29675
rect 20750 -29825 20900 -27250
rect 20500 -32525 20650 -30050
rect 21000 -30175 21150 -27200
rect 21250 -30375 21400 -27100
rect 21500 -30200 21650 -27000
rect 21750 -29975 21900 -26875
rect 22000 -29700 22150 -26700
rect 22250 -29425 22400 -26400
rect 22500 -29100 22650 -26075
rect 22750 -28750 22900 -25800
rect 23000 -28425 23150 -25750
rect 23250 -28075 23400 -25725
rect 23500 -27600 23650 -25675
rect 23750 -27200 23900 -25600
rect 24000 -26625 24150 -25475
rect 21000 -30875 21150 -30600
rect 21250 -31750 21400 -30625
rect 20750 -32500 20900 -32075
rect 21500 -32500 21650 -30450
rect 21750 -32475 21900 -30250
rect 22000 -32475 22150 -30000
rect 22250 -32475 22400 -29725
rect 22500 -32550 22650 -29400
rect 22750 -32675 22900 -29050
rect 23000 -31150 23150 -28725
rect 23250 -31000 23400 -28375
rect 23500 -29400 23650 -27975
rect 23750 -29025 23900 -27500
rect 24000 -27700 24150 -27475
rect 24250 -27525 24400 -25325
rect 24500 -27225 24650 -25175
rect 24750 -26800 24900 -24975
rect 25000 -26375 25150 -24750
rect 25250 -25950 25400 -24475
rect 25500 -25500 25650 -24100
rect 25750 -25025 25900 -23475
rect 26000 -24550 26150 -21800
rect 26250 -24050 26400 -21350
rect 26500 -23525 26650 -20350
rect 26750 -22875 26900 -19650
rect 27000 -22175 27150 -19675
rect 26750 -24325 26900 -23700
rect 27000 -24100 27150 -22950
rect 27250 -23925 27400 -17650
rect 27500 -23700 27650 -12400
rect 29000 -12425 29150 -11625
rect 29250 -12475 29400 -11725
rect 29500 -12500 29650 -11750
rect 29750 -12525 29900 -11800
rect 27750 -23500 27900 -12550
rect 28000 -16625 28150 -12550
rect 28000 -17050 28150 -16900
rect 28000 -23275 28150 -17200
rect 28250 -17300 28400 -12550
rect 28250 -23025 28400 -17700
rect 28500 -18000 28650 -12550
rect 28500 -18450 28650 -18300
rect 28500 -22750 28650 -18600
rect 28750 -18875 28900 -12575
rect 28750 -19175 28900 -19025
rect 29000 -19100 29150 -12600
rect 29250 -18775 29400 -12625
rect 30000 -12650 30150 -11850
rect 30250 -12625 30400 -11875
rect 29500 -18300 29650 -12650
rect 30500 -12675 30650 -11950
rect 29750 -18100 29900 -12675
rect 30750 -12750 30900 -12000
rect 30000 -17950 30150 -12800
rect 30250 -17725 30400 -12800
rect 31000 -12825 31150 -12075
rect 30500 -17525 30650 -12850
rect 31250 -12900 31400 -12150
rect 30750 -17300 30900 -12900
rect 31500 -13000 31650 -12225
rect 31000 -17125 31150 -13000
rect 31250 -17000 31400 -13075
rect 31750 -13125 31900 -12325
rect 31500 -16825 31650 -13200
rect 32000 -13250 32150 -12425
rect 31750 -16650 31900 -13300
rect 32250 -13350 32400 -12525
rect 32000 -16500 32150 -13425
rect 32500 -13450 32650 -12650
rect 32250 -16375 32400 -13550
rect 32750 -13575 32900 -12750
rect 32500 -16250 32650 -13675
rect 33000 -13750 33150 -12875
rect 32750 -16125 32900 -13825
rect 33250 -13850 33400 -12975
rect 33000 -15950 33150 -13925
rect 33500 -13975 33650 -13100
rect 33750 -14050 33900 -13200
rect 33250 -15850 33400 -14050
rect 34000 -14150 34150 -13300
rect 33500 -15750 33650 -14150
rect 34250 -14225 34400 -13375
rect 33750 -15650 33900 -14250
rect 34500 -14300 34650 -13450
rect 34000 -15575 34150 -14325
rect 34750 -14375 34900 -13525
rect 35000 -14425 35150 -13575
rect 34250 -15450 34400 -14425
rect 35250 -14450 35400 -13625
rect 35500 -14475 35650 -13675
rect 34500 -15300 34650 -14475
rect 35750 -14500 35900 -13725
rect 36000 -14525 36150 -13775
rect 36250 -14475 36400 -13800
rect 36500 -14425 36650 -13875
rect 36750 -14450 36900 -13950
rect 34750 -15200 34900 -14550
rect 35000 -15050 35150 -14600
rect 35250 -14925 35400 -14675
rect 35500 -14850 35650 -14700
rect 30500 -17925 30650 -17775
rect 30750 -17950 30900 -17550
rect 31000 -18050 31150 -17350
rect 28750 -20100 28900 -19950
rect 28750 -22325 28900 -20275
rect 29000 -20475 29150 -19450
rect 29250 -19950 29400 -19075
rect 29500 -20025 29650 -18750
rect 29750 -20100 29900 -18425
rect 30000 -19025 30150 -18200
rect 30250 -18850 30400 -18150
rect 30500 -18650 30650 -18100
rect 30750 -18425 30900 -18125
rect 30000 -20050 30150 -19200
rect 30500 -19375 30650 -18850
rect 30250 -19950 30400 -19375
rect 30500 -19825 30650 -19600
rect 30750 -19650 30900 -18675
rect 29250 -20575 29400 -20150
rect 29250 -21100 29400 -20825
rect 29500 -21000 29650 -20275
rect 29750 -20925 29900 -20250
rect 30000 -20850 30150 -20225
rect 30250 -20575 30400 -20125
rect 30500 -20500 30650 -20000
rect 30750 -20400 30900 -19875
rect 31000 -20225 31150 -18450
rect 31250 -20050 31400 -17175
rect 31500 -19850 31650 -17000
rect 31750 -19625 31900 -16850
rect 32000 -19425 32150 -16725
rect 32250 -19200 32400 -16550
rect 32500 -18950 32650 -16425
rect 32750 -18700 32900 -16300
rect 33000 -18450 33150 -16175
rect 33250 -18200 33400 -16025
rect 33500 -17925 33650 -15925
rect 33750 -17675 33900 -15825
rect 34000 -17375 34150 -15725
rect 34250 -17075 34400 -15600
rect 34500 -16800 34650 -15500
rect 34750 -16525 34900 -15400
rect 35000 -16225 35150 -15275
rect 35250 -15800 35400 -15175
rect 35500 -15525 35650 -15075
rect 35750 -15275 35900 -14700
rect 36000 -15025 36150 -14700
rect 26500 -24500 26650 -24325
rect 26000 -25400 26150 -25250
rect 24000 -28775 24150 -27850
rect 24250 -28575 24400 -27975
rect 24500 -28425 24650 -27575
rect 24750 -28275 24900 -27125
rect 25000 -28050 25150 -26750
rect 25250 -27750 25400 -26300
rect 25500 -27350 25650 -25825
rect 25750 -26925 25900 -25400
rect 26000 -26525 26150 -25575
rect 26250 -26200 26400 -25075
rect 26500 -25900 26650 -24800
rect 26750 -25650 26900 -24550
rect 27000 -25375 27150 -24350
rect 27250 -25125 27400 -24125
rect 27500 -24900 27650 -23925
rect 27750 -24700 27900 -23725
rect 28000 -24475 28150 -23525
rect 28250 -24250 28400 -23300
rect 28500 -24050 28650 -22975
rect 28750 -23800 28900 -22750
rect 29000 -23525 29150 -21875
rect 29250 -23225 29400 -21275
rect 29500 -22750 29650 -21200
rect 29750 -22250 29900 -21100
rect 30000 -21925 30150 -21025
rect 30250 -21725 30400 -20900
rect 30500 -21600 30650 -20775
rect 30750 -21450 30900 -20625
rect 31000 -21325 31150 -20475
rect 31250 -21175 31400 -20275
rect 31500 -21000 31650 -20075
rect 31750 -20850 31900 -19875
rect 32000 -20600 32150 -19650
rect 32250 -20425 32400 -19425
rect 32500 -20200 32650 -19200
rect 32750 -19975 32900 -18975
rect 33000 -19750 33150 -18725
rect 33250 -19525 33400 -18450
rect 33500 -19275 33650 -18175
rect 33750 -19025 33900 -17925
rect 34000 -18750 34150 -17650
rect 34250 -18500 34400 -17350
rect 34500 -18175 34650 -17025
rect 34750 -17925 34900 -16800
rect 35000 -17625 35150 -16600
rect 35250 -17375 35400 -16275
rect 35500 -17100 35650 -15900
rect 35750 -16825 35900 -15600
rect 36000 -16500 36150 -15350
rect 36250 -16225 36400 -15100
rect 36500 -15900 36650 -14900
rect 36750 -15625 36900 -14725
rect 37000 -15300 37150 -14150
rect 23500 -30850 23650 -29850
rect 23750 -30700 23900 -29775
rect 24000 -30575 24150 -29650
rect 24250 -30425 24400 -29525
rect 24500 -30300 24650 -29400
rect 24750 -30150 24900 -29250
rect 25000 -30000 25150 -29125
rect 25250 -29850 25400 -29000
rect 25500 -29700 25650 -28900
rect 25750 -29575 25900 -28800
rect 26000 -29425 26150 -28750
rect 26250 -29300 26400 -28750
rect 26500 -29300 26650 -28775
rect 17500 -33550 17650 -33400
rect 17500 -33875 17650 -33700
rect 16000 -34400 16150 -34075
rect 16000 -35700 16150 -34550
rect 16250 -35725 16400 -34250
rect 16500 -35725 16650 -34100
rect 16750 -35750 16900 -33925
rect 17000 -35650 17150 -33975
rect 17250 -35475 17400 -33975
rect 17500 -35275 17650 -34125
rect 17750 -34475 17900 -33300
rect 18250 -33500 18400 -33075
rect 18500 -33800 18650 -32775
rect 19250 -32900 19400 -32750
rect 19500 -32900 19650 -32750
rect 19750 -32900 19900 -32750
rect 20000 -32900 20150 -32700
rect 20250 -32900 20400 -32750
rect 18750 -33700 18900 -33100
rect 19000 -33325 19150 -33175
rect 19250 -33275 19400 -33050
rect 18000 -34425 18150 -34050
rect 12750 -36650 12900 -36225
rect 13250 -36275 13400 -36025
rect 13500 -36350 13650 -36000
rect 13000 -36525 13150 -36350
rect 13750 -36400 13900 -35950
rect 11500 -37750 11650 -37575
rect 11750 -37725 11900 -37575
rect 12250 -37900 12400 -37475
rect 9500 -38625 9650 -38475
rect 9500 -39050 9650 -38825
rect 9750 -38900 9900 -38325
rect 2250 -42750 2400 -42250
rect 2000 -43700 2150 -42750
rect 2500 -42850 2650 -42100
rect 2250 -43375 2400 -42900
rect 2750 -43000 2900 -41950
rect 2500 -43150 2650 -43000
rect 1250 -44725 1400 -44575
rect 0 -49525 150 -48225
rect 250 -49600 400 -46850
rect 500 -49700 650 -46150
rect 750 -49750 900 -45850
rect 1000 -49800 1150 -45450
rect 1250 -49375 1400 -44950
rect 1500 -49375 1650 -44600
rect 1750 -49450 1900 -44300
rect 2000 -49500 2150 -43975
rect 2250 -49525 2400 -43750
rect 1250 -49850 1400 -49525
rect 1500 -49850 1650 -49525
rect 2500 -49600 2650 -43525
rect 2750 -49600 2900 -43300
rect 1750 -49900 1900 -49600
rect 3000 -49650 3150 -41825
rect 2000 -49925 2150 -49650
rect 3250 -49725 3400 -41700
rect 3500 -49725 3650 -41600
rect 3750 -49700 3900 -41500
rect 4000 -49725 4150 -41425
rect 4250 -49700 4400 -41400
rect 4500 -49700 4650 -41350
rect 4750 -49650 4900 -41275
rect 5000 -49600 5150 -41225
rect 5250 -49600 5400 -41150
rect 5500 -49625 5650 -41100
rect 5750 -49775 5900 -41025
rect 7750 -43725 7900 -40125
rect 8000 -42950 8150 -39950
rect 8250 -42375 8400 -39775
rect 8500 -41950 8650 -39600
rect 8750 -41450 8900 -39450
rect 7750 -44950 7900 -44050
rect 8000 -44950 8150 -43125
rect 8250 -44850 8400 -42550
rect 8500 -44775 8650 -42125
rect 8750 -44700 8900 -41700
rect 9000 -44775 9150 -39350
rect 8750 -49825 8900 -44850
rect 9000 -49175 9150 -45025
rect 9250 -45775 9400 -39275
rect 9250 -46075 9400 -45925
rect 9000 -49600 9150 -49325
rect 9250 -49475 9400 -46225
rect 9500 -46425 9650 -39250
rect 9500 -49275 9650 -46725
rect 9750 -46875 9900 -39150
rect 9750 -49075 9900 -47125
rect 10000 -47225 10150 -38250
rect 10000 -48850 10150 -47475
rect 10250 -47550 10400 -38150
rect 10500 -38500 10650 -38250
rect 10750 -38600 10900 -38125
rect 10250 -48575 10400 -47775
rect 10500 -47800 10650 -38650
rect 10750 -48050 10900 -38750
rect 10500 -48425 10650 -48050
rect 11000 -48175 11150 -37975
rect 11250 -38250 11400 -37925
rect 12500 -37950 12650 -37300
rect 12750 -37900 12900 -37125
rect 13000 -37900 13150 -36975
rect 11250 -43125 11400 -38525
rect 11500 -42025 11650 -38275
rect 11750 -41050 11900 -37975
rect 12000 -39775 12150 -37975
rect 12250 -39250 12400 -38050
rect 12500 -38625 12650 -38100
rect 12000 -40175 12150 -40025
rect 11500 -42350 11650 -42175
rect 11500 -43275 11650 -42650
rect 11250 -48075 11400 -43275
rect 11750 -43400 11900 -41425
rect 11500 -47950 11650 -43450
rect 12000 -43525 12150 -40350
rect 11750 -47800 11900 -43550
rect 12250 -43625 12400 -39650
rect 12000 -47650 12150 -43675
rect 12500 -43750 12650 -39175
rect 12250 -47475 12400 -43800
rect 12750 -43850 12900 -38800
rect 12500 -46825 12650 -43925
rect 13000 -43950 13150 -38250
rect 12750 -46625 12900 -44025
rect 13250 -44050 13400 -36850
rect 13000 -46425 13150 -44100
rect 13500 -44125 13650 -36750
rect 13750 -44200 13900 -36625
rect 13250 -46200 13400 -44200
rect 14000 -44275 14150 -35950
rect 13500 -46075 13650 -44300
rect 14250 -44350 14400 -35950
rect 14500 -44350 14650 -35900
rect 14750 -44300 14900 -35900
rect 15000 -44225 15150 -35950
rect 15250 -44200 15400 -35900
rect 15500 -44125 15650 -35925
rect 15750 -44075 15900 -35950
rect 16000 -44025 16150 -36000
rect 16250 -43950 16400 -36075
rect 16500 -43850 16650 -36050
rect 16750 -43725 16900 -36025
rect 17000 -43750 17150 -35900
rect 17250 -43775 17400 -35700
rect 17500 -43850 17650 -35500
rect 17750 -43900 17900 -35275
rect 18000 -43900 18150 -34950
rect 18250 -43850 18400 -34450
rect 18500 -43750 18650 -34325
rect 18750 -43775 18900 -33900
rect 19000 -43750 19150 -33850
rect 19250 -43650 19400 -33800
rect 19500 -43575 19650 -33475
rect 19750 -43475 19900 -33500
rect 20000 -43400 20150 -33300
rect 20250 -43275 20400 -33125
rect 20500 -43175 20650 -32950
rect 20750 -43050 20900 -32850
rect 21000 -42925 21150 -32775
rect 21250 -42800 21400 -32750
rect 21500 -42675 21650 -32750
rect 23000 -32825 23150 -31400
rect 23250 -31650 23400 -31175
rect 21750 -34975 21900 -32825
rect 22000 -34950 22150 -32850
rect 22250 -34925 22400 -32950
rect 23250 -32975 23400 -31850
rect 23500 -32250 23650 -31025
rect 22500 -34900 22650 -33000
rect 23500 -33100 23650 -32675
rect 23750 -32850 23900 -30900
rect 22750 -34700 22900 -33200
rect 23000 -33275 23150 -33125
rect 23000 -33575 23150 -33425
rect 23000 -34875 23150 -33725
rect 23250 -34525 23400 -33250
rect 24000 -33450 24150 -30750
rect 23500 -34400 23650 -33625
rect 23750 -33750 23900 -33525
rect 24000 -33800 24150 -33625
rect 23250 -35225 23400 -35075
rect 23500 -35200 23650 -34900
rect 21750 -42500 21900 -35375
rect 22000 -38825 22150 -35250
rect 22250 -38675 22400 -35225
rect 22500 -38575 22650 -35225
rect 22750 -38450 22900 -35225
rect 23000 -38275 23150 -35250
rect 23750 -35275 23900 -34000
rect 24000 -34100 24150 -33950
rect 24250 -34100 24400 -30600
rect 24500 -31550 24650 -30475
rect 24750 -31425 24900 -30325
rect 25000 -31300 25150 -30175
rect 25250 -31175 25400 -30025
rect 25500 -31025 25650 -29875
rect 25750 -31025 25900 -29750
rect 25000 -31700 25150 -31450
rect 25250 -31575 25400 -31325
rect 25500 -31475 25650 -31325
rect 26000 -31450 26150 -29600
rect 24000 -34750 24150 -34450
rect 24000 -35350 24150 -35075
rect 23250 -38125 23400 -35375
rect 23500 -37775 23650 -35350
rect 23750 -37275 23900 -35450
rect 24250 -35475 24400 -34450
rect 24500 -34700 24650 -31950
rect 25000 -32275 25150 -32125
rect 24750 -34800 24900 -32300
rect 25000 -32575 25150 -32425
rect 25250 -32525 25400 -31725
rect 25500 -32925 25650 -31675
rect 25750 -32475 25900 -31650
rect 26000 -32400 26150 -32000
rect 26250 -32075 26400 -29500
rect 26750 -29775 26900 -28875
rect 25750 -32775 25900 -32625
rect 25000 -34675 25150 -33075
rect 25250 -34550 25400 -33275
rect 25500 -34400 25650 -33200
rect 25750 -34275 25900 -33075
rect 26000 -34150 26150 -32950
rect 26250 -34025 26400 -32850
rect 26500 -33900 26650 -29850
rect 27000 -30400 27150 -29000
rect 26750 -33775 26900 -30475
rect 27250 -31000 27400 -29225
rect 27000 -33650 27150 -31075
rect 27500 -31450 27650 -29350
rect 27750 -30700 27900 -29350
rect 28000 -30225 28150 -29250
rect 28250 -29925 28400 -29150
rect 28500 -29750 28650 -29050
rect 28750 -29650 28900 -29000
rect 29000 -29625 29150 -28975
rect 29250 -29625 29400 -29000
rect 29500 -29700 29650 -29025
rect 27750 -31025 27900 -30875
rect 27250 -33525 27400 -31650
rect 27750 -32200 27900 -31300
rect 27500 -33400 27650 -32300
rect 28000 -32850 28150 -30500
rect 27750 -33250 27900 -32975
rect 24000 -36700 24150 -35525
rect 24250 -35950 24400 -35675
rect 24000 -37700 24150 -37000
rect 23500 -38350 23650 -38075
rect 23250 -38850 23400 -38425
rect 23500 -38850 23650 -38700
rect 22000 -42325 22150 -38975
rect 22250 -42100 22400 -38900
rect 23750 -38950 23900 -37825
rect 22500 -41900 22650 -38950
rect 22750 -41650 22900 -38950
rect 23000 -41450 23150 -38950
rect 23250 -41250 23400 -39075
rect 24000 -39150 24150 -38675
rect 23500 -41075 23650 -39175
rect 24250 -39275 24400 -36275
rect 23750 -40800 23900 -39275
rect 24000 -40500 24150 -39350
rect 24500 -39450 24650 -35000
rect 24250 -40250 24400 -39450
rect 24750 -39775 24900 -35050
rect 24500 -40000 24650 -39800
rect 23500 -41425 23650 -41275
rect 23000 -42225 23150 -41650
rect 23500 -41925 23650 -41600
rect 23750 -42025 23900 -41025
rect 24000 -41900 24150 -40725
rect 24250 -41725 24400 -40475
rect 24500 -41575 24650 -40225
rect 24750 -41375 24900 -39975
rect 25000 -41200 25150 -35000
rect 25250 -41000 25400 -34850
rect 25500 -40725 25650 -34700
rect 25750 -40350 25900 -34575
rect 26000 -34600 26150 -34450
rect 26250 -34650 26400 -34325
rect 26000 -40025 26150 -34750
rect 26500 -34850 26650 -34225
rect 26250 -39550 26400 -34925
rect 26750 -35000 26900 -34100
rect 26500 -38950 26650 -35100
rect 27000 -35150 27150 -33975
rect 26750 -38350 26900 -35325
rect 27250 -35550 27400 -33850
rect 27500 -35425 27650 -33700
rect 27750 -34925 27900 -33600
rect 28000 -33775 28150 -33450
rect 28000 -34925 28150 -34075
rect 28250 -34150 28400 -30175
rect 28500 -34200 28650 -29950
rect 28750 -32375 28900 -29800
rect 29000 -32100 29150 -29775
rect 29250 -32075 29400 -29775
rect 29750 -29875 29900 -29100
rect 29500 -32175 29650 -29900
rect 30000 -30100 30150 -29225
rect 27000 -37600 27150 -35575
rect 27500 -35725 27650 -35575
rect 27500 -38050 27650 -36350
rect 24750 -42375 24900 -41925
rect 25000 -42300 25150 -41675
rect 25250 -41750 25400 -41600
rect 13750 -46150 13900 -44375
rect 14000 -45850 14150 -44425
rect 14250 -45575 14400 -44500
rect 14500 -45375 14650 -44500
rect 13500 -46375 13650 -46225
rect 12500 -47350 12650 -46975
rect 12750 -47175 12900 -46825
rect 13000 -46950 13150 -46625
rect 13250 -46725 13400 -46450
rect 13750 -46650 13900 -46425
rect 14000 -46900 14150 -46175
rect 14250 -46975 14400 -45900
rect 14500 -46425 14650 -45525
rect 14750 -46150 14900 -44450
rect 15000 -45950 15150 -44400
rect 15250 -45750 15400 -44350
rect 15500 -45550 15650 -44300
rect 15750 -45350 15900 -44250
rect 16000 -45150 16150 -44200
rect 16250 -44950 16400 -44100
rect 16500 -44750 16650 -44050
rect 16750 -44550 16900 -43950
rect 17000 -44275 17150 -43925
rect 14750 -47200 14900 -46350
rect 15000 -47050 15150 -46150
rect 15250 -46900 15400 -45950
rect 15500 -46700 15650 -45750
rect 15750 -46525 15900 -45550
rect 16000 -46325 16150 -45350
rect 16250 -46150 16400 -45175
rect 16500 -46000 16650 -44975
rect 16750 -45825 16900 -44750
rect 17000 -45625 17150 -44525
rect 17250 -44600 17400 -44250
rect 17750 -44850 17900 -44425
rect 18500 -44775 18650 -44575
rect 18750 -44700 18900 -44375
rect 19250 -44525 19400 -44075
rect 19500 -44475 19650 -44000
rect 19750 -44450 19900 -43875
rect 20000 -44350 20150 -43800
rect 20250 -44350 20400 -43725
rect 20500 -44350 20650 -43500
rect 17250 -45425 17400 -44950
rect 17500 -45975 17650 -45725
rect 17750 -45850 17900 -45600
rect 18000 -45725 18150 -45350
rect 18250 -45600 18400 -45075
rect 18500 -45500 18650 -44975
rect 18750 -45400 18900 -44850
rect 19000 -45300 19150 -44750
rect 19250 -45225 19400 -44675
rect 19500 -44775 19650 -44625
rect 19750 -44775 19900 -44625
rect 19500 -45125 19650 -44925
rect 19750 -45075 19900 -44925
rect 20000 -44975 20150 -44500
rect 20250 -44875 20400 -44500
rect 20500 -44775 20650 -44500
rect 20750 -44625 20900 -43350
rect 21000 -44550 21150 -43250
rect 21250 -44425 21400 -43125
rect 21500 -44350 21650 -42975
rect 21750 -44300 21900 -42775
rect 22000 -44225 22150 -42875
rect 22250 -43075 22400 -42450
rect 22250 -43525 22400 -43375
rect 22500 -43525 22650 -42400
rect 22250 -44175 22400 -43675
rect 22750 -44075 22900 -42550
rect 24500 -42600 24650 -42450
rect 23000 -44100 23150 -42750
rect 23250 -44050 23400 -42950
rect 24250 -43000 24400 -42825
rect 23500 -44050 23650 -43200
rect 23750 -44000 23900 -43100
rect 24000 -43925 24150 -43225
rect 24250 -43450 24400 -43300
rect 24250 -44000 24400 -43850
rect 24500 -43950 24650 -43100
rect 24750 -43800 24900 -42800
rect 25000 -43850 25150 -42500
rect 25250 -43275 25400 -42275
rect 25750 -42625 25900 -40850
rect 26000 -40900 26150 -40475
rect 26250 -40500 26400 -40075
rect 26500 -40175 26650 -39650
rect 26750 -39875 26900 -39050
rect 27000 -39575 27150 -38250
rect 27250 -39325 27400 -38050
rect 27500 -39100 27650 -38400
rect 27750 -38500 27900 -35100
rect 27750 -38900 27900 -38750
rect 28000 -38825 28150 -35100
rect 26000 -41200 26150 -41050
rect 26250 -41100 26400 -40750
rect 26500 -40950 26650 -40400
rect 26750 -40900 26900 -40100
rect 26000 -41975 26150 -41425
rect 26250 -41525 26400 -41275
rect 25500 -43050 25650 -42900
rect 25500 -43750 25650 -43600
rect 25750 -43925 25900 -42775
rect 26000 -44100 26150 -42250
rect 26250 -44125 26400 -41850
rect 26500 -44050 26650 -41400
rect 26750 -43950 26900 -41100
rect 27000 -43850 27150 -39850
rect 27250 -41350 27400 -39575
rect 27500 -40925 27650 -39325
rect 27750 -40600 27900 -39100
rect 28000 -40350 28150 -38975
rect 27500 -41375 27650 -41225
rect 27750 -41350 27900 -40850
rect 28000 -41300 28150 -40525
rect 27250 -43800 27400 -41600
rect 27500 -43750 27650 -41550
rect 27750 -43700 27900 -41500
rect 28000 -41700 28150 -41550
rect 28000 -42250 28150 -41850
rect 28000 -42575 28150 -42425
rect 28000 -43650 28150 -42725
rect 28250 -43125 28400 -34325
rect 28500 -36525 28650 -34550
rect 28750 -35050 28900 -32650
rect 29000 -35375 29150 -32300
rect 28750 -35750 28900 -35375
rect 29000 -35700 29150 -35550
rect 28500 -37900 28650 -36750
rect 28500 -38200 28650 -38050
rect 28500 -43300 28650 -38350
rect 28750 -38900 28900 -35975
rect 28750 -43300 28900 -39150
rect 29000 -39425 29150 -35850
rect 29000 -43275 29150 -39725
rect 29250 -39850 29400 -32225
rect 29500 -36125 29650 -32450
rect 29750 -32500 29900 -30125
rect 29750 -36325 29900 -32775
rect 30000 -32850 30150 -30350
rect 30250 -30375 30400 -29400
rect 30000 -35850 30150 -33125
rect 30250 -33225 30400 -30600
rect 30500 -30625 30650 -29600
rect 30250 -35875 30400 -33500
rect 30500 -33575 30650 -30850
rect 30750 -30900 30900 -29825
rect 30500 -36050 30650 -33850
rect 30750 -33975 30900 -31125
rect 31000 -31225 31150 -30100
rect 30750 -35850 30900 -34250
rect 31000 -34425 31150 -31550
rect 31250 -31700 31400 -30325
rect 31500 -31750 31650 -30500
rect 31750 -31425 31900 -30625
rect 32000 -31300 32150 -30675
rect 32250 -31300 32400 -30725
rect 31000 -35450 31150 -34875
rect 31250 -35175 31400 -32150
rect 31500 -35375 31650 -32200
rect 30750 -36150 30900 -36000
rect 31000 -36075 31150 -35725
rect 31250 -35875 31400 -35725
rect 29250 -43200 29400 -40050
rect 29500 -40100 29650 -36325
rect 30000 -36500 30150 -36175
rect 29500 -43250 29650 -40275
rect 29750 -43275 29900 -36500
rect 30250 -36725 30400 -36325
rect 30000 -43250 30150 -36725
rect 30500 -36900 30650 -36350
rect 30750 -36725 30900 -36575
rect 30250 -41100 30400 -36925
rect 30500 -41100 30650 -37125
rect 30750 -37150 30900 -36875
rect 31000 -37375 31150 -36275
rect 30750 -41100 30900 -37375
rect 31000 -40950 31150 -37600
rect 31250 -37625 31400 -36025
rect 31500 -37875 31650 -35575
rect 31750 -35675 31900 -31625
rect 31750 -38225 31900 -35975
rect 32000 -36175 32150 -31450
rect 31250 -40600 31400 -38375
rect 31500 -40075 31650 -38400
rect 31750 -39225 31900 -38500
rect 32000 -39175 32150 -36525
rect 32250 -36825 32400 -31550
rect 32500 -31650 32650 -30850
rect 32250 -38775 32400 -37025
rect 32500 -37650 32650 -31975
rect 32750 -32250 32900 -30975
rect 32500 -38300 32650 -38100
rect 32500 -38600 32650 -38450
rect 32750 -38725 32900 -32500
rect 33000 -32950 33150 -31200
rect 32250 -39300 32400 -39000
rect 31500 -40375 31650 -40225
rect 30250 -41450 30400 -41300
rect 30500 -41400 30650 -41250
rect 30250 -43200 30400 -41600
rect 30500 -43150 30650 -41600
rect 30750 -43100 30900 -41250
rect 31000 -43050 31150 -41100
rect 31250 -43050 31400 -40850
rect 31500 -43050 31650 -40525
rect 31750 -43025 31900 -39375
rect 32000 -41000 32150 -39325
rect 32000 -43000 32150 -41300
rect 32250 -41325 32400 -39750
rect 32500 -41450 32650 -39250
rect 32750 -41450 32900 -38950
rect 33000 -41325 33150 -33300
rect 33250 -33850 33400 -31525
rect 33250 -35700 33400 -34350
rect 33500 -35450 33650 -32025
rect 33250 -41100 33400 -35850
rect 33750 -35900 33900 -32700
rect 34000 -35725 34150 -33650
rect 34250 -35600 34400 -34550
rect 34500 -35500 34650 -34800
rect 34750 -35500 34900 -34925
rect 33500 -38675 33650 -36475
rect 33500 -40825 33650 -38850
rect 33750 -38875 33900 -36400
rect 33750 -39725 33900 -39275
rect 33750 -40100 33900 -39950
rect 32250 -43000 32400 -41500
rect 32500 -43000 32650 -41600
rect 32750 -42850 32900 -41600
rect 33000 -42575 33150 -41500
rect 33250 -42525 33400 -41325
rect 33500 -42300 33650 -41000
rect 33750 -41925 33900 -40350
rect 34000 -41625 34150 -35900
rect 34250 -41050 34400 -35750
rect 34500 -41275 34650 -35675
rect 34750 -40625 34900 -35700
rect 35000 -35925 35150 -35050
rect 35000 -36375 35150 -36175
rect 35000 -38850 35150 -36775
rect 35000 -39575 35150 -39250
rect 35000 -39875 35150 -39725
rect 33500 -42975 33650 -42575
rect 33750 -43025 33900 -42350
rect 34000 -43050 34150 -42400
rect 34250 -43050 34400 -42075
rect 34500 -43000 34650 -41625
rect 34750 -42925 34900 -40775
rect 35000 -42800 35150 -40025
rect 35250 -42625 35400 -35200
rect 35500 -42425 35650 -35500
rect 35750 -40075 35900 -36025
rect 35750 -42250 35900 -40875
rect 36000 -42025 36150 -40875
rect 36250 -41825 36400 -40750
rect 36500 -41600 36650 -40575
rect 36750 -41300 36900 -40425
rect 37000 -41125 37150 -40225
rect 37250 -41000 37400 -40050
rect 37500 -40800 37650 -39850
rect 37750 -40600 37900 -39675
rect 38000 -40425 38150 -39450
rect 38250 -40225 38400 -39250
rect 38500 -40025 38650 -39050
rect 38750 -39800 38900 -38850
rect 39000 -39625 39150 -38650
rect 39250 -39400 39400 -38450
rect 39500 -39200 39650 -38300
rect 39750 -39000 39900 -38200
rect 40000 -38775 40150 -38125
rect 40250 -38525 40400 -38125
rect 28250 -43600 28400 -43375
rect 15750 -47500 15900 -46725
rect 11250 -48400 11400 -48250
rect 11500 -48275 11650 -48125
rect 10500 -49900 10650 -48700
rect 10750 -49775 10900 -48500
rect 11000 -49650 11150 -48550
rect 16000 -48675 16150 -46550
rect 16000 -49100 16150 -48825
rect 23500 -49925 23650 -44300
rect 24750 -44350 24900 -44200
rect 23750 -49575 23900 -44425
rect 24000 -49200 24150 -44400
rect 24250 -48825 24400 -44675
rect 24500 -47525 24650 -44550
rect 24750 -47425 24900 -44875
rect 25250 -45050 25400 -44900
rect 25000 -47275 25150 -45050
rect 25250 -46900 25400 -45900
rect 25500 -45950 25650 -44750
rect 25500 -47300 25650 -46200
rect 24500 -48500 24650 -47675
rect 24750 -48175 24900 -47575
rect 24250 -49600 24400 -49100
rect 24500 -49275 24650 -48725
rect 25000 -49225 25150 -48875
rect 25250 -49150 25400 -48000
rect 25500 -49050 25650 -47800
rect 25750 -48950 25900 -44700
rect 26000 -48800 26150 -44425
rect 26250 -48675 26400 -44325
rect 26500 -48525 26650 -44225
rect 26750 -48400 26900 -44125
rect 27000 -48225 27150 -44050
rect 27250 -48050 27400 -43950
rect 27500 -47875 27650 -43900
rect 27750 -47650 27900 -43850
rect 28000 -47425 28150 -43800
rect 28250 -47200 28400 -43750
rect 28500 -46975 28650 -43700
rect 28750 -46775 28900 -43700
rect 29000 -46575 29150 -43650
rect 29250 -46375 29400 -43575
rect 29500 -46200 29650 -43550
rect 29750 -45975 29900 -43475
rect 30000 -45775 30150 -43425
rect 30250 -45600 30400 -43350
rect 30500 -45400 30650 -43300
rect 30750 -45200 30900 -43300
rect 31000 -45025 31150 -43250
rect 31250 -44800 31400 -43225
rect 31500 -44625 31650 -43200
rect 31750 -44425 31900 -43175
rect 32000 -44150 32150 -43150
rect 32250 -43900 32400 -43150
rect 32500 -43725 32650 -43150
rect 32750 -43550 32900 -43150
rect 33000 -43350 33150 -43150
rect 34000 -43600 34150 -43325
rect 34250 -43450 34400 -43300
rect 36000 -48575 36150 -42350
rect 36250 -48950 36400 -42175
rect 36500 -48475 36650 -41950
rect 36750 -48450 36900 -41675
rect 37000 -48450 37150 -41425
rect 37250 -48450 37400 -41200
rect 37500 -48450 37650 -41100
rect 37750 -48450 37900 -40925
rect 38000 -48475 38150 -40600
rect 38250 -45900 38400 -40425
rect 38500 -45825 38650 -40225
rect 38250 -48575 38400 -46225
rect 38750 -47350 38900 -40050
rect 38500 -48150 38650 -47400
rect 38500 -48500 38650 -48300
rect 38750 -48550 38900 -47500
rect 36500 -49200 36650 -48625
rect 36750 -49350 36900 -48600
rect 37000 -49525 37150 -48600
rect 37250 -49700 37400 -48600
rect 37500 -49800 37650 -48600
rect 37750 -49900 37900 -48600
rect 39000 -48725 39150 -39825
rect 39250 -49000 39400 -39600
rect 39500 -47125 39650 -39400
rect 39750 -45700 39900 -39200
rect 39500 -47425 39650 -47275
rect 39500 -47850 39650 -47650
rect 39500 -48250 39650 -48050
rect 39750 -48700 39900 -46425
rect 40000 -46450 40150 -38975
rect 40500 -39625 40650 -38175
rect 40500 -40200 40650 -39775
rect 40750 -40125 40900 -38300
rect 41000 -40175 41150 -38550
rect 41250 -40150 41400 -38875
rect 41500 -40125 41650 -39125
rect 41750 -40050 41900 -39225
rect 42000 -40025 42150 -39250
rect 42250 -40000 42400 -39250
rect 42500 -39975 42650 -39200
rect 42750 -39950 42900 -39200
rect 43000 -39950 43150 -39175
rect 43250 -39925 43400 -39150
rect 43500 -39875 43650 -39125
rect 43750 -39850 43900 -39100
rect 44000 -39825 44150 -39075
rect 44250 -39800 44400 -39050
rect 44500 -39800 44650 -39025
rect 44750 -39775 44900 -39000
rect 45000 -39775 45150 -39000
rect 45250 -39775 45400 -39000
rect 45500 -39775 45650 -39000
rect 45750 -39775 45900 -39000
rect 46000 -39775 46150 -38975
rect 46250 -39750 46400 -38950
rect 46500 -39750 46650 -38950
rect 46750 -39750 46900 -38950
rect 47000 -39750 47150 -38950
rect 47250 -39750 47400 -38950
rect 47500 -39750 47650 -38950
rect 47750 -39725 47900 -38925
rect 48000 -39700 48150 -38900
rect 48250 -39650 48400 -38850
rect 48500 -39600 48650 -38800
rect 48750 -39550 48900 -38775
rect 49250 -39425 49400 -38625
rect 49500 -39350 49650 -38550
rect 49750 -39300 49900 -38475
rect 40750 -40525 40900 -40350
rect 41000 -40525 41150 -40375
rect 40000 -46975 40150 -46725
rect 40000 -48650 40150 -47250
rect 39000 -49200 39150 -49050
rect 39250 -49650 39400 -49250
<< end >>
