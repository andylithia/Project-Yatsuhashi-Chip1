magic
tech sky130A
timestamp 1659233347
<< metal1 >>
rect -100 550 500 600
rect -100 50 -50 550
rect 450 450 500 550
rect 50 400 500 450
rect 50 50 100 400
rect -100 0 100 50
<< via1 >>
rect -50 450 450 550
rect -50 50 50 450
<< metal2 >>
rect -100 550 500 600
rect -100 50 -50 550
rect 450 450 500 550
rect 50 400 500 450
rect 50 50 100 400
rect -100 0 100 50
<< via2 >>
rect -50 450 450 550
rect -50 50 50 450
<< metal3 >>
rect -100 550 500 600
rect -100 50 -50 550
rect 450 450 500 550
rect 50 400 500 450
rect 50 50 100 400
rect -100 0 100 50
<< via3 >>
rect -50 450 450 550
rect -50 50 50 450
<< metal4 >>
rect -100 550 500 600
rect -100 50 -50 550
rect 450 450 500 550
rect 150 400 500 450
rect 150 350 200 400
rect 50 300 200 350
rect 50 50 100 300
rect -100 0 100 50
<< via4 >>
rect -50 450 150 550
rect -50 350 50 450
rect 50 350 150 450
<< metal5 >>
rect -100 550 500 600
rect -100 350 -50 550
rect 150 400 500 550
rect 150 350 200 400
rect -100 300 200 350
rect -100 0 100 300
<< end >>
