magic
tech sky130A
magscale 1 2
timestamp 1620310959
