magic
tech sky130B
magscale 1 2
timestamp 1660524083
<< metal4 >>
rect -35900 -22112 -27500 -22000
rect -35900 -23888 -29388 -22112
rect -27612 -23888 -27500 -22112
rect -35900 -24000 -27500 -23888
<< via4 >>
rect -29388 -23888 -27612 -22112
<< metal5 >>
tri -31012 -8675 -28337 -6000 se
rect -28337 -8000 -14263 -6000
tri -14263 -8000 -12263 -6000 sw
rect -28337 -8675 -28184 -8000
tri -28184 -8675 -27509 -8000 nw
tri -15091 -8600 -14491 -8000 ne
rect -14491 -8600 -12263 -8000
tri -27336 -8675 -27261 -8600 se
rect -27261 -8675 -15339 -8600
tri -32700 -10363 -31012 -8675 se
rect -31012 -9523 -29032 -8675
tri -29032 -9523 -28184 -8675 nw
tri -28184 -9523 -27336 -8675 se
rect -27336 -9448 -15339 -8675
tri -15339 -9448 -14491 -8600 sw
tri -14491 -9448 -13643 -8600 ne
rect -13643 -9448 -12263 -8600
rect -27336 -9523 -14491 -9448
rect -31012 -10363 -29880 -9523
tri -32928 -10591 -32700 -10363 se
rect -32700 -10371 -29880 -10363
tri -29880 -10371 -29032 -9523 nw
tri -29032 -10371 -28184 -9523 se
rect -28184 -9752 -14491 -9523
tri -14491 -9752 -14187 -9448 sw
tri -13643 -9752 -13339 -9448 ne
rect -13339 -9752 -12263 -9448
rect -28184 -10371 -14187 -9752
rect -32700 -10591 -30109 -10371
tri -35528 -13191 -32928 -10591 se
rect -32928 -10600 -30109 -10591
tri -30109 -10600 -29880 -10371 nw
tri -29261 -10600 -29032 -10371 se
rect -29032 -10600 -14187 -10371
tri -14187 -10600 -13339 -9752 sw
tri -13339 -10600 -12491 -9752 ne
rect -12491 -10600 -12263 -9752
tri -12263 -10600 -9663 -8000 sw
rect -32928 -11439 -30948 -10600
tri -30948 -11439 -30109 -10600 nw
tri -30100 -11439 -29261 -10600 se
rect -29261 -11200 -27032 -10600
tri -27032 -11200 -26432 -10600 nw
tri -16168 -11200 -15568 -10600 ne
rect -15568 -11200 -13339 -10600
rect -29261 -11439 -27880 -11200
rect -32928 -12287 -31796 -11439
tri -31796 -12287 -30948 -11439 nw
tri -30948 -12287 -30100 -11439 se
rect -30100 -12048 -27880 -11439
tri -27880 -12048 -27032 -11200 nw
tri -27032 -12048 -26184 -11200 se
rect -26184 -12048 -16416 -11200
tri -16416 -12048 -15568 -11200 sw
tri -15568 -12048 -14720 -11200 ne
rect -14720 -11448 -13339 -11200
tri -13339 -11448 -12491 -10600 sw
tri -12491 -11448 -11643 -10600 ne
rect -11643 -11448 -9663 -10600
rect -14720 -11504 -12491 -11448
tri -12491 -11504 -12435 -11448 sw
tri -11643 -11504 -11587 -11448 ne
rect -11587 -11504 -9663 -11448
rect -14720 -12048 -12435 -11504
rect -30100 -12287 -28184 -12048
rect -32928 -12352 -31861 -12287
tri -31861 -12352 -31796 -12287 nw
tri -31013 -12352 -30948 -12287 se
rect -30948 -12352 -28184 -12287
tri -28184 -12352 -27880 -12048 nw
tri -27336 -12352 -27032 -12048 se
rect -27032 -12352 -15568 -12048
tri -15568 -12352 -15264 -12048 sw
tri -14720 -12352 -14416 -12048 ne
rect -14416 -12352 -12435 -12048
tri -12435 -12352 -11587 -11504 sw
tri -11587 -12352 -10739 -11504 ne
rect -10739 -12352 -9663 -11504
rect -32928 -13191 -32700 -12352
tri -32700 -13191 -31861 -12352 nw
tri -31852 -13191 -31013 -12352 se
rect -31013 -13191 -29032 -12352
tri -37300 -14963 -35528 -13191 se
rect -35528 -14039 -33548 -13191
tri -33548 -14039 -32700 -13191 nw
tri -32700 -14039 -31852 -13191 se
rect -31852 -13200 -29032 -13191
tri -29032 -13200 -28184 -12352 nw
tri -28184 -13200 -27336 -12352 se
rect -27336 -13200 -15264 -12352
tri -15264 -13200 -14416 -12352 sw
tri -14416 -13200 -13568 -12352 ne
rect -13568 -13200 -11587 -12352
tri -11587 -13200 -10739 -12352 sw
tri -10739 -13200 -9891 -12352 ne
rect -9891 -13200 -9663 -12352
tri -9663 -13200 -7063 -10600 sw
rect -31852 -14039 -29880 -13200
rect -35528 -14268 -33777 -14039
tri -33777 -14268 -33548 -14039 nw
tri -32929 -14268 -32700 -14039 se
rect -32700 -14048 -29880 -14039
tri -29880 -14048 -29032 -13200 nw
tri -29032 -14048 -28184 -13200 se
rect -32700 -14268 -30100 -14048
tri -30100 -14268 -29880 -14048 nw
tri -29252 -14268 -29032 -14048 se
rect -29032 -14268 -28184 -14048
rect -35528 -14963 -34625 -14268
rect -37300 -15116 -34625 -14963
tri -34625 -15116 -33777 -14268 nw
tri -33777 -15116 -32929 -14268 se
rect -32929 -15116 -30948 -14268
tri -30948 -15116 -30100 -14268 nw
tri -30100 -15116 -29252 -14268 se
rect -29252 -15116 -28184 -14268
rect -37300 -16000 -35300 -15116
tri -35300 -15791 -34625 -15116 nw
tri -34452 -15791 -33777 -15116 se
rect -33777 -15791 -31796 -15116
rect -39300 -18000 -35300 -16000
tri -34700 -16039 -34452 -15791 se
rect -34452 -15964 -31796 -15791
tri -31796 -15964 -30948 -15116 nw
tri -30948 -15964 -30100 -15116 se
rect -30100 -15964 -28184 -15116
rect -34452 -16039 -32100 -15964
rect -34700 -16268 -32100 -16039
tri -32100 -16268 -31796 -15964 nw
tri -31252 -16268 -30948 -15964 se
rect -30948 -16029 -28184 -15964
tri -28184 -16029 -25355 -13200 nw
tri -17245 -16029 -14416 -13200 ne
tri -14416 -14048 -13568 -13200 sw
tri -13568 -14048 -12720 -13200 ne
rect -12720 -14048 -10739 -13200
tri -10739 -14048 -9891 -13200 sw
tri -9891 -14048 -9043 -13200 ne
rect -9043 -14048 -7063 -13200
rect -14416 -14268 -13568 -14048
tri -13568 -14268 -13348 -14048 sw
tri -12720 -14268 -12500 -14048 ne
rect -12500 -14268 -9891 -14048
tri -9891 -14268 -9671 -14048 sw
tri -9043 -14268 -8823 -14048 ne
rect -8823 -14268 -7063 -14048
rect -14416 -15116 -13348 -14268
tri -13348 -15116 -12500 -14268 sw
tri -12500 -15116 -11652 -14268 ne
rect -11652 -15116 -9671 -14268
tri -9671 -15116 -8823 -14268 sw
tri -8823 -15116 -7975 -14268 ne
rect -7975 -14963 -7063 -14268
tri -7063 -14963 -5300 -13200 sw
rect -7975 -15116 -5300 -14963
rect -14416 -15964 -12500 -15116
tri -12500 -15964 -11652 -15116 sw
tri -11652 -15964 -10804 -15116 ne
rect -10804 -15791 -8823 -15116
tri -8823 -15791 -8148 -15116 sw
tri -7975 -15791 -7300 -15116 ne
rect -10804 -15964 -8148 -15791
rect -14416 -16029 -11652 -15964
rect -30948 -16268 -30100 -16029
rect -34700 -25571 -32700 -16268
tri -32700 -16868 -32100 -16268 nw
tri -32100 -17116 -31252 -16268 se
rect -31252 -17116 -30100 -16268
rect -32100 -24494 -30100 -17116
tri -30100 -17945 -28184 -16029 nw
tri -14416 -17945 -12500 -16029 ne
rect -12500 -16268 -11652 -16029
tri -11652 -16268 -11348 -15964 sw
tri -10804 -16268 -10500 -15964 ne
rect -10500 -16039 -8148 -15964
tri -8148 -16039 -7900 -15791 sw
rect -10500 -16268 -7900 -16039
rect -12500 -17116 -11348 -16268
tri -11348 -17116 -10500 -16268 sw
tri -10500 -16868 -9900 -16268 ne
rect -29500 -22112 -27500 -22000
rect -29500 -23888 -29388 -22112
rect -27612 -23888 -27500 -22112
tri -30100 -24494 -29500 -23894 sw
rect -29500 -24000 -27500 -23888
rect -32100 -24722 -29500 -24494
tri -32700 -25571 -32100 -24971 sw
tri -32100 -25571 -31251 -24722 ne
rect -31251 -24796 -29500 -24722
tri -29500 -24796 -29198 -24494 sw
tri -29145 -24796 -28349 -24000 ne
rect -28349 -24796 -27500 -24000
rect -31251 -25571 -29198 -24796
rect -34700 -25645 -32100 -25571
tri -32100 -25645 -32026 -25571 sw
tri -31251 -25645 -31177 -25571 ne
rect -31177 -25645 -29198 -25571
tri -29198 -25645 -28349 -24796 sw
tri -28349 -25645 -27500 -24796 ne
tri -27500 -25645 -24672 -22817 sw
tri -13655 -23972 -12500 -22817 se
rect -12500 -23645 -10500 -17116
rect -12500 -23972 -11349 -23645
tri -15328 -25645 -13655 -23972 se
rect -13655 -24494 -11349 -23972
tri -11349 -24494 -10500 -23645 nw
tri -10500 -24494 -9900 -23894 se
rect -9900 -24494 -7900 -16268
rect -13655 -24796 -11651 -24494
tri -11651 -24796 -11349 -24494 nw
tri -10802 -24796 -10500 -24494 se
rect -10500 -24722 -7900 -24494
rect -10500 -24796 -8749 -24722
rect -13655 -25645 -12500 -24796
tri -12500 -25645 -11651 -24796 nw
tri -11651 -25645 -10802 -24796 se
rect -10802 -25571 -8749 -24796
tri -8749 -25571 -7900 -24722 nw
tri -7900 -25571 -7300 -24971 se
rect -7300 -25571 -5300 -15116
rect -10802 -25645 -8823 -25571
tri -8823 -25645 -8749 -25571 nw
tri -7974 -25645 -7900 -25571 se
rect -7900 -25645 -5300 -25571
rect -34700 -25799 -32026 -25645
tri -34700 -26800 -33699 -25799 ne
rect -33699 -26494 -32026 -25799
tri -32026 -26494 -31177 -25645 sw
tri -31177 -26494 -30328 -25645 ne
rect -30328 -26494 -28349 -25645
tri -28349 -26494 -27500 -25645 sw
tri -27500 -26494 -26651 -25645 ne
rect -26651 -26494 -24672 -25645
rect -33699 -26800 -31177 -26494
tri -31177 -26800 -30871 -26494 sw
tri -30328 -26800 -30022 -26494 ne
rect -30022 -26800 -27500 -26494
tri -27500 -26800 -27194 -26494 sw
tri -26651 -26800 -26345 -26494 ne
rect -26345 -26800 -24672 -26494
tri -24672 -26800 -23517 -25645 sw
tri -16483 -26800 -15328 -25645 se
rect -15328 -26494 -13349 -25645
tri -13349 -26494 -12500 -25645 nw
tri -12500 -26494 -11651 -25645 se
rect -11651 -26494 -9672 -25645
tri -9672 -26494 -8823 -25645 nw
tri -8823 -26494 -7974 -25645 se
rect -7974 -25799 -5300 -25645
rect -7974 -26494 -7300 -25799
rect -15328 -26800 -13655 -26494
tri -13655 -26800 -13349 -26494 nw
tri -12806 -26800 -12500 -26494 se
rect -12500 -26722 -9900 -26494
tri -9900 -26722 -9672 -26494 nw
tri -9051 -26722 -8823 -26494 se
rect -8823 -26722 -7300 -26494
rect -12500 -26800 -10749 -26722
tri -33699 -29400 -31099 -26800 ne
rect -31099 -27649 -30871 -26800
tri -30871 -27649 -30022 -26800 sw
tri -30022 -27649 -29173 -26800 ne
rect -29173 -27649 -27194 -26800
tri -27194 -27649 -26345 -26800 sw
tri -26345 -27649 -25496 -26800 ne
rect -25496 -27649 -14504 -26800
tri -14504 -27649 -13655 -26800 nw
tri -13655 -27649 -12806 -26800 se
rect -12806 -27571 -10749 -26800
tri -10749 -27571 -9900 -26722 nw
tri -9900 -27571 -9051 -26722 se
rect -9051 -27571 -7300 -26722
rect -12806 -27649 -10827 -27571
tri -10827 -27649 -10749 -27571 nw
tri -9978 -27649 -9900 -27571 se
rect -9900 -27649 -7300 -27571
rect -31099 -28498 -30022 -27649
tri -30022 -28498 -29173 -27649 sw
tri -29173 -28498 -28324 -27649 ne
rect -28324 -27951 -26345 -27649
tri -26345 -27951 -26043 -27649 sw
tri -25496 -27951 -25194 -27649 ne
rect -25194 -27951 -14806 -27649
tri -14806 -27951 -14504 -27649 nw
tri -13957 -27951 -13655 -27649 se
rect -13655 -27951 -11651 -27649
rect -28324 -28498 -26043 -27951
rect -31099 -28551 -29173 -28498
tri -29173 -28551 -29120 -28498 sw
tri -28324 -28551 -28271 -28498 ne
rect -28271 -28551 -26043 -28498
rect -31099 -29400 -29120 -28551
tri -29120 -29400 -28271 -28551 sw
tri -28271 -29400 -27422 -28551 ne
rect -27422 -28800 -26043 -28551
tri -26043 -28800 -25194 -27951 sw
tri -25194 -28800 -24345 -27951 ne
rect -24345 -28800 -15655 -27951
tri -15655 -28800 -14806 -27951 nw
tri -14806 -28800 -13957 -27951 se
rect -13957 -28473 -11651 -27951
tri -11651 -28473 -10827 -27649 nw
tri -10802 -28473 -9978 -27649 se
rect -9978 -27799 -7300 -27649
tri -7300 -27799 -5300 -25799 nw
rect -9978 -28473 -9900 -27799
rect -13957 -28800 -12500 -28473
rect -27422 -29400 -25194 -28800
tri -25194 -29400 -24594 -28800 sw
tri -15406 -29400 -14806 -28800 se
rect -14806 -29322 -12500 -28800
tri -12500 -29322 -11651 -28473 nw
tri -11651 -29322 -10802 -28473 se
rect -10802 -29322 -9900 -28473
rect -14806 -29400 -13349 -29322
tri -31099 -32000 -28499 -29400 ne
rect -28499 -30249 -28271 -29400
tri -28271 -30249 -27422 -29400 sw
tri -27422 -30249 -26573 -29400 ne
rect -26573 -30171 -13349 -29400
tri -13349 -30171 -12500 -29322 nw
tri -12500 -30171 -11651 -29322 se
rect -11651 -30171 -9900 -29322
rect -26573 -30249 -13655 -30171
rect -28499 -30551 -27422 -30249
tri -27422 -30551 -27120 -30249 sw
tri -26573 -30551 -26271 -30249 ne
rect -26271 -30477 -13655 -30249
tri -13655 -30477 -13349 -30171 nw
tri -12806 -30477 -12500 -30171 se
rect -12500 -30399 -9900 -30171
tri -9900 -30399 -7300 -27799 nw
rect -26271 -30551 -14504 -30477
rect -28499 -31400 -27120 -30551
tri -27120 -31400 -26271 -30551 sw
tri -26271 -31400 -25422 -30551 ne
rect -25422 -31326 -14504 -30551
tri -14504 -31326 -13655 -30477 nw
tri -13655 -31326 -12806 -30477 se
rect -12806 -31326 -12500 -30477
rect -25422 -31400 -14578 -31326
tri -14578 -31400 -14504 -31326 nw
rect -28499 -32000 -26271 -31400
tri -26271 -32000 -25671 -31400 sw
tri -14329 -32000 -13655 -31326 se
rect -13655 -32000 -12500 -31326
tri -28499 -34000 -26499 -32000 ne
rect -26499 -32999 -12500 -32000
tri -12500 -32999 -9900 -30399 nw
rect -26499 -34000 -13501 -32999
tri -13501 -34000 -12500 -32999 nw
<< end >>
