magic
tech sky130B
timestamp 1660789662
<< metal1 >>
rect 200 840 500 850
rect 200 760 260 840
rect 440 760 500 840
rect 200 700 500 760
rect 850 840 1150 900
rect 850 760 910 840
rect 1090 760 1150 840
rect 850 700 1150 760
rect 1500 850 1900 900
rect 1500 840 1800 850
rect 1500 760 1560 840
rect 1740 760 1800 840
rect 1500 700 1800 760
rect 200 -860 500 -850
rect 200 -940 260 -860
rect 440 -940 500 -860
rect 200 -1000 500 -940
rect 850 -860 1150 -850
rect 850 -940 910 -860
rect 1090 -940 1150 -860
rect 850 -1000 1150 -940
rect 1500 -860 1800 -800
rect 1500 -940 1560 -860
rect 1740 -940 1800 -860
rect 1500 -1000 1800 -940
<< via1 >>
rect 260 760 440 840
rect 910 760 1090 840
rect 1560 760 1740 840
rect 260 -940 440 -860
rect 910 -940 1090 -860
rect 1560 -940 1740 -860
<< metal2 >>
rect 0 890 200 900
rect 0 760 10 890
rect 90 850 200 890
rect 500 890 850 900
rect 500 850 610 890
rect 90 760 100 850
rect 0 750 100 760
rect 250 840 450 850
rect 250 760 260 840
rect 440 760 450 840
rect 250 750 450 760
rect 600 760 610 850
rect 740 850 850 890
rect 1150 890 1500 900
rect 1150 850 1260 890
rect 740 760 750 850
rect 600 750 750 760
rect 900 840 1100 850
rect 900 760 910 840
rect 1090 760 1100 840
rect 900 750 1100 760
rect 1250 760 1260 850
rect 1390 850 1500 890
rect 1800 890 2050 900
rect 1800 850 1910 890
rect 1390 760 1400 850
rect 1250 750 1400 760
rect 1550 840 1750 850
rect 1550 760 1560 840
rect 1740 760 1750 840
rect 1550 750 1750 760
rect 1900 750 1910 850
rect 2040 750 2050 890
rect 0 710 200 750
rect 500 710 850 750
rect 1150 710 1500 750
rect 1800 710 2050 750
rect 0 700 210 710
rect 80 690 210 700
rect 490 700 870 710
rect 490 690 620 700
rect 710 690 870 700
rect 1130 690 1520 710
rect 1780 690 2050 710
rect 0 -850 200 -800
rect 500 -850 850 -800
rect 1150 -850 1500 -800
rect 1800 -850 2050 -800
rect 0 -860 100 -850
rect 0 -1000 10 -860
rect 90 -950 100 -860
rect 250 -860 450 -850
rect 250 -940 260 -860
rect 440 -940 450 -860
rect 250 -950 450 -940
rect 600 -860 750 -850
rect 600 -950 610 -860
rect 90 -990 200 -950
rect 500 -990 610 -950
rect 90 -1000 220 -990
rect 0 -1010 220 -1000
rect 480 -1000 610 -990
rect 740 -950 750 -860
rect 900 -860 1100 -850
rect 900 -940 910 -860
rect 1090 -940 1100 -860
rect 900 -950 1100 -940
rect 1250 -860 1400 -850
rect 1250 -950 1260 -860
rect 740 -990 850 -950
rect 1150 -990 1260 -950
rect 740 -1000 870 -990
rect 480 -1010 870 -1000
rect 1130 -1000 1260 -990
rect 1390 -950 1400 -860
rect 1550 -860 1750 -850
rect 1550 -940 1560 -860
rect 1740 -940 1750 -860
rect 1550 -950 1750 -940
rect 1900 -860 2050 -850
rect 1900 -950 1910 -860
rect 1390 -990 1500 -950
rect 1800 -990 1910 -950
rect 1390 -1000 1520 -990
rect 1130 -1010 1520 -1000
rect 1780 -1000 1910 -990
rect 2040 -1000 2050 -860
rect 1780 -1010 2050 -1000
<< via2 >>
rect 10 760 90 890
rect 260 760 440 840
rect 610 760 740 890
rect 910 760 1090 840
rect 1260 760 1390 890
rect 1560 760 1740 840
rect 1910 750 2040 890
rect 10 -1000 90 -860
rect 260 -940 440 -860
rect 610 -1000 740 -860
rect 910 -940 1090 -860
rect 1260 -1000 1390 -860
rect 1560 -940 1740 -860
rect 1910 -1000 2040 -860
<< metal3 >>
rect 0 900 100 910
rect 0 760 10 900
rect 90 760 100 900
rect 600 900 750 910
rect 0 750 100 760
rect 250 840 450 850
rect 250 760 260 840
rect 440 760 450 840
rect 250 700 450 760
rect 600 760 610 900
rect 740 760 750 900
rect 1250 900 1400 910
rect 600 750 750 760
rect 900 840 1100 850
rect 900 760 910 840
rect 1090 760 1100 840
rect 900 700 1100 760
rect 1250 760 1260 900
rect 1390 760 1400 900
rect 1900 890 2050 900
rect 1250 750 1400 760
rect 1550 840 1750 850
rect 1550 760 1560 840
rect 1740 760 1750 840
rect 1550 700 1750 760
rect 1900 750 1910 890
rect 2040 750 2050 890
rect 1900 740 2050 750
rect -200 500 1750 700
rect -200 -600 0 500
rect -200 -800 1750 -600
rect 0 -860 100 -850
rect 0 -1000 10 -860
rect 90 -1000 100 -860
rect 250 -860 450 -800
rect 250 -940 260 -860
rect 440 -940 450 -860
rect 250 -950 450 -940
rect 600 -860 750 -850
rect 0 -1010 100 -1000
rect 600 -1000 610 -860
rect 740 -1000 750 -860
rect 900 -860 1100 -800
rect 900 -940 910 -860
rect 1090 -940 1100 -860
rect 900 -950 1100 -940
rect 1250 -860 1400 -850
rect 600 -1010 750 -1000
rect 1250 -1000 1260 -860
rect 1390 -1000 1400 -860
rect 1550 -860 1750 -800
rect 1550 -940 1560 -860
rect 1740 -940 1750 -860
rect 1550 -950 1750 -940
rect 1900 -860 2050 -850
rect 1250 -1010 1400 -1000
rect 1900 -1000 1910 -860
rect 2040 -1000 2050 -860
rect 1900 -1010 2050 -1000
<< via3 >>
rect 220 1530 280 1760
rect 470 1530 530 1760
rect 720 1530 780 1760
rect 970 1530 1030 1760
rect 1220 1530 1280 1760
rect 1470 1530 1530 1760
rect 1720 1530 1780 1760
rect 10 890 90 900
rect 10 760 90 890
rect 610 890 740 900
rect 610 760 740 890
rect 1260 890 1390 900
rect 1260 760 1390 890
rect 1910 750 2040 890
rect 470 -170 530 50
rect 720 -170 780 50
rect 970 -170 1030 50
rect 1220 -170 1280 50
rect 1470 -170 1530 50
rect 10 -1000 90 -860
rect 610 -1000 740 -860
rect 1260 -1000 1390 -860
rect 1910 -1000 2040 -860
rect 220 -1880 280 -1650
rect 470 -1880 530 -1650
rect 720 -1880 780 -1650
rect 970 -1880 1030 -1650
rect 1220 -1880 1280 -1650
rect 1470 -1880 1530 -1650
rect 1720 -1880 1780 -1650
<< metal4 >>
rect 210 1760 1790 1770
rect 210 1530 220 1760
rect 280 1530 430 1760
rect 570 1530 680 1760
rect 820 1530 970 1760
rect 1030 1530 1180 1760
rect 1320 1530 1430 1760
rect 1570 1530 1720 1760
rect 1780 1530 1790 1760
rect 210 1520 1790 1530
rect 0 900 2200 910
rect 0 760 10 900
rect 90 760 610 900
rect 740 760 1260 900
rect 1390 890 2200 900
rect 1390 760 1910 890
rect 0 750 1910 760
rect 2040 750 2200 890
rect 1900 740 2200 750
rect 420 60 480 70
rect 1520 60 1580 70
rect 420 -170 430 60
rect 570 -170 680 60
rect 820 50 1180 60
rect 820 -170 970 50
rect 1030 -170 1180 50
rect 1320 -170 1430 60
rect 1570 -170 1580 60
rect 420 -180 1580 -170
rect 2050 -850 2200 740
rect 0 -860 2200 -850
rect 0 -1000 10 -860
rect 90 -1000 610 -860
rect 740 -1000 1260 -860
rect 1390 -1000 1910 -860
rect 2040 -1000 2200 -860
rect 0 -1010 2200 -1000
rect 210 -1650 1790 -1640
rect 210 -1880 220 -1650
rect 280 -1880 430 -1650
rect 570 -1880 680 -1650
rect 820 -1880 970 -1650
rect 1030 -1880 1180 -1650
rect 1320 -1880 1430 -1650
rect 1570 -1880 1720 -1650
rect 1780 -1880 1790 -1650
rect 210 -1890 1790 -1880
<< via4 >>
rect 430 1530 470 1760
rect 470 1530 530 1760
rect 530 1530 570 1760
rect 680 1530 720 1760
rect 720 1530 780 1760
rect 780 1530 820 1760
rect 1180 1530 1220 1760
rect 1220 1530 1280 1760
rect 1280 1530 1320 1760
rect 1430 1530 1470 1760
rect 1470 1530 1530 1760
rect 1530 1530 1570 1760
rect 430 50 570 60
rect 430 -170 470 50
rect 470 -170 530 50
rect 530 -170 570 50
rect 680 50 820 60
rect 1180 50 1320 60
rect 680 -170 720 50
rect 720 -170 780 50
rect 780 -170 820 50
rect 1180 -170 1220 50
rect 1220 -170 1280 50
rect 1280 -170 1320 50
rect 1430 50 1570 60
rect 1430 -170 1470 50
rect 1470 -170 1530 50
rect 1530 -170 1570 50
rect 430 -1880 470 -1650
rect 470 -1880 530 -1650
rect 530 -1880 570 -1650
rect 680 -1880 720 -1650
rect 720 -1880 780 -1650
rect 780 -1880 820 -1650
rect 1180 -1880 1220 -1650
rect 1220 -1880 1280 -1650
rect 1280 -1880 1320 -1650
rect 1430 -1880 1470 -1650
rect 1470 -1880 1530 -1650
rect 1530 -1880 1570 -1650
<< metal5 >>
rect 0 1760 2000 1780
rect 0 1530 430 1760
rect 570 1530 680 1760
rect 820 1530 1180 1760
rect 1320 1530 1430 1760
rect 1570 1530 2000 1760
rect 0 1520 2000 1530
rect 410 60 840 1520
rect 410 -170 430 60
rect 570 -170 680 60
rect 820 -170 840 60
rect 410 -1640 840 -170
rect 1160 60 1590 1520
rect 1160 -170 1180 60
rect 1320 -170 1430 60
rect 1570 -170 1590 60
rect 1160 -1640 1590 -170
rect 0 -1650 2000 -1640
rect 0 -1880 430 -1650
rect 570 -1880 680 -1650
rect 820 -1880 1180 -1650
rect 1320 -1880 1430 -1650
rect 1570 -1880 2000 -1650
rect 0 -1900 2000 -1880
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659929390
transform 1 0 253 0 1 -1055
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_1
timestamp 1659929390
transform 1 0 253 0 -1 940
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_2
timestamp 1659929390
transform 1 0 253 0 -1 2640
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_3
timestamp 1659929390
transform 1 0 253 0 1 -2755
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_4
timestamp 1659929390
transform -1 0 1080 0 1 -2755
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_5
timestamp 1659929390
transform -1 0 1080 0 -1 2640
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_6
timestamp 1659929390
transform -1 0 1080 0 1 -1055
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_7
timestamp 1659929390
transform -1 0 1080 0 -1 940
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_8
timestamp 1659929390
transform 1 0 1543 0 1 -2755
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_9
timestamp 1659929390
transform 1 0 1543 0 -1 2640
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_10
timestamp 1659929390
transform 1 0 1543 0 1 -1055
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_11
timestamp 1659929390
transform 1 0 1543 0 -1 940
box -253 1105 435 1790
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660275339
transform 1 0 -50 0 1 2070
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_1
timestamp 1660275339
transform 1 0 200 0 1 2070
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_2
timestamp 1660275339
transform 1 0 450 0 1 2070
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_3
timestamp 1660275339
transform 1 0 700 0 1 2070
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_4
timestamp 1660275339
transform 1 0 950 0 1 2070
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_5
timestamp 1660275339
transform 1 0 1200 0 1 2070
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_6
timestamp 1660275339
transform 1 0 1450 0 1 2070
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_7
timestamp 1660275339
transform 1 0 1700 0 1 2070
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_8
timestamp 1660275339
transform 1 0 1700 0 1 -1340
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_9
timestamp 1660275339
transform 1 0 -50 0 1 -1340
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_10
timestamp 1660275339
transform 1 0 200 0 1 -1340
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_11
timestamp 1660275339
transform 1 0 450 0 1 -1340
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_12
timestamp 1660275339
transform 1 0 950 0 1 -1340
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_13
timestamp 1660275339
transform 1 0 700 0 1 -1340
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_14
timestamp 1660275339
transform 1 0 1200 0 1 -1340
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_15
timestamp 1660275339
transform 1 0 1450 0 1 -1340
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_17
timestamp 1660275339
transform 1 0 200 0 1 370
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_18
timestamp 1660275339
transform 1 0 450 0 1 370
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_19
timestamp 1660275339
transform 1 0 700 0 1 370
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_20
timestamp 1660275339
transform 1 0 950 0 1 370
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_21
timestamp 1660275339
transform 1 0 1200 0 1 370
box 50 -550 300 -300
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_22
timestamp 1660275339
transform 1 0 1450 0 1 370
box 50 -550 300 -300
<< labels >>
rlabel metal3 -200 -800 0 700 1 G
rlabel metal5 0 1520 2000 1780 1 SG
rlabel metal4 2050 -1010 2200 910 1 D
<< end >>
