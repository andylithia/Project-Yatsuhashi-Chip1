magic
tech sky130B
magscale 1 2
timestamp 1659146707
<< pwell >>
rect 0 66 676 1128
<< nmos >>
rect 194 92 224 1102
rect 280 92 310 1102
rect 366 92 396 1102
rect 452 92 482 1102
<< ndiff >>
rect 138 1090 194 1102
rect 138 1056 149 1090
rect 183 1056 194 1090
rect 138 1022 194 1056
rect 138 988 149 1022
rect 183 988 194 1022
rect 138 954 194 988
rect 138 920 149 954
rect 183 920 194 954
rect 138 886 194 920
rect 138 852 149 886
rect 183 852 194 886
rect 138 818 194 852
rect 138 784 149 818
rect 183 784 194 818
rect 138 750 194 784
rect 138 716 149 750
rect 183 716 194 750
rect 138 682 194 716
rect 138 648 149 682
rect 183 648 194 682
rect 138 614 194 648
rect 138 580 149 614
rect 183 580 194 614
rect 138 546 194 580
rect 138 512 149 546
rect 183 512 194 546
rect 138 478 194 512
rect 138 444 149 478
rect 183 444 194 478
rect 138 410 194 444
rect 138 376 149 410
rect 183 376 194 410
rect 138 342 194 376
rect 138 308 149 342
rect 183 308 194 342
rect 138 274 194 308
rect 138 240 149 274
rect 183 240 194 274
rect 138 206 194 240
rect 138 172 149 206
rect 183 172 194 206
rect 138 138 194 172
rect 138 104 149 138
rect 183 104 194 138
rect 138 92 194 104
rect 224 1090 280 1102
rect 224 1056 235 1090
rect 269 1056 280 1090
rect 224 1022 280 1056
rect 224 988 235 1022
rect 269 988 280 1022
rect 224 954 280 988
rect 224 920 235 954
rect 269 920 280 954
rect 224 886 280 920
rect 224 852 235 886
rect 269 852 280 886
rect 224 818 280 852
rect 224 784 235 818
rect 269 784 280 818
rect 224 750 280 784
rect 224 716 235 750
rect 269 716 280 750
rect 224 682 280 716
rect 224 648 235 682
rect 269 648 280 682
rect 224 614 280 648
rect 224 580 235 614
rect 269 580 280 614
rect 224 546 280 580
rect 224 512 235 546
rect 269 512 280 546
rect 224 478 280 512
rect 224 444 235 478
rect 269 444 280 478
rect 224 410 280 444
rect 224 376 235 410
rect 269 376 280 410
rect 224 342 280 376
rect 224 308 235 342
rect 269 308 280 342
rect 224 274 280 308
rect 224 240 235 274
rect 269 240 280 274
rect 224 206 280 240
rect 224 172 235 206
rect 269 172 280 206
rect 224 138 280 172
rect 224 104 235 138
rect 269 104 280 138
rect 224 92 280 104
rect 310 1090 366 1102
rect 310 1056 321 1090
rect 355 1056 366 1090
rect 310 1022 366 1056
rect 310 988 321 1022
rect 355 988 366 1022
rect 310 954 366 988
rect 310 920 321 954
rect 355 920 366 954
rect 310 886 366 920
rect 310 852 321 886
rect 355 852 366 886
rect 310 818 366 852
rect 310 784 321 818
rect 355 784 366 818
rect 310 750 366 784
rect 310 716 321 750
rect 355 716 366 750
rect 310 682 366 716
rect 310 648 321 682
rect 355 648 366 682
rect 310 614 366 648
rect 310 580 321 614
rect 355 580 366 614
rect 310 546 366 580
rect 310 512 321 546
rect 355 512 366 546
rect 310 478 366 512
rect 310 444 321 478
rect 355 444 366 478
rect 310 410 366 444
rect 310 376 321 410
rect 355 376 366 410
rect 310 342 366 376
rect 310 308 321 342
rect 355 308 366 342
rect 310 274 366 308
rect 310 240 321 274
rect 355 240 366 274
rect 310 206 366 240
rect 310 172 321 206
rect 355 172 366 206
rect 310 138 366 172
rect 310 104 321 138
rect 355 104 366 138
rect 310 92 366 104
rect 396 1090 452 1102
rect 396 1056 407 1090
rect 441 1056 452 1090
rect 396 1022 452 1056
rect 396 988 407 1022
rect 441 988 452 1022
rect 396 954 452 988
rect 396 920 407 954
rect 441 920 452 954
rect 396 886 452 920
rect 396 852 407 886
rect 441 852 452 886
rect 396 818 452 852
rect 396 784 407 818
rect 441 784 452 818
rect 396 750 452 784
rect 396 716 407 750
rect 441 716 452 750
rect 396 682 452 716
rect 396 648 407 682
rect 441 648 452 682
rect 396 614 452 648
rect 396 580 407 614
rect 441 580 452 614
rect 396 546 452 580
rect 396 512 407 546
rect 441 512 452 546
rect 396 478 452 512
rect 396 444 407 478
rect 441 444 452 478
rect 396 410 452 444
rect 396 376 407 410
rect 441 376 452 410
rect 396 342 452 376
rect 396 308 407 342
rect 441 308 452 342
rect 396 274 452 308
rect 396 240 407 274
rect 441 240 452 274
rect 396 206 452 240
rect 396 172 407 206
rect 441 172 452 206
rect 396 138 452 172
rect 396 104 407 138
rect 441 104 452 138
rect 396 92 452 104
rect 482 1090 538 1102
rect 482 1056 493 1090
rect 527 1056 538 1090
rect 482 1022 538 1056
rect 482 988 493 1022
rect 527 988 538 1022
rect 482 954 538 988
rect 482 920 493 954
rect 527 920 538 954
rect 482 886 538 920
rect 482 852 493 886
rect 527 852 538 886
rect 482 818 538 852
rect 482 784 493 818
rect 527 784 538 818
rect 482 750 538 784
rect 482 716 493 750
rect 527 716 538 750
rect 482 682 538 716
rect 482 648 493 682
rect 527 648 538 682
rect 482 614 538 648
rect 482 580 493 614
rect 527 580 538 614
rect 482 546 538 580
rect 482 512 493 546
rect 527 512 538 546
rect 482 478 538 512
rect 482 444 493 478
rect 527 444 538 478
rect 482 410 538 444
rect 482 376 493 410
rect 527 376 538 410
rect 482 342 538 376
rect 482 308 493 342
rect 527 308 538 342
rect 482 274 538 308
rect 482 240 493 274
rect 527 240 538 274
rect 482 206 538 240
rect 482 172 493 206
rect 527 172 538 206
rect 482 138 538 172
rect 482 104 493 138
rect 527 104 538 138
rect 482 92 538 104
<< ndiffc >>
rect 149 1056 183 1090
rect 149 988 183 1022
rect 149 920 183 954
rect 149 852 183 886
rect 149 784 183 818
rect 149 716 183 750
rect 149 648 183 682
rect 149 580 183 614
rect 149 512 183 546
rect 149 444 183 478
rect 149 376 183 410
rect 149 308 183 342
rect 149 240 183 274
rect 149 172 183 206
rect 149 104 183 138
rect 235 1056 269 1090
rect 235 988 269 1022
rect 235 920 269 954
rect 235 852 269 886
rect 235 784 269 818
rect 235 716 269 750
rect 235 648 269 682
rect 235 580 269 614
rect 235 512 269 546
rect 235 444 269 478
rect 235 376 269 410
rect 235 308 269 342
rect 235 240 269 274
rect 235 172 269 206
rect 235 104 269 138
rect 321 1056 355 1090
rect 321 988 355 1022
rect 321 920 355 954
rect 321 852 355 886
rect 321 784 355 818
rect 321 716 355 750
rect 321 648 355 682
rect 321 580 355 614
rect 321 512 355 546
rect 321 444 355 478
rect 321 376 355 410
rect 321 308 355 342
rect 321 240 355 274
rect 321 172 355 206
rect 321 104 355 138
rect 407 1056 441 1090
rect 407 988 441 1022
rect 407 920 441 954
rect 407 852 441 886
rect 407 784 441 818
rect 407 716 441 750
rect 407 648 441 682
rect 407 580 441 614
rect 407 512 441 546
rect 407 444 441 478
rect 407 376 441 410
rect 407 308 441 342
rect 407 240 441 274
rect 407 172 441 206
rect 407 104 441 138
rect 493 1056 527 1090
rect 493 988 527 1022
rect 493 920 527 954
rect 493 852 527 886
rect 493 784 527 818
rect 493 716 527 750
rect 493 648 527 682
rect 493 580 527 614
rect 493 512 527 546
rect 493 444 527 478
rect 493 376 527 410
rect 493 308 527 342
rect 493 240 527 274
rect 493 172 527 206
rect 493 104 527 138
<< psubdiff >>
rect 26 1056 84 1102
rect 26 1022 38 1056
rect 72 1022 84 1056
rect 26 988 84 1022
rect 26 954 38 988
rect 72 954 84 988
rect 26 920 84 954
rect 26 886 38 920
rect 72 886 84 920
rect 26 852 84 886
rect 26 818 38 852
rect 72 818 84 852
rect 26 784 84 818
rect 26 750 38 784
rect 72 750 84 784
rect 26 716 84 750
rect 26 682 38 716
rect 72 682 84 716
rect 26 648 84 682
rect 26 614 38 648
rect 72 614 84 648
rect 26 580 84 614
rect 26 546 38 580
rect 72 546 84 580
rect 26 512 84 546
rect 26 478 38 512
rect 72 478 84 512
rect 26 444 84 478
rect 26 410 38 444
rect 72 410 84 444
rect 26 376 84 410
rect 26 342 38 376
rect 72 342 84 376
rect 26 308 84 342
rect 26 274 38 308
rect 72 274 84 308
rect 26 240 84 274
rect 26 206 38 240
rect 72 206 84 240
rect 26 172 84 206
rect 26 138 38 172
rect 72 138 84 172
rect 26 92 84 138
rect 592 1056 650 1102
rect 592 1022 604 1056
rect 638 1022 650 1056
rect 592 988 650 1022
rect 592 954 604 988
rect 638 954 650 988
rect 592 920 650 954
rect 592 886 604 920
rect 638 886 650 920
rect 592 852 650 886
rect 592 818 604 852
rect 638 818 650 852
rect 592 784 650 818
rect 592 750 604 784
rect 638 750 650 784
rect 592 716 650 750
rect 592 682 604 716
rect 638 682 650 716
rect 592 648 650 682
rect 592 614 604 648
rect 638 614 650 648
rect 592 580 650 614
rect 592 546 604 580
rect 638 546 650 580
rect 592 512 650 546
rect 592 478 604 512
rect 638 478 650 512
rect 592 444 650 478
rect 592 410 604 444
rect 638 410 650 444
rect 592 376 650 410
rect 592 342 604 376
rect 638 342 650 376
rect 592 308 650 342
rect 592 274 604 308
rect 638 274 650 308
rect 592 240 650 274
rect 592 206 604 240
rect 638 206 650 240
rect 592 172 650 206
rect 592 138 604 172
rect 638 138 650 172
rect 592 92 650 138
<< psubdiffcont >>
rect 38 1022 72 1056
rect 38 954 72 988
rect 38 886 72 920
rect 38 818 72 852
rect 38 750 72 784
rect 38 682 72 716
rect 38 614 72 648
rect 38 546 72 580
rect 38 478 72 512
rect 38 410 72 444
rect 38 342 72 376
rect 38 274 72 308
rect 38 206 72 240
rect 38 138 72 172
rect 604 1022 638 1056
rect 604 954 638 988
rect 604 886 638 920
rect 604 818 638 852
rect 604 750 638 784
rect 604 682 638 716
rect 604 614 638 648
rect 604 546 638 580
rect 604 478 638 512
rect 604 410 638 444
rect 604 342 638 376
rect 604 274 638 308
rect 604 206 638 240
rect 604 138 638 172
<< poly >>
rect 169 1174 507 1194
rect 169 1140 185 1174
rect 219 1140 253 1174
rect 287 1140 321 1174
rect 355 1140 389 1174
rect 423 1140 457 1174
rect 491 1140 507 1174
rect 169 1124 507 1140
rect 194 1102 224 1124
rect 280 1102 310 1124
rect 366 1102 396 1124
rect 452 1102 482 1124
rect 194 70 224 92
rect 280 70 310 92
rect 366 70 396 92
rect 452 70 482 92
rect 169 54 507 70
rect 169 20 185 54
rect 219 20 253 54
rect 287 20 321 54
rect 355 20 389 54
rect 423 20 457 54
rect 491 20 507 54
rect 169 0 507 20
<< polycont >>
rect 185 1140 219 1174
rect 253 1140 287 1174
rect 321 1140 355 1174
rect 389 1140 423 1174
rect 457 1140 491 1174
rect 185 20 219 54
rect 253 20 287 54
rect 321 20 355 54
rect 389 20 423 54
rect 457 20 491 54
<< locali >>
rect 169 1140 177 1174
rect 219 1140 249 1174
rect 287 1140 321 1174
rect 355 1140 389 1174
rect 427 1140 457 1174
rect 499 1140 507 1174
rect 149 1090 183 1106
rect 38 1010 72 1022
rect 38 938 72 954
rect 38 866 72 886
rect 38 794 72 818
rect 38 722 72 750
rect 38 650 72 682
rect 38 580 72 614
rect 38 512 72 544
rect 38 444 72 472
rect 38 376 72 400
rect 38 308 72 328
rect 38 240 72 256
rect 38 172 72 184
rect 149 1022 183 1048
rect 149 954 183 976
rect 149 886 183 904
rect 149 818 183 832
rect 149 750 183 760
rect 149 682 183 688
rect 149 614 183 616
rect 149 578 183 580
rect 149 506 183 512
rect 149 434 183 444
rect 149 362 183 376
rect 149 290 183 308
rect 149 218 183 240
rect 149 146 183 172
rect 149 88 183 104
rect 235 1090 269 1106
rect 235 1022 269 1048
rect 235 954 269 976
rect 235 886 269 904
rect 235 818 269 832
rect 235 750 269 760
rect 235 682 269 688
rect 235 614 269 616
rect 235 578 269 580
rect 235 506 269 512
rect 235 434 269 444
rect 235 362 269 376
rect 235 290 269 308
rect 235 218 269 240
rect 235 146 269 172
rect 235 88 269 104
rect 321 1090 355 1106
rect 321 1022 355 1048
rect 321 954 355 976
rect 321 886 355 904
rect 321 818 355 832
rect 321 750 355 760
rect 321 682 355 688
rect 321 614 355 616
rect 321 578 355 580
rect 321 506 355 512
rect 321 434 355 444
rect 321 362 355 376
rect 321 290 355 308
rect 321 218 355 240
rect 321 146 355 172
rect 321 88 355 104
rect 407 1090 441 1106
rect 407 1022 441 1048
rect 407 954 441 976
rect 407 886 441 904
rect 407 818 441 832
rect 407 750 441 760
rect 407 682 441 688
rect 407 614 441 616
rect 407 578 441 580
rect 407 506 441 512
rect 407 434 441 444
rect 407 362 441 376
rect 407 290 441 308
rect 407 218 441 240
rect 407 146 441 172
rect 407 88 441 104
rect 493 1090 527 1106
rect 493 1022 527 1048
rect 493 954 527 976
rect 493 886 527 904
rect 493 818 527 832
rect 493 750 527 760
rect 493 682 527 688
rect 493 614 527 616
rect 493 578 527 580
rect 493 506 527 512
rect 493 434 527 444
rect 493 362 527 376
rect 493 290 527 308
rect 493 218 527 240
rect 493 146 527 172
rect 604 1010 638 1022
rect 604 938 638 954
rect 604 866 638 886
rect 604 794 638 818
rect 604 722 638 750
rect 604 650 638 682
rect 604 580 638 614
rect 604 512 638 544
rect 604 444 638 472
rect 604 376 638 400
rect 604 308 638 328
rect 604 240 638 256
rect 604 172 638 184
rect 493 88 527 104
rect 169 20 177 54
rect 219 20 249 54
rect 287 20 321 54
rect 355 20 389 54
rect 427 20 457 54
rect 499 20 507 54
<< viali >>
rect 177 1140 185 1174
rect 185 1140 211 1174
rect 249 1140 253 1174
rect 253 1140 283 1174
rect 321 1140 355 1174
rect 393 1140 423 1174
rect 423 1140 427 1174
rect 465 1140 491 1174
rect 491 1140 499 1174
rect 38 1056 72 1082
rect 38 1048 72 1056
rect 38 988 72 1010
rect 38 976 72 988
rect 38 920 72 938
rect 38 904 72 920
rect 38 852 72 866
rect 38 832 72 852
rect 38 784 72 794
rect 38 760 72 784
rect 38 716 72 722
rect 38 688 72 716
rect 38 648 72 650
rect 38 616 72 648
rect 38 546 72 578
rect 38 544 72 546
rect 38 478 72 506
rect 38 472 72 478
rect 38 410 72 434
rect 38 400 72 410
rect 38 342 72 362
rect 38 328 72 342
rect 38 274 72 290
rect 38 256 72 274
rect 38 206 72 218
rect 38 184 72 206
rect 38 138 72 146
rect 38 112 72 138
rect 149 1056 183 1082
rect 149 1048 183 1056
rect 149 988 183 1010
rect 149 976 183 988
rect 149 920 183 938
rect 149 904 183 920
rect 149 852 183 866
rect 149 832 183 852
rect 149 784 183 794
rect 149 760 183 784
rect 149 716 183 722
rect 149 688 183 716
rect 149 648 183 650
rect 149 616 183 648
rect 149 546 183 578
rect 149 544 183 546
rect 149 478 183 506
rect 149 472 183 478
rect 149 410 183 434
rect 149 400 183 410
rect 149 342 183 362
rect 149 328 183 342
rect 149 274 183 290
rect 149 256 183 274
rect 149 206 183 218
rect 149 184 183 206
rect 149 138 183 146
rect 149 112 183 138
rect 235 1056 269 1082
rect 235 1048 269 1056
rect 235 988 269 1010
rect 235 976 269 988
rect 235 920 269 938
rect 235 904 269 920
rect 235 852 269 866
rect 235 832 269 852
rect 235 784 269 794
rect 235 760 269 784
rect 235 716 269 722
rect 235 688 269 716
rect 235 648 269 650
rect 235 616 269 648
rect 235 546 269 578
rect 235 544 269 546
rect 235 478 269 506
rect 235 472 269 478
rect 235 410 269 434
rect 235 400 269 410
rect 235 342 269 362
rect 235 328 269 342
rect 235 274 269 290
rect 235 256 269 274
rect 235 206 269 218
rect 235 184 269 206
rect 235 138 269 146
rect 235 112 269 138
rect 321 1056 355 1082
rect 321 1048 355 1056
rect 321 988 355 1010
rect 321 976 355 988
rect 321 920 355 938
rect 321 904 355 920
rect 321 852 355 866
rect 321 832 355 852
rect 321 784 355 794
rect 321 760 355 784
rect 321 716 355 722
rect 321 688 355 716
rect 321 648 355 650
rect 321 616 355 648
rect 321 546 355 578
rect 321 544 355 546
rect 321 478 355 506
rect 321 472 355 478
rect 321 410 355 434
rect 321 400 355 410
rect 321 342 355 362
rect 321 328 355 342
rect 321 274 355 290
rect 321 256 355 274
rect 321 206 355 218
rect 321 184 355 206
rect 321 138 355 146
rect 321 112 355 138
rect 407 1056 441 1082
rect 407 1048 441 1056
rect 407 988 441 1010
rect 407 976 441 988
rect 407 920 441 938
rect 407 904 441 920
rect 407 852 441 866
rect 407 832 441 852
rect 407 784 441 794
rect 407 760 441 784
rect 407 716 441 722
rect 407 688 441 716
rect 407 648 441 650
rect 407 616 441 648
rect 407 546 441 578
rect 407 544 441 546
rect 407 478 441 506
rect 407 472 441 478
rect 407 410 441 434
rect 407 400 441 410
rect 407 342 441 362
rect 407 328 441 342
rect 407 274 441 290
rect 407 256 441 274
rect 407 206 441 218
rect 407 184 441 206
rect 407 138 441 146
rect 407 112 441 138
rect 493 1056 527 1082
rect 493 1048 527 1056
rect 493 988 527 1010
rect 493 976 527 988
rect 493 920 527 938
rect 493 904 527 920
rect 493 852 527 866
rect 493 832 527 852
rect 493 784 527 794
rect 493 760 527 784
rect 493 716 527 722
rect 493 688 527 716
rect 493 648 527 650
rect 493 616 527 648
rect 493 546 527 578
rect 493 544 527 546
rect 493 478 527 506
rect 493 472 527 478
rect 493 410 527 434
rect 493 400 527 410
rect 493 342 527 362
rect 493 328 527 342
rect 493 274 527 290
rect 493 256 527 274
rect 493 206 527 218
rect 493 184 527 206
rect 493 138 527 146
rect 493 112 527 138
rect 604 1056 638 1082
rect 604 1048 638 1056
rect 604 988 638 1010
rect 604 976 638 988
rect 604 920 638 938
rect 604 904 638 920
rect 604 852 638 866
rect 604 832 638 852
rect 604 784 638 794
rect 604 760 638 784
rect 604 716 638 722
rect 604 688 638 716
rect 604 648 638 650
rect 604 616 638 648
rect 604 546 638 578
rect 604 544 638 546
rect 604 478 638 506
rect 604 472 638 478
rect 604 410 638 434
rect 604 400 638 410
rect 604 342 638 362
rect 604 328 638 342
rect 604 274 638 290
rect 604 256 638 274
rect 604 206 638 218
rect 604 184 638 206
rect 604 138 638 146
rect 604 112 638 138
rect 177 20 185 54
rect 185 20 211 54
rect 249 20 253 54
rect 253 20 283 54
rect 321 20 355 54
rect 393 20 423 54
rect 423 20 427 54
rect 465 20 491 54
rect 491 20 499 54
<< metal1 >>
rect 165 1174 511 1194
rect 165 1140 177 1174
rect 211 1140 249 1174
rect 283 1140 321 1174
rect 355 1140 393 1174
rect 427 1140 465 1174
rect 499 1140 511 1174
rect 165 1128 511 1140
rect 26 1082 84 1094
rect 26 1048 38 1082
rect 72 1048 84 1082
rect 26 1010 84 1048
rect 26 976 38 1010
rect 72 976 84 1010
rect 26 938 84 976
rect 26 904 38 938
rect 72 904 84 938
rect 26 866 84 904
rect 26 832 38 866
rect 72 832 84 866
rect 26 794 84 832
rect 26 760 38 794
rect 72 760 84 794
rect 26 722 84 760
rect 26 688 38 722
rect 72 688 84 722
rect 26 650 84 688
rect 26 616 38 650
rect 72 616 84 650
rect 26 578 84 616
rect 26 544 38 578
rect 72 544 84 578
rect 26 506 84 544
rect 26 472 38 506
rect 72 472 84 506
rect 26 434 84 472
rect 26 400 38 434
rect 72 400 84 434
rect 26 362 84 400
rect 26 328 38 362
rect 72 328 84 362
rect 26 290 84 328
rect 26 256 38 290
rect 72 256 84 290
rect 26 218 84 256
rect 26 184 38 218
rect 72 184 84 218
rect 26 146 84 184
rect 26 112 38 146
rect 72 112 84 146
rect 26 100 84 112
rect 140 1082 192 1094
rect 140 1054 149 1082
rect 183 1054 192 1082
rect 140 990 149 1002
rect 183 990 192 1002
rect 140 926 149 938
rect 183 926 192 938
rect 140 866 192 874
rect 140 862 149 866
rect 183 862 192 866
rect 140 798 192 810
rect 140 734 192 746
rect 140 670 192 682
rect 140 616 149 618
rect 183 616 192 618
rect 140 606 192 616
rect 140 544 149 554
rect 183 544 192 554
rect 140 542 192 544
rect 140 478 149 490
rect 183 478 192 490
rect 140 414 149 426
rect 183 414 192 426
rect 140 350 149 362
rect 183 350 192 362
rect 140 290 192 298
rect 140 286 149 290
rect 183 286 192 290
rect 140 222 192 234
rect 140 158 192 170
rect 140 100 192 106
rect 226 1088 278 1094
rect 226 1024 278 1036
rect 226 960 278 972
rect 226 904 235 908
rect 269 904 278 908
rect 226 896 278 904
rect 226 832 235 844
rect 269 832 278 844
rect 226 768 235 780
rect 269 768 278 780
rect 226 704 235 716
rect 269 704 278 716
rect 226 650 278 652
rect 226 640 235 650
rect 269 640 278 650
rect 226 578 278 588
rect 226 576 235 578
rect 269 576 278 578
rect 226 512 278 524
rect 226 448 278 460
rect 226 384 278 396
rect 226 328 235 332
rect 269 328 278 332
rect 226 320 278 328
rect 226 256 235 268
rect 269 256 278 268
rect 226 192 235 204
rect 269 192 278 204
rect 226 112 235 140
rect 269 112 278 140
rect 226 100 278 112
rect 312 1082 364 1094
rect 312 1054 321 1082
rect 355 1054 364 1082
rect 312 990 321 1002
rect 355 990 364 1002
rect 312 926 321 938
rect 355 926 364 938
rect 312 866 364 874
rect 312 862 321 866
rect 355 862 364 866
rect 312 798 364 810
rect 312 734 364 746
rect 312 670 364 682
rect 312 616 321 618
rect 355 616 364 618
rect 312 606 364 616
rect 312 544 321 554
rect 355 544 364 554
rect 312 542 364 544
rect 312 478 321 490
rect 355 478 364 490
rect 312 414 321 426
rect 355 414 364 426
rect 312 350 321 362
rect 355 350 364 362
rect 312 290 364 298
rect 312 286 321 290
rect 355 286 364 290
rect 312 222 364 234
rect 312 158 364 170
rect 312 100 364 106
rect 398 1088 450 1094
rect 398 1024 450 1036
rect 398 960 450 972
rect 398 904 407 908
rect 441 904 450 908
rect 398 896 450 904
rect 398 832 407 844
rect 441 832 450 844
rect 398 768 407 780
rect 441 768 450 780
rect 398 704 407 716
rect 441 704 450 716
rect 398 650 450 652
rect 398 640 407 650
rect 441 640 450 650
rect 398 578 450 588
rect 398 576 407 578
rect 441 576 450 578
rect 398 512 450 524
rect 398 448 450 460
rect 398 384 450 396
rect 398 328 407 332
rect 441 328 450 332
rect 398 320 450 328
rect 398 256 407 268
rect 441 256 450 268
rect 398 192 407 204
rect 441 192 450 204
rect 398 112 407 140
rect 441 112 450 140
rect 398 100 450 112
rect 484 1082 536 1094
rect 484 1054 493 1082
rect 527 1054 536 1082
rect 484 990 493 1002
rect 527 990 536 1002
rect 484 926 493 938
rect 527 926 536 938
rect 484 866 536 874
rect 484 862 493 866
rect 527 862 536 866
rect 484 798 536 810
rect 484 734 536 746
rect 484 670 536 682
rect 484 616 493 618
rect 527 616 536 618
rect 484 606 536 616
rect 484 544 493 554
rect 527 544 536 554
rect 484 542 536 544
rect 484 478 493 490
rect 527 478 536 490
rect 484 414 493 426
rect 527 414 536 426
rect 484 350 493 362
rect 527 350 536 362
rect 484 290 536 298
rect 484 286 493 290
rect 527 286 536 290
rect 484 222 536 234
rect 484 158 536 170
rect 484 100 536 106
rect 592 1082 650 1094
rect 592 1048 604 1082
rect 638 1048 650 1082
rect 592 1010 650 1048
rect 592 976 604 1010
rect 638 976 650 1010
rect 592 938 650 976
rect 592 904 604 938
rect 638 904 650 938
rect 592 866 650 904
rect 592 832 604 866
rect 638 832 650 866
rect 592 794 650 832
rect 592 760 604 794
rect 638 760 650 794
rect 592 722 650 760
rect 592 688 604 722
rect 638 688 650 722
rect 592 650 650 688
rect 592 616 604 650
rect 638 616 650 650
rect 592 578 650 616
rect 592 544 604 578
rect 638 544 650 578
rect 592 506 650 544
rect 592 472 604 506
rect 638 472 650 506
rect 592 434 650 472
rect 592 400 604 434
rect 638 400 650 434
rect 592 362 650 400
rect 592 328 604 362
rect 638 328 650 362
rect 592 290 650 328
rect 592 256 604 290
rect 638 256 650 290
rect 592 218 650 256
rect 592 184 604 218
rect 638 184 650 218
rect 592 146 650 184
rect 592 112 604 146
rect 638 112 650 146
rect 592 100 650 112
rect 165 54 511 66
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 465 54
rect 499 20 511 54
rect 165 0 511 20
<< via1 >>
rect 140 1048 149 1054
rect 149 1048 183 1054
rect 183 1048 192 1054
rect 140 1010 192 1048
rect 140 1002 149 1010
rect 149 1002 183 1010
rect 183 1002 192 1010
rect 140 976 149 990
rect 149 976 183 990
rect 183 976 192 990
rect 140 938 192 976
rect 140 904 149 926
rect 149 904 183 926
rect 183 904 192 926
rect 140 874 192 904
rect 140 832 149 862
rect 149 832 183 862
rect 183 832 192 862
rect 140 810 192 832
rect 140 794 192 798
rect 140 760 149 794
rect 149 760 183 794
rect 183 760 192 794
rect 140 746 192 760
rect 140 722 192 734
rect 140 688 149 722
rect 149 688 183 722
rect 183 688 192 722
rect 140 682 192 688
rect 140 650 192 670
rect 140 618 149 650
rect 149 618 183 650
rect 183 618 192 650
rect 140 578 192 606
rect 140 554 149 578
rect 149 554 183 578
rect 183 554 192 578
rect 140 506 192 542
rect 140 490 149 506
rect 149 490 183 506
rect 183 490 192 506
rect 140 472 149 478
rect 149 472 183 478
rect 183 472 192 478
rect 140 434 192 472
rect 140 426 149 434
rect 149 426 183 434
rect 183 426 192 434
rect 140 400 149 414
rect 149 400 183 414
rect 183 400 192 414
rect 140 362 192 400
rect 140 328 149 350
rect 149 328 183 350
rect 183 328 192 350
rect 140 298 192 328
rect 140 256 149 286
rect 149 256 183 286
rect 183 256 192 286
rect 140 234 192 256
rect 140 218 192 222
rect 140 184 149 218
rect 149 184 183 218
rect 183 184 192 218
rect 140 170 192 184
rect 140 146 192 158
rect 140 112 149 146
rect 149 112 183 146
rect 183 112 192 146
rect 140 106 192 112
rect 226 1082 278 1088
rect 226 1048 235 1082
rect 235 1048 269 1082
rect 269 1048 278 1082
rect 226 1036 278 1048
rect 226 1010 278 1024
rect 226 976 235 1010
rect 235 976 269 1010
rect 269 976 278 1010
rect 226 972 278 976
rect 226 938 278 960
rect 226 908 235 938
rect 235 908 269 938
rect 269 908 278 938
rect 226 866 278 896
rect 226 844 235 866
rect 235 844 269 866
rect 269 844 278 866
rect 226 794 278 832
rect 226 780 235 794
rect 235 780 269 794
rect 269 780 278 794
rect 226 760 235 768
rect 235 760 269 768
rect 269 760 278 768
rect 226 722 278 760
rect 226 716 235 722
rect 235 716 269 722
rect 269 716 278 722
rect 226 688 235 704
rect 235 688 269 704
rect 269 688 278 704
rect 226 652 278 688
rect 226 616 235 640
rect 235 616 269 640
rect 269 616 278 640
rect 226 588 278 616
rect 226 544 235 576
rect 235 544 269 576
rect 269 544 278 576
rect 226 524 278 544
rect 226 506 278 512
rect 226 472 235 506
rect 235 472 269 506
rect 269 472 278 506
rect 226 460 278 472
rect 226 434 278 448
rect 226 400 235 434
rect 235 400 269 434
rect 269 400 278 434
rect 226 396 278 400
rect 226 362 278 384
rect 226 332 235 362
rect 235 332 269 362
rect 269 332 278 362
rect 226 290 278 320
rect 226 268 235 290
rect 235 268 269 290
rect 269 268 278 290
rect 226 218 278 256
rect 226 204 235 218
rect 235 204 269 218
rect 269 204 278 218
rect 226 184 235 192
rect 235 184 269 192
rect 269 184 278 192
rect 226 146 278 184
rect 226 140 235 146
rect 235 140 269 146
rect 269 140 278 146
rect 312 1048 321 1054
rect 321 1048 355 1054
rect 355 1048 364 1054
rect 312 1010 364 1048
rect 312 1002 321 1010
rect 321 1002 355 1010
rect 355 1002 364 1010
rect 312 976 321 990
rect 321 976 355 990
rect 355 976 364 990
rect 312 938 364 976
rect 312 904 321 926
rect 321 904 355 926
rect 355 904 364 926
rect 312 874 364 904
rect 312 832 321 862
rect 321 832 355 862
rect 355 832 364 862
rect 312 810 364 832
rect 312 794 364 798
rect 312 760 321 794
rect 321 760 355 794
rect 355 760 364 794
rect 312 746 364 760
rect 312 722 364 734
rect 312 688 321 722
rect 321 688 355 722
rect 355 688 364 722
rect 312 682 364 688
rect 312 650 364 670
rect 312 618 321 650
rect 321 618 355 650
rect 355 618 364 650
rect 312 578 364 606
rect 312 554 321 578
rect 321 554 355 578
rect 355 554 364 578
rect 312 506 364 542
rect 312 490 321 506
rect 321 490 355 506
rect 355 490 364 506
rect 312 472 321 478
rect 321 472 355 478
rect 355 472 364 478
rect 312 434 364 472
rect 312 426 321 434
rect 321 426 355 434
rect 355 426 364 434
rect 312 400 321 414
rect 321 400 355 414
rect 355 400 364 414
rect 312 362 364 400
rect 312 328 321 350
rect 321 328 355 350
rect 355 328 364 350
rect 312 298 364 328
rect 312 256 321 286
rect 321 256 355 286
rect 355 256 364 286
rect 312 234 364 256
rect 312 218 364 222
rect 312 184 321 218
rect 321 184 355 218
rect 355 184 364 218
rect 312 170 364 184
rect 312 146 364 158
rect 312 112 321 146
rect 321 112 355 146
rect 355 112 364 146
rect 312 106 364 112
rect 398 1082 450 1088
rect 398 1048 407 1082
rect 407 1048 441 1082
rect 441 1048 450 1082
rect 398 1036 450 1048
rect 398 1010 450 1024
rect 398 976 407 1010
rect 407 976 441 1010
rect 441 976 450 1010
rect 398 972 450 976
rect 398 938 450 960
rect 398 908 407 938
rect 407 908 441 938
rect 441 908 450 938
rect 398 866 450 896
rect 398 844 407 866
rect 407 844 441 866
rect 441 844 450 866
rect 398 794 450 832
rect 398 780 407 794
rect 407 780 441 794
rect 441 780 450 794
rect 398 760 407 768
rect 407 760 441 768
rect 441 760 450 768
rect 398 722 450 760
rect 398 716 407 722
rect 407 716 441 722
rect 441 716 450 722
rect 398 688 407 704
rect 407 688 441 704
rect 441 688 450 704
rect 398 652 450 688
rect 398 616 407 640
rect 407 616 441 640
rect 441 616 450 640
rect 398 588 450 616
rect 398 544 407 576
rect 407 544 441 576
rect 441 544 450 576
rect 398 524 450 544
rect 398 506 450 512
rect 398 472 407 506
rect 407 472 441 506
rect 441 472 450 506
rect 398 460 450 472
rect 398 434 450 448
rect 398 400 407 434
rect 407 400 441 434
rect 441 400 450 434
rect 398 396 450 400
rect 398 362 450 384
rect 398 332 407 362
rect 407 332 441 362
rect 441 332 450 362
rect 398 290 450 320
rect 398 268 407 290
rect 407 268 441 290
rect 441 268 450 290
rect 398 218 450 256
rect 398 204 407 218
rect 407 204 441 218
rect 441 204 450 218
rect 398 184 407 192
rect 407 184 441 192
rect 441 184 450 192
rect 398 146 450 184
rect 398 140 407 146
rect 407 140 441 146
rect 441 140 450 146
rect 484 1048 493 1054
rect 493 1048 527 1054
rect 527 1048 536 1054
rect 484 1010 536 1048
rect 484 1002 493 1010
rect 493 1002 527 1010
rect 527 1002 536 1010
rect 484 976 493 990
rect 493 976 527 990
rect 527 976 536 990
rect 484 938 536 976
rect 484 904 493 926
rect 493 904 527 926
rect 527 904 536 926
rect 484 874 536 904
rect 484 832 493 862
rect 493 832 527 862
rect 527 832 536 862
rect 484 810 536 832
rect 484 794 536 798
rect 484 760 493 794
rect 493 760 527 794
rect 527 760 536 794
rect 484 746 536 760
rect 484 722 536 734
rect 484 688 493 722
rect 493 688 527 722
rect 527 688 536 722
rect 484 682 536 688
rect 484 650 536 670
rect 484 618 493 650
rect 493 618 527 650
rect 527 618 536 650
rect 484 578 536 606
rect 484 554 493 578
rect 493 554 527 578
rect 527 554 536 578
rect 484 506 536 542
rect 484 490 493 506
rect 493 490 527 506
rect 527 490 536 506
rect 484 472 493 478
rect 493 472 527 478
rect 527 472 536 478
rect 484 434 536 472
rect 484 426 493 434
rect 493 426 527 434
rect 527 426 536 434
rect 484 400 493 414
rect 493 400 527 414
rect 527 400 536 414
rect 484 362 536 400
rect 484 328 493 350
rect 493 328 527 350
rect 527 328 536 350
rect 484 298 536 328
rect 484 256 493 286
rect 493 256 527 286
rect 527 256 536 286
rect 484 234 536 256
rect 484 218 536 222
rect 484 184 493 218
rect 493 184 527 218
rect 527 184 536 218
rect 484 170 536 184
rect 484 146 536 158
rect 484 112 493 146
rect 493 112 527 146
rect 527 112 536 146
rect 484 106 536 112
<< metal2 >>
rect 138 1202 538 1258
rect 138 1054 194 1202
rect 138 1002 140 1054
rect 192 1002 194 1054
rect 138 990 194 1002
rect 138 938 140 990
rect 192 938 194 990
rect 138 926 194 938
rect 138 874 140 926
rect 192 874 194 926
rect 138 862 194 874
rect 138 810 140 862
rect 192 810 194 862
rect 138 798 194 810
rect 138 746 140 798
rect 192 746 194 798
rect 138 734 194 746
rect 138 682 140 734
rect 192 682 194 734
rect 138 670 194 682
rect 138 618 140 670
rect 192 618 194 670
rect 138 606 194 618
rect 138 554 140 606
rect 192 554 194 606
rect 138 542 194 554
rect 138 490 140 542
rect 192 490 194 542
rect 138 478 194 490
rect 138 426 140 478
rect 192 426 194 478
rect 138 414 194 426
rect 138 362 140 414
rect 192 362 194 414
rect 138 350 194 362
rect 138 298 140 350
rect 192 298 194 350
rect 138 286 194 298
rect 138 234 140 286
rect 192 234 194 286
rect 138 222 194 234
rect 138 170 140 222
rect 192 170 194 222
rect 138 158 194 170
rect 138 106 140 158
rect 192 106 194 158
rect 138 92 194 106
rect 224 1088 280 1102
rect 224 1036 226 1088
rect 278 1036 280 1088
rect 224 1024 280 1036
rect 224 972 226 1024
rect 278 972 280 1024
rect 224 960 280 972
rect 224 908 226 960
rect 278 908 280 960
rect 224 896 280 908
rect 224 844 226 896
rect 278 844 280 896
rect 224 832 280 844
rect 224 780 226 832
rect 278 780 280 832
rect 224 768 280 780
rect 224 716 226 768
rect 278 716 280 768
rect 224 704 280 716
rect 224 652 226 704
rect 278 652 280 704
rect 224 640 280 652
rect 224 588 226 640
rect 278 588 280 640
rect 224 576 280 588
rect 224 524 226 576
rect 278 524 280 576
rect 224 512 280 524
rect 224 460 226 512
rect 278 460 280 512
rect 224 448 280 460
rect 224 396 226 448
rect 278 396 280 448
rect 224 384 280 396
rect 224 332 226 384
rect 278 332 280 384
rect 224 320 280 332
rect 224 268 226 320
rect 278 268 280 320
rect 224 256 280 268
rect 224 204 226 256
rect 278 204 280 256
rect 224 192 280 204
rect 224 140 226 192
rect 278 140 280 192
rect 224 -8 280 140
rect 310 1054 366 1202
rect 310 1002 312 1054
rect 364 1002 366 1054
rect 310 990 366 1002
rect 310 938 312 990
rect 364 938 366 990
rect 310 926 366 938
rect 310 874 312 926
rect 364 874 366 926
rect 310 862 366 874
rect 310 810 312 862
rect 364 810 366 862
rect 310 798 366 810
rect 310 746 312 798
rect 364 746 366 798
rect 310 734 366 746
rect 310 682 312 734
rect 364 682 366 734
rect 310 670 366 682
rect 310 618 312 670
rect 364 618 366 670
rect 310 606 366 618
rect 310 554 312 606
rect 364 554 366 606
rect 310 542 366 554
rect 310 490 312 542
rect 364 490 366 542
rect 310 478 366 490
rect 310 426 312 478
rect 364 426 366 478
rect 310 414 366 426
rect 310 362 312 414
rect 364 362 366 414
rect 310 350 366 362
rect 310 298 312 350
rect 364 298 366 350
rect 310 286 366 298
rect 310 234 312 286
rect 364 234 366 286
rect 310 222 366 234
rect 310 170 312 222
rect 364 170 366 222
rect 310 158 366 170
rect 310 106 312 158
rect 364 106 366 158
rect 310 92 366 106
rect 396 1088 452 1102
rect 396 1036 398 1088
rect 450 1036 452 1088
rect 396 1024 452 1036
rect 396 972 398 1024
rect 450 972 452 1024
rect 396 960 452 972
rect 396 908 398 960
rect 450 908 452 960
rect 396 896 452 908
rect 396 844 398 896
rect 450 844 452 896
rect 396 832 452 844
rect 396 780 398 832
rect 450 780 452 832
rect 396 768 452 780
rect 396 716 398 768
rect 450 716 452 768
rect 396 704 452 716
rect 396 652 398 704
rect 450 652 452 704
rect 396 640 452 652
rect 396 588 398 640
rect 450 588 452 640
rect 396 576 452 588
rect 396 524 398 576
rect 450 524 452 576
rect 396 512 452 524
rect 396 460 398 512
rect 450 460 452 512
rect 396 448 452 460
rect 396 396 398 448
rect 450 396 452 448
rect 396 384 452 396
rect 396 332 398 384
rect 450 332 452 384
rect 396 320 452 332
rect 396 268 398 320
rect 450 268 452 320
rect 396 256 452 268
rect 396 204 398 256
rect 450 204 452 256
rect 396 192 452 204
rect 396 140 398 192
rect 450 140 452 192
rect 396 -8 452 140
rect 482 1054 538 1202
rect 482 1002 484 1054
rect 536 1002 538 1054
rect 482 990 538 1002
rect 482 938 484 990
rect 536 938 538 990
rect 482 926 538 938
rect 482 874 484 926
rect 536 874 538 926
rect 482 862 538 874
rect 482 810 484 862
rect 536 810 538 862
rect 482 798 538 810
rect 482 746 484 798
rect 536 746 538 798
rect 482 734 538 746
rect 482 682 484 734
rect 536 682 538 734
rect 482 670 538 682
rect 482 618 484 670
rect 536 618 538 670
rect 482 606 538 618
rect 482 554 484 606
rect 536 554 538 606
rect 482 542 538 554
rect 482 490 484 542
rect 536 490 538 542
rect 482 478 538 490
rect 482 426 484 478
rect 536 426 538 478
rect 482 414 538 426
rect 482 362 484 414
rect 536 362 538 414
rect 482 350 538 362
rect 482 298 484 350
rect 536 298 538 350
rect 482 286 538 298
rect 482 234 484 286
rect 536 234 538 286
rect 482 222 538 234
rect 482 170 484 222
rect 536 170 538 222
rect 482 158 538 170
rect 482 106 484 158
rect 536 106 538 158
rect 482 92 538 106
rect 224 -64 452 -8
<< labels >>
rlabel metal2 138 1202 538 1258 1 D
rlabel metal2 224 -64 452 -8 1 S
rlabel metal1 25 100 84 1094 1 B
rlabel metal1 592 99 651 1093 1 B
rlabel metal1 165 -1 511 66 1 G
<< end >>
