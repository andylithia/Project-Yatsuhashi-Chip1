magic
tech sky130B
timestamp 1659501637
<< metal1 >>
rect 0 1990 2000 2000
rect 0 1955 75 1990
rect 175 1955 325 1990
rect 425 1955 575 1990
rect 675 1955 825 1990
rect 925 1955 1075 1990
rect 1175 1955 1325 1990
rect 1425 1955 1575 1990
rect 1675 1955 1825 1990
rect 1925 1955 2000 1990
rect 0 1950 2000 1955
rect 0 1940 60 1950
rect 190 1940 310 1950
rect 440 1940 560 1950
rect 690 1940 810 1950
rect 940 1940 1060 1950
rect 1190 1940 1310 1950
rect 1440 1940 1560 1950
rect 1690 1940 1810 1950
rect 1940 1940 2000 1950
rect 0 1925 50 1940
rect 0 1825 10 1925
rect 45 1825 50 1925
rect 0 1810 50 1825
rect 200 1925 300 1940
rect 200 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 300 1925
rect 200 1810 300 1825
rect 450 1925 550 1940
rect 450 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 550 1925
rect 450 1810 550 1825
rect 700 1925 800 1940
rect 700 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 800 1925
rect 700 1810 800 1825
rect 950 1925 1050 1940
rect 950 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1050 1925
rect 950 1810 1050 1825
rect 1200 1925 1300 1940
rect 1200 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1300 1925
rect 1200 1810 1300 1825
rect 1450 1925 1550 1940
rect 1450 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1550 1925
rect 1450 1810 1550 1825
rect 1700 1925 1800 1940
rect 1700 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1800 1925
rect 1700 1810 1800 1825
rect 1950 1925 2000 1940
rect 1950 1825 1955 1925
rect 1990 1825 2000 1925
rect 1950 1810 2000 1825
rect 0 1800 60 1810
rect 190 1800 310 1810
rect 440 1800 560 1810
rect 690 1800 810 1810
rect 940 1800 1060 1810
rect 1190 1800 1310 1810
rect 1440 1800 1560 1810
rect 1690 1800 1810 1810
rect 1940 1800 2000 1810
rect 0 1795 2000 1800
rect 0 1760 75 1795
rect 175 1760 325 1795
rect 425 1760 575 1795
rect 675 1760 825 1795
rect 925 1760 1075 1795
rect 1175 1760 1325 1795
rect 1425 1760 1575 1795
rect 1675 1760 1825 1795
rect 1925 1760 2000 1795
rect 0 1740 2000 1760
rect 0 1705 75 1740
rect 175 1705 325 1740
rect 425 1705 575 1740
rect 675 1705 825 1740
rect 925 1705 1075 1740
rect 1175 1705 1325 1740
rect 1425 1705 1575 1740
rect 1675 1705 1825 1740
rect 1925 1705 2000 1740
rect 0 1700 2000 1705
rect 0 1690 60 1700
rect 190 1690 310 1700
rect 440 1690 560 1700
rect 690 1690 810 1700
rect 940 1690 1060 1700
rect 1190 1690 1310 1700
rect 1440 1690 1560 1700
rect 1690 1690 1810 1700
rect 1940 1690 2000 1700
rect 0 1675 50 1690
rect 0 1575 10 1675
rect 45 1575 50 1675
rect 0 1560 50 1575
rect 200 1675 300 1690
rect 200 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 300 1675
rect 200 1560 300 1575
rect 450 1675 550 1690
rect 450 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 550 1675
rect 450 1560 550 1575
rect 700 1675 800 1690
rect 700 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 800 1675
rect 700 1560 800 1575
rect 950 1675 1050 1690
rect 950 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1050 1675
rect 950 1560 1050 1575
rect 1200 1675 1300 1690
rect 1200 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1300 1675
rect 1200 1560 1300 1575
rect 1450 1675 1550 1690
rect 1450 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1550 1675
rect 1450 1560 1550 1575
rect 1700 1675 1800 1690
rect 1700 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1800 1675
rect 1700 1560 1800 1575
rect 1950 1675 2000 1690
rect 1950 1575 1955 1675
rect 1990 1575 2000 1675
rect 1950 1560 2000 1575
rect 0 1550 60 1560
rect 190 1550 310 1560
rect 440 1550 560 1560
rect 690 1550 810 1560
rect 940 1550 1060 1560
rect 1190 1550 1310 1560
rect 1440 1550 1560 1560
rect 1690 1550 1810 1560
rect 1940 1550 2000 1560
rect 0 1545 2000 1550
rect 0 1510 75 1545
rect 175 1510 325 1545
rect 425 1510 575 1545
rect 675 1510 825 1545
rect 925 1510 1075 1545
rect 1175 1510 1325 1545
rect 1425 1510 1575 1545
rect 1675 1510 1825 1545
rect 1925 1510 2000 1545
rect 0 1490 2000 1510
rect 0 1455 75 1490
rect 175 1455 325 1490
rect 425 1455 575 1490
rect 675 1455 825 1490
rect 925 1455 1075 1490
rect 1175 1455 1325 1490
rect 1425 1455 1575 1490
rect 1675 1455 1825 1490
rect 1925 1455 2000 1490
rect 0 1450 2000 1455
rect 0 1440 60 1450
rect 190 1440 310 1450
rect 440 1440 560 1450
rect 690 1440 810 1450
rect 940 1440 1060 1450
rect 1190 1440 1310 1450
rect 1440 1440 1560 1450
rect 1690 1440 1810 1450
rect 1940 1440 2000 1450
rect 0 1425 50 1440
rect 0 1325 10 1425
rect 45 1325 50 1425
rect 0 1310 50 1325
rect 200 1425 300 1440
rect 200 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 300 1425
rect 200 1310 300 1325
rect 450 1425 550 1440
rect 450 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 550 1425
rect 450 1310 550 1325
rect 700 1425 800 1440
rect 700 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 800 1425
rect 700 1310 800 1325
rect 950 1425 1050 1440
rect 950 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1050 1425
rect 950 1310 1050 1325
rect 1200 1425 1300 1440
rect 1200 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1300 1425
rect 1200 1310 1300 1325
rect 1450 1425 1550 1440
rect 1450 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1550 1425
rect 1450 1310 1550 1325
rect 1700 1425 1800 1440
rect 1700 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1800 1425
rect 1700 1310 1800 1325
rect 1950 1425 2000 1440
rect 1950 1325 1955 1425
rect 1990 1325 2000 1425
rect 1950 1310 2000 1325
rect 0 1300 60 1310
rect 190 1300 310 1310
rect 440 1300 560 1310
rect 690 1300 810 1310
rect 940 1300 1060 1310
rect 1190 1300 1310 1310
rect 1440 1300 1560 1310
rect 1690 1300 1810 1310
rect 1940 1300 2000 1310
rect 0 1295 2000 1300
rect 0 1260 75 1295
rect 175 1260 325 1295
rect 425 1260 575 1295
rect 675 1260 825 1295
rect 925 1260 1075 1295
rect 1175 1260 1325 1295
rect 1425 1260 1575 1295
rect 1675 1260 1825 1295
rect 1925 1260 2000 1295
rect 0 1240 2000 1260
rect 0 1205 75 1240
rect 175 1205 325 1240
rect 425 1205 575 1240
rect 675 1205 825 1240
rect 925 1205 1075 1240
rect 1175 1205 1325 1240
rect 1425 1205 1575 1240
rect 1675 1205 1825 1240
rect 1925 1205 2000 1240
rect 0 1200 2000 1205
rect 0 1190 60 1200
rect 190 1190 310 1200
rect 440 1190 560 1200
rect 690 1190 810 1200
rect 940 1190 1060 1200
rect 1190 1190 1310 1200
rect 1440 1190 1560 1200
rect 1690 1190 1810 1200
rect 1940 1190 2000 1200
rect 0 1175 50 1190
rect 0 1075 10 1175
rect 45 1075 50 1175
rect 0 1060 50 1075
rect 200 1175 300 1190
rect 200 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 300 1175
rect 200 1060 300 1075
rect 450 1175 550 1190
rect 450 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 550 1175
rect 450 1060 550 1075
rect 700 1175 800 1190
rect 700 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 800 1175
rect 700 1060 800 1075
rect 950 1175 1050 1190
rect 950 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1050 1175
rect 950 1060 1050 1075
rect 1200 1175 1300 1190
rect 1200 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1300 1175
rect 1200 1060 1300 1075
rect 1450 1175 1550 1190
rect 1450 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1550 1175
rect 1450 1060 1550 1075
rect 1700 1175 1800 1190
rect 1700 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1800 1175
rect 1700 1060 1800 1075
rect 1950 1175 2000 1190
rect 1950 1075 1955 1175
rect 1990 1075 2000 1175
rect 1950 1060 2000 1075
rect 0 1050 60 1060
rect 190 1050 310 1060
rect 440 1050 560 1060
rect 690 1050 810 1060
rect 940 1050 1060 1060
rect 1190 1050 1310 1060
rect 1440 1050 1560 1060
rect 1690 1050 1810 1060
rect 1940 1050 2000 1060
rect 0 1045 2000 1050
rect 0 1010 75 1045
rect 175 1010 325 1045
rect 425 1010 575 1045
rect 675 1010 825 1045
rect 925 1010 1075 1045
rect 1175 1010 1325 1045
rect 1425 1010 1575 1045
rect 1675 1010 1825 1045
rect 1925 1010 2000 1045
rect 0 990 2000 1010
rect 0 955 75 990
rect 175 955 325 990
rect 425 955 575 990
rect 675 955 825 990
rect 925 955 1075 990
rect 1175 955 1325 990
rect 1425 955 1575 990
rect 1675 955 1825 990
rect 1925 955 2000 990
rect 0 950 2000 955
rect 0 940 60 950
rect 190 940 310 950
rect 440 940 560 950
rect 690 940 810 950
rect 940 940 1060 950
rect 1190 940 1310 950
rect 1440 940 1560 950
rect 1690 940 1810 950
rect 1940 940 2000 950
rect 0 925 50 940
rect 0 825 10 925
rect 45 825 50 925
rect 0 810 50 825
rect 200 925 300 940
rect 200 825 205 925
rect 240 825 260 925
rect 295 825 300 925
rect 200 810 300 825
rect 450 925 550 940
rect 450 825 455 925
rect 490 825 510 925
rect 545 825 550 925
rect 450 810 550 825
rect 700 925 800 940
rect 700 825 705 925
rect 740 825 760 925
rect 795 825 800 925
rect 700 810 800 825
rect 950 925 1050 940
rect 950 825 955 925
rect 990 825 1010 925
rect 1045 825 1050 925
rect 950 810 1050 825
rect 1200 925 1300 940
rect 1200 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1300 925
rect 1200 810 1300 825
rect 1450 925 1550 940
rect 1450 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1550 925
rect 1450 810 1550 825
rect 1700 925 1800 940
rect 1700 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1800 925
rect 1700 810 1800 825
rect 1950 925 2000 940
rect 1950 825 1955 925
rect 1990 825 2000 925
rect 1950 810 2000 825
rect 0 800 60 810
rect 190 800 310 810
rect 440 800 560 810
rect 690 800 810 810
rect 940 800 1060 810
rect 1190 800 1310 810
rect 1440 800 1560 810
rect 1690 800 1810 810
rect 1940 800 2000 810
rect 0 795 2000 800
rect 0 760 75 795
rect 175 760 325 795
rect 425 760 575 795
rect 675 760 825 795
rect 925 760 1075 795
rect 1175 760 1325 795
rect 1425 760 1575 795
rect 1675 760 1825 795
rect 1925 760 2000 795
rect 0 740 2000 760
rect 0 705 75 740
rect 175 705 325 740
rect 425 705 575 740
rect 675 705 825 740
rect 925 705 1075 740
rect 1175 705 1325 740
rect 1425 705 1575 740
rect 1675 705 1825 740
rect 1925 705 2000 740
rect 0 700 2000 705
rect 0 690 60 700
rect 190 690 310 700
rect 440 690 560 700
rect 690 690 810 700
rect 940 690 1060 700
rect 1190 690 1310 700
rect 1440 690 1560 700
rect 1690 690 1810 700
rect 1940 690 2000 700
rect 0 675 50 690
rect 0 575 10 675
rect 45 575 50 675
rect 0 560 50 575
rect 200 675 300 690
rect 200 575 205 675
rect 240 575 260 675
rect 295 575 300 675
rect 200 560 300 575
rect 450 675 550 690
rect 450 575 455 675
rect 490 575 510 675
rect 545 575 550 675
rect 450 560 550 575
rect 700 675 800 690
rect 700 575 705 675
rect 740 575 760 675
rect 795 575 800 675
rect 700 560 800 575
rect 950 675 1050 690
rect 950 575 955 675
rect 990 575 1010 675
rect 1045 575 1050 675
rect 950 560 1050 575
rect 1200 675 1300 690
rect 1200 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1300 675
rect 1200 560 1300 575
rect 1450 675 1550 690
rect 1450 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1550 675
rect 1450 560 1550 575
rect 1700 675 1800 690
rect 1700 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1800 675
rect 1700 560 1800 575
rect 1950 675 2000 690
rect 1950 575 1955 675
rect 1990 575 2000 675
rect 1950 560 2000 575
rect 0 550 60 560
rect 190 550 310 560
rect 440 550 560 560
rect 690 550 810 560
rect 940 550 1060 560
rect 1190 550 1310 560
rect 1440 550 1560 560
rect 1690 550 1810 560
rect 1940 550 2000 560
rect 0 545 2000 550
rect 0 510 75 545
rect 175 510 325 545
rect 425 510 575 545
rect 675 510 825 545
rect 925 510 1075 545
rect 1175 510 1325 545
rect 1425 510 1575 545
rect 1675 510 1825 545
rect 1925 510 2000 545
rect 0 490 2000 510
rect 0 455 75 490
rect 175 455 325 490
rect 425 455 575 490
rect 675 455 825 490
rect 925 455 1075 490
rect 1175 455 1325 490
rect 1425 455 1575 490
rect 1675 455 1825 490
rect 1925 455 2000 490
rect 0 450 2000 455
rect 0 440 60 450
rect 190 440 310 450
rect 440 440 560 450
rect 690 440 810 450
rect 940 440 1060 450
rect 1190 440 1310 450
rect 1440 440 1560 450
rect 1690 440 1810 450
rect 1940 440 2000 450
rect 0 425 50 440
rect 0 325 10 425
rect 45 325 50 425
rect 0 310 50 325
rect 200 425 300 440
rect 200 325 205 425
rect 240 325 260 425
rect 295 325 300 425
rect 200 310 300 325
rect 450 425 550 440
rect 450 325 455 425
rect 490 325 510 425
rect 545 325 550 425
rect 450 310 550 325
rect 700 425 800 440
rect 700 325 705 425
rect 740 325 760 425
rect 795 325 800 425
rect 700 310 800 325
rect 950 425 1050 440
rect 950 325 955 425
rect 990 325 1010 425
rect 1045 325 1050 425
rect 950 310 1050 325
rect 1200 425 1300 440
rect 1200 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1300 425
rect 1200 310 1300 325
rect 1450 425 1550 440
rect 1450 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1550 425
rect 1450 310 1550 325
rect 1700 425 1800 440
rect 1700 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1800 425
rect 1700 310 1800 325
rect 1950 425 2000 440
rect 1950 325 1955 425
rect 1990 325 2000 425
rect 1950 310 2000 325
rect 0 300 60 310
rect 190 300 310 310
rect 440 300 560 310
rect 690 300 810 310
rect 940 300 1060 310
rect 1190 300 1310 310
rect 1440 300 1560 310
rect 1690 300 1810 310
rect 1940 300 2000 310
rect 0 295 2000 300
rect 0 260 75 295
rect 175 260 325 295
rect 425 260 575 295
rect 675 260 825 295
rect 925 260 1075 295
rect 1175 260 1325 295
rect 1425 260 1575 295
rect 1675 260 1825 295
rect 1925 260 2000 295
rect 0 240 2000 260
rect 0 205 75 240
rect 175 205 325 240
rect 425 205 575 240
rect 675 205 825 240
rect 925 205 1075 240
rect 1175 205 1325 240
rect 1425 205 1575 240
rect 1675 205 1825 240
rect 1925 205 2000 240
rect 0 200 2000 205
rect 0 190 60 200
rect 190 190 310 200
rect 440 190 560 200
rect 690 190 810 200
rect 940 190 1060 200
rect 1190 190 1310 200
rect 1440 190 1560 200
rect 1690 190 1810 200
rect 1940 190 2000 200
rect 0 175 50 190
rect 0 75 10 175
rect 45 75 50 175
rect 0 60 50 75
rect 200 175 300 190
rect 200 75 205 175
rect 240 75 260 175
rect 295 75 300 175
rect 200 60 300 75
rect 450 175 550 190
rect 450 75 455 175
rect 490 75 510 175
rect 545 75 550 175
rect 450 60 550 75
rect 700 175 800 190
rect 700 75 705 175
rect 740 75 760 175
rect 795 75 800 175
rect 700 60 800 75
rect 950 175 1050 190
rect 950 75 955 175
rect 990 75 1010 175
rect 1045 75 1050 175
rect 950 60 1050 75
rect 1200 175 1300 190
rect 1200 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1300 175
rect 1200 60 1300 75
rect 1450 175 1550 190
rect 1450 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1550 175
rect 1450 60 1550 75
rect 1700 175 1800 190
rect 1700 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1800 175
rect 1700 60 1800 75
rect 1950 175 2000 190
rect 1950 75 1955 175
rect 1990 75 2000 175
rect 1950 60 2000 75
rect 0 50 60 60
rect 190 50 310 60
rect 440 50 560 60
rect 690 50 810 60
rect 940 50 1060 60
rect 1190 50 1310 60
rect 1440 50 1560 60
rect 1690 50 1810 60
rect 1940 50 2000 60
rect 0 45 2000 50
rect 0 10 75 45
rect 175 10 325 45
rect 425 10 575 45
rect 675 10 825 45
rect 925 10 1075 45
rect 1175 10 1325 45
rect 1425 10 1575 45
rect 1675 10 1825 45
rect 1925 10 2000 45
rect 0 0 2000 10
<< via1 >>
rect 75 1955 175 1990
rect 325 1955 425 1990
rect 575 1955 675 1990
rect 825 1955 925 1990
rect 1075 1955 1175 1990
rect 1325 1955 1425 1990
rect 1575 1955 1675 1990
rect 1825 1955 1925 1990
rect 10 1825 45 1925
rect 205 1825 240 1925
rect 260 1825 295 1925
rect 455 1825 490 1925
rect 510 1825 545 1925
rect 705 1825 740 1925
rect 760 1825 795 1925
rect 955 1825 990 1925
rect 1010 1825 1045 1925
rect 1205 1825 1240 1925
rect 1260 1825 1295 1925
rect 1455 1825 1490 1925
rect 1510 1825 1545 1925
rect 1705 1825 1740 1925
rect 1760 1825 1795 1925
rect 1955 1825 1990 1925
rect 75 1760 175 1795
rect 325 1760 425 1795
rect 575 1760 675 1795
rect 825 1760 925 1795
rect 1075 1760 1175 1795
rect 1325 1760 1425 1795
rect 1575 1760 1675 1795
rect 1825 1760 1925 1795
rect 75 1705 175 1740
rect 325 1705 425 1740
rect 575 1705 675 1740
rect 825 1705 925 1740
rect 1075 1705 1175 1740
rect 1325 1705 1425 1740
rect 1575 1705 1675 1740
rect 1825 1705 1925 1740
rect 10 1575 45 1675
rect 205 1575 240 1675
rect 260 1575 295 1675
rect 455 1575 490 1675
rect 510 1575 545 1675
rect 705 1575 740 1675
rect 760 1575 795 1675
rect 955 1575 990 1675
rect 1010 1575 1045 1675
rect 1205 1575 1240 1675
rect 1260 1575 1295 1675
rect 1455 1575 1490 1675
rect 1510 1575 1545 1675
rect 1705 1575 1740 1675
rect 1760 1575 1795 1675
rect 1955 1575 1990 1675
rect 75 1510 175 1545
rect 325 1510 425 1545
rect 575 1510 675 1545
rect 825 1510 925 1545
rect 1075 1510 1175 1545
rect 1325 1510 1425 1545
rect 1575 1510 1675 1545
rect 1825 1510 1925 1545
rect 75 1455 175 1490
rect 325 1455 425 1490
rect 575 1455 675 1490
rect 825 1455 925 1490
rect 1075 1455 1175 1490
rect 1325 1455 1425 1490
rect 1575 1455 1675 1490
rect 1825 1455 1925 1490
rect 10 1325 45 1425
rect 205 1325 240 1425
rect 260 1325 295 1425
rect 455 1325 490 1425
rect 510 1325 545 1425
rect 705 1325 740 1425
rect 760 1325 795 1425
rect 955 1325 990 1425
rect 1010 1325 1045 1425
rect 1205 1325 1240 1425
rect 1260 1325 1295 1425
rect 1455 1325 1490 1425
rect 1510 1325 1545 1425
rect 1705 1325 1740 1425
rect 1760 1325 1795 1425
rect 1955 1325 1990 1425
rect 75 1260 175 1295
rect 325 1260 425 1295
rect 575 1260 675 1295
rect 825 1260 925 1295
rect 1075 1260 1175 1295
rect 1325 1260 1425 1295
rect 1575 1260 1675 1295
rect 1825 1260 1925 1295
rect 75 1205 175 1240
rect 325 1205 425 1240
rect 575 1205 675 1240
rect 825 1205 925 1240
rect 1075 1205 1175 1240
rect 1325 1205 1425 1240
rect 1575 1205 1675 1240
rect 1825 1205 1925 1240
rect 10 1075 45 1175
rect 205 1075 240 1175
rect 260 1075 295 1175
rect 455 1075 490 1175
rect 510 1075 545 1175
rect 705 1075 740 1175
rect 760 1075 795 1175
rect 955 1075 990 1175
rect 1010 1075 1045 1175
rect 1205 1075 1240 1175
rect 1260 1075 1295 1175
rect 1455 1075 1490 1175
rect 1510 1075 1545 1175
rect 1705 1075 1740 1175
rect 1760 1075 1795 1175
rect 1955 1075 1990 1175
rect 75 1010 175 1045
rect 325 1010 425 1045
rect 575 1010 675 1045
rect 825 1010 925 1045
rect 1075 1010 1175 1045
rect 1325 1010 1425 1045
rect 1575 1010 1675 1045
rect 1825 1010 1925 1045
rect 75 955 175 990
rect 325 955 425 990
rect 575 955 675 990
rect 825 955 925 990
rect 1075 955 1175 990
rect 1325 955 1425 990
rect 1575 955 1675 990
rect 1825 955 1925 990
rect 10 825 45 925
rect 205 825 240 925
rect 260 825 295 925
rect 455 825 490 925
rect 510 825 545 925
rect 705 825 740 925
rect 760 825 795 925
rect 955 825 990 925
rect 1010 825 1045 925
rect 1205 825 1240 925
rect 1260 825 1295 925
rect 1455 825 1490 925
rect 1510 825 1545 925
rect 1705 825 1740 925
rect 1760 825 1795 925
rect 1955 825 1990 925
rect 75 760 175 795
rect 325 760 425 795
rect 575 760 675 795
rect 825 760 925 795
rect 1075 760 1175 795
rect 1325 760 1425 795
rect 1575 760 1675 795
rect 1825 760 1925 795
rect 75 705 175 740
rect 325 705 425 740
rect 575 705 675 740
rect 825 705 925 740
rect 1075 705 1175 740
rect 1325 705 1425 740
rect 1575 705 1675 740
rect 1825 705 1925 740
rect 10 575 45 675
rect 205 575 240 675
rect 260 575 295 675
rect 455 575 490 675
rect 510 575 545 675
rect 705 575 740 675
rect 760 575 795 675
rect 955 575 990 675
rect 1010 575 1045 675
rect 1205 575 1240 675
rect 1260 575 1295 675
rect 1455 575 1490 675
rect 1510 575 1545 675
rect 1705 575 1740 675
rect 1760 575 1795 675
rect 1955 575 1990 675
rect 75 510 175 545
rect 325 510 425 545
rect 575 510 675 545
rect 825 510 925 545
rect 1075 510 1175 545
rect 1325 510 1425 545
rect 1575 510 1675 545
rect 1825 510 1925 545
rect 75 455 175 490
rect 325 455 425 490
rect 575 455 675 490
rect 825 455 925 490
rect 1075 455 1175 490
rect 1325 455 1425 490
rect 1575 455 1675 490
rect 1825 455 1925 490
rect 10 325 45 425
rect 205 325 240 425
rect 260 325 295 425
rect 455 325 490 425
rect 510 325 545 425
rect 705 325 740 425
rect 760 325 795 425
rect 955 325 990 425
rect 1010 325 1045 425
rect 1205 325 1240 425
rect 1260 325 1295 425
rect 1455 325 1490 425
rect 1510 325 1545 425
rect 1705 325 1740 425
rect 1760 325 1795 425
rect 1955 325 1990 425
rect 75 260 175 295
rect 325 260 425 295
rect 575 260 675 295
rect 825 260 925 295
rect 1075 260 1175 295
rect 1325 260 1425 295
rect 1575 260 1675 295
rect 1825 260 1925 295
rect 75 205 175 240
rect 325 205 425 240
rect 575 205 675 240
rect 825 205 925 240
rect 1075 205 1175 240
rect 1325 205 1425 240
rect 1575 205 1675 240
rect 1825 205 1925 240
rect 10 75 45 175
rect 205 75 240 175
rect 260 75 295 175
rect 455 75 490 175
rect 510 75 545 175
rect 705 75 740 175
rect 760 75 795 175
rect 955 75 990 175
rect 1010 75 1045 175
rect 1205 75 1240 175
rect 1260 75 1295 175
rect 1455 75 1490 175
rect 1510 75 1545 175
rect 1705 75 1740 175
rect 1760 75 1795 175
rect 1955 75 1990 175
rect 75 10 175 45
rect 325 10 425 45
rect 575 10 675 45
rect 825 10 925 45
rect 1075 10 1175 45
rect 1325 10 1425 45
rect 1575 10 1675 45
rect 1825 10 1925 45
<< metal2 >>
rect 70 1990 180 2000
rect 70 1955 75 1990
rect 175 1955 180 1990
rect 70 1930 180 1955
rect 320 1990 430 2000
rect 320 1955 325 1990
rect 425 1955 430 1990
rect 320 1930 430 1955
rect 570 1990 680 2000
rect 570 1955 575 1990
rect 675 1955 680 1990
rect 570 1930 680 1955
rect 820 1990 930 2000
rect 820 1955 825 1990
rect 925 1955 930 1990
rect 820 1930 930 1955
rect 1070 1990 1180 2000
rect 1070 1955 1075 1990
rect 1175 1955 1180 1990
rect 1070 1930 1180 1955
rect 1320 1990 1430 2000
rect 1320 1955 1325 1990
rect 1425 1955 1430 1990
rect 1320 1930 1430 1955
rect 1570 1990 1680 2000
rect 1570 1955 1575 1990
rect 1675 1955 1680 1990
rect 1570 1930 1680 1955
rect 1820 1990 1930 2000
rect 1820 1955 1825 1990
rect 1925 1955 1930 1990
rect 1820 1930 1930 1955
rect 0 1925 2000 1930
rect 0 1825 10 1925
rect 45 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1955 1925
rect 1990 1825 2000 1925
rect 0 1820 2000 1825
rect 70 1795 180 1820
rect 70 1760 75 1795
rect 175 1760 180 1795
rect 70 1740 180 1760
rect 70 1705 75 1740
rect 175 1705 180 1740
rect 70 1680 180 1705
rect 320 1795 430 1820
rect 320 1760 325 1795
rect 425 1760 430 1795
rect 320 1740 430 1760
rect 320 1705 325 1740
rect 425 1705 430 1740
rect 320 1680 430 1705
rect 570 1795 680 1820
rect 570 1760 575 1795
rect 675 1760 680 1795
rect 570 1740 680 1760
rect 570 1705 575 1740
rect 675 1705 680 1740
rect 570 1680 680 1705
rect 820 1795 930 1820
rect 820 1760 825 1795
rect 925 1760 930 1795
rect 820 1740 930 1760
rect 820 1705 825 1740
rect 925 1705 930 1740
rect 820 1680 930 1705
rect 1070 1795 1180 1820
rect 1070 1760 1075 1795
rect 1175 1760 1180 1795
rect 1070 1740 1180 1760
rect 1070 1705 1075 1740
rect 1175 1705 1180 1740
rect 1070 1680 1180 1705
rect 1320 1795 1430 1820
rect 1320 1760 1325 1795
rect 1425 1760 1430 1795
rect 1320 1740 1430 1760
rect 1320 1705 1325 1740
rect 1425 1705 1430 1740
rect 1320 1680 1430 1705
rect 1570 1795 1680 1820
rect 1570 1760 1575 1795
rect 1675 1760 1680 1795
rect 1570 1740 1680 1760
rect 1570 1705 1575 1740
rect 1675 1705 1680 1740
rect 1570 1680 1680 1705
rect 1820 1795 1930 1820
rect 1820 1760 1825 1795
rect 1925 1760 1930 1795
rect 1820 1740 1930 1760
rect 1820 1705 1825 1740
rect 1925 1705 1930 1740
rect 1820 1680 1930 1705
rect 0 1675 2000 1680
rect 0 1575 10 1675
rect 45 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1955 1675
rect 1990 1575 2000 1675
rect 0 1570 2000 1575
rect 70 1545 180 1570
rect 70 1510 75 1545
rect 175 1510 180 1545
rect 70 1490 180 1510
rect 70 1455 75 1490
rect 175 1455 180 1490
rect 70 1430 180 1455
rect 320 1545 430 1570
rect 320 1510 325 1545
rect 425 1510 430 1545
rect 320 1490 430 1510
rect 320 1455 325 1490
rect 425 1455 430 1490
rect 320 1430 430 1455
rect 570 1545 680 1570
rect 570 1510 575 1545
rect 675 1510 680 1545
rect 570 1490 680 1510
rect 570 1455 575 1490
rect 675 1455 680 1490
rect 570 1430 680 1455
rect 820 1545 930 1570
rect 820 1510 825 1545
rect 925 1510 930 1545
rect 820 1490 930 1510
rect 820 1455 825 1490
rect 925 1455 930 1490
rect 820 1430 930 1455
rect 1070 1545 1180 1570
rect 1070 1510 1075 1545
rect 1175 1510 1180 1545
rect 1070 1490 1180 1510
rect 1070 1455 1075 1490
rect 1175 1455 1180 1490
rect 1070 1430 1180 1455
rect 1320 1545 1430 1570
rect 1320 1510 1325 1545
rect 1425 1510 1430 1545
rect 1320 1490 1430 1510
rect 1320 1455 1325 1490
rect 1425 1455 1430 1490
rect 1320 1430 1430 1455
rect 1570 1545 1680 1570
rect 1570 1510 1575 1545
rect 1675 1510 1680 1545
rect 1570 1490 1680 1510
rect 1570 1455 1575 1490
rect 1675 1455 1680 1490
rect 1570 1430 1680 1455
rect 1820 1545 1930 1570
rect 1820 1510 1825 1545
rect 1925 1510 1930 1545
rect 1820 1490 1930 1510
rect 1820 1455 1825 1490
rect 1925 1455 1930 1490
rect 1820 1430 1930 1455
rect 0 1425 2000 1430
rect 0 1325 10 1425
rect 45 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1955 1425
rect 1990 1325 2000 1425
rect 0 1320 2000 1325
rect 70 1295 180 1320
rect 70 1260 75 1295
rect 175 1260 180 1295
rect 70 1240 180 1260
rect 70 1205 75 1240
rect 175 1205 180 1240
rect 70 1180 180 1205
rect 320 1295 430 1320
rect 320 1260 325 1295
rect 425 1260 430 1295
rect 320 1240 430 1260
rect 320 1205 325 1240
rect 425 1205 430 1240
rect 320 1180 430 1205
rect 570 1295 680 1320
rect 570 1260 575 1295
rect 675 1260 680 1295
rect 570 1240 680 1260
rect 570 1205 575 1240
rect 675 1205 680 1240
rect 570 1180 680 1205
rect 820 1295 930 1320
rect 820 1260 825 1295
rect 925 1260 930 1295
rect 820 1240 930 1260
rect 820 1205 825 1240
rect 925 1205 930 1240
rect 820 1180 930 1205
rect 1070 1295 1180 1320
rect 1070 1260 1075 1295
rect 1175 1260 1180 1295
rect 1070 1240 1180 1260
rect 1070 1205 1075 1240
rect 1175 1205 1180 1240
rect 1070 1180 1180 1205
rect 1320 1295 1430 1320
rect 1320 1260 1325 1295
rect 1425 1260 1430 1295
rect 1320 1240 1430 1260
rect 1320 1205 1325 1240
rect 1425 1205 1430 1240
rect 1320 1180 1430 1205
rect 1570 1295 1680 1320
rect 1570 1260 1575 1295
rect 1675 1260 1680 1295
rect 1570 1240 1680 1260
rect 1570 1205 1575 1240
rect 1675 1205 1680 1240
rect 1570 1180 1680 1205
rect 1820 1295 1930 1320
rect 1820 1260 1825 1295
rect 1925 1260 1930 1295
rect 1820 1240 1930 1260
rect 1820 1205 1825 1240
rect 1925 1205 1930 1240
rect 1820 1180 1930 1205
rect 0 1175 2000 1180
rect 0 1075 10 1175
rect 45 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1955 1175
rect 1990 1075 2000 1175
rect 0 1070 2000 1075
rect 70 1045 180 1070
rect 70 1010 75 1045
rect 175 1010 180 1045
rect 70 990 180 1010
rect 70 955 75 990
rect 175 955 180 990
rect 70 930 180 955
rect 320 1045 430 1070
rect 320 1010 325 1045
rect 425 1010 430 1045
rect 320 990 430 1010
rect 320 955 325 990
rect 425 955 430 990
rect 320 930 430 955
rect 570 1045 680 1070
rect 570 1010 575 1045
rect 675 1010 680 1045
rect 570 990 680 1010
rect 570 955 575 990
rect 675 955 680 990
rect 570 930 680 955
rect 820 1045 930 1070
rect 820 1010 825 1045
rect 925 1010 930 1045
rect 820 990 930 1010
rect 820 955 825 990
rect 925 955 930 990
rect 820 930 930 955
rect 1070 1045 1180 1070
rect 1070 1010 1075 1045
rect 1175 1010 1180 1045
rect 1070 990 1180 1010
rect 1070 955 1075 990
rect 1175 955 1180 990
rect 1070 930 1180 955
rect 1320 1045 1430 1070
rect 1320 1010 1325 1045
rect 1425 1010 1430 1045
rect 1320 990 1430 1010
rect 1320 955 1325 990
rect 1425 955 1430 990
rect 1320 930 1430 955
rect 1570 1045 1680 1070
rect 1570 1010 1575 1045
rect 1675 1010 1680 1045
rect 1570 990 1680 1010
rect 1570 955 1575 990
rect 1675 955 1680 990
rect 1570 930 1680 955
rect 1820 1045 1930 1070
rect 1820 1010 1825 1045
rect 1925 1010 1930 1045
rect 1820 990 1930 1010
rect 1820 955 1825 990
rect 1925 955 1930 990
rect 1820 930 1930 955
rect 0 925 2000 930
rect 0 825 10 925
rect 45 825 205 925
rect 240 825 260 925
rect 295 825 455 925
rect 490 825 510 925
rect 545 825 705 925
rect 740 825 760 925
rect 795 825 955 925
rect 990 825 1010 925
rect 1045 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1955 925
rect 1990 825 2000 925
rect 0 820 2000 825
rect 70 795 180 820
rect 70 760 75 795
rect 175 760 180 795
rect 70 740 180 760
rect 70 705 75 740
rect 175 705 180 740
rect 70 680 180 705
rect 320 795 430 820
rect 320 760 325 795
rect 425 760 430 795
rect 320 740 430 760
rect 320 705 325 740
rect 425 705 430 740
rect 320 680 430 705
rect 570 795 680 820
rect 570 760 575 795
rect 675 760 680 795
rect 570 740 680 760
rect 570 705 575 740
rect 675 705 680 740
rect 570 680 680 705
rect 820 795 930 820
rect 820 760 825 795
rect 925 760 930 795
rect 820 740 930 760
rect 820 705 825 740
rect 925 705 930 740
rect 820 680 930 705
rect 1070 795 1180 820
rect 1070 760 1075 795
rect 1175 760 1180 795
rect 1070 740 1180 760
rect 1070 705 1075 740
rect 1175 705 1180 740
rect 1070 680 1180 705
rect 1320 795 1430 820
rect 1320 760 1325 795
rect 1425 760 1430 795
rect 1320 740 1430 760
rect 1320 705 1325 740
rect 1425 705 1430 740
rect 1320 680 1430 705
rect 1570 795 1680 820
rect 1570 760 1575 795
rect 1675 760 1680 795
rect 1570 740 1680 760
rect 1570 705 1575 740
rect 1675 705 1680 740
rect 1570 680 1680 705
rect 1820 795 1930 820
rect 1820 760 1825 795
rect 1925 760 1930 795
rect 1820 740 1930 760
rect 1820 705 1825 740
rect 1925 705 1930 740
rect 1820 680 1930 705
rect 0 675 2000 680
rect 0 575 10 675
rect 45 575 205 675
rect 240 575 260 675
rect 295 575 455 675
rect 490 575 510 675
rect 545 575 705 675
rect 740 575 760 675
rect 795 575 955 675
rect 990 575 1010 675
rect 1045 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1955 675
rect 1990 575 2000 675
rect 0 570 2000 575
rect 70 545 180 570
rect 70 510 75 545
rect 175 510 180 545
rect 70 490 180 510
rect 70 455 75 490
rect 175 455 180 490
rect 70 430 180 455
rect 320 545 430 570
rect 320 510 325 545
rect 425 510 430 545
rect 320 490 430 510
rect 320 455 325 490
rect 425 455 430 490
rect 320 430 430 455
rect 570 545 680 570
rect 570 510 575 545
rect 675 510 680 545
rect 570 490 680 510
rect 570 455 575 490
rect 675 455 680 490
rect 570 430 680 455
rect 820 545 930 570
rect 820 510 825 545
rect 925 510 930 545
rect 820 490 930 510
rect 820 455 825 490
rect 925 455 930 490
rect 820 430 930 455
rect 1070 545 1180 570
rect 1070 510 1075 545
rect 1175 510 1180 545
rect 1070 490 1180 510
rect 1070 455 1075 490
rect 1175 455 1180 490
rect 1070 430 1180 455
rect 1320 545 1430 570
rect 1320 510 1325 545
rect 1425 510 1430 545
rect 1320 490 1430 510
rect 1320 455 1325 490
rect 1425 455 1430 490
rect 1320 430 1430 455
rect 1570 545 1680 570
rect 1570 510 1575 545
rect 1675 510 1680 545
rect 1570 490 1680 510
rect 1570 455 1575 490
rect 1675 455 1680 490
rect 1570 430 1680 455
rect 1820 545 1930 570
rect 1820 510 1825 545
rect 1925 510 1930 545
rect 1820 490 1930 510
rect 1820 455 1825 490
rect 1925 455 1930 490
rect 1820 430 1930 455
rect 0 425 2000 430
rect 0 325 10 425
rect 45 325 205 425
rect 240 325 260 425
rect 295 325 455 425
rect 490 325 510 425
rect 545 325 705 425
rect 740 325 760 425
rect 795 325 955 425
rect 990 325 1010 425
rect 1045 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1955 425
rect 1990 325 2000 425
rect 0 320 2000 325
rect 70 295 180 320
rect 70 260 75 295
rect 175 260 180 295
rect 70 240 180 260
rect 70 205 75 240
rect 175 205 180 240
rect 70 180 180 205
rect 320 295 430 320
rect 320 260 325 295
rect 425 260 430 295
rect 320 240 430 260
rect 320 205 325 240
rect 425 205 430 240
rect 320 180 430 205
rect 570 295 680 320
rect 570 260 575 295
rect 675 260 680 295
rect 570 240 680 260
rect 570 205 575 240
rect 675 205 680 240
rect 570 180 680 205
rect 820 295 930 320
rect 820 260 825 295
rect 925 260 930 295
rect 820 240 930 260
rect 820 205 825 240
rect 925 205 930 240
rect 820 180 930 205
rect 1070 295 1180 320
rect 1070 260 1075 295
rect 1175 260 1180 295
rect 1070 240 1180 260
rect 1070 205 1075 240
rect 1175 205 1180 240
rect 1070 180 1180 205
rect 1320 295 1430 320
rect 1320 260 1325 295
rect 1425 260 1430 295
rect 1320 240 1430 260
rect 1320 205 1325 240
rect 1425 205 1430 240
rect 1320 180 1430 205
rect 1570 295 1680 320
rect 1570 260 1575 295
rect 1675 260 1680 295
rect 1570 240 1680 260
rect 1570 205 1575 240
rect 1675 205 1680 240
rect 1570 180 1680 205
rect 1820 295 1930 320
rect 1820 260 1825 295
rect 1925 260 1930 295
rect 1820 240 1930 260
rect 1820 205 1825 240
rect 1925 205 1930 240
rect 1820 180 1930 205
rect 0 175 2000 180
rect 0 75 10 175
rect 45 75 205 175
rect 240 75 260 175
rect 295 75 455 175
rect 490 75 510 175
rect 545 75 705 175
rect 740 75 760 175
rect 795 75 955 175
rect 990 75 1010 175
rect 1045 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1955 175
rect 1990 75 2000 175
rect 0 70 2000 75
rect 70 45 180 70
rect 70 10 75 45
rect 175 10 180 45
rect 70 0 180 10
rect 320 45 430 70
rect 320 10 325 45
rect 425 10 430 45
rect 320 0 430 10
rect 570 45 680 70
rect 570 10 575 45
rect 675 10 680 45
rect 570 0 680 10
rect 820 45 930 70
rect 820 10 825 45
rect 925 10 930 45
rect 820 0 930 10
rect 1070 45 1180 70
rect 1070 10 1075 45
rect 1175 10 1180 45
rect 1070 0 1180 10
rect 1320 45 1430 70
rect 1320 10 1325 45
rect 1425 10 1430 45
rect 1320 0 1430 10
rect 1570 45 1680 70
rect 1570 10 1575 45
rect 1675 10 1680 45
rect 1570 0 1680 10
rect 1820 45 1930 70
rect 1820 10 1825 45
rect 1925 10 1930 45
rect 1820 0 1930 10
<< via2 >>
rect 75 1955 175 1990
rect 325 1955 425 1990
rect 575 1955 675 1990
rect 825 1955 925 1990
rect 1075 1955 1175 1990
rect 1325 1955 1425 1990
rect 1575 1955 1675 1990
rect 1825 1955 1925 1990
rect 10 1825 45 1925
rect 205 1825 240 1925
rect 260 1825 295 1925
rect 455 1825 490 1925
rect 510 1825 545 1925
rect 705 1825 740 1925
rect 760 1825 795 1925
rect 955 1825 990 1925
rect 1010 1825 1045 1925
rect 1205 1825 1240 1925
rect 1260 1825 1295 1925
rect 1455 1825 1490 1925
rect 1510 1825 1545 1925
rect 1705 1825 1740 1925
rect 1760 1825 1795 1925
rect 1955 1825 1990 1925
rect 75 1760 175 1795
rect 75 1705 175 1740
rect 325 1760 425 1795
rect 325 1705 425 1740
rect 575 1760 675 1795
rect 575 1705 675 1740
rect 825 1760 925 1795
rect 825 1705 925 1740
rect 1075 1760 1175 1795
rect 1075 1705 1175 1740
rect 1325 1760 1425 1795
rect 1325 1705 1425 1740
rect 1575 1760 1675 1795
rect 1575 1705 1675 1740
rect 1825 1760 1925 1795
rect 1825 1705 1925 1740
rect 10 1575 45 1675
rect 205 1575 240 1675
rect 260 1575 295 1675
rect 455 1575 490 1675
rect 510 1575 545 1675
rect 705 1575 740 1675
rect 760 1575 795 1675
rect 955 1575 990 1675
rect 1010 1575 1045 1675
rect 1205 1575 1240 1675
rect 1260 1575 1295 1675
rect 1455 1575 1490 1675
rect 1510 1575 1545 1675
rect 1705 1575 1740 1675
rect 1760 1575 1795 1675
rect 1955 1575 1990 1675
rect 75 1510 175 1545
rect 75 1455 175 1490
rect 325 1510 425 1545
rect 325 1455 425 1490
rect 575 1510 675 1545
rect 575 1455 675 1490
rect 825 1510 925 1545
rect 825 1455 925 1490
rect 1075 1510 1175 1545
rect 1075 1455 1175 1490
rect 1325 1510 1425 1545
rect 1325 1455 1425 1490
rect 1575 1510 1675 1545
rect 1575 1455 1675 1490
rect 1825 1510 1925 1545
rect 1825 1455 1925 1490
rect 10 1325 45 1425
rect 205 1325 240 1425
rect 260 1325 295 1425
rect 455 1325 490 1425
rect 510 1325 545 1425
rect 705 1325 740 1425
rect 760 1325 795 1425
rect 955 1325 990 1425
rect 1010 1325 1045 1425
rect 1205 1325 1240 1425
rect 1260 1325 1295 1425
rect 1455 1325 1490 1425
rect 1510 1325 1545 1425
rect 1705 1325 1740 1425
rect 1760 1325 1795 1425
rect 1955 1325 1990 1425
rect 75 1260 175 1295
rect 75 1205 175 1240
rect 325 1260 425 1295
rect 325 1205 425 1240
rect 575 1260 675 1295
rect 575 1205 675 1240
rect 825 1260 925 1295
rect 825 1205 925 1240
rect 1075 1260 1175 1295
rect 1075 1205 1175 1240
rect 1325 1260 1425 1295
rect 1325 1205 1425 1240
rect 1575 1260 1675 1295
rect 1575 1205 1675 1240
rect 1825 1260 1925 1295
rect 1825 1205 1925 1240
rect 10 1075 45 1175
rect 205 1075 240 1175
rect 260 1075 295 1175
rect 455 1075 490 1175
rect 510 1075 545 1175
rect 705 1075 740 1175
rect 760 1075 795 1175
rect 955 1075 990 1175
rect 1010 1075 1045 1175
rect 1205 1075 1240 1175
rect 1260 1075 1295 1175
rect 1455 1075 1490 1175
rect 1510 1075 1545 1175
rect 1705 1075 1740 1175
rect 1760 1075 1795 1175
rect 1955 1075 1990 1175
rect 75 1010 175 1045
rect 75 955 175 990
rect 325 1010 425 1045
rect 325 955 425 990
rect 575 1010 675 1045
rect 575 955 675 990
rect 825 1010 925 1045
rect 825 955 925 990
rect 1075 1010 1175 1045
rect 1075 955 1175 990
rect 1325 1010 1425 1045
rect 1325 955 1425 990
rect 1575 1010 1675 1045
rect 1575 955 1675 990
rect 1825 1010 1925 1045
rect 1825 955 1925 990
rect 10 825 45 925
rect 205 825 240 925
rect 260 825 295 925
rect 455 825 490 925
rect 510 825 545 925
rect 705 825 740 925
rect 760 825 795 925
rect 955 825 990 925
rect 1010 825 1045 925
rect 1205 825 1240 925
rect 1260 825 1295 925
rect 1455 825 1490 925
rect 1510 825 1545 925
rect 1705 825 1740 925
rect 1760 825 1795 925
rect 1955 825 1990 925
rect 75 760 175 795
rect 75 705 175 740
rect 325 760 425 795
rect 325 705 425 740
rect 575 760 675 795
rect 575 705 675 740
rect 825 760 925 795
rect 825 705 925 740
rect 1075 760 1175 795
rect 1075 705 1175 740
rect 1325 760 1425 795
rect 1325 705 1425 740
rect 1575 760 1675 795
rect 1575 705 1675 740
rect 1825 760 1925 795
rect 1825 705 1925 740
rect 10 575 45 675
rect 205 575 240 675
rect 260 575 295 675
rect 455 575 490 675
rect 510 575 545 675
rect 705 575 740 675
rect 760 575 795 675
rect 955 575 990 675
rect 1010 575 1045 675
rect 1205 575 1240 675
rect 1260 575 1295 675
rect 1455 575 1490 675
rect 1510 575 1545 675
rect 1705 575 1740 675
rect 1760 575 1795 675
rect 1955 575 1990 675
rect 75 510 175 545
rect 75 455 175 490
rect 325 510 425 545
rect 325 455 425 490
rect 575 510 675 545
rect 575 455 675 490
rect 825 510 925 545
rect 825 455 925 490
rect 1075 510 1175 545
rect 1075 455 1175 490
rect 1325 510 1425 545
rect 1325 455 1425 490
rect 1575 510 1675 545
rect 1575 455 1675 490
rect 1825 510 1925 545
rect 1825 455 1925 490
rect 10 325 45 425
rect 205 325 240 425
rect 260 325 295 425
rect 455 325 490 425
rect 510 325 545 425
rect 705 325 740 425
rect 760 325 795 425
rect 955 325 990 425
rect 1010 325 1045 425
rect 1205 325 1240 425
rect 1260 325 1295 425
rect 1455 325 1490 425
rect 1510 325 1545 425
rect 1705 325 1740 425
rect 1760 325 1795 425
rect 1955 325 1990 425
rect 75 260 175 295
rect 75 205 175 240
rect 325 260 425 295
rect 325 205 425 240
rect 575 260 675 295
rect 575 205 675 240
rect 825 260 925 295
rect 825 205 925 240
rect 1075 260 1175 295
rect 1075 205 1175 240
rect 1325 260 1425 295
rect 1325 205 1425 240
rect 1575 260 1675 295
rect 1575 205 1675 240
rect 1825 260 1925 295
rect 1825 205 1925 240
rect 10 75 45 175
rect 205 75 240 175
rect 260 75 295 175
rect 455 75 490 175
rect 510 75 545 175
rect 705 75 740 175
rect 760 75 795 175
rect 955 75 990 175
rect 1010 75 1045 175
rect 1205 75 1240 175
rect 1260 75 1295 175
rect 1455 75 1490 175
rect 1510 75 1545 175
rect 1705 75 1740 175
rect 1760 75 1795 175
rect 1955 75 1990 175
rect 75 10 175 45
rect 325 10 425 45
rect 575 10 675 45
rect 825 10 925 45
rect 1075 10 1175 45
rect 1325 10 1425 45
rect 1575 10 1675 45
rect 1825 10 1925 45
<< metal3 >>
rect 0 1990 2000 2000
rect 0 1955 75 1990
rect 175 1955 325 1990
rect 425 1955 575 1990
rect 675 1955 825 1990
rect 925 1955 1075 1990
rect 1175 1955 1325 1990
rect 1425 1955 1575 1990
rect 1675 1955 1825 1990
rect 1925 1955 2000 1990
rect 0 1950 2000 1955
rect 0 1940 60 1950
rect 190 1940 310 1950
rect 440 1940 560 1950
rect 690 1940 810 1950
rect 940 1940 1060 1950
rect 1190 1940 1310 1950
rect 1440 1940 1560 1950
rect 1690 1940 1810 1950
rect 1940 1940 2000 1950
rect 0 1925 50 1940
rect 0 1825 10 1925
rect 45 1825 50 1925
rect 0 1810 50 1825
rect 200 1925 300 1940
rect 200 1825 205 1925
rect 240 1825 260 1925
rect 295 1825 300 1925
rect 200 1810 300 1825
rect 450 1925 550 1940
rect 450 1825 455 1925
rect 490 1825 510 1925
rect 545 1825 550 1925
rect 450 1810 550 1825
rect 700 1925 800 1940
rect 700 1825 705 1925
rect 740 1825 760 1925
rect 795 1825 800 1925
rect 700 1810 800 1825
rect 950 1925 1050 1940
rect 950 1825 955 1925
rect 990 1825 1010 1925
rect 1045 1825 1050 1925
rect 950 1810 1050 1825
rect 1200 1925 1300 1940
rect 1200 1825 1205 1925
rect 1240 1825 1260 1925
rect 1295 1825 1300 1925
rect 1200 1810 1300 1825
rect 1450 1925 1550 1940
rect 1450 1825 1455 1925
rect 1490 1825 1510 1925
rect 1545 1825 1550 1925
rect 1450 1810 1550 1825
rect 1700 1925 1800 1940
rect 1700 1825 1705 1925
rect 1740 1825 1760 1925
rect 1795 1825 1800 1925
rect 1700 1810 1800 1825
rect 1950 1925 2000 1940
rect 1950 1825 1955 1925
rect 1990 1825 2000 1925
rect 1950 1810 2000 1825
rect 0 1800 60 1810
rect 190 1800 310 1810
rect 440 1800 560 1810
rect 690 1800 810 1810
rect 940 1800 1060 1810
rect 1190 1800 1310 1810
rect 1440 1800 1560 1810
rect 1690 1800 1810 1810
rect 1940 1800 2000 1810
rect 0 1795 200 1800
rect 0 1760 75 1795
rect 175 1760 200 1795
rect 0 1740 200 1760
rect 0 1705 75 1740
rect 175 1705 200 1740
rect 0 1700 200 1705
rect 300 1795 450 1800
rect 300 1760 325 1795
rect 425 1760 450 1795
rect 300 1740 450 1760
rect 300 1705 325 1740
rect 425 1705 450 1740
rect 300 1700 450 1705
rect 550 1795 700 1800
rect 550 1760 575 1795
rect 675 1760 700 1795
rect 550 1740 700 1760
rect 550 1705 575 1740
rect 675 1705 700 1740
rect 550 1700 700 1705
rect 800 1795 1200 1800
rect 800 1760 825 1795
rect 925 1760 1075 1795
rect 1175 1760 1200 1795
rect 800 1740 1200 1760
rect 800 1705 825 1740
rect 925 1705 1075 1740
rect 1175 1705 1200 1740
rect 800 1700 1200 1705
rect 1300 1795 1450 1800
rect 1300 1760 1325 1795
rect 1425 1760 1450 1795
rect 1300 1740 1450 1760
rect 1300 1705 1325 1740
rect 1425 1705 1450 1740
rect 1300 1700 1450 1705
rect 1550 1795 1700 1800
rect 1550 1760 1575 1795
rect 1675 1760 1700 1795
rect 1550 1740 1700 1760
rect 1550 1705 1575 1740
rect 1675 1705 1700 1740
rect 1550 1700 1700 1705
rect 1800 1795 2000 1800
rect 1800 1760 1825 1795
rect 1925 1760 2000 1795
rect 1800 1740 2000 1760
rect 1800 1705 1825 1740
rect 1925 1705 2000 1740
rect 1800 1700 2000 1705
rect 0 1690 60 1700
rect 190 1690 310 1700
rect 440 1690 560 1700
rect 690 1690 810 1700
rect 940 1690 1060 1700
rect 1190 1690 1310 1700
rect 1440 1690 1560 1700
rect 1690 1690 1810 1700
rect 1940 1690 2000 1700
rect 0 1675 50 1690
rect 0 1575 10 1675
rect 45 1575 50 1675
rect 0 1560 50 1575
rect 200 1675 300 1690
rect 200 1575 205 1675
rect 240 1575 260 1675
rect 295 1575 300 1675
rect 200 1560 300 1575
rect 450 1675 550 1690
rect 450 1575 455 1675
rect 490 1575 510 1675
rect 545 1575 550 1675
rect 450 1560 550 1575
rect 700 1675 800 1690
rect 700 1575 705 1675
rect 740 1575 760 1675
rect 795 1575 800 1675
rect 700 1560 800 1575
rect 950 1675 1050 1690
rect 950 1575 955 1675
rect 990 1575 1010 1675
rect 1045 1575 1050 1675
rect 950 1560 1050 1575
rect 1200 1675 1300 1690
rect 1200 1575 1205 1675
rect 1240 1575 1260 1675
rect 1295 1575 1300 1675
rect 1200 1560 1300 1575
rect 1450 1675 1550 1690
rect 1450 1575 1455 1675
rect 1490 1575 1510 1675
rect 1545 1575 1550 1675
rect 1450 1560 1550 1575
rect 1700 1675 1800 1690
rect 1700 1575 1705 1675
rect 1740 1575 1760 1675
rect 1795 1575 1800 1675
rect 1700 1560 1800 1575
rect 1950 1675 2000 1690
rect 1950 1575 1955 1675
rect 1990 1575 2000 1675
rect 1950 1560 2000 1575
rect 0 1550 60 1560
rect 190 1550 310 1560
rect 440 1550 560 1560
rect 690 1550 810 1560
rect 940 1550 1060 1560
rect 1190 1550 1310 1560
rect 1440 1550 1560 1560
rect 1690 1550 1810 1560
rect 1940 1550 2000 1560
rect 0 1545 200 1550
rect 0 1510 75 1545
rect 175 1510 200 1545
rect 0 1490 200 1510
rect 0 1455 75 1490
rect 175 1455 200 1490
rect 0 1450 200 1455
rect 300 1545 450 1550
rect 300 1510 325 1545
rect 425 1510 450 1545
rect 300 1490 450 1510
rect 300 1455 325 1490
rect 425 1455 450 1490
rect 300 1450 450 1455
rect 550 1545 700 1550
rect 550 1510 575 1545
rect 675 1510 700 1545
rect 550 1490 700 1510
rect 550 1455 575 1490
rect 675 1455 700 1490
rect 550 1450 700 1455
rect 800 1545 950 1550
rect 800 1510 825 1545
rect 925 1510 950 1545
rect 800 1490 950 1510
rect 800 1455 825 1490
rect 925 1455 950 1490
rect 800 1450 950 1455
rect 1050 1545 1200 1550
rect 1050 1510 1075 1545
rect 1175 1510 1200 1545
rect 1050 1490 1200 1510
rect 1050 1455 1075 1490
rect 1175 1455 1200 1490
rect 1050 1450 1200 1455
rect 1300 1545 1450 1550
rect 1300 1510 1325 1545
rect 1425 1510 1450 1545
rect 1300 1490 1450 1510
rect 1300 1455 1325 1490
rect 1425 1455 1450 1490
rect 1300 1450 1450 1455
rect 1550 1545 1700 1550
rect 1550 1510 1575 1545
rect 1675 1510 1700 1545
rect 1550 1490 1700 1510
rect 1550 1455 1575 1490
rect 1675 1455 1700 1490
rect 1550 1450 1700 1455
rect 1800 1545 2000 1550
rect 1800 1510 1825 1545
rect 1925 1510 2000 1545
rect 1800 1490 2000 1510
rect 1800 1455 1825 1490
rect 1925 1455 2000 1490
rect 1800 1450 2000 1455
rect 0 1440 60 1450
rect 190 1440 310 1450
rect 440 1440 560 1450
rect 690 1440 810 1450
rect 940 1440 1060 1450
rect 1190 1440 1310 1450
rect 1440 1440 1560 1450
rect 1690 1440 1810 1450
rect 1940 1440 2000 1450
rect 0 1425 50 1440
rect 0 1325 10 1425
rect 45 1325 50 1425
rect 0 1310 50 1325
rect 200 1425 300 1440
rect 200 1325 205 1425
rect 240 1325 260 1425
rect 295 1325 300 1425
rect 200 1310 300 1325
rect 450 1425 550 1440
rect 450 1325 455 1425
rect 490 1325 510 1425
rect 545 1325 550 1425
rect 450 1310 550 1325
rect 700 1425 800 1440
rect 700 1325 705 1425
rect 740 1325 760 1425
rect 795 1325 800 1425
rect 700 1310 800 1325
rect 950 1425 1050 1440
rect 950 1325 955 1425
rect 990 1325 1010 1425
rect 1045 1325 1050 1425
rect 950 1310 1050 1325
rect 1200 1425 1300 1440
rect 1200 1325 1205 1425
rect 1240 1325 1260 1425
rect 1295 1325 1300 1425
rect 1200 1310 1300 1325
rect 1450 1425 1550 1440
rect 1450 1325 1455 1425
rect 1490 1325 1510 1425
rect 1545 1325 1550 1425
rect 1450 1310 1550 1325
rect 1700 1425 1800 1440
rect 1700 1325 1705 1425
rect 1740 1325 1760 1425
rect 1795 1325 1800 1425
rect 1700 1310 1800 1325
rect 1950 1425 2000 1440
rect 1950 1325 1955 1425
rect 1990 1325 2000 1425
rect 1950 1310 2000 1325
rect 0 1300 60 1310
rect 190 1300 310 1310
rect 440 1300 560 1310
rect 690 1300 810 1310
rect 940 1300 1060 1310
rect 1190 1300 1310 1310
rect 1440 1300 1560 1310
rect 1690 1300 1810 1310
rect 1940 1300 2000 1310
rect 0 1295 200 1300
rect 0 1260 75 1295
rect 175 1260 200 1295
rect 0 1240 200 1260
rect 0 1205 75 1240
rect 175 1205 200 1240
rect 0 1200 200 1205
rect 300 1295 450 1300
rect 300 1260 325 1295
rect 425 1260 450 1295
rect 300 1240 450 1260
rect 300 1205 325 1240
rect 425 1205 450 1240
rect 300 1200 450 1205
rect 550 1295 700 1300
rect 550 1260 575 1295
rect 675 1260 700 1295
rect 550 1240 700 1260
rect 550 1205 575 1240
rect 675 1205 700 1240
rect 550 1200 700 1205
rect 800 1295 1200 1300
rect 800 1260 825 1295
rect 925 1260 1075 1295
rect 1175 1260 1200 1295
rect 800 1240 1200 1260
rect 800 1205 825 1240
rect 925 1205 1075 1240
rect 1175 1205 1200 1240
rect 800 1200 1200 1205
rect 1300 1295 1450 1300
rect 1300 1260 1325 1295
rect 1425 1260 1450 1295
rect 1300 1240 1450 1260
rect 1300 1205 1325 1240
rect 1425 1205 1450 1240
rect 1300 1200 1450 1205
rect 1550 1295 1700 1300
rect 1550 1260 1575 1295
rect 1675 1260 1700 1295
rect 1550 1240 1700 1260
rect 1550 1205 1575 1240
rect 1675 1205 1700 1240
rect 1550 1200 1700 1205
rect 1800 1295 2000 1300
rect 1800 1260 1825 1295
rect 1925 1260 2000 1295
rect 1800 1240 2000 1260
rect 1800 1205 1825 1240
rect 1925 1205 2000 1240
rect 1800 1200 2000 1205
rect 0 1190 60 1200
rect 190 1190 310 1200
rect 440 1190 560 1200
rect 690 1190 810 1200
rect 940 1190 1060 1200
rect 1190 1190 1310 1200
rect 1440 1190 1560 1200
rect 1690 1190 1810 1200
rect 1940 1190 2000 1200
rect 0 1175 50 1190
rect 0 1075 10 1175
rect 45 1075 50 1175
rect 0 1060 50 1075
rect 200 1175 300 1190
rect 200 1075 205 1175
rect 240 1075 260 1175
rect 295 1075 300 1175
rect 200 1060 300 1075
rect 450 1175 550 1190
rect 450 1075 455 1175
rect 490 1075 510 1175
rect 545 1075 550 1175
rect 450 1060 550 1075
rect 700 1175 800 1190
rect 700 1075 705 1175
rect 740 1075 760 1175
rect 795 1075 800 1175
rect 700 1060 800 1075
rect 950 1175 1050 1190
rect 950 1075 955 1175
rect 990 1075 1010 1175
rect 1045 1075 1050 1175
rect 950 1060 1050 1075
rect 1200 1175 1300 1190
rect 1200 1075 1205 1175
rect 1240 1075 1260 1175
rect 1295 1075 1300 1175
rect 1200 1060 1300 1075
rect 1450 1175 1550 1190
rect 1450 1075 1455 1175
rect 1490 1075 1510 1175
rect 1545 1075 1550 1175
rect 1450 1060 1550 1075
rect 1700 1175 1800 1190
rect 1700 1075 1705 1175
rect 1740 1075 1760 1175
rect 1795 1075 1800 1175
rect 1700 1060 1800 1075
rect 1950 1175 2000 1190
rect 1950 1075 1955 1175
rect 1990 1075 2000 1175
rect 1950 1060 2000 1075
rect 0 1050 60 1060
rect 190 1050 310 1060
rect 440 1050 560 1060
rect 690 1050 810 1060
rect 940 1050 1060 1060
rect 1190 1050 1310 1060
rect 1440 1050 1560 1060
rect 1690 1050 1810 1060
rect 1940 1050 2000 1060
rect 0 1045 450 1050
rect 0 1010 75 1045
rect 175 1010 325 1045
rect 425 1010 450 1045
rect 0 990 450 1010
rect 0 955 75 990
rect 175 955 325 990
rect 425 955 450 990
rect 0 950 450 955
rect 550 1045 1450 1050
rect 550 1010 575 1045
rect 675 1010 825 1045
rect 925 1010 1075 1045
rect 1175 1010 1325 1045
rect 1425 1010 1450 1045
rect 550 990 1450 1010
rect 550 955 575 990
rect 675 955 825 990
rect 925 955 1075 990
rect 1175 955 1325 990
rect 1425 955 1450 990
rect 550 950 1450 955
rect 1550 1045 2000 1050
rect 1550 1010 1575 1045
rect 1675 1010 1825 1045
rect 1925 1010 2000 1045
rect 1550 990 2000 1010
rect 1550 955 1575 990
rect 1675 955 1825 990
rect 1925 955 2000 990
rect 1550 950 2000 955
rect 0 940 60 950
rect 190 940 310 950
rect 440 940 560 950
rect 690 940 810 950
rect 940 940 1060 950
rect 1190 940 1310 950
rect 1440 940 1560 950
rect 1690 940 1810 950
rect 1940 940 2000 950
rect 0 925 50 940
rect 0 825 10 925
rect 45 825 50 925
rect 0 810 50 825
rect 200 925 300 940
rect 200 825 205 925
rect 240 825 260 925
rect 295 825 300 925
rect 200 810 300 825
rect 450 925 550 940
rect 450 825 455 925
rect 490 825 510 925
rect 545 825 550 925
rect 450 810 550 825
rect 700 925 800 940
rect 700 825 705 925
rect 740 825 760 925
rect 795 825 800 925
rect 700 810 800 825
rect 950 925 1050 940
rect 950 825 955 925
rect 990 825 1010 925
rect 1045 825 1050 925
rect 950 810 1050 825
rect 1200 925 1300 940
rect 1200 825 1205 925
rect 1240 825 1260 925
rect 1295 825 1300 925
rect 1200 810 1300 825
rect 1450 925 1550 940
rect 1450 825 1455 925
rect 1490 825 1510 925
rect 1545 825 1550 925
rect 1450 810 1550 825
rect 1700 925 1800 940
rect 1700 825 1705 925
rect 1740 825 1760 925
rect 1795 825 1800 925
rect 1700 810 1800 825
rect 1950 925 2000 940
rect 1950 825 1955 925
rect 1990 825 2000 925
rect 1950 810 2000 825
rect 0 800 60 810
rect 190 800 310 810
rect 440 800 560 810
rect 690 800 810 810
rect 940 800 1060 810
rect 1190 800 1310 810
rect 1440 800 1560 810
rect 1690 800 1810 810
rect 1940 800 2000 810
rect 0 795 200 800
rect 0 760 75 795
rect 175 760 200 795
rect 0 740 200 760
rect 0 705 75 740
rect 175 705 200 740
rect 0 700 200 705
rect 300 795 450 800
rect 300 760 325 795
rect 425 760 450 795
rect 300 740 450 760
rect 300 705 325 740
rect 425 705 450 740
rect 300 700 450 705
rect 550 795 700 800
rect 550 760 575 795
rect 675 760 700 795
rect 550 740 700 760
rect 550 705 575 740
rect 675 705 700 740
rect 550 700 700 705
rect 800 795 1200 800
rect 800 760 825 795
rect 925 760 1075 795
rect 1175 760 1200 795
rect 800 740 1200 760
rect 800 705 825 740
rect 925 705 1075 740
rect 1175 705 1200 740
rect 800 700 1200 705
rect 1300 795 1450 800
rect 1300 760 1325 795
rect 1425 760 1450 795
rect 1300 740 1450 760
rect 1300 705 1325 740
rect 1425 705 1450 740
rect 1300 700 1450 705
rect 1550 795 1700 800
rect 1550 760 1575 795
rect 1675 760 1700 795
rect 1550 740 1700 760
rect 1550 705 1575 740
rect 1675 705 1700 740
rect 1550 700 1700 705
rect 1800 795 2000 800
rect 1800 760 1825 795
rect 1925 760 2000 795
rect 1800 740 2000 760
rect 1800 705 1825 740
rect 1925 705 2000 740
rect 1800 700 2000 705
rect 0 690 60 700
rect 190 690 310 700
rect 440 690 560 700
rect 690 690 810 700
rect 940 690 1060 700
rect 1190 690 1310 700
rect 1440 690 1560 700
rect 1690 690 1810 700
rect 1940 690 2000 700
rect 0 675 50 690
rect 0 575 10 675
rect 45 575 50 675
rect 0 560 50 575
rect 200 675 300 690
rect 200 575 205 675
rect 240 575 260 675
rect 295 575 300 675
rect 200 560 300 575
rect 450 675 550 690
rect 450 575 455 675
rect 490 575 510 675
rect 545 575 550 675
rect 450 560 550 575
rect 700 675 800 690
rect 700 575 705 675
rect 740 575 760 675
rect 795 575 800 675
rect 700 560 800 575
rect 950 675 1050 690
rect 950 575 955 675
rect 990 575 1010 675
rect 1045 575 1050 675
rect 950 560 1050 575
rect 1200 675 1300 690
rect 1200 575 1205 675
rect 1240 575 1260 675
rect 1295 575 1300 675
rect 1200 560 1300 575
rect 1450 675 1550 690
rect 1450 575 1455 675
rect 1490 575 1510 675
rect 1545 575 1550 675
rect 1450 560 1550 575
rect 1700 675 1800 690
rect 1700 575 1705 675
rect 1740 575 1760 675
rect 1795 575 1800 675
rect 1700 560 1800 575
rect 1950 675 2000 690
rect 1950 575 1955 675
rect 1990 575 2000 675
rect 1950 560 2000 575
rect 0 550 60 560
rect 190 550 310 560
rect 440 550 560 560
rect 690 550 810 560
rect 940 550 1060 560
rect 1190 550 1310 560
rect 1440 550 1560 560
rect 1690 550 1810 560
rect 1940 550 2000 560
rect 0 545 200 550
rect 0 510 75 545
rect 175 510 200 545
rect 0 490 200 510
rect 0 455 75 490
rect 175 455 200 490
rect 0 450 200 455
rect 300 545 450 550
rect 300 510 325 545
rect 425 510 450 545
rect 300 490 450 510
rect 300 455 325 490
rect 425 455 450 490
rect 300 450 450 455
rect 550 545 700 550
rect 550 510 575 545
rect 675 510 700 545
rect 550 490 700 510
rect 550 455 575 490
rect 675 455 700 490
rect 550 450 700 455
rect 800 545 950 550
rect 800 510 825 545
rect 925 510 950 545
rect 800 490 950 510
rect 800 455 825 490
rect 925 455 950 490
rect 800 450 950 455
rect 1050 545 1200 550
rect 1050 510 1075 545
rect 1175 510 1200 545
rect 1050 490 1200 510
rect 1050 455 1075 490
rect 1175 455 1200 490
rect 1050 450 1200 455
rect 1300 545 1450 550
rect 1300 510 1325 545
rect 1425 510 1450 545
rect 1300 490 1450 510
rect 1300 455 1325 490
rect 1425 455 1450 490
rect 1300 450 1450 455
rect 1550 545 1700 550
rect 1550 510 1575 545
rect 1675 510 1700 545
rect 1550 490 1700 510
rect 1550 455 1575 490
rect 1675 455 1700 490
rect 1550 450 1700 455
rect 1800 545 2000 550
rect 1800 510 1825 545
rect 1925 510 2000 545
rect 1800 490 2000 510
rect 1800 455 1825 490
rect 1925 455 2000 490
rect 1800 450 2000 455
rect 0 440 60 450
rect 190 440 310 450
rect 440 440 560 450
rect 690 440 810 450
rect 940 440 1060 450
rect 1190 440 1310 450
rect 1440 440 1560 450
rect 1690 440 1810 450
rect 1940 440 2000 450
rect 0 425 50 440
rect 0 325 10 425
rect 45 325 50 425
rect 0 310 50 325
rect 200 425 300 440
rect 200 325 205 425
rect 240 325 260 425
rect 295 325 300 425
rect 200 310 300 325
rect 450 425 550 440
rect 450 325 455 425
rect 490 325 510 425
rect 545 325 550 425
rect 450 310 550 325
rect 700 425 800 440
rect 700 325 705 425
rect 740 325 760 425
rect 795 325 800 425
rect 700 310 800 325
rect 950 425 1050 440
rect 950 325 955 425
rect 990 325 1010 425
rect 1045 325 1050 425
rect 950 310 1050 325
rect 1200 425 1300 440
rect 1200 325 1205 425
rect 1240 325 1260 425
rect 1295 325 1300 425
rect 1200 310 1300 325
rect 1450 425 1550 440
rect 1450 325 1455 425
rect 1490 325 1510 425
rect 1545 325 1550 425
rect 1450 310 1550 325
rect 1700 425 1800 440
rect 1700 325 1705 425
rect 1740 325 1760 425
rect 1795 325 1800 425
rect 1700 310 1800 325
rect 1950 425 2000 440
rect 1950 325 1955 425
rect 1990 325 2000 425
rect 1950 310 2000 325
rect 0 300 60 310
rect 190 300 310 310
rect 440 300 560 310
rect 690 300 810 310
rect 940 300 1060 310
rect 1190 300 1310 310
rect 1440 300 1560 310
rect 1690 300 1810 310
rect 1940 300 2000 310
rect 0 295 200 300
rect 0 260 75 295
rect 175 260 200 295
rect 0 240 200 260
rect 0 205 75 240
rect 175 205 200 240
rect 0 200 200 205
rect 300 295 450 300
rect 300 260 325 295
rect 425 260 450 295
rect 300 240 450 260
rect 300 205 325 240
rect 425 205 450 240
rect 300 200 450 205
rect 550 295 700 300
rect 550 260 575 295
rect 675 260 700 295
rect 550 240 700 260
rect 550 205 575 240
rect 675 205 700 240
rect 550 200 700 205
rect 800 295 1200 300
rect 800 260 825 295
rect 925 260 1075 295
rect 1175 260 1200 295
rect 800 240 1200 260
rect 800 205 825 240
rect 925 205 1075 240
rect 1175 205 1200 240
rect 800 200 1200 205
rect 1300 295 1450 300
rect 1300 260 1325 295
rect 1425 260 1450 295
rect 1300 240 1450 260
rect 1300 205 1325 240
rect 1425 205 1450 240
rect 1300 200 1450 205
rect 1550 295 1700 300
rect 1550 260 1575 295
rect 1675 260 1700 295
rect 1550 240 1700 260
rect 1550 205 1575 240
rect 1675 205 1700 240
rect 1550 200 1700 205
rect 1800 295 2000 300
rect 1800 260 1825 295
rect 1925 260 2000 295
rect 1800 240 2000 260
rect 1800 205 1825 240
rect 1925 205 2000 240
rect 1800 200 2000 205
rect 0 190 60 200
rect 190 190 310 200
rect 440 190 560 200
rect 690 190 810 200
rect 940 190 1060 200
rect 1190 190 1310 200
rect 1440 190 1560 200
rect 1690 190 1810 200
rect 1940 190 2000 200
rect 0 175 50 190
rect 0 75 10 175
rect 45 75 50 175
rect 0 60 50 75
rect 200 175 300 190
rect 200 75 205 175
rect 240 75 260 175
rect 295 75 300 175
rect 200 60 300 75
rect 450 175 550 190
rect 450 75 455 175
rect 490 75 510 175
rect 545 75 550 175
rect 450 60 550 75
rect 700 175 800 190
rect 700 75 705 175
rect 740 75 760 175
rect 795 75 800 175
rect 700 60 800 75
rect 950 175 1050 190
rect 950 75 955 175
rect 990 75 1010 175
rect 1045 75 1050 175
rect 950 60 1050 75
rect 1200 175 1300 190
rect 1200 75 1205 175
rect 1240 75 1260 175
rect 1295 75 1300 175
rect 1200 60 1300 75
rect 1450 175 1550 190
rect 1450 75 1455 175
rect 1490 75 1510 175
rect 1545 75 1550 175
rect 1450 60 1550 75
rect 1700 175 1800 190
rect 1700 75 1705 175
rect 1740 75 1760 175
rect 1795 75 1800 175
rect 1700 60 1800 75
rect 1950 175 2000 190
rect 1950 75 1955 175
rect 1990 75 2000 175
rect 1950 60 2000 75
rect 0 50 60 60
rect 190 50 310 60
rect 440 50 560 60
rect 690 50 810 60
rect 940 50 1060 60
rect 1190 50 1310 60
rect 1440 50 1560 60
rect 1690 50 1810 60
rect 1940 50 2000 60
rect 0 45 2000 50
rect 0 10 75 45
rect 175 10 325 45
rect 425 10 575 45
rect 675 10 825 45
rect 925 10 1075 45
rect 1175 10 1325 45
rect 1425 10 1575 45
rect 1675 10 1825 45
rect 1925 10 2000 45
rect 0 0 2000 10
<< via3 >>
rect 200 1700 300 1800
rect 450 1700 550 1800
rect 700 1700 800 1800
rect 1200 1700 1300 1800
rect 1450 1700 1550 1800
rect 1700 1700 1800 1800
rect 200 1450 300 1550
rect 450 1450 550 1550
rect 700 1450 800 1550
rect 950 1450 1050 1550
rect 1200 1450 1300 1550
rect 1450 1450 1550 1550
rect 1700 1450 1800 1550
rect 200 1200 300 1300
rect 450 1200 550 1300
rect 700 1200 800 1300
rect 1200 1200 1300 1300
rect 1450 1200 1550 1300
rect 1700 1200 1800 1300
rect 450 950 550 1050
rect 1450 950 1550 1050
rect 200 700 300 800
rect 450 700 550 800
rect 700 700 800 800
rect 1200 700 1300 800
rect 1450 700 1550 800
rect 1700 700 1800 800
rect 200 450 300 550
rect 450 450 550 550
rect 700 450 800 550
rect 950 450 1050 550
rect 1200 450 1300 550
rect 1450 450 1550 550
rect 1700 450 1800 550
rect 200 200 300 300
rect 450 200 550 300
rect 700 200 800 300
rect 1200 200 1300 300
rect 1450 200 1550 300
rect 1700 200 1800 300
<< metal4 >>
rect 260 1820 740 2000
rect 1260 1820 1740 2000
rect 180 1800 820 1820
rect 180 1740 200 1800
rect 0 1700 200 1740
rect 300 1700 450 1800
rect 550 1700 700 1800
rect 800 1740 820 1800
rect 1180 1800 1820 1820
rect 1180 1740 1200 1800
rect 800 1700 1200 1740
rect 1300 1700 1450 1800
rect 1550 1700 1700 1800
rect 1800 1740 1820 1800
rect 1800 1700 2000 1740
rect 0 1550 2000 1700
rect 0 1450 200 1550
rect 300 1450 450 1550
rect 550 1450 700 1550
rect 800 1450 950 1550
rect 1050 1450 1200 1550
rect 1300 1450 1450 1550
rect 1550 1450 1700 1550
rect 1800 1450 2000 1550
rect 0 1300 2000 1450
rect 0 1260 200 1300
rect 180 1200 200 1260
rect 300 1200 450 1300
rect 550 1200 700 1300
rect 800 1260 1200 1300
rect 800 1200 820 1260
rect 180 1180 820 1200
rect 1180 1200 1200 1260
rect 1300 1200 1450 1300
rect 1550 1200 1700 1300
rect 1800 1260 2000 1300
rect 1800 1200 1820 1260
rect 1180 1180 1820 1200
rect 260 1050 740 1180
rect 260 950 450 1050
rect 550 950 740 1050
rect 260 820 740 950
rect 1260 1050 1740 1180
rect 1260 950 1450 1050
rect 1550 950 1740 1050
rect 1260 820 1740 950
rect 180 800 820 820
rect 180 740 200 800
rect 0 700 200 740
rect 300 700 450 800
rect 550 700 700 800
rect 800 740 820 800
rect 1180 800 1820 820
rect 1180 740 1200 800
rect 800 700 1200 740
rect 1300 700 1450 800
rect 1550 700 1700 800
rect 1800 740 1820 800
rect 1800 700 2000 740
rect 0 550 2000 700
rect 0 450 200 550
rect 300 450 450 550
rect 550 450 700 550
rect 800 450 950 550
rect 1050 450 1200 550
rect 1300 450 1450 550
rect 1550 450 1700 550
rect 1800 450 2000 550
rect 0 300 2000 450
rect 0 260 200 300
rect 180 200 200 260
rect 300 200 450 300
rect 550 200 700 300
rect 800 260 1200 300
rect 800 200 820 260
rect 180 180 820 200
rect 1180 200 1200 260
rect 1300 200 1450 300
rect 1550 200 1700 300
rect 1800 260 2000 300
rect 1800 200 1820 260
rect 1180 180 1820 200
rect 260 0 740 180
rect 1260 0 1740 180
<< end >>
