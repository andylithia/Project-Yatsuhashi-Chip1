magic
tech sky130B
magscale 1 2
timestamp 1662473609
<< nwell >>
rect 1060 -80 3880 1180
<< nsubdiff >>
rect 1100 1080 1180 1120
rect 1100 1040 1120 1080
rect 1160 1040 1180 1080
rect 1100 1000 1180 1040
rect 1100 960 1120 1000
rect 1160 960 1180 1000
rect 1100 920 1180 960
rect 1100 880 1120 920
rect 1160 880 1180 920
rect 1100 840 1180 880
rect 1100 800 1120 840
rect 1160 800 1180 840
rect 1100 760 1180 800
rect 1100 720 1120 760
rect 1160 720 1180 760
rect 1100 680 1180 720
rect 1100 640 1120 680
rect 1160 640 1180 680
rect 1100 600 1180 640
rect 1100 560 1120 600
rect 1160 560 1180 600
rect 1100 520 1180 560
rect 1100 480 1120 520
rect 1160 480 1180 520
rect 1100 440 1180 480
rect 1100 400 1120 440
rect 1160 400 1180 440
rect 1100 360 1180 400
rect 1100 320 1120 360
rect 1160 320 1180 360
rect 1100 280 1180 320
rect 1100 240 1120 280
rect 1160 240 1180 280
rect 1100 200 1180 240
rect 1100 160 1120 200
rect 1160 160 1180 200
rect 1100 60 1180 160
rect 3760 1080 3840 1120
rect 3760 1040 3780 1080
rect 3820 1040 3840 1080
rect 3760 1000 3840 1040
rect 3760 960 3780 1000
rect 3820 960 3840 1000
rect 3760 920 3840 960
rect 3760 880 3780 920
rect 3820 880 3840 920
rect 3760 840 3840 880
rect 3760 800 3780 840
rect 3820 800 3840 840
rect 3760 760 3840 800
rect 3760 720 3780 760
rect 3820 720 3840 760
rect 3760 680 3840 720
rect 3760 640 3780 680
rect 3820 640 3840 680
rect 3760 600 3840 640
rect 3760 560 3780 600
rect 3820 560 3840 600
rect 3760 520 3840 560
rect 3760 480 3780 520
rect 3820 480 3840 520
rect 3760 440 3840 480
rect 3760 400 3780 440
rect 3820 400 3840 440
rect 3760 360 3840 400
rect 3760 320 3780 360
rect 3820 320 3840 360
rect 3760 280 3840 320
rect 3760 240 3780 280
rect 3820 240 3840 280
rect 3760 200 3840 240
rect 3760 160 3780 200
rect 3820 160 3840 200
rect 3760 60 3840 160
rect 1100 40 3840 60
rect 1100 0 1300 40
rect 1340 0 1380 40
rect 1420 0 1460 40
rect 1500 0 1540 40
rect 1580 0 1620 40
rect 1660 0 1700 40
rect 1740 0 1780 40
rect 1820 0 1860 40
rect 1900 0 1940 40
rect 1980 0 2020 40
rect 2060 0 2100 40
rect 2140 0 2180 40
rect 2220 0 2260 40
rect 2300 0 2340 40
rect 2380 0 2420 40
rect 2460 0 2500 40
rect 2540 0 2580 40
rect 2620 0 2660 40
rect 2700 0 2740 40
rect 2780 0 2820 40
rect 2860 0 2900 40
rect 2940 0 2980 40
rect 3020 0 3060 40
rect 3100 0 3140 40
rect 3180 0 3220 40
rect 3260 0 3300 40
rect 3340 0 3380 40
rect 3420 0 3460 40
rect 3500 0 3540 40
rect 3580 0 3620 40
rect 3660 0 3840 40
rect 1100 -20 3840 0
<< nsubdiffcont >>
rect 1120 1040 1160 1080
rect 1120 960 1160 1000
rect 1120 880 1160 920
rect 1120 800 1160 840
rect 1120 720 1160 760
rect 1120 640 1160 680
rect 1120 560 1160 600
rect 1120 480 1160 520
rect 1120 400 1160 440
rect 1120 320 1160 360
rect 1120 240 1160 280
rect 1120 160 1160 200
rect 3780 1040 3820 1080
rect 3780 960 3820 1000
rect 3780 880 3820 920
rect 3780 800 3820 840
rect 3780 720 3820 760
rect 3780 640 3820 680
rect 3780 560 3820 600
rect 3780 480 3820 520
rect 3780 400 3820 440
rect 3780 320 3820 360
rect 3780 240 3820 280
rect 3780 160 3820 200
rect 1300 0 1340 40
rect 1380 0 1420 40
rect 1460 0 1500 40
rect 1540 0 1580 40
rect 1620 0 1660 40
rect 1700 0 1740 40
rect 1780 0 1820 40
rect 1860 0 1900 40
rect 1940 0 1980 40
rect 2020 0 2060 40
rect 2100 0 2140 40
rect 2180 0 2220 40
rect 2260 0 2300 40
rect 2340 0 2380 40
rect 2420 0 2460 40
rect 2500 0 2540 40
rect 2580 0 2620 40
rect 2660 0 2700 40
rect 2740 0 2780 40
rect 2820 0 2860 40
rect 2900 0 2940 40
rect 2980 0 3020 40
rect 3060 0 3100 40
rect 3140 0 3180 40
rect 3220 0 3260 40
rect 3300 0 3340 40
rect 3380 0 3420 40
rect 3460 0 3500 40
rect 3540 0 3580 40
rect 3620 0 3660 40
<< locali >>
rect 1120 1100 1200 1120
rect 1120 1080 1140 1100
rect 1120 1000 1140 1040
rect 1120 920 1140 960
rect 1120 840 1140 880
rect 1120 760 1140 800
rect 1120 680 1140 720
rect 1120 600 1140 640
rect 1120 520 1140 560
rect 1120 440 1140 480
rect 1120 360 1140 400
rect 1120 280 1140 320
rect 1120 200 1140 240
rect 1180 160 1200 1100
rect 1120 140 1200 160
rect 3740 1100 3820 1120
rect 3740 160 3760 1100
rect 3800 1080 3820 1100
rect 3800 1000 3820 1040
rect 3800 920 3820 960
rect 3800 840 3820 880
rect 3800 760 3820 800
rect 3800 680 3820 720
rect 3800 600 3820 640
rect 3800 520 3820 560
rect 3800 440 3820 480
rect 3800 360 3820 400
rect 3800 280 3820 320
rect 3800 200 3820 240
rect 3740 140 3820 160
rect 1240 40 3700 60
rect 1240 0 1260 40
rect 3680 0 3700 40
rect 1240 -20 3700 0
<< viali >>
rect 1140 1080 1180 1100
rect 1140 1040 1160 1080
rect 1160 1040 1180 1080
rect 1140 1000 1180 1040
rect 1140 960 1160 1000
rect 1160 960 1180 1000
rect 1140 920 1180 960
rect 1140 880 1160 920
rect 1160 880 1180 920
rect 1140 840 1180 880
rect 1140 800 1160 840
rect 1160 800 1180 840
rect 1140 760 1180 800
rect 1140 720 1160 760
rect 1160 720 1180 760
rect 1140 680 1180 720
rect 1140 640 1160 680
rect 1160 640 1180 680
rect 1140 600 1180 640
rect 1140 560 1160 600
rect 1160 560 1180 600
rect 1140 520 1180 560
rect 1140 480 1160 520
rect 1160 480 1180 520
rect 1140 440 1180 480
rect 1140 400 1160 440
rect 1160 400 1180 440
rect 1140 360 1180 400
rect 1140 320 1160 360
rect 1160 320 1180 360
rect 1140 280 1180 320
rect 1140 240 1160 280
rect 1160 240 1180 280
rect 1140 200 1180 240
rect 1140 160 1160 200
rect 1160 160 1180 200
rect 3760 1080 3800 1100
rect 3760 1040 3780 1080
rect 3780 1040 3800 1080
rect 3760 1000 3800 1040
rect 3760 960 3780 1000
rect 3780 960 3800 1000
rect 3760 920 3800 960
rect 3760 880 3780 920
rect 3780 880 3800 920
rect 3760 840 3800 880
rect 3760 800 3780 840
rect 3780 800 3800 840
rect 3760 760 3800 800
rect 3760 720 3780 760
rect 3780 720 3800 760
rect 3760 680 3800 720
rect 3760 640 3780 680
rect 3780 640 3800 680
rect 3760 600 3800 640
rect 3760 560 3780 600
rect 3780 560 3800 600
rect 3760 520 3800 560
rect 3760 480 3780 520
rect 3780 480 3800 520
rect 3760 440 3800 480
rect 3760 400 3780 440
rect 3780 400 3800 440
rect 3760 360 3800 400
rect 3760 320 3780 360
rect 3780 320 3800 360
rect 3760 280 3800 320
rect 3760 240 3780 280
rect 3780 240 3800 280
rect 3760 200 3800 240
rect 3760 160 3780 200
rect 3780 160 3800 200
rect 1260 0 1300 40
rect 1300 0 1340 40
rect 1340 0 1380 40
rect 1380 0 1420 40
rect 1420 0 1460 40
rect 1460 0 1500 40
rect 1500 0 1540 40
rect 1540 0 1580 40
rect 1580 0 1620 40
rect 1620 0 1660 40
rect 1660 0 1700 40
rect 1700 0 1740 40
rect 1740 0 1780 40
rect 1780 0 1820 40
rect 1820 0 1860 40
rect 1860 0 1900 40
rect 1900 0 1940 40
rect 1940 0 1980 40
rect 1980 0 2020 40
rect 2020 0 2060 40
rect 2060 0 2100 40
rect 2100 0 2140 40
rect 2140 0 2180 40
rect 2180 0 2220 40
rect 2220 0 2260 40
rect 2260 0 2300 40
rect 2300 0 2340 40
rect 2340 0 2380 40
rect 2380 0 2420 40
rect 2420 0 2460 40
rect 2460 0 2500 40
rect 2500 0 2540 40
rect 2540 0 2580 40
rect 2580 0 2620 40
rect 2620 0 2660 40
rect 2660 0 2700 40
rect 2700 0 2740 40
rect 2740 0 2780 40
rect 2780 0 2820 40
rect 2820 0 2860 40
rect 2860 0 2900 40
rect 2900 0 2940 40
rect 2940 0 2980 40
rect 2980 0 3020 40
rect 3020 0 3060 40
rect 3060 0 3100 40
rect 3100 0 3140 40
rect 3140 0 3180 40
rect 3180 0 3220 40
rect 3220 0 3260 40
rect 3260 0 3300 40
rect 3300 0 3340 40
rect 3340 0 3380 40
rect 3380 0 3420 40
rect 3420 0 3460 40
rect 3460 0 3500 40
rect 3500 0 3540 40
rect 3540 0 3580 40
rect 3580 0 3620 40
rect 3620 0 3660 40
rect 3660 0 3680 40
<< metal1 >>
rect 1289 1170 3634 1386
rect 1120 1100 1280 1120
rect 1120 160 1140 1100
rect 1180 160 1280 1100
rect 1120 140 1280 160
rect 3660 1100 3820 1120
rect 3660 160 3760 1100
rect 3800 160 3820 1100
rect 3660 140 3820 160
rect 1240 0 1260 40
rect 3680 0 3700 40
rect 1240 -40 3700 0
rect 2380 -100 2440 -40
<< metal3 >>
rect 980 1060 3600 1120
use sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1660669191
transform 1 0 1200 0 1 97
box 0 -97 466 1135
use sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15_1
timestamp 1660669191
transform -1 0 2010 0 1 97
box 0 -97 466 1135
use sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15_2
timestamp 1660669191
transform 1 0 1888 0 1 97
box 0 -97 466 1135
use sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15_3
timestamp 1660669191
transform -1 0 2698 0 1 97
box 0 -97 466 1135
use sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15_4
timestamp 1660669191
transform 1 0 2920 0 1 97
box 0 -97 466 1135
use sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15_5
timestamp 1660669191
transform -1 0 3730 0 1 97
box 0 -97 466 1135
use sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF04W5p00L0p15_6
timestamp 1660669191
transform -1 0 3042 0 1 97
box 0 -97 466 1135
<< labels >>
rlabel metal1 1300 1320 1560 1380 1 G
rlabel metal3 980 1060 1020 1120 1 SD
rlabel metal1 2380 -100 2440 -80 1 S
<< end >>
