magic
tech sky130B
magscale 1 2
timestamp 1662238829
<< nwell >>
rect -296 -40349 296 40349
<< pmos >>
rect -100 38130 100 40130
rect -100 35894 100 37894
rect -100 33658 100 35658
rect -100 31422 100 33422
rect -100 29186 100 31186
rect -100 26950 100 28950
rect -100 24714 100 26714
rect -100 22478 100 24478
rect -100 20242 100 22242
rect -100 18006 100 20006
rect -100 15770 100 17770
rect -100 13534 100 15534
rect -100 11298 100 13298
rect -100 9062 100 11062
rect -100 6826 100 8826
rect -100 4590 100 6590
rect -100 2354 100 4354
rect -100 118 100 2118
rect -100 -2118 100 -118
rect -100 -4354 100 -2354
rect -100 -6590 100 -4590
rect -100 -8826 100 -6826
rect -100 -11062 100 -9062
rect -100 -13298 100 -11298
rect -100 -15534 100 -13534
rect -100 -17770 100 -15770
rect -100 -20006 100 -18006
rect -100 -22242 100 -20242
rect -100 -24478 100 -22478
rect -100 -26714 100 -24714
rect -100 -28950 100 -26950
rect -100 -31186 100 -29186
rect -100 -33422 100 -31422
rect -100 -35658 100 -33658
rect -100 -37894 100 -35894
rect -100 -40130 100 -38130
<< pdiff >>
rect -158 40118 -100 40130
rect -158 38142 -146 40118
rect -112 38142 -100 40118
rect -158 38130 -100 38142
rect 100 40118 158 40130
rect 100 38142 112 40118
rect 146 38142 158 40118
rect 100 38130 158 38142
rect -158 37882 -100 37894
rect -158 35906 -146 37882
rect -112 35906 -100 37882
rect -158 35894 -100 35906
rect 100 37882 158 37894
rect 100 35906 112 37882
rect 146 35906 158 37882
rect 100 35894 158 35906
rect -158 35646 -100 35658
rect -158 33670 -146 35646
rect -112 33670 -100 35646
rect -158 33658 -100 33670
rect 100 35646 158 35658
rect 100 33670 112 35646
rect 146 33670 158 35646
rect 100 33658 158 33670
rect -158 33410 -100 33422
rect -158 31434 -146 33410
rect -112 31434 -100 33410
rect -158 31422 -100 31434
rect 100 33410 158 33422
rect 100 31434 112 33410
rect 146 31434 158 33410
rect 100 31422 158 31434
rect -158 31174 -100 31186
rect -158 29198 -146 31174
rect -112 29198 -100 31174
rect -158 29186 -100 29198
rect 100 31174 158 31186
rect 100 29198 112 31174
rect 146 29198 158 31174
rect 100 29186 158 29198
rect -158 28938 -100 28950
rect -158 26962 -146 28938
rect -112 26962 -100 28938
rect -158 26950 -100 26962
rect 100 28938 158 28950
rect 100 26962 112 28938
rect 146 26962 158 28938
rect 100 26950 158 26962
rect -158 26702 -100 26714
rect -158 24726 -146 26702
rect -112 24726 -100 26702
rect -158 24714 -100 24726
rect 100 26702 158 26714
rect 100 24726 112 26702
rect 146 24726 158 26702
rect 100 24714 158 24726
rect -158 24466 -100 24478
rect -158 22490 -146 24466
rect -112 22490 -100 24466
rect -158 22478 -100 22490
rect 100 24466 158 24478
rect 100 22490 112 24466
rect 146 22490 158 24466
rect 100 22478 158 22490
rect -158 22230 -100 22242
rect -158 20254 -146 22230
rect -112 20254 -100 22230
rect -158 20242 -100 20254
rect 100 22230 158 22242
rect 100 20254 112 22230
rect 146 20254 158 22230
rect 100 20242 158 20254
rect -158 19994 -100 20006
rect -158 18018 -146 19994
rect -112 18018 -100 19994
rect -158 18006 -100 18018
rect 100 19994 158 20006
rect 100 18018 112 19994
rect 146 18018 158 19994
rect 100 18006 158 18018
rect -158 17758 -100 17770
rect -158 15782 -146 17758
rect -112 15782 -100 17758
rect -158 15770 -100 15782
rect 100 17758 158 17770
rect 100 15782 112 17758
rect 146 15782 158 17758
rect 100 15770 158 15782
rect -158 15522 -100 15534
rect -158 13546 -146 15522
rect -112 13546 -100 15522
rect -158 13534 -100 13546
rect 100 15522 158 15534
rect 100 13546 112 15522
rect 146 13546 158 15522
rect 100 13534 158 13546
rect -158 13286 -100 13298
rect -158 11310 -146 13286
rect -112 11310 -100 13286
rect -158 11298 -100 11310
rect 100 13286 158 13298
rect 100 11310 112 13286
rect 146 11310 158 13286
rect 100 11298 158 11310
rect -158 11050 -100 11062
rect -158 9074 -146 11050
rect -112 9074 -100 11050
rect -158 9062 -100 9074
rect 100 11050 158 11062
rect 100 9074 112 11050
rect 146 9074 158 11050
rect 100 9062 158 9074
rect -158 8814 -100 8826
rect -158 6838 -146 8814
rect -112 6838 -100 8814
rect -158 6826 -100 6838
rect 100 8814 158 8826
rect 100 6838 112 8814
rect 146 6838 158 8814
rect 100 6826 158 6838
rect -158 6578 -100 6590
rect -158 4602 -146 6578
rect -112 4602 -100 6578
rect -158 4590 -100 4602
rect 100 6578 158 6590
rect 100 4602 112 6578
rect 146 4602 158 6578
rect 100 4590 158 4602
rect -158 4342 -100 4354
rect -158 2366 -146 4342
rect -112 2366 -100 4342
rect -158 2354 -100 2366
rect 100 4342 158 4354
rect 100 2366 112 4342
rect 146 2366 158 4342
rect 100 2354 158 2366
rect -158 2106 -100 2118
rect -158 130 -146 2106
rect -112 130 -100 2106
rect -158 118 -100 130
rect 100 2106 158 2118
rect 100 130 112 2106
rect 146 130 158 2106
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -2106 -146 -130
rect -112 -2106 -100 -130
rect -158 -2118 -100 -2106
rect 100 -130 158 -118
rect 100 -2106 112 -130
rect 146 -2106 158 -130
rect 100 -2118 158 -2106
rect -158 -2366 -100 -2354
rect -158 -4342 -146 -2366
rect -112 -4342 -100 -2366
rect -158 -4354 -100 -4342
rect 100 -2366 158 -2354
rect 100 -4342 112 -2366
rect 146 -4342 158 -2366
rect 100 -4354 158 -4342
rect -158 -4602 -100 -4590
rect -158 -6578 -146 -4602
rect -112 -6578 -100 -4602
rect -158 -6590 -100 -6578
rect 100 -4602 158 -4590
rect 100 -6578 112 -4602
rect 146 -6578 158 -4602
rect 100 -6590 158 -6578
rect -158 -6838 -100 -6826
rect -158 -8814 -146 -6838
rect -112 -8814 -100 -6838
rect -158 -8826 -100 -8814
rect 100 -6838 158 -6826
rect 100 -8814 112 -6838
rect 146 -8814 158 -6838
rect 100 -8826 158 -8814
rect -158 -9074 -100 -9062
rect -158 -11050 -146 -9074
rect -112 -11050 -100 -9074
rect -158 -11062 -100 -11050
rect 100 -9074 158 -9062
rect 100 -11050 112 -9074
rect 146 -11050 158 -9074
rect 100 -11062 158 -11050
rect -158 -11310 -100 -11298
rect -158 -13286 -146 -11310
rect -112 -13286 -100 -11310
rect -158 -13298 -100 -13286
rect 100 -11310 158 -11298
rect 100 -13286 112 -11310
rect 146 -13286 158 -11310
rect 100 -13298 158 -13286
rect -158 -13546 -100 -13534
rect -158 -15522 -146 -13546
rect -112 -15522 -100 -13546
rect -158 -15534 -100 -15522
rect 100 -13546 158 -13534
rect 100 -15522 112 -13546
rect 146 -15522 158 -13546
rect 100 -15534 158 -15522
rect -158 -15782 -100 -15770
rect -158 -17758 -146 -15782
rect -112 -17758 -100 -15782
rect -158 -17770 -100 -17758
rect 100 -15782 158 -15770
rect 100 -17758 112 -15782
rect 146 -17758 158 -15782
rect 100 -17770 158 -17758
rect -158 -18018 -100 -18006
rect -158 -19994 -146 -18018
rect -112 -19994 -100 -18018
rect -158 -20006 -100 -19994
rect 100 -18018 158 -18006
rect 100 -19994 112 -18018
rect 146 -19994 158 -18018
rect 100 -20006 158 -19994
rect -158 -20254 -100 -20242
rect -158 -22230 -146 -20254
rect -112 -22230 -100 -20254
rect -158 -22242 -100 -22230
rect 100 -20254 158 -20242
rect 100 -22230 112 -20254
rect 146 -22230 158 -20254
rect 100 -22242 158 -22230
rect -158 -22490 -100 -22478
rect -158 -24466 -146 -22490
rect -112 -24466 -100 -22490
rect -158 -24478 -100 -24466
rect 100 -22490 158 -22478
rect 100 -24466 112 -22490
rect 146 -24466 158 -22490
rect 100 -24478 158 -24466
rect -158 -24726 -100 -24714
rect -158 -26702 -146 -24726
rect -112 -26702 -100 -24726
rect -158 -26714 -100 -26702
rect 100 -24726 158 -24714
rect 100 -26702 112 -24726
rect 146 -26702 158 -24726
rect 100 -26714 158 -26702
rect -158 -26962 -100 -26950
rect -158 -28938 -146 -26962
rect -112 -28938 -100 -26962
rect -158 -28950 -100 -28938
rect 100 -26962 158 -26950
rect 100 -28938 112 -26962
rect 146 -28938 158 -26962
rect 100 -28950 158 -28938
rect -158 -29198 -100 -29186
rect -158 -31174 -146 -29198
rect -112 -31174 -100 -29198
rect -158 -31186 -100 -31174
rect 100 -29198 158 -29186
rect 100 -31174 112 -29198
rect 146 -31174 158 -29198
rect 100 -31186 158 -31174
rect -158 -31434 -100 -31422
rect -158 -33410 -146 -31434
rect -112 -33410 -100 -31434
rect -158 -33422 -100 -33410
rect 100 -31434 158 -31422
rect 100 -33410 112 -31434
rect 146 -33410 158 -31434
rect 100 -33422 158 -33410
rect -158 -33670 -100 -33658
rect -158 -35646 -146 -33670
rect -112 -35646 -100 -33670
rect -158 -35658 -100 -35646
rect 100 -33670 158 -33658
rect 100 -35646 112 -33670
rect 146 -35646 158 -33670
rect 100 -35658 158 -35646
rect -158 -35906 -100 -35894
rect -158 -37882 -146 -35906
rect -112 -37882 -100 -35906
rect -158 -37894 -100 -37882
rect 100 -35906 158 -35894
rect 100 -37882 112 -35906
rect 146 -37882 158 -35906
rect 100 -37894 158 -37882
rect -158 -38142 -100 -38130
rect -158 -40118 -146 -38142
rect -112 -40118 -100 -38142
rect -158 -40130 -100 -40118
rect 100 -38142 158 -38130
rect 100 -40118 112 -38142
rect 146 -40118 158 -38142
rect 100 -40130 158 -40118
<< pdiffc >>
rect -146 38142 -112 40118
rect 112 38142 146 40118
rect -146 35906 -112 37882
rect 112 35906 146 37882
rect -146 33670 -112 35646
rect 112 33670 146 35646
rect -146 31434 -112 33410
rect 112 31434 146 33410
rect -146 29198 -112 31174
rect 112 29198 146 31174
rect -146 26962 -112 28938
rect 112 26962 146 28938
rect -146 24726 -112 26702
rect 112 24726 146 26702
rect -146 22490 -112 24466
rect 112 22490 146 24466
rect -146 20254 -112 22230
rect 112 20254 146 22230
rect -146 18018 -112 19994
rect 112 18018 146 19994
rect -146 15782 -112 17758
rect 112 15782 146 17758
rect -146 13546 -112 15522
rect 112 13546 146 15522
rect -146 11310 -112 13286
rect 112 11310 146 13286
rect -146 9074 -112 11050
rect 112 9074 146 11050
rect -146 6838 -112 8814
rect 112 6838 146 8814
rect -146 4602 -112 6578
rect 112 4602 146 6578
rect -146 2366 -112 4342
rect 112 2366 146 4342
rect -146 130 -112 2106
rect 112 130 146 2106
rect -146 -2106 -112 -130
rect 112 -2106 146 -130
rect -146 -4342 -112 -2366
rect 112 -4342 146 -2366
rect -146 -6578 -112 -4602
rect 112 -6578 146 -4602
rect -146 -8814 -112 -6838
rect 112 -8814 146 -6838
rect -146 -11050 -112 -9074
rect 112 -11050 146 -9074
rect -146 -13286 -112 -11310
rect 112 -13286 146 -11310
rect -146 -15522 -112 -13546
rect 112 -15522 146 -13546
rect -146 -17758 -112 -15782
rect 112 -17758 146 -15782
rect -146 -19994 -112 -18018
rect 112 -19994 146 -18018
rect -146 -22230 -112 -20254
rect 112 -22230 146 -20254
rect -146 -24466 -112 -22490
rect 112 -24466 146 -22490
rect -146 -26702 -112 -24726
rect 112 -26702 146 -24726
rect -146 -28938 -112 -26962
rect 112 -28938 146 -26962
rect -146 -31174 -112 -29198
rect 112 -31174 146 -29198
rect -146 -33410 -112 -31434
rect 112 -33410 146 -31434
rect -146 -35646 -112 -33670
rect 112 -35646 146 -33670
rect -146 -37882 -112 -35906
rect 112 -37882 146 -35906
rect -146 -40118 -112 -38142
rect 112 -40118 146 -38142
<< nsubdiff >>
rect -260 40279 -164 40313
rect 164 40279 260 40313
rect -260 40217 -226 40279
rect 226 40217 260 40279
rect -260 -40279 -226 -40217
rect 226 -40279 260 -40217
rect -260 -40313 -164 -40279
rect 164 -40313 260 -40279
<< nsubdiffcont >>
rect -164 40279 164 40313
rect -260 -40217 -226 40217
rect 226 -40217 260 40217
rect -164 -40313 164 -40279
<< poly >>
rect -100 40211 100 40227
rect -100 40177 -84 40211
rect 84 40177 100 40211
rect -100 40130 100 40177
rect -100 38083 100 38130
rect -100 38049 -84 38083
rect 84 38049 100 38083
rect -100 38033 100 38049
rect -100 37975 100 37991
rect -100 37941 -84 37975
rect 84 37941 100 37975
rect -100 37894 100 37941
rect -100 35847 100 35894
rect -100 35813 -84 35847
rect 84 35813 100 35847
rect -100 35797 100 35813
rect -100 35739 100 35755
rect -100 35705 -84 35739
rect 84 35705 100 35739
rect -100 35658 100 35705
rect -100 33611 100 33658
rect -100 33577 -84 33611
rect 84 33577 100 33611
rect -100 33561 100 33577
rect -100 33503 100 33519
rect -100 33469 -84 33503
rect 84 33469 100 33503
rect -100 33422 100 33469
rect -100 31375 100 31422
rect -100 31341 -84 31375
rect 84 31341 100 31375
rect -100 31325 100 31341
rect -100 31267 100 31283
rect -100 31233 -84 31267
rect 84 31233 100 31267
rect -100 31186 100 31233
rect -100 29139 100 29186
rect -100 29105 -84 29139
rect 84 29105 100 29139
rect -100 29089 100 29105
rect -100 29031 100 29047
rect -100 28997 -84 29031
rect 84 28997 100 29031
rect -100 28950 100 28997
rect -100 26903 100 26950
rect -100 26869 -84 26903
rect 84 26869 100 26903
rect -100 26853 100 26869
rect -100 26795 100 26811
rect -100 26761 -84 26795
rect 84 26761 100 26795
rect -100 26714 100 26761
rect -100 24667 100 24714
rect -100 24633 -84 24667
rect 84 24633 100 24667
rect -100 24617 100 24633
rect -100 24559 100 24575
rect -100 24525 -84 24559
rect 84 24525 100 24559
rect -100 24478 100 24525
rect -100 22431 100 22478
rect -100 22397 -84 22431
rect 84 22397 100 22431
rect -100 22381 100 22397
rect -100 22323 100 22339
rect -100 22289 -84 22323
rect 84 22289 100 22323
rect -100 22242 100 22289
rect -100 20195 100 20242
rect -100 20161 -84 20195
rect 84 20161 100 20195
rect -100 20145 100 20161
rect -100 20087 100 20103
rect -100 20053 -84 20087
rect 84 20053 100 20087
rect -100 20006 100 20053
rect -100 17959 100 18006
rect -100 17925 -84 17959
rect 84 17925 100 17959
rect -100 17909 100 17925
rect -100 17851 100 17867
rect -100 17817 -84 17851
rect 84 17817 100 17851
rect -100 17770 100 17817
rect -100 15723 100 15770
rect -100 15689 -84 15723
rect 84 15689 100 15723
rect -100 15673 100 15689
rect -100 15615 100 15631
rect -100 15581 -84 15615
rect 84 15581 100 15615
rect -100 15534 100 15581
rect -100 13487 100 13534
rect -100 13453 -84 13487
rect 84 13453 100 13487
rect -100 13437 100 13453
rect -100 13379 100 13395
rect -100 13345 -84 13379
rect 84 13345 100 13379
rect -100 13298 100 13345
rect -100 11251 100 11298
rect -100 11217 -84 11251
rect 84 11217 100 11251
rect -100 11201 100 11217
rect -100 11143 100 11159
rect -100 11109 -84 11143
rect 84 11109 100 11143
rect -100 11062 100 11109
rect -100 9015 100 9062
rect -100 8981 -84 9015
rect 84 8981 100 9015
rect -100 8965 100 8981
rect -100 8907 100 8923
rect -100 8873 -84 8907
rect 84 8873 100 8907
rect -100 8826 100 8873
rect -100 6779 100 6826
rect -100 6745 -84 6779
rect 84 6745 100 6779
rect -100 6729 100 6745
rect -100 6671 100 6687
rect -100 6637 -84 6671
rect 84 6637 100 6671
rect -100 6590 100 6637
rect -100 4543 100 4590
rect -100 4509 -84 4543
rect 84 4509 100 4543
rect -100 4493 100 4509
rect -100 4435 100 4451
rect -100 4401 -84 4435
rect 84 4401 100 4435
rect -100 4354 100 4401
rect -100 2307 100 2354
rect -100 2273 -84 2307
rect 84 2273 100 2307
rect -100 2257 100 2273
rect -100 2199 100 2215
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect -100 2118 100 2165
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -2165 100 -2118
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect -100 -2215 100 -2199
rect -100 -2273 100 -2257
rect -100 -2307 -84 -2273
rect 84 -2307 100 -2273
rect -100 -2354 100 -2307
rect -100 -4401 100 -4354
rect -100 -4435 -84 -4401
rect 84 -4435 100 -4401
rect -100 -4451 100 -4435
rect -100 -4509 100 -4493
rect -100 -4543 -84 -4509
rect 84 -4543 100 -4509
rect -100 -4590 100 -4543
rect -100 -6637 100 -6590
rect -100 -6671 -84 -6637
rect 84 -6671 100 -6637
rect -100 -6687 100 -6671
rect -100 -6745 100 -6729
rect -100 -6779 -84 -6745
rect 84 -6779 100 -6745
rect -100 -6826 100 -6779
rect -100 -8873 100 -8826
rect -100 -8907 -84 -8873
rect 84 -8907 100 -8873
rect -100 -8923 100 -8907
rect -100 -8981 100 -8965
rect -100 -9015 -84 -8981
rect 84 -9015 100 -8981
rect -100 -9062 100 -9015
rect -100 -11109 100 -11062
rect -100 -11143 -84 -11109
rect 84 -11143 100 -11109
rect -100 -11159 100 -11143
rect -100 -11217 100 -11201
rect -100 -11251 -84 -11217
rect 84 -11251 100 -11217
rect -100 -11298 100 -11251
rect -100 -13345 100 -13298
rect -100 -13379 -84 -13345
rect 84 -13379 100 -13345
rect -100 -13395 100 -13379
rect -100 -13453 100 -13437
rect -100 -13487 -84 -13453
rect 84 -13487 100 -13453
rect -100 -13534 100 -13487
rect -100 -15581 100 -15534
rect -100 -15615 -84 -15581
rect 84 -15615 100 -15581
rect -100 -15631 100 -15615
rect -100 -15689 100 -15673
rect -100 -15723 -84 -15689
rect 84 -15723 100 -15689
rect -100 -15770 100 -15723
rect -100 -17817 100 -17770
rect -100 -17851 -84 -17817
rect 84 -17851 100 -17817
rect -100 -17867 100 -17851
rect -100 -17925 100 -17909
rect -100 -17959 -84 -17925
rect 84 -17959 100 -17925
rect -100 -18006 100 -17959
rect -100 -20053 100 -20006
rect -100 -20087 -84 -20053
rect 84 -20087 100 -20053
rect -100 -20103 100 -20087
rect -100 -20161 100 -20145
rect -100 -20195 -84 -20161
rect 84 -20195 100 -20161
rect -100 -20242 100 -20195
rect -100 -22289 100 -22242
rect -100 -22323 -84 -22289
rect 84 -22323 100 -22289
rect -100 -22339 100 -22323
rect -100 -22397 100 -22381
rect -100 -22431 -84 -22397
rect 84 -22431 100 -22397
rect -100 -22478 100 -22431
rect -100 -24525 100 -24478
rect -100 -24559 -84 -24525
rect 84 -24559 100 -24525
rect -100 -24575 100 -24559
rect -100 -24633 100 -24617
rect -100 -24667 -84 -24633
rect 84 -24667 100 -24633
rect -100 -24714 100 -24667
rect -100 -26761 100 -26714
rect -100 -26795 -84 -26761
rect 84 -26795 100 -26761
rect -100 -26811 100 -26795
rect -100 -26869 100 -26853
rect -100 -26903 -84 -26869
rect 84 -26903 100 -26869
rect -100 -26950 100 -26903
rect -100 -28997 100 -28950
rect -100 -29031 -84 -28997
rect 84 -29031 100 -28997
rect -100 -29047 100 -29031
rect -100 -29105 100 -29089
rect -100 -29139 -84 -29105
rect 84 -29139 100 -29105
rect -100 -29186 100 -29139
rect -100 -31233 100 -31186
rect -100 -31267 -84 -31233
rect 84 -31267 100 -31233
rect -100 -31283 100 -31267
rect -100 -31341 100 -31325
rect -100 -31375 -84 -31341
rect 84 -31375 100 -31341
rect -100 -31422 100 -31375
rect -100 -33469 100 -33422
rect -100 -33503 -84 -33469
rect 84 -33503 100 -33469
rect -100 -33519 100 -33503
rect -100 -33577 100 -33561
rect -100 -33611 -84 -33577
rect 84 -33611 100 -33577
rect -100 -33658 100 -33611
rect -100 -35705 100 -35658
rect -100 -35739 -84 -35705
rect 84 -35739 100 -35705
rect -100 -35755 100 -35739
rect -100 -35813 100 -35797
rect -100 -35847 -84 -35813
rect 84 -35847 100 -35813
rect -100 -35894 100 -35847
rect -100 -37941 100 -37894
rect -100 -37975 -84 -37941
rect 84 -37975 100 -37941
rect -100 -37991 100 -37975
rect -100 -38049 100 -38033
rect -100 -38083 -84 -38049
rect 84 -38083 100 -38049
rect -100 -38130 100 -38083
rect -100 -40177 100 -40130
rect -100 -40211 -84 -40177
rect 84 -40211 100 -40177
rect -100 -40227 100 -40211
<< polycont >>
rect -84 40177 84 40211
rect -84 38049 84 38083
rect -84 37941 84 37975
rect -84 35813 84 35847
rect -84 35705 84 35739
rect -84 33577 84 33611
rect -84 33469 84 33503
rect -84 31341 84 31375
rect -84 31233 84 31267
rect -84 29105 84 29139
rect -84 28997 84 29031
rect -84 26869 84 26903
rect -84 26761 84 26795
rect -84 24633 84 24667
rect -84 24525 84 24559
rect -84 22397 84 22431
rect -84 22289 84 22323
rect -84 20161 84 20195
rect -84 20053 84 20087
rect -84 17925 84 17959
rect -84 17817 84 17851
rect -84 15689 84 15723
rect -84 15581 84 15615
rect -84 13453 84 13487
rect -84 13345 84 13379
rect -84 11217 84 11251
rect -84 11109 84 11143
rect -84 8981 84 9015
rect -84 8873 84 8907
rect -84 6745 84 6779
rect -84 6637 84 6671
rect -84 4509 84 4543
rect -84 4401 84 4435
rect -84 2273 84 2307
rect -84 2165 84 2199
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -2199 84 -2165
rect -84 -2307 84 -2273
rect -84 -4435 84 -4401
rect -84 -4543 84 -4509
rect -84 -6671 84 -6637
rect -84 -6779 84 -6745
rect -84 -8907 84 -8873
rect -84 -9015 84 -8981
rect -84 -11143 84 -11109
rect -84 -11251 84 -11217
rect -84 -13379 84 -13345
rect -84 -13487 84 -13453
rect -84 -15615 84 -15581
rect -84 -15723 84 -15689
rect -84 -17851 84 -17817
rect -84 -17959 84 -17925
rect -84 -20087 84 -20053
rect -84 -20195 84 -20161
rect -84 -22323 84 -22289
rect -84 -22431 84 -22397
rect -84 -24559 84 -24525
rect -84 -24667 84 -24633
rect -84 -26795 84 -26761
rect -84 -26903 84 -26869
rect -84 -29031 84 -28997
rect -84 -29139 84 -29105
rect -84 -31267 84 -31233
rect -84 -31375 84 -31341
rect -84 -33503 84 -33469
rect -84 -33611 84 -33577
rect -84 -35739 84 -35705
rect -84 -35847 84 -35813
rect -84 -37975 84 -37941
rect -84 -38083 84 -38049
rect -84 -40211 84 -40177
<< locali >>
rect -260 40279 -164 40313
rect 164 40279 260 40313
rect -260 40217 -226 40279
rect 226 40217 260 40279
rect -100 40177 -84 40211
rect 84 40177 100 40211
rect -146 40118 -112 40134
rect -146 38126 -112 38142
rect 112 40118 146 40134
rect 112 38126 146 38142
rect -100 38049 -84 38083
rect 84 38049 100 38083
rect -100 37941 -84 37975
rect 84 37941 100 37975
rect -146 37882 -112 37898
rect -146 35890 -112 35906
rect 112 37882 146 37898
rect 112 35890 146 35906
rect -100 35813 -84 35847
rect 84 35813 100 35847
rect -100 35705 -84 35739
rect 84 35705 100 35739
rect -146 35646 -112 35662
rect -146 33654 -112 33670
rect 112 35646 146 35662
rect 112 33654 146 33670
rect -100 33577 -84 33611
rect 84 33577 100 33611
rect -100 33469 -84 33503
rect 84 33469 100 33503
rect -146 33410 -112 33426
rect -146 31418 -112 31434
rect 112 33410 146 33426
rect 112 31418 146 31434
rect -100 31341 -84 31375
rect 84 31341 100 31375
rect -100 31233 -84 31267
rect 84 31233 100 31267
rect -146 31174 -112 31190
rect -146 29182 -112 29198
rect 112 31174 146 31190
rect 112 29182 146 29198
rect -100 29105 -84 29139
rect 84 29105 100 29139
rect -100 28997 -84 29031
rect 84 28997 100 29031
rect -146 28938 -112 28954
rect -146 26946 -112 26962
rect 112 28938 146 28954
rect 112 26946 146 26962
rect -100 26869 -84 26903
rect 84 26869 100 26903
rect -100 26761 -84 26795
rect 84 26761 100 26795
rect -146 26702 -112 26718
rect -146 24710 -112 24726
rect 112 26702 146 26718
rect 112 24710 146 24726
rect -100 24633 -84 24667
rect 84 24633 100 24667
rect -100 24525 -84 24559
rect 84 24525 100 24559
rect -146 24466 -112 24482
rect -146 22474 -112 22490
rect 112 24466 146 24482
rect 112 22474 146 22490
rect -100 22397 -84 22431
rect 84 22397 100 22431
rect -100 22289 -84 22323
rect 84 22289 100 22323
rect -146 22230 -112 22246
rect -146 20238 -112 20254
rect 112 22230 146 22246
rect 112 20238 146 20254
rect -100 20161 -84 20195
rect 84 20161 100 20195
rect -100 20053 -84 20087
rect 84 20053 100 20087
rect -146 19994 -112 20010
rect -146 18002 -112 18018
rect 112 19994 146 20010
rect 112 18002 146 18018
rect -100 17925 -84 17959
rect 84 17925 100 17959
rect -100 17817 -84 17851
rect 84 17817 100 17851
rect -146 17758 -112 17774
rect -146 15766 -112 15782
rect 112 17758 146 17774
rect 112 15766 146 15782
rect -100 15689 -84 15723
rect 84 15689 100 15723
rect -100 15581 -84 15615
rect 84 15581 100 15615
rect -146 15522 -112 15538
rect -146 13530 -112 13546
rect 112 15522 146 15538
rect 112 13530 146 13546
rect -100 13453 -84 13487
rect 84 13453 100 13487
rect -100 13345 -84 13379
rect 84 13345 100 13379
rect -146 13286 -112 13302
rect -146 11294 -112 11310
rect 112 13286 146 13302
rect 112 11294 146 11310
rect -100 11217 -84 11251
rect 84 11217 100 11251
rect -100 11109 -84 11143
rect 84 11109 100 11143
rect -146 11050 -112 11066
rect -146 9058 -112 9074
rect 112 11050 146 11066
rect 112 9058 146 9074
rect -100 8981 -84 9015
rect 84 8981 100 9015
rect -100 8873 -84 8907
rect 84 8873 100 8907
rect -146 8814 -112 8830
rect -146 6822 -112 6838
rect 112 8814 146 8830
rect 112 6822 146 6838
rect -100 6745 -84 6779
rect 84 6745 100 6779
rect -100 6637 -84 6671
rect 84 6637 100 6671
rect -146 6578 -112 6594
rect -146 4586 -112 4602
rect 112 6578 146 6594
rect 112 4586 146 4602
rect -100 4509 -84 4543
rect 84 4509 100 4543
rect -100 4401 -84 4435
rect 84 4401 100 4435
rect -146 4342 -112 4358
rect -146 2350 -112 2366
rect 112 4342 146 4358
rect 112 2350 146 2366
rect -100 2273 -84 2307
rect 84 2273 100 2307
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect -146 2106 -112 2122
rect -146 114 -112 130
rect 112 2106 146 2122
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -2122 -112 -2106
rect 112 -130 146 -114
rect 112 -2122 146 -2106
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect -100 -2307 -84 -2273
rect 84 -2307 100 -2273
rect -146 -2366 -112 -2350
rect -146 -4358 -112 -4342
rect 112 -2366 146 -2350
rect 112 -4358 146 -4342
rect -100 -4435 -84 -4401
rect 84 -4435 100 -4401
rect -100 -4543 -84 -4509
rect 84 -4543 100 -4509
rect -146 -4602 -112 -4586
rect -146 -6594 -112 -6578
rect 112 -4602 146 -4586
rect 112 -6594 146 -6578
rect -100 -6671 -84 -6637
rect 84 -6671 100 -6637
rect -100 -6779 -84 -6745
rect 84 -6779 100 -6745
rect -146 -6838 -112 -6822
rect -146 -8830 -112 -8814
rect 112 -6838 146 -6822
rect 112 -8830 146 -8814
rect -100 -8907 -84 -8873
rect 84 -8907 100 -8873
rect -100 -9015 -84 -8981
rect 84 -9015 100 -8981
rect -146 -9074 -112 -9058
rect -146 -11066 -112 -11050
rect 112 -9074 146 -9058
rect 112 -11066 146 -11050
rect -100 -11143 -84 -11109
rect 84 -11143 100 -11109
rect -100 -11251 -84 -11217
rect 84 -11251 100 -11217
rect -146 -11310 -112 -11294
rect -146 -13302 -112 -13286
rect 112 -11310 146 -11294
rect 112 -13302 146 -13286
rect -100 -13379 -84 -13345
rect 84 -13379 100 -13345
rect -100 -13487 -84 -13453
rect 84 -13487 100 -13453
rect -146 -13546 -112 -13530
rect -146 -15538 -112 -15522
rect 112 -13546 146 -13530
rect 112 -15538 146 -15522
rect -100 -15615 -84 -15581
rect 84 -15615 100 -15581
rect -100 -15723 -84 -15689
rect 84 -15723 100 -15689
rect -146 -15782 -112 -15766
rect -146 -17774 -112 -17758
rect 112 -15782 146 -15766
rect 112 -17774 146 -17758
rect -100 -17851 -84 -17817
rect 84 -17851 100 -17817
rect -100 -17959 -84 -17925
rect 84 -17959 100 -17925
rect -146 -18018 -112 -18002
rect -146 -20010 -112 -19994
rect 112 -18018 146 -18002
rect 112 -20010 146 -19994
rect -100 -20087 -84 -20053
rect 84 -20087 100 -20053
rect -100 -20195 -84 -20161
rect 84 -20195 100 -20161
rect -146 -20254 -112 -20238
rect -146 -22246 -112 -22230
rect 112 -20254 146 -20238
rect 112 -22246 146 -22230
rect -100 -22323 -84 -22289
rect 84 -22323 100 -22289
rect -100 -22431 -84 -22397
rect 84 -22431 100 -22397
rect -146 -22490 -112 -22474
rect -146 -24482 -112 -24466
rect 112 -22490 146 -22474
rect 112 -24482 146 -24466
rect -100 -24559 -84 -24525
rect 84 -24559 100 -24525
rect -100 -24667 -84 -24633
rect 84 -24667 100 -24633
rect -146 -24726 -112 -24710
rect -146 -26718 -112 -26702
rect 112 -24726 146 -24710
rect 112 -26718 146 -26702
rect -100 -26795 -84 -26761
rect 84 -26795 100 -26761
rect -100 -26903 -84 -26869
rect 84 -26903 100 -26869
rect -146 -26962 -112 -26946
rect -146 -28954 -112 -28938
rect 112 -26962 146 -26946
rect 112 -28954 146 -28938
rect -100 -29031 -84 -28997
rect 84 -29031 100 -28997
rect -100 -29139 -84 -29105
rect 84 -29139 100 -29105
rect -146 -29198 -112 -29182
rect -146 -31190 -112 -31174
rect 112 -29198 146 -29182
rect 112 -31190 146 -31174
rect -100 -31267 -84 -31233
rect 84 -31267 100 -31233
rect -100 -31375 -84 -31341
rect 84 -31375 100 -31341
rect -146 -31434 -112 -31418
rect -146 -33426 -112 -33410
rect 112 -31434 146 -31418
rect 112 -33426 146 -33410
rect -100 -33503 -84 -33469
rect 84 -33503 100 -33469
rect -100 -33611 -84 -33577
rect 84 -33611 100 -33577
rect -146 -33670 -112 -33654
rect -146 -35662 -112 -35646
rect 112 -33670 146 -33654
rect 112 -35662 146 -35646
rect -100 -35739 -84 -35705
rect 84 -35739 100 -35705
rect -100 -35847 -84 -35813
rect 84 -35847 100 -35813
rect -146 -35906 -112 -35890
rect -146 -37898 -112 -37882
rect 112 -35906 146 -35890
rect 112 -37898 146 -37882
rect -100 -37975 -84 -37941
rect 84 -37975 100 -37941
rect -100 -38083 -84 -38049
rect 84 -38083 100 -38049
rect -146 -38142 -112 -38126
rect -146 -40134 -112 -40118
rect 112 -38142 146 -38126
rect 112 -40134 146 -40118
rect -100 -40211 -84 -40177
rect 84 -40211 100 -40177
rect -260 -40279 -226 -40217
rect 226 -40279 260 -40217
rect -260 -40313 -164 -40279
rect 164 -40313 260 -40279
<< viali >>
rect -84 40177 84 40211
rect -146 38142 -112 40118
rect 112 38142 146 40118
rect -84 38049 84 38083
rect -84 37941 84 37975
rect -146 35906 -112 37882
rect 112 35906 146 37882
rect -84 35813 84 35847
rect -84 35705 84 35739
rect -146 33670 -112 35646
rect 112 33670 146 35646
rect -84 33577 84 33611
rect -84 33469 84 33503
rect -146 31434 -112 33410
rect 112 31434 146 33410
rect -84 31341 84 31375
rect -84 31233 84 31267
rect -146 29198 -112 31174
rect 112 29198 146 31174
rect -84 29105 84 29139
rect -84 28997 84 29031
rect -146 26962 -112 28938
rect 112 26962 146 28938
rect -84 26869 84 26903
rect -84 26761 84 26795
rect -146 24726 -112 26702
rect 112 24726 146 26702
rect -84 24633 84 24667
rect -84 24525 84 24559
rect -146 22490 -112 24466
rect 112 22490 146 24466
rect -84 22397 84 22431
rect -84 22289 84 22323
rect -146 20254 -112 22230
rect 112 20254 146 22230
rect -84 20161 84 20195
rect -84 20053 84 20087
rect -146 18018 -112 19994
rect 112 18018 146 19994
rect -84 17925 84 17959
rect -84 17817 84 17851
rect -146 15782 -112 17758
rect 112 15782 146 17758
rect -84 15689 84 15723
rect -84 15581 84 15615
rect -146 13546 -112 15522
rect 112 13546 146 15522
rect -84 13453 84 13487
rect -84 13345 84 13379
rect -146 11310 -112 13286
rect 112 11310 146 13286
rect -84 11217 84 11251
rect -84 11109 84 11143
rect -146 9074 -112 11050
rect 112 9074 146 11050
rect -84 8981 84 9015
rect -84 8873 84 8907
rect -146 6838 -112 8814
rect 112 6838 146 8814
rect -84 6745 84 6779
rect -84 6637 84 6671
rect -146 4602 -112 6578
rect 112 4602 146 6578
rect -84 4509 84 4543
rect -84 4401 84 4435
rect -146 2366 -112 4342
rect 112 2366 146 4342
rect -84 2273 84 2307
rect -84 2165 84 2199
rect -146 130 -112 2106
rect 112 130 146 2106
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -2106 -112 -130
rect 112 -2106 146 -130
rect -84 -2199 84 -2165
rect -84 -2307 84 -2273
rect -146 -4342 -112 -2366
rect 112 -4342 146 -2366
rect -84 -4435 84 -4401
rect -84 -4543 84 -4509
rect -146 -6578 -112 -4602
rect 112 -6578 146 -4602
rect -84 -6671 84 -6637
rect -84 -6779 84 -6745
rect -146 -8814 -112 -6838
rect 112 -8814 146 -6838
rect -84 -8907 84 -8873
rect -84 -9015 84 -8981
rect -146 -11050 -112 -9074
rect 112 -11050 146 -9074
rect -84 -11143 84 -11109
rect -84 -11251 84 -11217
rect -146 -13286 -112 -11310
rect 112 -13286 146 -11310
rect -84 -13379 84 -13345
rect -84 -13487 84 -13453
rect -146 -15522 -112 -13546
rect 112 -15522 146 -13546
rect -84 -15615 84 -15581
rect -84 -15723 84 -15689
rect -146 -17758 -112 -15782
rect 112 -17758 146 -15782
rect -84 -17851 84 -17817
rect -84 -17959 84 -17925
rect -146 -19994 -112 -18018
rect 112 -19994 146 -18018
rect -84 -20087 84 -20053
rect -84 -20195 84 -20161
rect -146 -22230 -112 -20254
rect 112 -22230 146 -20254
rect -84 -22323 84 -22289
rect -84 -22431 84 -22397
rect -146 -24466 -112 -22490
rect 112 -24466 146 -22490
rect -84 -24559 84 -24525
rect -84 -24667 84 -24633
rect -146 -26702 -112 -24726
rect 112 -26702 146 -24726
rect -84 -26795 84 -26761
rect -84 -26903 84 -26869
rect -146 -28938 -112 -26962
rect 112 -28938 146 -26962
rect -84 -29031 84 -28997
rect -84 -29139 84 -29105
rect -146 -31174 -112 -29198
rect 112 -31174 146 -29198
rect -84 -31267 84 -31233
rect -84 -31375 84 -31341
rect -146 -33410 -112 -31434
rect 112 -33410 146 -31434
rect -84 -33503 84 -33469
rect -84 -33611 84 -33577
rect -146 -35646 -112 -33670
rect 112 -35646 146 -33670
rect -84 -35739 84 -35705
rect -84 -35847 84 -35813
rect -146 -37882 -112 -35906
rect 112 -37882 146 -35906
rect -84 -37975 84 -37941
rect -84 -38083 84 -38049
rect -146 -40118 -112 -38142
rect 112 -40118 146 -38142
rect -84 -40211 84 -40177
<< metal1 >>
rect -96 40211 96 40217
rect -96 40177 -84 40211
rect 84 40177 96 40211
rect -96 40171 96 40177
rect -152 40118 -106 40130
rect -152 38142 -146 40118
rect -112 38142 -106 40118
rect -152 38130 -106 38142
rect 106 40118 152 40130
rect 106 38142 112 40118
rect 146 38142 152 40118
rect 106 38130 152 38142
rect -96 38083 96 38089
rect -96 38049 -84 38083
rect 84 38049 96 38083
rect -96 38043 96 38049
rect -96 37975 96 37981
rect -96 37941 -84 37975
rect 84 37941 96 37975
rect -96 37935 96 37941
rect -152 37882 -106 37894
rect -152 35906 -146 37882
rect -112 35906 -106 37882
rect -152 35894 -106 35906
rect 106 37882 152 37894
rect 106 35906 112 37882
rect 146 35906 152 37882
rect 106 35894 152 35906
rect -96 35847 96 35853
rect -96 35813 -84 35847
rect 84 35813 96 35847
rect -96 35807 96 35813
rect -96 35739 96 35745
rect -96 35705 -84 35739
rect 84 35705 96 35739
rect -96 35699 96 35705
rect -152 35646 -106 35658
rect -152 33670 -146 35646
rect -112 33670 -106 35646
rect -152 33658 -106 33670
rect 106 35646 152 35658
rect 106 33670 112 35646
rect 146 33670 152 35646
rect 106 33658 152 33670
rect -96 33611 96 33617
rect -96 33577 -84 33611
rect 84 33577 96 33611
rect -96 33571 96 33577
rect -96 33503 96 33509
rect -96 33469 -84 33503
rect 84 33469 96 33503
rect -96 33463 96 33469
rect -152 33410 -106 33422
rect -152 31434 -146 33410
rect -112 31434 -106 33410
rect -152 31422 -106 31434
rect 106 33410 152 33422
rect 106 31434 112 33410
rect 146 31434 152 33410
rect 106 31422 152 31434
rect -96 31375 96 31381
rect -96 31341 -84 31375
rect 84 31341 96 31375
rect -96 31335 96 31341
rect -96 31267 96 31273
rect -96 31233 -84 31267
rect 84 31233 96 31267
rect -96 31227 96 31233
rect -152 31174 -106 31186
rect -152 29198 -146 31174
rect -112 29198 -106 31174
rect -152 29186 -106 29198
rect 106 31174 152 31186
rect 106 29198 112 31174
rect 146 29198 152 31174
rect 106 29186 152 29198
rect -96 29139 96 29145
rect -96 29105 -84 29139
rect 84 29105 96 29139
rect -96 29099 96 29105
rect -96 29031 96 29037
rect -96 28997 -84 29031
rect 84 28997 96 29031
rect -96 28991 96 28997
rect -152 28938 -106 28950
rect -152 26962 -146 28938
rect -112 26962 -106 28938
rect -152 26950 -106 26962
rect 106 28938 152 28950
rect 106 26962 112 28938
rect 146 26962 152 28938
rect 106 26950 152 26962
rect -96 26903 96 26909
rect -96 26869 -84 26903
rect 84 26869 96 26903
rect -96 26863 96 26869
rect -96 26795 96 26801
rect -96 26761 -84 26795
rect 84 26761 96 26795
rect -96 26755 96 26761
rect -152 26702 -106 26714
rect -152 24726 -146 26702
rect -112 24726 -106 26702
rect -152 24714 -106 24726
rect 106 26702 152 26714
rect 106 24726 112 26702
rect 146 24726 152 26702
rect 106 24714 152 24726
rect -96 24667 96 24673
rect -96 24633 -84 24667
rect 84 24633 96 24667
rect -96 24627 96 24633
rect -96 24559 96 24565
rect -96 24525 -84 24559
rect 84 24525 96 24559
rect -96 24519 96 24525
rect -152 24466 -106 24478
rect -152 22490 -146 24466
rect -112 22490 -106 24466
rect -152 22478 -106 22490
rect 106 24466 152 24478
rect 106 22490 112 24466
rect 146 22490 152 24466
rect 106 22478 152 22490
rect -96 22431 96 22437
rect -96 22397 -84 22431
rect 84 22397 96 22431
rect -96 22391 96 22397
rect -96 22323 96 22329
rect -96 22289 -84 22323
rect 84 22289 96 22323
rect -96 22283 96 22289
rect -152 22230 -106 22242
rect -152 20254 -146 22230
rect -112 20254 -106 22230
rect -152 20242 -106 20254
rect 106 22230 152 22242
rect 106 20254 112 22230
rect 146 20254 152 22230
rect 106 20242 152 20254
rect -96 20195 96 20201
rect -96 20161 -84 20195
rect 84 20161 96 20195
rect -96 20155 96 20161
rect -96 20087 96 20093
rect -96 20053 -84 20087
rect 84 20053 96 20087
rect -96 20047 96 20053
rect -152 19994 -106 20006
rect -152 18018 -146 19994
rect -112 18018 -106 19994
rect -152 18006 -106 18018
rect 106 19994 152 20006
rect 106 18018 112 19994
rect 146 18018 152 19994
rect 106 18006 152 18018
rect -96 17959 96 17965
rect -96 17925 -84 17959
rect 84 17925 96 17959
rect -96 17919 96 17925
rect -96 17851 96 17857
rect -96 17817 -84 17851
rect 84 17817 96 17851
rect -96 17811 96 17817
rect -152 17758 -106 17770
rect -152 15782 -146 17758
rect -112 15782 -106 17758
rect -152 15770 -106 15782
rect 106 17758 152 17770
rect 106 15782 112 17758
rect 146 15782 152 17758
rect 106 15770 152 15782
rect -96 15723 96 15729
rect -96 15689 -84 15723
rect 84 15689 96 15723
rect -96 15683 96 15689
rect -96 15615 96 15621
rect -96 15581 -84 15615
rect 84 15581 96 15615
rect -96 15575 96 15581
rect -152 15522 -106 15534
rect -152 13546 -146 15522
rect -112 13546 -106 15522
rect -152 13534 -106 13546
rect 106 15522 152 15534
rect 106 13546 112 15522
rect 146 13546 152 15522
rect 106 13534 152 13546
rect -96 13487 96 13493
rect -96 13453 -84 13487
rect 84 13453 96 13487
rect -96 13447 96 13453
rect -96 13379 96 13385
rect -96 13345 -84 13379
rect 84 13345 96 13379
rect -96 13339 96 13345
rect -152 13286 -106 13298
rect -152 11310 -146 13286
rect -112 11310 -106 13286
rect -152 11298 -106 11310
rect 106 13286 152 13298
rect 106 11310 112 13286
rect 146 11310 152 13286
rect 106 11298 152 11310
rect -96 11251 96 11257
rect -96 11217 -84 11251
rect 84 11217 96 11251
rect -96 11211 96 11217
rect -96 11143 96 11149
rect -96 11109 -84 11143
rect 84 11109 96 11143
rect -96 11103 96 11109
rect -152 11050 -106 11062
rect -152 9074 -146 11050
rect -112 9074 -106 11050
rect -152 9062 -106 9074
rect 106 11050 152 11062
rect 106 9074 112 11050
rect 146 9074 152 11050
rect 106 9062 152 9074
rect -96 9015 96 9021
rect -96 8981 -84 9015
rect 84 8981 96 9015
rect -96 8975 96 8981
rect -96 8907 96 8913
rect -96 8873 -84 8907
rect 84 8873 96 8907
rect -96 8867 96 8873
rect -152 8814 -106 8826
rect -152 6838 -146 8814
rect -112 6838 -106 8814
rect -152 6826 -106 6838
rect 106 8814 152 8826
rect 106 6838 112 8814
rect 146 6838 152 8814
rect 106 6826 152 6838
rect -96 6779 96 6785
rect -96 6745 -84 6779
rect 84 6745 96 6779
rect -96 6739 96 6745
rect -96 6671 96 6677
rect -96 6637 -84 6671
rect 84 6637 96 6671
rect -96 6631 96 6637
rect -152 6578 -106 6590
rect -152 4602 -146 6578
rect -112 4602 -106 6578
rect -152 4590 -106 4602
rect 106 6578 152 6590
rect 106 4602 112 6578
rect 146 4602 152 6578
rect 106 4590 152 4602
rect -96 4543 96 4549
rect -96 4509 -84 4543
rect 84 4509 96 4543
rect -96 4503 96 4509
rect -96 4435 96 4441
rect -96 4401 -84 4435
rect 84 4401 96 4435
rect -96 4395 96 4401
rect -152 4342 -106 4354
rect -152 2366 -146 4342
rect -112 2366 -106 4342
rect -152 2354 -106 2366
rect 106 4342 152 4354
rect 106 2366 112 4342
rect 146 2366 152 4342
rect 106 2354 152 2366
rect -96 2307 96 2313
rect -96 2273 -84 2307
rect 84 2273 96 2307
rect -96 2267 96 2273
rect -96 2199 96 2205
rect -96 2165 -84 2199
rect 84 2165 96 2199
rect -96 2159 96 2165
rect -152 2106 -106 2118
rect -152 130 -146 2106
rect -112 130 -106 2106
rect -152 118 -106 130
rect 106 2106 152 2118
rect 106 130 112 2106
rect 146 130 152 2106
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -2106 -146 -130
rect -112 -2106 -106 -130
rect -152 -2118 -106 -2106
rect 106 -130 152 -118
rect 106 -2106 112 -130
rect 146 -2106 152 -130
rect 106 -2118 152 -2106
rect -96 -2165 96 -2159
rect -96 -2199 -84 -2165
rect 84 -2199 96 -2165
rect -96 -2205 96 -2199
rect -96 -2273 96 -2267
rect -96 -2307 -84 -2273
rect 84 -2307 96 -2273
rect -96 -2313 96 -2307
rect -152 -2366 -106 -2354
rect -152 -4342 -146 -2366
rect -112 -4342 -106 -2366
rect -152 -4354 -106 -4342
rect 106 -2366 152 -2354
rect 106 -4342 112 -2366
rect 146 -4342 152 -2366
rect 106 -4354 152 -4342
rect -96 -4401 96 -4395
rect -96 -4435 -84 -4401
rect 84 -4435 96 -4401
rect -96 -4441 96 -4435
rect -96 -4509 96 -4503
rect -96 -4543 -84 -4509
rect 84 -4543 96 -4509
rect -96 -4549 96 -4543
rect -152 -4602 -106 -4590
rect -152 -6578 -146 -4602
rect -112 -6578 -106 -4602
rect -152 -6590 -106 -6578
rect 106 -4602 152 -4590
rect 106 -6578 112 -4602
rect 146 -6578 152 -4602
rect 106 -6590 152 -6578
rect -96 -6637 96 -6631
rect -96 -6671 -84 -6637
rect 84 -6671 96 -6637
rect -96 -6677 96 -6671
rect -96 -6745 96 -6739
rect -96 -6779 -84 -6745
rect 84 -6779 96 -6745
rect -96 -6785 96 -6779
rect -152 -6838 -106 -6826
rect -152 -8814 -146 -6838
rect -112 -8814 -106 -6838
rect -152 -8826 -106 -8814
rect 106 -6838 152 -6826
rect 106 -8814 112 -6838
rect 146 -8814 152 -6838
rect 106 -8826 152 -8814
rect -96 -8873 96 -8867
rect -96 -8907 -84 -8873
rect 84 -8907 96 -8873
rect -96 -8913 96 -8907
rect -96 -8981 96 -8975
rect -96 -9015 -84 -8981
rect 84 -9015 96 -8981
rect -96 -9021 96 -9015
rect -152 -9074 -106 -9062
rect -152 -11050 -146 -9074
rect -112 -11050 -106 -9074
rect -152 -11062 -106 -11050
rect 106 -9074 152 -9062
rect 106 -11050 112 -9074
rect 146 -11050 152 -9074
rect 106 -11062 152 -11050
rect -96 -11109 96 -11103
rect -96 -11143 -84 -11109
rect 84 -11143 96 -11109
rect -96 -11149 96 -11143
rect -96 -11217 96 -11211
rect -96 -11251 -84 -11217
rect 84 -11251 96 -11217
rect -96 -11257 96 -11251
rect -152 -11310 -106 -11298
rect -152 -13286 -146 -11310
rect -112 -13286 -106 -11310
rect -152 -13298 -106 -13286
rect 106 -11310 152 -11298
rect 106 -13286 112 -11310
rect 146 -13286 152 -11310
rect 106 -13298 152 -13286
rect -96 -13345 96 -13339
rect -96 -13379 -84 -13345
rect 84 -13379 96 -13345
rect -96 -13385 96 -13379
rect -96 -13453 96 -13447
rect -96 -13487 -84 -13453
rect 84 -13487 96 -13453
rect -96 -13493 96 -13487
rect -152 -13546 -106 -13534
rect -152 -15522 -146 -13546
rect -112 -15522 -106 -13546
rect -152 -15534 -106 -15522
rect 106 -13546 152 -13534
rect 106 -15522 112 -13546
rect 146 -15522 152 -13546
rect 106 -15534 152 -15522
rect -96 -15581 96 -15575
rect -96 -15615 -84 -15581
rect 84 -15615 96 -15581
rect -96 -15621 96 -15615
rect -96 -15689 96 -15683
rect -96 -15723 -84 -15689
rect 84 -15723 96 -15689
rect -96 -15729 96 -15723
rect -152 -15782 -106 -15770
rect -152 -17758 -146 -15782
rect -112 -17758 -106 -15782
rect -152 -17770 -106 -17758
rect 106 -15782 152 -15770
rect 106 -17758 112 -15782
rect 146 -17758 152 -15782
rect 106 -17770 152 -17758
rect -96 -17817 96 -17811
rect -96 -17851 -84 -17817
rect 84 -17851 96 -17817
rect -96 -17857 96 -17851
rect -96 -17925 96 -17919
rect -96 -17959 -84 -17925
rect 84 -17959 96 -17925
rect -96 -17965 96 -17959
rect -152 -18018 -106 -18006
rect -152 -19994 -146 -18018
rect -112 -19994 -106 -18018
rect -152 -20006 -106 -19994
rect 106 -18018 152 -18006
rect 106 -19994 112 -18018
rect 146 -19994 152 -18018
rect 106 -20006 152 -19994
rect -96 -20053 96 -20047
rect -96 -20087 -84 -20053
rect 84 -20087 96 -20053
rect -96 -20093 96 -20087
rect -96 -20161 96 -20155
rect -96 -20195 -84 -20161
rect 84 -20195 96 -20161
rect -96 -20201 96 -20195
rect -152 -20254 -106 -20242
rect -152 -22230 -146 -20254
rect -112 -22230 -106 -20254
rect -152 -22242 -106 -22230
rect 106 -20254 152 -20242
rect 106 -22230 112 -20254
rect 146 -22230 152 -20254
rect 106 -22242 152 -22230
rect -96 -22289 96 -22283
rect -96 -22323 -84 -22289
rect 84 -22323 96 -22289
rect -96 -22329 96 -22323
rect -96 -22397 96 -22391
rect -96 -22431 -84 -22397
rect 84 -22431 96 -22397
rect -96 -22437 96 -22431
rect -152 -22490 -106 -22478
rect -152 -24466 -146 -22490
rect -112 -24466 -106 -22490
rect -152 -24478 -106 -24466
rect 106 -22490 152 -22478
rect 106 -24466 112 -22490
rect 146 -24466 152 -22490
rect 106 -24478 152 -24466
rect -96 -24525 96 -24519
rect -96 -24559 -84 -24525
rect 84 -24559 96 -24525
rect -96 -24565 96 -24559
rect -96 -24633 96 -24627
rect -96 -24667 -84 -24633
rect 84 -24667 96 -24633
rect -96 -24673 96 -24667
rect -152 -24726 -106 -24714
rect -152 -26702 -146 -24726
rect -112 -26702 -106 -24726
rect -152 -26714 -106 -26702
rect 106 -24726 152 -24714
rect 106 -26702 112 -24726
rect 146 -26702 152 -24726
rect 106 -26714 152 -26702
rect -96 -26761 96 -26755
rect -96 -26795 -84 -26761
rect 84 -26795 96 -26761
rect -96 -26801 96 -26795
rect -96 -26869 96 -26863
rect -96 -26903 -84 -26869
rect 84 -26903 96 -26869
rect -96 -26909 96 -26903
rect -152 -26962 -106 -26950
rect -152 -28938 -146 -26962
rect -112 -28938 -106 -26962
rect -152 -28950 -106 -28938
rect 106 -26962 152 -26950
rect 106 -28938 112 -26962
rect 146 -28938 152 -26962
rect 106 -28950 152 -28938
rect -96 -28997 96 -28991
rect -96 -29031 -84 -28997
rect 84 -29031 96 -28997
rect -96 -29037 96 -29031
rect -96 -29105 96 -29099
rect -96 -29139 -84 -29105
rect 84 -29139 96 -29105
rect -96 -29145 96 -29139
rect -152 -29198 -106 -29186
rect -152 -31174 -146 -29198
rect -112 -31174 -106 -29198
rect -152 -31186 -106 -31174
rect 106 -29198 152 -29186
rect 106 -31174 112 -29198
rect 146 -31174 152 -29198
rect 106 -31186 152 -31174
rect -96 -31233 96 -31227
rect -96 -31267 -84 -31233
rect 84 -31267 96 -31233
rect -96 -31273 96 -31267
rect -96 -31341 96 -31335
rect -96 -31375 -84 -31341
rect 84 -31375 96 -31341
rect -96 -31381 96 -31375
rect -152 -31434 -106 -31422
rect -152 -33410 -146 -31434
rect -112 -33410 -106 -31434
rect -152 -33422 -106 -33410
rect 106 -31434 152 -31422
rect 106 -33410 112 -31434
rect 146 -33410 152 -31434
rect 106 -33422 152 -33410
rect -96 -33469 96 -33463
rect -96 -33503 -84 -33469
rect 84 -33503 96 -33469
rect -96 -33509 96 -33503
rect -96 -33577 96 -33571
rect -96 -33611 -84 -33577
rect 84 -33611 96 -33577
rect -96 -33617 96 -33611
rect -152 -33670 -106 -33658
rect -152 -35646 -146 -33670
rect -112 -35646 -106 -33670
rect -152 -35658 -106 -35646
rect 106 -33670 152 -33658
rect 106 -35646 112 -33670
rect 146 -35646 152 -33670
rect 106 -35658 152 -35646
rect -96 -35705 96 -35699
rect -96 -35739 -84 -35705
rect 84 -35739 96 -35705
rect -96 -35745 96 -35739
rect -96 -35813 96 -35807
rect -96 -35847 -84 -35813
rect 84 -35847 96 -35813
rect -96 -35853 96 -35847
rect -152 -35906 -106 -35894
rect -152 -37882 -146 -35906
rect -112 -37882 -106 -35906
rect -152 -37894 -106 -37882
rect 106 -35906 152 -35894
rect 106 -37882 112 -35906
rect 146 -37882 152 -35906
rect 106 -37894 152 -37882
rect -96 -37941 96 -37935
rect -96 -37975 -84 -37941
rect 84 -37975 96 -37941
rect -96 -37981 96 -37975
rect -96 -38049 96 -38043
rect -96 -38083 -84 -38049
rect 84 -38083 96 -38049
rect -96 -38089 96 -38083
rect -152 -38142 -106 -38130
rect -152 -40118 -146 -38142
rect -112 -40118 -106 -38142
rect -152 -40130 -106 -40118
rect 106 -38142 152 -38130
rect 106 -40118 112 -38142
rect 146 -40118 152 -38142
rect 106 -40130 152 -40118
rect -96 -40177 96 -40171
rect -96 -40211 -84 -40177
rect 84 -40211 96 -40177
rect -96 -40217 96 -40211
<< properties >>
string FIXED_BBOX -243 -40296 243 40296
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 1 m 36 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
