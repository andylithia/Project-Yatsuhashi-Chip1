magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< pwell >>
rect -26 -26 392 362
<< scnmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
<< ndiff >>
rect 0 0 60 336
rect 90 0 168 336
rect 198 0 276 336
rect 306 0 366 336
<< poly >>
rect 60 362 306 392
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
<< locali >>
rect 112 235 358 269
rect 8 135 42 201
rect 112 168 146 235
rect 220 135 254 201
rect 324 168 358 235
use sky130_sram_1r1w_24x128_8_contact_10  sky130_sram_1r1w_24x128_8_contact_10_0
timestamp 1661296025
transform 1 0 316 0 1 135
box -26 -22 76 88
use sky130_sram_1r1w_24x128_8_contact_10  sky130_sram_1r1w_24x128_8_contact_10_1
timestamp 1661296025
transform 1 0 212 0 1 135
box -26 -22 76 88
use sky130_sram_1r1w_24x128_8_contact_10  sky130_sram_1r1w_24x128_8_contact_10_2
timestamp 1661296025
transform 1 0 104 0 1 135
box -26 -22 76 88
use sky130_sram_1r1w_24x128_8_contact_10  sky130_sram_1r1w_24x128_8_contact_10_3
timestamp 1661296025
transform 1 0 0 0 1 135
box -26 -22 76 88
<< labels >>
rlabel poly s 183 377 183 377 4 G
port 1 nsew
rlabel locali s 237 168 237 168 4 S
port 2 nsew
rlabel locali s 25 168 25 168 4 S
port 2 nsew
rlabel locali s 235 252 235 252 4 D
port 3 nsew
<< properties >>
string FIXED_BBOX -25 -26 391 392
<< end >>
