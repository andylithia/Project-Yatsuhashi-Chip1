magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< locali >>
rect 3470 8467 5718 8501
rect 5718 7053 10430 7087
rect 3817 6790 4036 6824
rect 4002 6308 4036 6790
rect 3470 5639 6598 5673
rect 4864 4225 10430 4259
rect 3470 2811 5232 2845
rect 3799 2541 3984 2575
rect 3799 2176 3833 2541
rect 3666 2142 3833 2176
rect 5232 1397 10430 1431
rect 3470 -17 10430 17
<< metal1 >>
rect 3438 8458 3502 8510
rect 2980 7800 3551 7828
rect 4870 7751 4934 7803
rect 10398 7044 10462 7096
rect 5964 6337 6028 6389
rect 2896 6160 3699 6188
rect 3064 5912 3599 5940
rect 3438 5630 3502 5682
rect 2896 5372 3566 5400
rect 2980 5248 3699 5276
rect 3316 5124 3832 5152
rect 4762 4923 4826 4975
rect 1553 4308 2896 4336
rect 10398 4216 10462 4268
rect 383 4148 3148 4176
rect 4338 3493 4402 3545
rect 3316 3332 3699 3360
rect 3148 3084 3599 3112
rect 3438 2802 3502 2854
rect 4035 2284 4099 2336
rect 3148 2145 3551 2173
rect 4706 2111 4770 2163
rect 10398 1388 10462 1440
rect 3519 643 3583 695
rect 8608 681 8672 733
rect 3438 -26 3502 26
<< metal2 >>
rect -57 17699 -29 17727
rect 1539 4322 1567 6401
rect 369 1414 397 4162
rect 1844 861 1900 909
rect 137 538 203 590
rect 2350 479 2406 527
rect 2798 0 2826 8524
rect 2882 0 2910 8524
rect 2966 0 2994 8524
rect 3050 0 3078 8524
rect 3134 0 3162 8524
rect 3218 0 3246 8524
rect 3302 0 3330 8524
rect 3442 8460 3498 8508
rect 4902 7763 10514 7791
rect 10402 7046 10458 7094
rect 5996 6349 10514 6377
rect 3442 5632 3498 5680
rect 4794 4935 10514 4963
rect 10402 4218 10458 4266
rect 4342 3495 4398 3543
rect 3442 2804 3498 2852
rect 4039 2286 4095 2334
rect 4724 1713 4752 2137
rect 10402 1390 10458 1438
rect 8640 707 10514 721
rect 8626 693 10514 707
rect 3537 655 3565 683
rect 8626 283 8654 693
rect 3442 -24 3498 24
<< metal3 >>
rect 3395 8452 3545 8516
rect 10355 7038 10505 7102
rect 3395 5624 3545 5688
rect 10355 4210 10505 4274
rect 3064 3489 4370 3549
rect 3395 2796 3545 2860
rect 3316 2280 4067 2340
rect 2980 1683 4738 1743
rect 1228 1365 1326 1463
rect 10355 1382 10505 1446
rect 1872 855 3316 915
rect 2378 473 3232 533
rect 3148 253 8640 313
rect 1228 -49 1326 49
rect 3395 -32 3545 32
<< metal4 >>
rect 335 5606 401 18415
rect 1439 5623 1505 18432
rect 3437 -33 3503 8517
rect 10397 1381 10463 7103
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 3441 0 1 8451
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 10401 0 1 7037
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_2
timestamp 1661296025
transform 1 0 3441 0 1 5623
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_3
timestamp 1661296025
transform 1 0 10401 0 1 7037
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_4
timestamp 1661296025
transform 1 0 3441 0 1 5623
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_5
timestamp 1661296025
transform 1 0 10401 0 1 4209
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_6
timestamp 1661296025
transform 1 0 3441 0 1 2795
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_7
timestamp 1661296025
transform 1 0 10401 0 1 4209
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_8
timestamp 1661296025
transform 1 0 3441 0 1 2795
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_9
timestamp 1661296025
transform 1 0 10401 0 1 1381
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_10
timestamp 1661296025
transform 1 0 3441 0 1 -33
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_11
timestamp 1661296025
transform 1 0 10401 0 1 1381
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_12
timestamp 1661296025
transform 1 0 4341 0 1 3486
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_13
timestamp 1661296025
transform 1 0 4341 0 1 3486
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_14
timestamp 1661296025
transform 1 0 3670 0 1 3313
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_15
timestamp 1661296025
transform 1 0 3570 0 1 3065
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_16
timestamp 1661296025
transform 1 0 4709 0 1 2104
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_17
timestamp 1661296025
transform 1 0 4038 0 1 2277
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_18
timestamp 1661296025
transform 1 0 4038 0 1 2277
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_19
timestamp 1661296025
transform 1 0 3522 0 1 2126
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_20
timestamp 1661296025
transform 1 0 8611 0 1 674
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_21
timestamp 1661296025
transform 1 0 8611 0 1 674
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_22
timestamp 1661296025
transform 1 0 3522 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_23
timestamp 1661296025
transform 1 0 5967 0 1 6330
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_24
timestamp 1661296025
transform 1 0 3670 0 1 6141
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_25
timestamp 1661296025
transform 1 0 3570 0 1 5893
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_26
timestamp 1661296025
transform 1 0 4765 0 1 4916
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_27
timestamp 1661296025
transform 1 0 3803 0 1 5105
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_28
timestamp 1661296025
transform 1 0 3670 0 1 5229
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_29
timestamp 1661296025
transform 1 0 3537 0 1 5353
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_30
timestamp 1661296025
transform 1 0 4873 0 1 7744
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_31
timestamp 1661296025
transform 1 0 3522 0 1 7781
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_0
timestamp 1661296025
transform 1 0 3438 0 1 8452
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_1
timestamp 1661296025
transform 1 0 10398 0 1 7038
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_2
timestamp 1661296025
transform 1 0 3438 0 1 5624
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_3
timestamp 1661296025
transform 1 0 10398 0 1 7038
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_4
timestamp 1661296025
transform 1 0 3438 0 1 5624
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_5
timestamp 1661296025
transform 1 0 10398 0 1 4210
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_6
timestamp 1661296025
transform 1 0 3438 0 1 2796
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_7
timestamp 1661296025
transform 1 0 10398 0 1 4210
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_8
timestamp 1661296025
transform 1 0 3438 0 1 2796
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_9
timestamp 1661296025
transform 1 0 10398 0 1 1382
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_10
timestamp 1661296025
transform 1 0 3438 0 1 -32
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_11
timestamp 1661296025
transform 1 0 10398 0 1 1382
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_12
timestamp 1661296025
transform 1 0 4338 0 1 3487
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_13
timestamp 1661296025
transform 1 0 4338 0 1 3487
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_14
timestamp 1661296025
transform 1 0 3284 0 1 3314
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_15
timestamp 1661296025
transform 1 0 3116 0 1 3066
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_16
timestamp 1661296025
transform 1 0 4706 0 1 2105
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_17
timestamp 1661296025
transform 1 0 4035 0 1 2278
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_18
timestamp 1661296025
transform 1 0 4035 0 1 2278
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_19
timestamp 1661296025
transform 1 0 3116 0 1 2127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_20
timestamp 1661296025
transform 1 0 8608 0 1 675
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_21
timestamp 1661296025
transform 1 0 8608 0 1 675
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_22
timestamp 1661296025
transform 1 0 3519 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_23
timestamp 1661296025
transform 1 0 5964 0 1 6331
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_24
timestamp 1661296025
transform 1 0 2864 0 1 6142
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_25
timestamp 1661296025
transform 1 0 3032 0 1 5894
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_26
timestamp 1661296025
transform 1 0 2864 0 1 4290
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_27
timestamp 1661296025
transform 1 0 1521 0 1 4290
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_28
timestamp 1661296025
transform 1 0 4762 0 1 4917
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_29
timestamp 1661296025
transform 1 0 3284 0 1 5106
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_30
timestamp 1661296025
transform 1 0 2948 0 1 5230
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_31
timestamp 1661296025
transform 1 0 2864 0 1 5354
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_32
timestamp 1661296025
transform 1 0 4870 0 1 7745
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_33
timestamp 1661296025
transform 1 0 2948 0 1 7782
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_34
timestamp 1661296025
transform 1 0 3116 0 1 4130
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_35
timestamp 1661296025
transform 1 0 351 0 1 4130
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_0
timestamp 1661296025
transform 1 0 3437 0 1 8447
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_1
timestamp 1661296025
transform 1 0 10397 0 1 7033
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_2
timestamp 1661296025
transform 1 0 3437 0 1 5619
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_3
timestamp 1661296025
transform 1 0 10397 0 1 7033
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_4
timestamp 1661296025
transform 1 0 3437 0 1 5619
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_5
timestamp 1661296025
transform 1 0 10397 0 1 4205
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_6
timestamp 1661296025
transform 1 0 3437 0 1 2791
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_7
timestamp 1661296025
transform 1 0 10397 0 1 4205
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_8
timestamp 1661296025
transform 1 0 3437 0 1 2791
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_9
timestamp 1661296025
transform 1 0 10397 0 1 1377
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_10
timestamp 1661296025
transform 1 0 3437 0 1 -37
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_11
timestamp 1661296025
transform 1 0 10397 0 1 1377
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_12
timestamp 1661296025
transform 1 0 4337 0 1 3482
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_13
timestamp 1661296025
transform 1 0 4034 0 1 2273
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_14
timestamp 1661296025
transform 1 0 4034 0 1 2273
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_15
timestamp 1661296025
transform 1 0 2345 0 1 466
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_16
timestamp 1661296025
transform 1 0 1839 0 1 848
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_0
timestamp 1661296025
transform 1 0 3432 0 1 8451
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_1
timestamp 1661296025
transform 1 0 10392 0 1 7037
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_2
timestamp 1661296025
transform 1 0 3432 0 1 5623
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_3
timestamp 1661296025
transform 1 0 10392 0 1 7037
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_4
timestamp 1661296025
transform 1 0 3432 0 1 5623
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_5
timestamp 1661296025
transform 1 0 10392 0 1 4209
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_6
timestamp 1661296025
transform 1 0 3432 0 1 2795
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_7
timestamp 1661296025
transform 1 0 10392 0 1 4209
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_8
timestamp 1661296025
transform 1 0 3432 0 1 2795
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_9
timestamp 1661296025
transform 1 0 10392 0 1 1381
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_10
timestamp 1661296025
transform 1 0 3432 0 1 -33
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_11
timestamp 1661296025
transform 1 0 10392 0 1 1381
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_0
timestamp 1661296025
transform 1 0 3031 0 1 3482
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_1
timestamp 1661296025
transform 1 0 2947 0 1 1676
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_2
timestamp 1661296025
transform 1 0 4705 0 1 1676
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_3
timestamp 1661296025
transform 1 0 3283 0 1 2273
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_4
timestamp 1661296025
transform 1 0 3115 0 1 246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_5
timestamp 1661296025
transform 1 0 8607 0 1 246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_6
timestamp 1661296025
transform 1 0 3199 0 1 466
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_32  sky130_sram_1r1w_24x128_8_contact_32_7
timestamp 1661296025
transform 1 0 3283 0 1 848
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_delay_chain  sky130_sram_1r1w_24x128_8_delay_chain_0
timestamp 1661296025
transform 1 0 0 0 -1 18382
box -75 -50 1876 12783
use sky130_sram_1r1w_24x128_8_dff_buf_array  sky130_sram_1r1w_24x128_8_dff_buf_array_0
timestamp 1661296025
transform 1 0 0 0 1 0
box -36 -49 2590 1471
use sky130_sram_1r1w_24x128_8_pand2  sky130_sram_1r1w_24x128_8_pand2_0
timestamp 1661296025
transform 1 0 3470 0 1 2828
box -36 -17 1430 1471
use sky130_sram_1r1w_24x128_8_pand2  sky130_sram_1r1w_24x128_8_pand2_1
timestamp 1661296025
transform 1 0 3838 0 -1 2828
box -36 -17 1430 1471
use sky130_sram_1r1w_24x128_8_pand3_0  sky130_sram_1r1w_24x128_8_pand3_0_0
timestamp 1661296025
transform 1 0 3470 0 -1 5656
box -36 -17 2178 1471
use sky130_sram_1r1w_24x128_8_pdriver_0  sky130_sram_1r1w_24x128_8_pdriver_0_0
timestamp 1661296025
transform 1 0 3470 0 1 0
box -36 -17 6996 1471
use sky130_sram_1r1w_24x128_8_pdriver_1  sky130_sram_1r1w_24x128_8_pdriver_1_0
timestamp 1661296025
transform 1 0 3470 0 -1 8484
box -36 -17 2284 1471
use sky130_sram_1r1w_24x128_8_pdriver_4  sky130_sram_1r1w_24x128_8_pdriver_4_0
timestamp 1661296025
transform 1 0 3938 0 1 5656
box -36 -17 2696 1471
use sky130_sram_1r1w_24x128_8_pinv  sky130_sram_1r1w_24x128_8_pinv_0
timestamp 1661296025
transform 1 0 3470 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pnand2_0  sky130_sram_1r1w_24x128_8_pnand2_0_0
timestamp 1661296025
transform 1 0 3470 0 1 5656
box -36 -17 504 1471
<< labels >>
rlabel metal2 s 137 538 203 590 4 csb
port 1 nsew
rlabel metal2 s 4902 7763 10514 7791 4 wl_en
port 2 nsew
rlabel metal2 s 4794 4935 10514 4963 4 s_en
port 3 nsew
rlabel metal2 s -57 17699 -29 17727 4 rbl_bl
port 4 nsew
rlabel metal2 s 5996 6349 10514 6377 4 p_en_bar
port 5 nsew
rlabel metal2 s 3537 655 3565 683 4 clk
port 6 nsew
rlabel metal2 s 8640 693 10514 721 4 clk_buf
port 7 nsew
rlabel metal3 s 1228 1365 1326 1463 4 vdd
port 8 nsew
rlabel metal4 s 10397 1381 10463 7103 4 vdd
port 8 nsew
rlabel metal4 s 335 5606 401 18415 4 vdd
port 8 nsew
rlabel metal4 s 1439 5623 1505 18432 4 gnd
port 9 nsew
rlabel metal4 s 3437 -33 3503 8517 4 gnd
port 9 nsew
rlabel metal3 s 1228 -49 1326 49 4 gnd
port 9 nsew
<< properties >>
string FIXED_BBOX 0 0 10514 18542
<< end >>
