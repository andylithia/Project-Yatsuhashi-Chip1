magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< error_p >>
rect 79 421 91 424
rect 38 420 91 421
rect 101 420 113 424
rect 151 420 163 424
rect 173 420 185 424
rect 38 412 80 420
rect 38 395 113 412
rect 114 400 125 412
rect 139 400 150 412
rect 42 378 76 395
rect 79 378 113 395
rect 42 299 46 333
rect 72 299 76 333
rect -25 262 25 264
rect 0 254 14 255
rect 0 253 17 254
rect 25 253 27 262
rect 0 246 38 253
rect 0 245 34 246
rect 0 229 8 245
rect 14 229 34 245
rect 0 228 34 229
rect 0 221 38 228
rect 14 220 17 221
rect 25 212 27 221
rect 42 192 45 282
rect 71 251 80 279
rect 69 213 80 251
rect 107 207 119 241
rect 129 213 143 241
rect 129 207 141 213
rect 42 141 46 175
rect 72 141 76 175
rect 42 94 76 98
rect 42 64 46 94
rect 72 64 76 94
rect 16 55 38 61
rect 80 55 102 61
rect 144 55 148 395
rect 151 378 156 412
rect 180 381 185 412
rect 186 400 197 412
rect 400 395 442 421
rect 174 373 246 381
rect 256 373 328 381
rect 332 379 336 395
rect 400 387 438 395
rect 400 380 408 387
rect 434 380 438 387
rect 388 379 454 380
rect 224 343 226 359
rect 196 335 226 343
rect 196 331 230 335
rect 196 301 204 331
rect 216 301 230 331
rect 224 254 226 301
rect 300 274 308 343
rect 332 341 342 379
rect 400 371 404 379
rect 454 365 504 367
rect 494 361 548 365
rect 494 356 514 361
rect 504 341 506 356
rect 336 329 342 341
rect 289 264 308 274
rect 300 258 308 264
rect 332 295 342 329
rect 400 333 404 341
rect 400 299 408 333
rect 434 299 438 333
rect 498 331 506 341
rect 514 331 515 351
rect 504 315 506 331
rect 525 322 528 356
rect 547 331 548 351
rect 557 331 564 341
rect 514 315 530 321
rect 532 315 548 321
rect 332 267 373 295
rect 332 261 351 267
rect 196 220 204 254
rect 216 220 230 254
rect 244 220 257 254
rect 278 224 291 258
rect 300 242 321 258
rect 336 251 351 261
rect 300 240 312 242
rect 300 224 321 240
rect 332 233 351 251
rect 361 233 375 267
rect 400 261 411 299
rect 562 262 612 264
rect 400 233 409 261
rect 466 253 497 255
rect 565 253 596 255
rect 442 246 500 253
rect 466 245 500 246
rect 565 245 599 253
rect 174 183 181 207
rect 224 173 226 220
rect 300 211 308 224
rect 289 208 305 210
rect 332 183 342 233
rect 400 213 404 233
rect 497 229 500 245
rect 596 229 599 245
rect 466 228 500 229
rect 442 221 500 228
rect 565 221 599 229
rect 612 212 614 262
rect 256 173 328 181
rect 336 175 342 183
rect 400 175 404 183
rect 196 143 204 173
rect 216 143 230 173
rect 196 139 230 143
rect 196 131 226 139
rect 224 115 226 131
rect 332 103 336 171
rect 400 141 408 175
rect 434 141 438 175
rect 454 159 504 161
rect 504 143 506 159
rect 514 153 530 159
rect 532 153 548 159
rect 525 143 548 152
rect 400 133 404 141
rect 498 133 506 143
rect 504 109 506 133
rect 514 123 515 143
rect 525 118 528 143
rect 547 123 548 143
rect 557 133 564 143
rect 514 109 548 113
rect 400 103 442 104
rect 174 93 246 101
rect 400 96 404 103
rect 295 62 300 96
rect 324 62 329 96
rect 367 62 438 96
rect 400 61 404 62
rect 378 55 404 61
rect 442 55 464 61
rect 38 39 80 55
rect 400 39 442 55
rect -25 25 25 27
rect 455 25 505 27
rect 557 25 607 27
rect 16 17 102 25
rect 378 17 464 25
rect 8 -17 17 17
rect 18 15 51 17
rect 80 15 100 17
rect 18 -17 100 15
rect 380 15 404 17
rect 429 15 438 17
rect 442 15 462 17
rect 16 -25 102 -17
rect 42 -41 76 -39
rect 16 -61 38 -55
rect 80 -61 102 -55
rect 144 -79 148 0
rect 332 -55 336 0
rect 380 -17 462 15
rect 463 -17 472 17
rect 480 -17 497 17
rect 378 -25 464 -17
rect 505 -25 507 25
rect 514 -17 548 17
rect 565 -17 582 17
rect 607 -25 609 25
rect 404 -41 438 -39
rect 378 -61 404 -55
rect 442 -61 464 -55
rect 400 -79 404 -61
rect 38 -105 80 -79
rect 400 -105 442 -79
<< nwell >>
rect 144 -79 336 395
<< pwell >>
rect 12 279 106 421
rect -26 195 106 279
rect 12 -105 106 195
rect 374 279 468 421
rect 374 195 650 279
rect 374 -105 468 195
<< npd >>
rect 38 341 80 371
rect 38 261 80 291
rect 38 183 80 213
rect 400 341 442 371
rect 400 261 442 291
rect 400 183 442 213
rect 38 103 80 133
rect 400 103 442 133
rect 38 39 80 55
rect 400 39 442 55
rect 38 -55 80 -39
rect 400 -55 442 -39
<< ppu >>
rect 196 343 224 359
rect 196 263 224 293
rect 196 181 224 211
rect 196 115 224 131
<< sramnvar >>
rect 278 343 306 359
rect 278 195 306 211
<< srampvar >>
rect 38 25 80 39
rect 400 25 442 39
rect 38 -39 80 -25
rect 400 -39 442 -25
<< ndiff >>
rect 38 378 42 395
rect 76 378 80 395
rect 38 371 80 378
rect 400 380 404 395
rect 438 380 442 395
rect 400 371 442 380
rect 38 333 80 341
rect 38 299 42 333
rect 76 299 80 333
rect 38 291 80 299
rect 38 253 80 261
rect 14 221 80 253
rect 38 213 80 221
rect 400 333 442 341
rect 400 299 404 333
rect 438 299 442 333
rect 400 291 442 299
rect 400 253 442 261
rect 400 221 466 253
rect 497 221 565 253
rect 596 221 624 253
rect 400 213 442 221
rect 38 175 80 183
rect 38 141 42 175
rect 76 141 80 175
rect 38 133 80 141
rect 400 175 442 183
rect 400 141 404 175
rect 438 141 442 175
rect 400 133 442 141
rect 38 94 80 103
rect 38 64 42 94
rect 76 64 80 94
rect 38 55 80 64
rect 400 96 442 103
rect 400 62 404 96
rect 438 62 442 96
rect 400 55 442 62
rect 38 -79 80 -55
rect 400 -79 442 -55
<< pdiff >>
rect 196 335 224 343
rect 196 293 224 301
rect 196 254 224 263
rect 196 211 224 220
rect 196 173 224 181
rect 196 131 224 139
<< ndiffc >>
rect 42 378 76 395
rect 404 380 438 395
rect 42 299 76 333
rect 0 221 14 253
rect 404 299 438 333
rect 466 221 497 253
rect 565 221 596 253
rect 42 141 76 175
rect 404 141 438 175
rect 42 64 76 94
rect 404 62 438 96
<< pdiffc >>
rect 196 301 224 335
rect 196 220 224 254
rect 196 139 224 173
<< psubdiff >>
rect 38 17 80 25
rect 38 -17 42 17
rect 76 -17 80 17
rect 38 -25 80 -17
rect 400 17 442 25
rect 400 -17 404 17
rect 438 -17 442 17
rect 400 -25 442 -17
<< nsubdiff >>
rect 278 258 306 343
rect 305 224 306 258
rect 278 211 306 224
<< psubdiffcont >>
rect 42 -17 76 17
rect 404 -17 438 17
<< nsubdiffcont >>
rect 278 224 305 258
<< poly >>
rect 127 371 353 373
rect 0 341 38 371
rect 80 359 400 371
rect 80 343 196 359
rect 224 343 278 359
rect 306 343 400 359
rect 80 341 138 343
rect 128 291 196 293
rect 16 261 38 291
rect 80 263 196 291
rect 224 263 256 293
rect 80 261 139 263
rect 109 241 139 261
rect 16 183 38 213
rect 80 207 107 213
rect 342 341 400 343
rect 442 365 624 371
rect 442 341 514 365
rect 505 331 514 341
rect 548 341 624 365
rect 548 331 557 341
rect 505 321 557 331
rect 341 267 400 291
rect 373 261 400 267
rect 442 261 464 291
rect 341 213 371 233
rect 341 211 400 213
rect 80 183 139 207
rect 174 181 196 211
rect 224 195 278 211
rect 306 195 400 211
rect 224 183 400 195
rect 442 183 464 213
rect 224 181 352 183
rect 0 103 38 133
rect 80 131 138 133
rect 505 143 557 153
rect 505 133 514 143
rect 342 131 400 133
rect 80 115 196 131
rect 224 115 400 131
rect 80 103 400 115
rect 442 109 514 133
rect 548 133 557 143
rect 548 109 624 133
rect 442 103 624 109
rect 127 101 353 103
rect 127 55 353 57
rect 0 25 38 55
rect 80 27 400 55
rect 80 25 138 27
rect 342 25 400 27
rect 442 25 624 55
rect 505 17 557 25
rect 505 -17 514 17
rect 548 -17 557 17
rect 505 -25 557 -17
rect 0 -55 38 -25
rect 80 -27 138 -25
rect 342 -27 400 -25
rect 80 -55 400 -27
rect 442 -55 624 -25
rect 127 -57 353 -55
<< polycont >>
rect 109 213 139 241
rect 107 207 139 213
rect 514 331 548 365
rect 341 261 373 267
rect 341 233 371 261
rect 514 109 548 143
rect 514 -17 548 17
<< corelocali >>
rect 14 412 118 420
rect 14 395 79 412
rect 14 378 42 395
rect 76 378 79 395
rect 113 378 118 412
rect 14 370 118 378
rect 146 412 382 420
rect 146 378 151 412
rect 185 410 382 412
rect 185 395 466 410
rect 185 380 404 395
rect 438 380 466 395
rect 185 378 382 380
rect 146 370 382 378
rect 494 365 568 377
rect 494 356 514 365
rect 14 335 373 336
rect 14 333 196 335
rect 14 301 42 333
rect 76 301 196 333
rect 224 301 373 335
rect 76 300 373 301
rect -14 254 14 273
rect -14 122 14 220
rect 42 175 76 299
rect 339 267 373 300
rect 42 122 76 141
rect 107 241 141 261
rect 107 213 109 241
rect 139 207 141 241
rect 172 258 308 264
rect 172 254 278 258
rect 172 220 196 254
rect 257 224 278 254
rect 305 224 308 258
rect 257 220 308 224
rect 172 210 308 220
rect 339 233 341 267
rect 371 233 373 261
rect 339 213 373 233
rect 404 333 438 352
rect 548 331 568 365
rect 528 322 568 331
rect 494 314 568 322
rect 107 174 141 207
rect 404 175 438 299
rect 466 254 596 270
rect 466 253 569 254
rect 497 221 565 253
rect 466 220 569 221
rect 466 204 596 220
rect 107 173 404 174
rect 107 139 196 173
rect 224 141 404 173
rect 438 141 466 173
rect 224 139 466 141
rect 107 138 466 139
rect 494 152 568 160
rect 528 143 568 152
rect 494 109 514 118
rect 548 109 568 143
rect 98 96 334 104
rect 98 94 295 96
rect 14 64 42 94
rect 76 64 295 94
rect 98 62 295 64
rect 329 62 334 96
rect 98 54 334 62
rect 362 96 466 104
rect 494 97 568 109
rect 362 62 367 96
rect 401 62 404 96
rect 438 62 466 96
rect 362 54 466 62
rect 480 18 582 26
rect -42 17 624 18
rect -42 -17 -17 17
rect 17 -17 42 17
rect 76 -17 404 17
rect 438 -17 463 17
rect 497 -17 514 17
rect 548 -17 565 17
rect 599 -17 624 17
rect -42 -18 624 -17
rect 480 -26 582 -18
<< viali >>
rect 79 378 113 412
rect 151 378 185 412
rect -17 253 17 254
rect -17 221 0 253
rect 0 221 14 253
rect 14 221 17 253
rect -17 220 17 221
rect 223 220 224 254
rect 224 220 257 254
rect 494 331 514 356
rect 514 331 528 356
rect 494 322 528 331
rect 569 253 603 254
rect 569 221 596 253
rect 596 221 603 253
rect 569 220 603 221
rect 494 143 528 152
rect 494 118 514 143
rect 514 118 528 143
rect 295 62 329 96
rect 367 62 401 96
rect -17 -17 17 17
rect 463 -17 497 17
rect 565 -17 599 17
<< metal1 >>
rect -42 262 42 420
rect -42 212 -25 262
rect 25 212 42 262
rect -42 25 42 212
rect -42 -25 -25 25
rect 25 -25 42 25
rect -42 -104 42 -25
rect 78 412 114 420
rect 78 378 79 412
rect 113 378 114 412
rect 78 -104 114 378
rect 150 412 186 420
rect 150 378 151 412
rect 185 378 186 412
rect 150 -104 186 378
rect 222 254 258 420
rect 222 220 223 254
rect 257 220 258 254
rect 222 -104 258 220
rect 294 96 330 420
rect 294 62 295 96
rect 329 62 330 96
rect 294 -104 330 62
rect 366 96 402 420
rect 438 365 531 377
rect 438 315 454 365
rect 504 356 531 365
rect 528 322 531 356
rect 504 315 531 322
rect 438 311 531 315
rect 438 295 515 311
tri 515 295 531 311 nw
rect 567 278 624 420
rect 550 262 624 278
rect 550 212 562 262
rect 612 212 624 262
rect 550 196 624 212
rect 438 163 515 179
tri 515 163 531 179 sw
rect 438 159 531 163
rect 438 109 454 159
rect 504 152 531 159
rect 528 118 531 152
rect 504 109 531 118
rect 438 97 531 109
rect 366 62 367 96
rect 401 62 402 96
rect 366 -104 402 62
rect 567 38 624 196
rect 438 25 624 38
rect 438 -25 455 25
rect 505 -25 557 25
rect 607 -25 624 25
rect 438 -38 624 -25
rect 567 -104 624 -38
<< via1 >>
rect -25 254 25 262
rect -25 220 -17 254
rect -17 220 17 254
rect 17 220 25 254
rect -25 212 25 220
rect -25 17 25 25
rect -25 -17 -17 17
rect -17 -17 17 17
rect 17 -17 25 17
rect -25 -25 25 -17
rect 454 356 504 365
rect 454 322 494 356
rect 494 322 504 356
rect 454 315 504 322
rect 562 254 612 262
rect 562 220 569 254
rect 569 220 603 254
rect 603 220 612 254
rect 562 212 612 220
rect 454 152 504 159
rect 454 118 494 152
rect 494 118 504 152
rect 454 109 504 118
rect 455 17 505 25
rect 455 -17 463 17
rect 463 -17 497 17
rect 497 -17 505 17
rect 455 -25 505 -17
rect 557 17 607 25
rect 557 -17 565 17
rect 565 -17 599 17
rect 599 -17 607 17
rect 557 -25 607 -17
<< metal2 >>
rect -42 365 624 371
rect -42 323 454 365
rect 438 315 454 323
rect 504 323 624 365
rect 504 315 520 323
rect 438 309 520 315
rect -42 262 404 275
rect -42 212 -25 262
rect 25 261 404 262
rect 554 262 624 275
rect 554 261 562 262
rect 25 213 562 261
rect 25 212 404 213
rect -42 199 404 212
rect 554 212 562 213
rect 612 212 624 262
rect 554 199 624 212
rect 438 159 520 165
rect 438 151 454 159
rect -42 109 454 151
rect 504 151 520 159
rect 504 109 624 151
rect -42 103 624 109
rect -42 25 624 55
rect -42 -25 -25 25
rect 25 -25 455 25
rect 505 -25 557 25
rect 607 -25 624 25
rect -42 -55 624 -25
<< labels >>
rlabel comment s 32 142 32 142 4 short li
rlabel comment s 40 159 40 159 4 no mcon
rlabel comment s 32 180 32 180 4 in cell
rlabel comment s 240 169 240 169 4 MAIN CELL
rlabel comment s 241 150 241 150 4 opt.1
rlabel comment s 45 57 45 57 4 short met1
rlabel comment s 43 259 43 259 4 short met1
rlabel comment s 32 174 32 174 4 short li
rlabel comment s 40 157 40 157 4 no mcon
rlabel comment s 32 136 32 136 4 in cell
rlabel comment s 45 57 45 57 4 short met1
rlabel comment s 43 259 43 259 4 short met1
rlabel comment s 32 174 32 174 4 short li
rlabel comment s 40 157 40 157 4 no mcon
rlabel comment s 32 136 32 136 4 in cell
rlabel comment s 45 57 45 57 4 short met1
rlabel comment s 43 259 43 259 4 short met1
rlabel comment s 32 174 32 174 4 short li
rlabel comment s 40 157 40 157 4 no mcon
rlabel comment s 32 136 32 136 4 in cell
rlabel comment s 45 57 45 57 4 short met1
rlabel comment s 43 259 43 259 4 short met1
rlabel comment s 32 174 32 174 4 short li
rlabel comment s 40 157 40 157 4 no mcon
rlabel comment s 32 136 32 136 4 in cell
rlabel metal2 s 186 199 294 275 4 GND
port 1 nsew
rlabel metal2 s 186 -55 294 55 4 GND
port 1 nsew
rlabel metal2 s 0 323 480 371 4 WL0
port 2 nsew
rlabel metal2 s 0 103 480 151 4 WL1
port 3 nsew
rlabel metal1 s 222 79 258 420 4 VDD
port 4 nsew
rlabel metal1 s 78 79 114 420 4 BL0
port 5 nsew
rlabel metal1 s 294 79 330 420 4 BL1
port 6 nsew
rlabel metal1 s 150 79 186 420 4 BR0
port 7 nsew
rlabel metal1 s 366 79 402 420 4 BR1
port 8 nsew
rlabel metal1 s 96 249 96 249 4 bl0
port 9 nsew
rlabel metal1 s 168 249 168 249 4 br0
port 10 nsew
rlabel metal1 s 312 249 312 249 4 bl1
port 11 nsew
rlabel metal1 s 384 249 384 249 4 br1
port 12 nsew
rlabel metal2 s 240 347 240 347 4 wl0
port 13 nsew
rlabel metal2 s 240 127 240 127 4 wl1
port 14 nsew
rlabel metal1 s 240 249 240 249 4 vdd
port 15 nsew
rlabel metal2 s 240 237 240 237 4 gnd
port 16 nsew
rlabel metal2 s 240 0 240 0 4 gnd
port 16 nsew
<< properties >>
string FIXED_BBOX 0 0 624 395
<< end >>
