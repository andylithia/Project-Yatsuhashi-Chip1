magic
tech sky130B
magscale 1 2
timestamp 1659923234
<< error_p >>
rect -23 1357 23 1369
rect -23 1317 -17 1357
rect -23 1305 23 1317
rect -23 583 23 595
rect -23 543 -17 583
rect -23 531 23 543
rect -23 407 23 419
rect -23 367 -17 407
rect -23 355 23 367
rect -23 -367 23 -355
rect -23 -407 -17 -367
rect -23 -419 23 -407
rect -23 -543 23 -531
rect -23 -583 -17 -543
rect -23 -595 23 -583
rect -23 -1317 23 -1305
rect -23 -1357 -17 -1317
rect -23 -1369 23 -1357
<< pwell >>
rect -199 -1539 199 1539
<< psubdiff >>
rect -163 1469 -67 1503
rect 67 1469 163 1503
rect -163 1407 -129 1469
rect 129 1407 163 1469
rect -163 -1469 -129 -1407
rect 129 -1469 163 -1407
rect -163 -1503 -67 -1469
rect 67 -1503 163 -1469
<< psubdiffcont >>
rect -67 1469 67 1503
rect -163 -1407 -129 1407
rect 129 -1407 163 1407
rect -67 -1503 67 -1469
<< poly >>
rect -33 1357 33 1373
rect -33 1323 -17 1357
rect 17 1323 33 1357
rect -33 1300 33 1323
rect -33 577 33 600
rect -33 543 -17 577
rect 17 543 33 577
rect -33 527 33 543
rect -33 407 33 423
rect -33 373 -17 407
rect 17 373 33 407
rect -33 350 33 373
rect -33 -373 33 -350
rect -33 -407 -17 -373
rect 17 -407 33 -373
rect -33 -423 33 -407
rect -33 -543 33 -527
rect -33 -577 -17 -543
rect 17 -577 33 -543
rect -33 -600 33 -577
rect -33 -1323 33 -1300
rect -33 -1357 -17 -1323
rect 17 -1357 33 -1323
rect -33 -1373 33 -1357
<< polycont >>
rect -17 1323 17 1357
rect -17 543 17 577
rect -17 373 17 407
rect -17 -407 17 -373
rect -17 -577 17 -543
rect -17 -1357 17 -1323
<< npolyres >>
rect -33 600 33 1300
rect -33 -350 33 350
rect -33 -1300 33 -600
<< locali >>
rect -163 1469 -67 1503
rect 67 1469 163 1503
rect -163 1407 -129 1469
rect 129 1407 163 1469
rect -33 1323 -17 1357
rect 17 1323 33 1357
rect -33 543 -17 577
rect 17 543 33 577
rect -33 373 -17 407
rect 17 373 33 407
rect -33 -407 -17 -373
rect 17 -407 33 -373
rect -33 -577 -17 -543
rect 17 -577 33 -543
rect -33 -1357 -17 -1323
rect 17 -1357 33 -1323
rect -163 -1469 -129 -1407
rect 129 -1469 163 -1407
rect -163 -1503 -67 -1469
rect 67 -1503 163 -1469
<< viali >>
rect -17 1323 17 1357
rect -17 1317 17 1323
rect -17 577 17 583
rect -17 543 17 577
rect -17 373 17 407
rect -17 367 17 373
rect -17 -373 17 -367
rect -17 -407 17 -373
rect -17 -577 17 -543
rect -17 -583 17 -577
rect -17 -1323 17 -1317
rect -17 -1357 17 -1323
<< metal1 >>
rect -23 1357 23 1369
rect -23 1317 -17 1357
rect 17 1317 23 1357
rect -23 1305 23 1317
rect -23 583 23 595
rect -23 543 -17 583
rect 17 543 23 583
rect -23 531 23 543
rect -23 407 23 419
rect -23 367 -17 407
rect 17 367 23 407
rect -23 355 23 367
rect -23 -367 23 -355
rect -23 -407 -17 -367
rect 17 -407 23 -367
rect -23 -419 23 -407
rect -23 -543 23 -531
rect -23 -583 -17 -543
rect 17 -583 23 -543
rect -23 -595 23 -583
rect -23 -1317 23 -1305
rect -23 -1357 -17 -1317
rect 17 -1357 23 -1317
rect -23 -1369 23 -1357
<< properties >>
string FIXED_BBOX -146 -1486 146 1486
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.33 l 3.5 m 3 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 511.212 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 1 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
