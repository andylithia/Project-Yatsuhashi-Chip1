magic
tech sky130B
magscale 1 2
timestamp 1661649517
<< metal4 >>
rect -6300 -11576 -2300 -11464
rect -6300 -15352 -6188 -11576
rect -2412 -15352 -2300 -11576
tri -7958 -18529 -6300 -16871 se
rect -6300 -18529 -2300 -15352
tri -10900 -21471 -7958 -18529 se
rect -7958 -21471 -6900 -18529
rect -10900 -24648 -6900 -21471
tri -6900 -23129 -2300 -18529 nw
rect -10900 -28424 -10788 -24648
rect -7012 -28424 -6900 -24648
rect -10900 -28536 -6900 -28424
<< via4 >>
rect -6188 -15352 -2412 -11576
rect -10788 -28424 -7012 -24648
<< metal5 >>
tri -34584 3500 -30584 7500 se
rect -30584 3500 -14016 7500
tri -14016 3500 -10016 7500 sw
tri -38300 -216 -34584 3500 se
rect -34584 2900 -29527 3500
tri -29527 2900 -28927 3500 nw
tri -15673 2900 -15073 3500 ne
rect -15073 2900 -10016 3500
rect -34584 2052 -30375 2900
tri -30375 2052 -29527 2900 nw
tri -29527 2052 -28679 2900 se
rect -28679 2052 -15921 2900
tri -15921 2052 -15073 2900 sw
tri -15073 2052 -14225 2900 ne
rect -14225 2052 -10016 2900
rect -34584 1204 -31223 2052
tri -31223 1204 -30375 2052 nw
tri -30375 1204 -29527 2052 se
rect -29527 1204 -15073 2052
tri -15073 1204 -14225 2052 sw
tri -14225 1204 -13377 2052 ne
rect -13377 1204 -10016 2052
rect -34584 632 -31795 1204
tri -31795 632 -31223 1204 nw
tri -30947 632 -30375 1204 se
rect -30375 632 -14225 1204
tri -14225 632 -13653 1204 sw
tri -13377 632 -12805 1204 ne
rect -12805 632 -10016 1204
rect -34584 -216 -32643 632
tri -32643 -216 -31795 632 nw
tri -31795 -216 -30947 632 se
rect -30947 -216 -13653 632
tri -13653 -216 -12805 632 sw
tri -12805 -216 -11957 632 ne
rect -11957 -216 -10016 632
tri -10016 -216 -6300 3500 sw
tri -40241 -2157 -38300 -216 se
rect -38300 -252 -32679 -216
tri -32679 -252 -32643 -216 nw
tri -31831 -252 -31795 -216 se
rect -31795 -252 -12805 -216
rect -38300 -1100 -33527 -252
tri -33527 -1100 -32679 -252 nw
tri -32679 -1100 -31831 -252 se
rect -31831 -1064 -12805 -252
tri -12805 -1064 -11957 -216 sw
tri -11957 -1064 -11109 -216 ne
rect -11109 -1064 -6300 -216
rect -31831 -1100 -11957 -1064
rect -38300 -1948 -34375 -1100
tri -34375 -1948 -33527 -1100 nw
tri -33527 -1948 -32679 -1100 se
rect -38300 -2157 -34584 -1948
tri -34584 -2157 -34375 -1948 nw
tri -33736 -2157 -33527 -1948 se
rect -33527 -2157 -32679 -1948
tri -42300 -4216 -40241 -2157 se
rect -40241 -3005 -35432 -2157
tri -35432 -3005 -34584 -2157 nw
tri -34584 -3005 -33736 -2157 se
rect -33736 -3005 -32679 -2157
rect -40241 -3853 -36280 -3005
tri -36280 -3853 -35432 -3005 nw
tri -35432 -3853 -34584 -3005 se
rect -34584 -3853 -32679 -3005
rect -40241 -4216 -36852 -3853
rect -42300 -4425 -36852 -4216
tri -36852 -4425 -36280 -3853 nw
tri -36004 -4425 -35432 -3853 se
rect -35432 -4425 -32679 -3853
rect -42300 -5273 -37700 -4425
tri -37700 -5273 -36852 -4425 nw
tri -36852 -5273 -36004 -4425 se
rect -36004 -5273 -32679 -4425
rect -42300 -11464 -38300 -5273
tri -38300 -5873 -37700 -5273 nw
rect -43322 -15464 -38300 -11464
tri -37700 -6121 -36852 -5273 se
rect -36852 -6121 -32679 -5273
rect -37700 -6757 -32679 -6121
tri -32679 -6757 -27022 -1100 nw
tri -17578 -5873 -12805 -1100 ne
rect -12805 -1273 -11957 -1100
tri -11957 -1273 -11748 -1064 sw
tri -11109 -1273 -10900 -1064 ne
rect -10900 -1273 -6300 -1064
rect -12805 -2121 -11748 -1273
tri -11748 -2121 -10900 -1273 sw
tri -10900 -2121 -10052 -1273 ne
rect -10052 -2121 -6300 -1273
rect -12805 -2969 -10900 -2121
tri -10900 -2969 -10052 -2121 sw
tri -10052 -2969 -9204 -2121 ne
rect -9204 -2969 -6300 -2121
rect -12805 -3817 -10052 -2969
tri -10052 -3817 -9204 -2969 sw
tri -9204 -3817 -8356 -2969 ne
rect -8356 -3817 -6300 -2969
rect -12805 -4425 -9204 -3817
tri -9204 -4425 -8596 -3817 sw
tri -8356 -4425 -7748 -3817 ne
rect -7748 -4216 -6300 -3817
tri -6300 -4216 -2300 -216 sw
rect -7748 -4425 -2300 -4216
rect -12805 -5273 -8596 -4425
tri -8596 -5273 -7748 -4425 sw
tri -7748 -5273 -6900 -4425 ne
rect -6900 -5273 -2300 -4425
rect -12805 -5873 -7748 -5273
rect -43322 -28536 -38300 -24536
rect -42300 -34727 -38300 -28536
rect -37700 -33879 -33700 -6757
tri -33700 -7778 -32679 -6757 nw
tri -12805 -7778 -10900 -5873 ne
rect -10900 -6121 -7748 -5873
tri -7748 -6121 -6900 -5273 sw
tri -6900 -5873 -6300 -5273 ne
rect -10900 -18529 -6900 -6121
rect -6300 -11576 -2300 -5273
rect -6300 -15352 -6188 -11576
rect -2412 -15352 -2300 -11576
rect -6300 -15464 -2300 -15352
tri -10900 -22529 -6900 -18529 ne
tri -6900 -21471 -2300 -16871 sw
rect -6900 -22529 -2300 -21471
tri -6900 -23129 -6300 -22529 ne
rect -10900 -24648 -6900 -24536
rect -10900 -28424 -10788 -24648
rect -7012 -28424 -6900 -24648
tri -38300 -34727 -37700 -34127 sw
tri -37700 -34727 -36852 -33879 ne
rect -36852 -34727 -33700 -33879
rect -42300 -35575 -37700 -34727
tri -37700 -35575 -36852 -34727 sw
tri -36852 -35575 -36004 -34727 ne
rect -36004 -35575 -33700 -34727
rect -42300 -35784 -36852 -35575
tri -42300 -39784 -38300 -35784 ne
rect -38300 -36147 -36852 -35784
tri -36852 -36147 -36280 -35575 sw
tri -36004 -36147 -35432 -35575 ne
rect -35432 -36147 -33700 -35575
rect -38300 -36995 -36280 -36147
tri -36280 -36995 -35432 -36147 sw
tri -35432 -36995 -34584 -36147 ne
rect -34584 -36995 -33700 -36147
rect -38300 -37843 -35432 -36995
tri -35432 -37843 -34584 -36995 sw
tri -34584 -37843 -33736 -36995 ne
rect -33736 -37843 -33700 -36995
tri -33700 -37843 -28079 -32222 sw
tri -11921 -33243 -10900 -32222 se
rect -10900 -33243 -6900 -28424
tri -12805 -34127 -11921 -33243 se
rect -11921 -33879 -6900 -33243
rect -11921 -34127 -7748 -33879
rect -38300 -38052 -34584 -37843
tri -34584 -38052 -34375 -37843 sw
tri -33736 -38052 -33527 -37843 ne
rect -33527 -38052 -28079 -37843
rect -38300 -38900 -34375 -38052
tri -34375 -38900 -33527 -38052 sw
tri -33527 -38900 -32679 -38052 ne
rect -32679 -38900 -28079 -38052
tri -28079 -38900 -27022 -37843 sw
tri -16557 -37879 -12805 -34127 se
rect -12805 -34727 -7748 -34127
tri -7748 -34727 -6900 -33879 nw
tri -6900 -34727 -6300 -34127 se
rect -6300 -34727 -2300 -22529
rect -12805 -35575 -8596 -34727
tri -8596 -35575 -7748 -34727 nw
tri -7748 -35575 -6900 -34727 se
rect -6900 -35575 -2300 -34727
rect -12805 -36183 -9204 -35575
tri -9204 -36183 -8596 -35575 nw
tri -8356 -36183 -7748 -35575 se
rect -7748 -35784 -2300 -35575
rect -7748 -36183 -6300 -35784
rect -12805 -37031 -10052 -36183
tri -10052 -37031 -9204 -36183 nw
tri -9204 -37031 -8356 -36183 se
rect -8356 -37031 -6300 -36183
rect -12805 -37879 -10900 -37031
tri -10900 -37879 -10052 -37031 nw
tri -10052 -37879 -9204 -37031 se
rect -9204 -37879 -6300 -37031
tri -17578 -38900 -16557 -37879 se
rect -16557 -38727 -11748 -37879
tri -11748 -38727 -10900 -37879 nw
tri -10900 -38727 -10052 -37879 se
rect -10052 -38727 -6300 -37879
rect -16557 -38900 -11957 -38727
rect -38300 -39748 -33527 -38900
tri -33527 -39748 -32679 -38900 sw
tri -32679 -39748 -31831 -38900 ne
rect -31831 -38936 -11957 -38900
tri -11957 -38936 -11748 -38727 nw
tri -11109 -38936 -10900 -38727 se
rect -10900 -38936 -6300 -38727
rect -31831 -39748 -12805 -38936
rect -38300 -39784 -32679 -39748
tri -32679 -39784 -32643 -39748 sw
tri -31831 -39784 -31795 -39748 ne
rect -31795 -39784 -12805 -39748
tri -12805 -39784 -11957 -38936 nw
tri -11957 -39784 -11109 -38936 se
rect -11109 -39784 -6300 -38936
tri -6300 -39784 -2300 -35784 nw
tri -38300 -43500 -34584 -39784 ne
rect -34584 -40632 -32643 -39784
tri -32643 -40632 -31795 -39784 sw
tri -31795 -40632 -30947 -39784 ne
rect -30947 -40632 -13653 -39784
tri -13653 -40632 -12805 -39784 nw
tri -12805 -40632 -11957 -39784 se
rect -11957 -40632 -10016 -39784
rect -34584 -41204 -31795 -40632
tri -31795 -41204 -31223 -40632 sw
tri -30947 -41204 -30375 -40632 ne
rect -30375 -41204 -14225 -40632
tri -14225 -41204 -13653 -40632 nw
tri -13377 -41204 -12805 -40632 se
rect -12805 -41204 -10016 -40632
rect -34584 -42052 -31223 -41204
tri -31223 -42052 -30375 -41204 sw
tri -30375 -42052 -29527 -41204 ne
rect -29527 -42052 -15073 -41204
tri -15073 -42052 -14225 -41204 nw
tri -14225 -42052 -13377 -41204 se
rect -13377 -42052 -10016 -41204
rect -34584 -42900 -30375 -42052
tri -30375 -42900 -29527 -42052 sw
tri -29527 -42900 -28679 -42052 ne
rect -28679 -42900 -15921 -42052
tri -15921 -42900 -15073 -42052 nw
tri -15073 -42900 -14225 -42052 se
rect -14225 -42900 -10016 -42052
rect -34584 -43500 -29527 -42900
tri -29527 -43500 -28927 -42900 sw
tri -15673 -43500 -15073 -42900 se
rect -15073 -43500 -10016 -42900
tri -10016 -43500 -6300 -39784 nw
tri -34584 -47500 -30584 -43500 ne
rect -30584 -47500 -14016 -43500
tri -14016 -47500 -10016 -43500 nw
<< end >>
