magic
tech sky130A
magscale 1 2
timestamp 1664897280
<< error_p >>
rect 29830 38650 30170 38684
<< error_s >>
rect -3370 38650 -3030 38684
rect 25280 24700 25400 24900
rect 25600 24700 25720 24900
rect 25280 23500 25400 24000
rect 25600 23800 25720 24000
<< pwell >>
rect 29802 38680 30200 40458
rect 30802 25480 31200 27258
rect 30798 12500 31200 14016
<< psubdiff >>
rect 29838 40388 29934 40422
rect 30068 40388 30164 40422
rect 29838 40326 29872 40388
rect 30130 40326 30164 40388
rect 29838 38750 29872 38812
rect 30130 38750 30164 38812
rect 29838 38716 29934 38750
rect 30068 38716 30164 38750
rect 30838 27188 30934 27222
rect 31068 27188 31164 27222
rect 30838 27126 30872 27188
rect 31130 27126 31164 27188
rect 30838 25550 30872 25612
rect 31130 25550 31164 25612
rect 30838 25516 30934 25550
rect 31068 25516 31164 25550
rect 30834 13946 30930 13980
rect 31068 13946 31164 13980
rect 30834 13884 30868 13946
rect 31130 13884 31164 13946
rect 30834 12570 30868 12632
rect 31130 12570 31164 12632
rect 30834 12536 30930 12570
rect 31068 12536 31164 12570
<< psubdiffcont >>
rect 29934 40388 30068 40422
rect 29838 38812 29872 40326
rect 30130 38812 30164 40326
rect 29934 38716 30068 38750
rect 30934 27188 31068 27222
rect 30838 25612 30872 27126
rect 31130 25612 31164 27126
rect 30934 25516 31068 25550
rect 30930 13946 31068 13980
rect 30834 12632 30868 13884
rect 31130 12632 31164 13884
rect 30930 12536 31068 12570
<< poly >>
rect 29968 40276 30034 40292
rect 29968 40242 29984 40276
rect 30018 40242 30034 40276
rect 29968 40219 30034 40242
rect 29968 38896 30034 38919
rect 29968 38862 29984 38896
rect 30018 38862 30034 38896
rect 29968 38846 30034 38862
rect 30968 27076 31034 27092
rect 30968 27042 30984 27076
rect 31018 27042 31034 27076
rect 30968 27019 31034 27042
rect 30968 25696 31034 25719
rect 30968 25662 30984 25696
rect 31018 25662 31034 25696
rect 30968 25646 31034 25662
<< polycont >>
rect 29984 40242 30018 40276
rect 29984 38862 30018 38896
rect 30984 27042 31018 27076
rect 30984 25662 31018 25696
<< xpolycontact >>
rect 30964 13418 31034 13850
rect 30964 12666 31034 13098
<< npolyres >>
rect 29968 38919 30034 40219
rect 30968 25719 31034 27019
<< ppolyres >>
rect 30964 13098 31034 13418
<< locali >>
rect 29838 40388 29934 40422
rect 30068 40388 30164 40422
rect 29838 40326 29872 40388
rect 30130 40326 30164 40388
rect 29968 40242 29984 40276
rect 30018 40242 30034 40276
rect 29968 38862 29984 38896
rect 30018 38862 30034 38896
rect 29838 38750 29872 38812
rect 30130 38750 30164 38812
rect 29838 38716 29934 38750
rect 30068 38716 30164 38750
rect 30838 27188 30934 27222
rect 31068 27188 31164 27222
rect 30838 27126 30872 27188
rect 31130 27126 31164 27188
rect 30968 27042 30984 27076
rect 31018 27042 31034 27076
rect 30968 25662 30984 25696
rect 31018 25662 31034 25696
rect 30838 25550 30872 25612
rect 31130 25550 31164 25612
rect 30838 25516 30934 25550
rect 31068 25516 31164 25550
rect 30834 13946 30930 13980
rect 31068 13946 31164 13980
rect 30834 13884 30868 13946
rect 31130 13884 31164 13946
rect 30834 12570 30868 12632
rect 31130 12570 31164 12632
rect 30834 12536 30930 12570
rect 31068 12536 31164 12570
<< viali >>
rect 29984 40242 30018 40276
rect 29984 40236 30018 40242
rect 29984 38896 30018 38902
rect 29984 38862 30018 38896
rect 30984 27042 31018 27076
rect 30984 27036 31018 27042
rect 30984 25696 31018 25702
rect 30984 25662 31018 25696
rect 30980 13435 31018 13832
rect 30980 12684 31018 13081
<< metal1 >>
rect -3300 40450 -3100 40460
rect -3300 40190 -3290 40450
rect -3110 40190 -3100 40450
rect -3300 40180 -3100 40190
rect 29900 40450 30100 40460
rect 29900 40190 29910 40450
rect 30090 40190 30100 40450
rect 29900 40180 30100 40190
rect -3300 38910 -3100 38920
rect -3300 38690 -3290 38910
rect -3110 38690 -3100 38910
rect -3300 38680 -3100 38690
rect 29900 38910 30100 38920
rect 29900 38690 29910 38910
rect 30090 38690 30100 38910
rect 29900 38680 30100 38690
rect -4300 27250 -4100 27260
rect -4300 27030 -4290 27250
rect -4110 27030 -4100 27250
rect -4300 27020 -4100 27030
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect -4300 25710 -4100 25720
rect -4300 25490 -4290 25710
rect -4110 25490 -4100 25710
rect -4300 25480 -4100 25490
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect -4300 13900 -4100 13910
rect -4300 13420 -4290 13900
rect -4110 13420 -4100 13900
rect -4300 13410 -4100 13420
rect 30900 13900 31100 13910
rect 30900 13420 30910 13900
rect 31090 13420 31100 13900
rect 30900 13410 31100 13420
rect -4300 13090 -4100 13100
rect -4300 12610 -4290 13090
rect -4110 12610 -4100 13090
rect -4300 12600 -4100 12610
rect 30900 13090 31100 13100
rect 30900 12610 30910 13090
rect 31090 12610 31100 13090
rect 30900 12600 31100 12610
<< via1 >>
rect -3290 40190 -3110 40450
rect 29910 40276 30090 40450
rect 29910 40236 29984 40276
rect 29984 40236 30018 40276
rect 30018 40236 30090 40276
rect 29910 40190 30090 40236
rect -3290 38690 -3110 38910
rect 29910 38902 30090 38910
rect 29910 38862 29984 38902
rect 29984 38862 30018 38902
rect 30018 38862 30090 38902
rect 29910 38690 30090 38862
rect -4290 27030 -4110 27250
rect 30910 27076 31090 27250
rect 30910 27036 30984 27076
rect 30984 27036 31018 27076
rect 31018 27036 31090 27076
rect 30910 27030 31090 27036
rect -4290 25490 -4110 25710
rect 30910 25702 31090 25710
rect 30910 25662 30984 25702
rect 30984 25662 31018 25702
rect 31018 25662 31090 25702
rect 30910 25490 31090 25662
rect -4290 13420 -4110 13900
rect 30910 13832 31090 13900
rect 30910 13435 30980 13832
rect 30980 13435 31018 13832
rect 31018 13435 31090 13832
rect 30910 13420 31090 13435
rect -4290 12610 -4110 13090
rect 30910 13081 31090 13090
rect 30910 12684 30980 13081
rect 30980 12684 31018 13081
rect 31018 12684 31090 13081
rect 30910 12610 31090 12684
<< metal2 >>
rect -3300 40450 -3100 40460
rect -3300 40190 -3290 40450
rect -3110 40190 -3100 40450
rect -3300 40180 -3100 40190
rect 29900 40450 30100 40460
rect 29900 40190 29910 40450
rect 30090 40190 30100 40450
rect 29900 40180 30100 40190
rect -3300 38910 -3100 38920
rect -3300 38690 -3290 38910
rect -3110 38690 -3100 38910
rect -3300 38680 -3100 38690
rect 29900 38910 30100 38920
rect 29900 38690 29910 38910
rect 30090 38690 30100 38910
rect 29900 38680 30100 38690
rect -4300 27250 -4100 27260
rect -4300 27030 -4290 27250
rect -4110 27030 -4100 27250
rect -4300 27020 -4100 27030
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect -4300 25710 -4100 25720
rect -4300 25490 -4290 25710
rect -4110 25490 -4100 25710
rect -4300 25480 -4100 25490
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect -4300 13900 -4100 13910
rect -4300 13420 -4290 13900
rect -4110 13420 -4100 13900
rect -4300 13410 -4100 13420
rect 30900 13900 31100 13910
rect 30900 13420 30910 13900
rect 31090 13420 31100 13900
rect 30900 13410 31100 13420
rect -4300 13090 -4100 13100
rect -4300 12610 -4290 13090
rect -4110 12610 -4100 13090
rect -4300 12600 -4100 12610
rect 30900 13090 31100 13100
rect 30900 12610 30910 13090
rect 31090 12610 31100 13090
rect 30900 12600 31100 12610
<< via2 >>
rect -3290 40190 -3110 40450
rect 29910 40190 30090 40450
rect -3290 38690 -3110 38910
rect 29910 38690 30090 38910
rect -4290 27030 -4110 27250
rect 30910 27030 31090 27250
rect -4290 25490 -4110 25710
rect 30910 25490 31090 25710
rect -4290 13420 -4110 13900
rect 30910 13420 31090 13900
rect -4290 12610 -4110 13090
rect 30910 12610 31090 13090
<< metal3 >>
rect -3400 40480 -3000 40500
rect -3400 40410 -3380 40480
rect -3400 40190 -3390 40410
rect -3020 40410 -3000 40480
rect -3010 40190 -3000 40410
rect -3400 40180 -3000 40190
rect 29800 40480 30200 40500
rect 29800 40410 29820 40480
rect 29800 40190 29810 40410
rect 30180 40410 30200 40480
rect 30190 40190 30200 40410
rect 29800 40180 30200 40190
rect -3400 38910 -3000 38920
rect -3400 38690 -3390 38910
rect -3010 38690 -3000 38910
rect -3400 38680 -3000 38690
rect 29800 38910 30200 38920
rect 29800 38690 29810 38910
rect 30190 38690 30200 38910
rect 29800 38680 30200 38690
rect -4400 31700 2800 31800
rect -4400 31100 1400 31700
rect 2700 31100 2800 31700
rect -4400 31000 2800 31100
rect 24000 31700 31200 31800
rect 24000 31100 24100 31700
rect 25400 31100 31200 31700
rect 24000 31000 31200 31100
rect -4400 27250 -3900 31000
rect -4400 27030 -4290 27250
rect -4110 27030 -3900 27250
rect -4400 27000 -3900 27030
rect 30700 27250 31200 31000
rect 30700 27030 30910 27250
rect 31090 27030 31200 27250
rect 30700 27000 31200 27030
rect -4400 25710 -4000 25720
rect -4400 25490 -4390 25710
rect -4010 25490 -4000 25710
rect -4400 25480 -4000 25490
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25480 31200 25490
rect -4400 14000 -4000 14010
rect -4400 13420 -4390 14000
rect -4010 13420 -4000 14000
rect -4400 13410 -4000 13420
rect 30800 14000 31200 14010
rect 30800 13420 30810 14000
rect 31190 13420 31200 14000
rect 30800 13410 31200 13420
rect -4400 13090 -4000 13100
rect -4400 12510 -4390 13090
rect -4010 12510 -4000 13090
rect -4400 12500 -4000 12510
rect 30800 13090 31200 13100
rect 30800 12510 30810 13090
rect 31190 12510 31200 13090
rect 30800 12500 31200 12510
<< via3 >>
rect -3380 40450 -3020 40480
rect -3380 40410 -3290 40450
rect -3390 40190 -3290 40410
rect -3290 40190 -3110 40450
rect -3110 40410 -3020 40450
rect -3110 40190 -3010 40410
rect 29820 40450 30180 40480
rect 29820 40410 29910 40450
rect 29810 40190 29910 40410
rect 29910 40190 30090 40450
rect 30090 40410 30180 40450
rect 30090 40190 30190 40410
rect -3390 38690 -3290 38910
rect -3290 38690 -3110 38910
rect -3110 38690 -3010 38910
rect 29810 38690 29910 38910
rect 29910 38690 30090 38910
rect 30090 38690 30190 38910
rect 1400 31100 2700 31700
rect 24100 31100 25400 31700
rect -4390 25490 -4290 25710
rect -4290 25490 -4110 25710
rect -4110 25490 -4010 25710
rect 30810 25490 30910 25710
rect 30910 25490 31090 25710
rect 31090 25490 31190 25710
rect -4390 13900 -4010 14000
rect -4390 13420 -4290 13900
rect -4290 13420 -4110 13900
rect -4110 13420 -4010 13900
rect 30810 13900 31190 14000
rect 30810 13420 30910 13900
rect 30910 13420 31090 13900
rect 31090 13420 31190 13900
rect -4390 12610 -4290 13090
rect -4290 12610 -4110 13090
rect -4110 12610 -4010 13090
rect -4390 12510 -4010 12610
rect 30810 12610 30910 13090
rect 30910 12610 31090 13090
rect 31090 12610 31190 13090
rect 30810 12510 31190 12610
<< metal4 >>
rect -3400 40800 800 46000
rect -3400 40480 -3000 40500
rect -3400 40410 -3380 40480
rect -3400 40190 -3390 40410
rect -3020 40410 -3000 40480
rect -3010 40190 -3000 40410
rect -3400 40100 -3000 40190
rect -1000 39100 800 40800
rect -3400 38910 -3000 38920
rect -3400 38690 -3390 38910
rect -3010 38700 -3000 38910
rect -3010 38690 -1600 38700
rect -3400 38650 -3370 38690
rect -3030 38650 -1600 38690
rect -3400 38600 -1600 38650
rect -3400 37600 -3300 38600
rect -1700 37600 -1600 38600
rect -3400 37500 -1600 37600
rect -4400 25710 -4000 25720
rect -4400 25490 -4390 25710
rect -4010 25490 -4000 25710
rect -4400 25450 -4370 25490
rect -4030 25450 -4000 25490
rect -4400 25430 -4000 25450
rect -3400 24900 -1600 37100
rect -6400 14300 -1600 24900
rect -1000 25500 -600 39100
rect 700 25500 800 39100
rect 26000 40800 30200 46000
rect 26000 40700 27800 40800
rect 26000 39900 26100 40700
rect 27700 39900 27800 40700
rect 29800 40480 30200 40500
rect 29800 40410 29820 40480
rect 29800 40190 29810 40410
rect 30180 40410 30200 40480
rect 30190 40190 30200 40410
rect 29800 40100 30200 40190
rect 26000 38100 27800 39900
rect 29800 38910 30200 38920
rect 29800 38700 29810 38910
rect -1000 23200 800 25500
rect -1000 18500 -600 23200
rect 700 18500 800 23200
rect -1000 17800 800 18500
rect -1000 16600 -900 17800
rect 700 16600 800 17800
rect -1000 16500 800 16600
rect 26000 25500 26100 38100
rect 27400 25500 27800 38100
rect 28400 38690 29810 38700
rect 30190 38690 30200 38910
rect 28400 38650 29830 38690
rect 30170 38650 30200 38690
rect 28400 38600 30200 38650
rect 28400 37600 28500 38600
rect 30100 37600 30200 38600
rect 28400 37500 30200 37600
rect 26000 23200 27800 25500
rect 26000 18500 26100 23200
rect 27400 18500 27800 23200
rect 26000 17800 27800 18500
rect 26000 16600 26100 17800
rect 27700 16600 27800 17800
rect 26000 16500 27800 16600
rect 28400 24900 30200 37100
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25450 30830 25490
rect 31170 25450 31200 25490
rect 30800 25430 31200 25450
rect -4400 14000 -4000 14010
rect -4400 13420 -4390 14000
rect -4010 13420 -4000 14000
rect -4400 13410 -4000 13420
rect -3400 13900 -1600 14300
rect 28400 14300 33200 24900
rect 28400 13900 30200 14300
rect -3400 13100 800 13900
rect -4400 13090 800 13100
rect -4400 12510 -4390 13090
rect -4010 12510 800 13090
rect -4400 12500 800 12510
rect -3400 12100 800 12500
rect -3400 11100 -600 12100
rect -1000 8000 -600 11100
rect 700 10100 800 12100
rect 200 10000 800 10100
rect 26000 13100 30200 13900
rect 30800 14000 31200 14010
rect 30800 13420 30810 14000
rect 31190 13420 31200 14000
rect 30800 13410 31200 13420
rect 26000 13090 31200 13100
rect 26000 12510 30810 13090
rect 31190 12510 31200 13090
rect 26000 12500 31200 12510
rect 26000 12100 30200 12500
rect 26000 10100 26100 12100
rect 27400 11100 30200 12100
rect 26000 10000 26600 10100
rect 200 8000 300 10000
rect -1000 7900 300 8000
rect 26500 8000 26600 10000
rect 27400 8000 27800 11100
rect 26500 7900 27800 8000
rect -1000 7400 800 7900
rect -7200 3600 800 7400
rect 26000 7400 27800 7900
rect 26000 3600 34000 7400
rect -7200 1200 2800 3600
rect -7200 400 -7100 1200
rect 2600 400 2800 1200
rect 24000 1200 34000 3600
rect 24000 400 25600 1200
rect 33900 400 34000 1200
rect -7200 200 2800 400
rect 25500 200 34000 400
<< via4 >>
rect -3370 40210 -3030 40450
rect -3370 38690 -3030 38890
rect -3370 38650 -3030 38690
rect -3300 37600 -1700 38600
rect -4370 25490 -4030 25690
rect -4370 25450 -4030 25490
rect -600 25500 700 39100
rect 26100 39900 27700 40700
rect 29830 40210 30170 40450
rect -600 18500 700 23200
rect -900 16600 700 17800
rect 26100 25500 27400 38100
rect 29830 38690 30170 38890
rect 29830 38650 30170 38690
rect 28500 37600 30100 38600
rect 26100 18500 27400 23200
rect 26100 16600 27700 17800
rect 30830 25490 31170 25690
rect 30830 25450 31170 25490
rect -4370 13440 -4030 13980
rect -600 10100 700 12100
rect -600 8000 200 10100
rect 30830 13440 31170 13980
rect 26100 10100 27400 12100
rect 26600 8000 27400 10100
rect -7100 400 2600 1200
rect 25600 400 33900 1200
<< mimcap2 >>
rect -3300 45800 700 45900
rect -3300 41000 -3200 45800
rect 600 41000 700 45800
rect -3300 40900 700 41000
rect 26100 45800 30100 45900
rect 26100 41000 26200 45800
rect 30000 41000 30100 45800
rect 26100 40900 30100 41000
rect -3300 36900 -1700 37000
rect -3300 26700 -3200 36900
rect -1800 26700 -1700 36900
rect -3300 26600 -1700 26700
rect 28500 36900 30100 37000
rect 28500 26700 28600 36900
rect 30000 26700 30100 36900
rect 28500 26600 30100 26700
rect -6300 24700 -1700 24800
rect -6300 14500 -6200 24700
rect -1800 14500 -1700 24700
rect -6300 14400 -1700 14500
rect 28500 24700 33100 24800
rect 28500 14500 28600 24700
rect 33000 14500 33100 24700
rect 28500 14400 33100 14500
rect -7100 7200 700 7300
rect -7100 2400 -7000 7200
rect 600 2400 700 7200
rect -7100 2300 700 2400
rect 26100 7200 33900 7300
rect 26100 2400 26200 7200
rect 33800 2400 33900 7200
rect 26100 2300 33900 2400
<< mimcap2contact >>
rect -3200 41000 600 45800
rect 26200 41000 30000 45800
rect -3200 26700 -1800 36900
rect 28600 26700 30000 36900
rect -6200 14500 -1800 24700
rect 28600 14500 33000 24700
rect -7000 2400 600 7200
rect 26200 2400 33800 7200
<< metal5 >>
rect 1300 48100 2800 48500
rect 24000 48100 25500 48500
rect -600 46700 1300 47600
rect 25500 46700 27400 47600
rect -600 46000 800 46700
rect -3400 45800 800 46000
rect -3400 41000 -3200 45800
rect 600 41000 800 45800
rect -3400 40800 800 41000
rect 26000 46000 27400 46700
rect 26000 45800 30200 46000
rect 26000 41000 26200 45800
rect 30000 41000 30200 45800
rect 26000 40800 30200 41000
rect -3400 40450 -3000 40800
rect -3400 40210 -3370 40450
rect -3030 40210 -3000 40450
rect -3400 40100 -3000 40210
rect 26000 40700 27800 40800
rect -2400 40100 1200 40200
rect -2500 40000 1200 40100
rect -2600 39900 1200 40000
rect -2700 39800 1200 39900
rect 26000 39900 26100 40700
rect 27700 39900 27800 40700
rect 29800 40450 30200 40800
rect 29800 40210 29830 40450
rect 30170 40210 30200 40450
rect 29800 40100 30200 40210
rect 26000 39800 27800 39900
rect -2800 39700 1200 39800
rect -2900 39600 -1400 39700
rect -3000 39500 -1500 39600
rect -3000 39000 -1600 39500
rect 25400 39200 29200 39300
rect -3400 38890 -1600 39000
rect -3400 38650 -3370 38890
rect -3030 38650 -1600 38890
rect -3400 38600 -1600 38650
rect -3400 37600 -3300 38600
rect -1700 37600 -1600 38600
rect -3400 36900 -1600 37600
rect -3400 26700 -3200 36900
rect -1800 26700 -1600 36900
rect -3400 26500 -1600 26700
rect -700 39100 800 39200
rect -4400 25690 -4000 25720
rect -4400 25450 -4370 25690
rect -4030 25450 -4000 25690
rect -4400 24900 -4000 25450
rect -700 25500 -600 39100
rect 700 25500 800 39100
rect 25400 39100 29300 39200
rect 25400 39000 29400 39100
rect 25400 38890 30200 39000
rect 25400 38800 29830 38890
rect 28200 38700 29830 38800
rect 28300 38650 29830 38700
rect 30170 38650 30200 38890
rect 28300 38600 30200 38650
rect -700 25400 800 25500
rect 26000 38100 27500 38200
rect 26000 25500 26100 38100
rect 27400 25500 27500 38100
rect 28400 37600 28500 38600
rect 30100 37600 30200 38600
rect 28400 36900 30200 37600
rect 28400 26700 28600 36900
rect 30000 26700 30200 36900
rect 28400 26500 30200 26700
rect 26000 25400 27500 25500
rect 30800 25690 31200 25720
rect 30800 25450 30830 25690
rect 31170 25450 31200 25690
rect 30800 24900 31200 25450
rect -6400 24700 1200 24900
rect 25600 24700 33200 24900
rect -6400 14500 -6200 24700
rect -1800 24000 2100 24700
rect 24700 24000 28600 24700
rect -1800 23800 1200 24000
rect 25600 23800 28600 24000
rect -1800 14500 -1600 23800
rect -700 23200 800 23300
rect -700 18500 -600 23200
rect 700 18500 800 23200
rect -700 18400 800 18500
rect 26000 23200 27500 23300
rect 26000 18500 26100 23200
rect 27400 18500 27500 23200
rect 26000 18400 27500 18500
rect -6400 14300 -1600 14500
rect -1200 17800 1300 17900
rect -1200 16600 -900 17800
rect 700 16600 1300 17800
rect -1200 16500 1300 16600
rect 25500 17800 28000 17900
rect 25500 16600 26100 17800
rect 27700 16600 28000 17800
rect 25500 16500 28000 16600
rect -4400 13980 -4000 14300
rect -4400 13440 -4370 13980
rect -4030 13440 -4000 13980
rect -1200 13900 0 16500
rect -4400 13410 -4000 13440
rect -3400 12600 0 13900
rect 26800 13900 28000 16500
rect 28400 14500 28600 23800
rect 33000 14500 33200 24700
rect 28400 14300 33200 14500
rect 30800 13980 31200 14300
rect 26800 12600 30200 13900
rect 30800 13440 30830 13980
rect 31170 13440 31200 13980
rect 30800 13410 31200 13440
rect -3400 7400 -1600 12600
rect -700 12100 800 12200
rect -700 8000 -600 12100
rect 700 10100 800 12100
rect 200 10000 800 10100
rect 26000 12100 27500 12200
rect 26000 10100 26100 12100
rect 26000 10000 26600 10100
rect 200 8000 300 10000
rect 700 9100 1200 9600
rect 25400 8200 25900 8700
rect -700 7900 300 8000
rect 26500 8000 26600 10000
rect 27400 8000 27500 12100
rect 26500 7900 27500 8000
rect 28400 7400 30200 12600
rect -7200 7200 800 7400
rect -7200 2400 -7000 7200
rect 600 2400 800 7200
rect -7200 2200 800 2400
rect 26000 7200 34000 7400
rect 26000 2400 26200 7200
rect 33800 2400 34000 7200
rect 26000 2200 34000 2400
rect -7200 1200 1400 1400
rect 25400 1200 34000 1400
rect -7200 400 -7100 1200
rect 24200 400 25600 1200
rect 33900 400 34000 1200
rect -7200 200 2800 400
rect 1300 0 2800 200
rect 24000 200 34000 400
rect 24000 0 25500 200
use cascode_1  cascode_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/CLASSE
timestamp 1664506494
transform 1 0 14700 0 1 -3700
box -14700 3700 10800 52200
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_1
timestamp 1664814488
transform 1 0 -4201 0 1 26369
box -199 -889 199 889
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_3
timestamp 1664814488
transform 1 0 -3201 0 1 39569
box -199 -889 199 889
use sky130_fd_pr__res_high_po_0p35_FFWWQH  sky130_fd_pr__res_high_po_0p35_FFWWQH_0
timestamp 1664805031
transform 1 0 -4199 0 1 13258
box -201 -758 201 758
<< labels >>
rlabel metal5 1300 48100 2800 48500 1 VDN
rlabel metal5 900 39700 1200 40200 1 VGN
rlabel metal3 800 31000 1000 31800 1 N2
rlabel metal5 900 16500 1200 17900 1 N
rlabel metal5 700 9100 1000 9600 1 VINN
rlabel metal5 1300 0 2800 400 1 VSS
rlabel metal5 800 23800 1000 24800 1 MIDGATE
rlabel metal5 24000 48300 25500 48500 1 VDP
rlabel metal3 25600 31100 25900 31700 1 P2
rlabel metal5 25600 16500 25900 17900 1 P
rlabel metal5 24000 0 25500 200 1 VSSH
rlabel metal5 25700 38800 25900 39300 1 VGP
rlabel metal5 25700 8200 25900 8700 1 VINP
<< end >>
