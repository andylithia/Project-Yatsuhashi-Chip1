magic
tech sky130B
magscale 1 2
timestamp 1661115194
<< nwell >>
rect 17438 6910 20258 8170
rect 17420 5020 20240 6280
<< pwell >>
rect 17444 9121 17468 9172
rect 19294 9121 19318 9172
rect 15970 8130 17330 8140
rect 15964 8116 16040 8130
rect 16050 8116 17340 8130
rect 15964 8090 17340 8116
rect 15964 8041 17302 8090
rect 17315 8041 17340 8090
rect 15964 6970 17340 8041
rect 15970 6948 17330 6970
rect 15970 6943 17233 6948
rect 15970 6940 17184 6943
rect 11636 5822 15708 6884
rect 15970 6217 17184 6220
rect 15970 6212 17233 6217
rect 15970 6190 17330 6212
rect 15964 5119 17340 6190
rect 15964 5070 17302 5119
rect 17315 5070 17340 5119
rect 15964 5044 17340 5070
rect 15964 5030 16040 5044
rect 16050 5030 17340 5044
rect 15970 5020 17330 5030
rect 17444 4071 17468 4122
rect 19294 4071 19318 4122
<< nmos >>
rect 16163 6969 16193 7979
rect 16249 6969 16279 7979
rect 16335 6969 16365 7979
rect 16421 6969 16451 7979
rect 16507 6969 16537 7979
rect 16593 6969 16623 7979
rect 16679 6969 16709 7979
rect 16765 6969 16795 7979
rect 16851 6969 16881 7979
rect 16937 6969 16967 7979
rect 17023 6969 17053 7979
rect 17109 6969 17139 7979
rect 11830 5848 11860 6858
rect 11916 5848 11946 6858
rect 12002 5848 12032 6858
rect 12088 5848 12118 6858
rect 12396 5848 12426 6858
rect 12482 5848 12512 6858
rect 12568 5848 12598 6858
rect 12654 5848 12684 6858
rect 12962 5848 12992 6858
rect 13048 5848 13078 6858
rect 13134 5848 13164 6858
rect 13220 5848 13250 6858
rect 13528 5848 13558 6858
rect 13614 5848 13644 6858
rect 13700 5848 13730 6858
rect 13786 5848 13816 6858
rect 14094 5848 14124 6858
rect 14180 5848 14210 6858
rect 14266 5848 14296 6858
rect 14352 5848 14382 6858
rect 14660 5848 14690 6858
rect 14746 5848 14776 6858
rect 14832 5848 14862 6858
rect 14918 5848 14948 6858
rect 15226 5848 15256 6858
rect 15312 5848 15342 6858
rect 15398 5848 15428 6858
rect 15484 5848 15514 6858
rect 16163 5181 16193 6191
rect 16249 5181 16279 6191
rect 16335 5181 16365 6191
rect 16421 5181 16451 6191
rect 16507 5181 16537 6191
rect 16593 5181 16623 6191
rect 16679 5181 16709 6191
rect 16765 5181 16795 6191
rect 16851 5181 16881 6191
rect 16937 5181 16967 6191
rect 17023 5181 17053 6191
rect 17109 5181 17139 6191
<< pmos >>
rect 17667 6957 17697 7957
rect 17753 6957 17783 7957
rect 17839 6957 17869 7957
rect 17925 6957 17955 7957
rect 18011 6957 18041 7957
rect 18097 6957 18127 7957
rect 18183 6957 18213 7957
rect 18269 6957 18299 7957
rect 18355 6957 18385 7957
rect 18441 6957 18471 7957
rect 18527 6957 18557 7957
rect 18613 6957 18643 7957
rect 18699 6957 18729 7957
rect 18785 6957 18815 7957
rect 18871 6957 18901 7957
rect 18957 6957 18987 7957
rect 19043 6957 19073 7957
rect 19129 6957 19159 7957
rect 19215 6957 19245 7957
rect 19301 6957 19331 7957
rect 19387 6957 19417 7957
rect 19473 6957 19503 7957
rect 19559 6957 19589 7957
rect 19645 6957 19675 7957
rect 19731 6957 19761 7957
rect 19817 6957 19847 7957
rect 19903 6957 19933 7957
rect 19989 6957 20019 7957
rect 17649 5233 17679 6233
rect 17735 5233 17765 6233
rect 17821 5233 17851 6233
rect 17907 5233 17937 6233
rect 17993 5233 18023 6233
rect 18079 5233 18109 6233
rect 18165 5233 18195 6233
rect 18251 5233 18281 6233
rect 18337 5233 18367 6233
rect 18423 5233 18453 6233
rect 18509 5233 18539 6233
rect 18595 5233 18625 6233
rect 18681 5233 18711 6233
rect 18767 5233 18797 6233
rect 18853 5233 18883 6233
rect 18939 5233 18969 6233
rect 19025 5233 19055 6233
rect 19111 5233 19141 6233
rect 19197 5233 19227 6233
rect 19283 5233 19313 6233
rect 19369 5233 19399 6233
rect 19455 5233 19485 6233
rect 19541 5233 19571 6233
rect 19627 5233 19657 6233
rect 19713 5233 19743 6233
rect 19799 5233 19829 6233
rect 19885 5233 19915 6233
rect 19971 5233 20001 6233
<< ndiff >>
rect 16107 7967 16163 7979
rect 16107 7933 16118 7967
rect 16152 7933 16163 7967
rect 16107 7899 16163 7933
rect 16107 7865 16118 7899
rect 16152 7865 16163 7899
rect 16107 7831 16163 7865
rect 16107 7797 16118 7831
rect 16152 7797 16163 7831
rect 16107 7763 16163 7797
rect 16107 7729 16118 7763
rect 16152 7729 16163 7763
rect 16107 7695 16163 7729
rect 16107 7661 16118 7695
rect 16152 7661 16163 7695
rect 16107 7627 16163 7661
rect 16107 7593 16118 7627
rect 16152 7593 16163 7627
rect 16107 7559 16163 7593
rect 16107 7525 16118 7559
rect 16152 7525 16163 7559
rect 16107 7491 16163 7525
rect 16107 7457 16118 7491
rect 16152 7457 16163 7491
rect 16107 7423 16163 7457
rect 16107 7389 16118 7423
rect 16152 7389 16163 7423
rect 16107 7355 16163 7389
rect 16107 7321 16118 7355
rect 16152 7321 16163 7355
rect 16107 7287 16163 7321
rect 16107 7253 16118 7287
rect 16152 7253 16163 7287
rect 16107 7219 16163 7253
rect 16107 7185 16118 7219
rect 16152 7185 16163 7219
rect 16107 7151 16163 7185
rect 16107 7117 16118 7151
rect 16152 7117 16163 7151
rect 16107 7083 16163 7117
rect 16107 7049 16118 7083
rect 16152 7049 16163 7083
rect 16107 7015 16163 7049
rect 16107 6981 16118 7015
rect 16152 6981 16163 7015
rect 16107 6969 16163 6981
rect 16193 7967 16249 7979
rect 16193 7933 16204 7967
rect 16238 7933 16249 7967
rect 16193 7899 16249 7933
rect 16193 7865 16204 7899
rect 16238 7865 16249 7899
rect 16193 7831 16249 7865
rect 16193 7797 16204 7831
rect 16238 7797 16249 7831
rect 16193 7763 16249 7797
rect 16193 7729 16204 7763
rect 16238 7729 16249 7763
rect 16193 7695 16249 7729
rect 16193 7661 16204 7695
rect 16238 7661 16249 7695
rect 16193 7627 16249 7661
rect 16193 7593 16204 7627
rect 16238 7593 16249 7627
rect 16193 7559 16249 7593
rect 16193 7525 16204 7559
rect 16238 7525 16249 7559
rect 16193 7491 16249 7525
rect 16193 7457 16204 7491
rect 16238 7457 16249 7491
rect 16193 7423 16249 7457
rect 16193 7389 16204 7423
rect 16238 7389 16249 7423
rect 16193 7355 16249 7389
rect 16193 7321 16204 7355
rect 16238 7321 16249 7355
rect 16193 7287 16249 7321
rect 16193 7253 16204 7287
rect 16238 7253 16249 7287
rect 16193 7219 16249 7253
rect 16193 7185 16204 7219
rect 16238 7185 16249 7219
rect 16193 7151 16249 7185
rect 16193 7117 16204 7151
rect 16238 7117 16249 7151
rect 16193 7083 16249 7117
rect 16193 7049 16204 7083
rect 16238 7049 16249 7083
rect 16193 7015 16249 7049
rect 16193 6981 16204 7015
rect 16238 6981 16249 7015
rect 16193 6969 16249 6981
rect 16279 7967 16335 7979
rect 16279 7933 16290 7967
rect 16324 7933 16335 7967
rect 16279 7899 16335 7933
rect 16279 7865 16290 7899
rect 16324 7865 16335 7899
rect 16279 7831 16335 7865
rect 16279 7797 16290 7831
rect 16324 7797 16335 7831
rect 16279 7763 16335 7797
rect 16279 7729 16290 7763
rect 16324 7729 16335 7763
rect 16279 7695 16335 7729
rect 16279 7661 16290 7695
rect 16324 7661 16335 7695
rect 16279 7627 16335 7661
rect 16279 7593 16290 7627
rect 16324 7593 16335 7627
rect 16279 7559 16335 7593
rect 16279 7525 16290 7559
rect 16324 7525 16335 7559
rect 16279 7491 16335 7525
rect 16279 7457 16290 7491
rect 16324 7457 16335 7491
rect 16279 7423 16335 7457
rect 16279 7389 16290 7423
rect 16324 7389 16335 7423
rect 16279 7355 16335 7389
rect 16279 7321 16290 7355
rect 16324 7321 16335 7355
rect 16279 7287 16335 7321
rect 16279 7253 16290 7287
rect 16324 7253 16335 7287
rect 16279 7219 16335 7253
rect 16279 7185 16290 7219
rect 16324 7185 16335 7219
rect 16279 7151 16335 7185
rect 16279 7117 16290 7151
rect 16324 7117 16335 7151
rect 16279 7083 16335 7117
rect 16279 7049 16290 7083
rect 16324 7049 16335 7083
rect 16279 7015 16335 7049
rect 16279 6981 16290 7015
rect 16324 6981 16335 7015
rect 16279 6969 16335 6981
rect 16365 7967 16421 7979
rect 16365 7933 16376 7967
rect 16410 7933 16421 7967
rect 16365 7899 16421 7933
rect 16365 7865 16376 7899
rect 16410 7865 16421 7899
rect 16365 7831 16421 7865
rect 16365 7797 16376 7831
rect 16410 7797 16421 7831
rect 16365 7763 16421 7797
rect 16365 7729 16376 7763
rect 16410 7729 16421 7763
rect 16365 7695 16421 7729
rect 16365 7661 16376 7695
rect 16410 7661 16421 7695
rect 16365 7627 16421 7661
rect 16365 7593 16376 7627
rect 16410 7593 16421 7627
rect 16365 7559 16421 7593
rect 16365 7525 16376 7559
rect 16410 7525 16421 7559
rect 16365 7491 16421 7525
rect 16365 7457 16376 7491
rect 16410 7457 16421 7491
rect 16365 7423 16421 7457
rect 16365 7389 16376 7423
rect 16410 7389 16421 7423
rect 16365 7355 16421 7389
rect 16365 7321 16376 7355
rect 16410 7321 16421 7355
rect 16365 7287 16421 7321
rect 16365 7253 16376 7287
rect 16410 7253 16421 7287
rect 16365 7219 16421 7253
rect 16365 7185 16376 7219
rect 16410 7185 16421 7219
rect 16365 7151 16421 7185
rect 16365 7117 16376 7151
rect 16410 7117 16421 7151
rect 16365 7083 16421 7117
rect 16365 7049 16376 7083
rect 16410 7049 16421 7083
rect 16365 7015 16421 7049
rect 16365 6981 16376 7015
rect 16410 6981 16421 7015
rect 16365 6969 16421 6981
rect 16451 7967 16507 7979
rect 16451 7933 16462 7967
rect 16496 7933 16507 7967
rect 16451 7899 16507 7933
rect 16451 7865 16462 7899
rect 16496 7865 16507 7899
rect 16451 7831 16507 7865
rect 16451 7797 16462 7831
rect 16496 7797 16507 7831
rect 16451 7763 16507 7797
rect 16451 7729 16462 7763
rect 16496 7729 16507 7763
rect 16451 7695 16507 7729
rect 16451 7661 16462 7695
rect 16496 7661 16507 7695
rect 16451 7627 16507 7661
rect 16451 7593 16462 7627
rect 16496 7593 16507 7627
rect 16451 7559 16507 7593
rect 16451 7525 16462 7559
rect 16496 7525 16507 7559
rect 16451 7491 16507 7525
rect 16451 7457 16462 7491
rect 16496 7457 16507 7491
rect 16451 7423 16507 7457
rect 16451 7389 16462 7423
rect 16496 7389 16507 7423
rect 16451 7355 16507 7389
rect 16451 7321 16462 7355
rect 16496 7321 16507 7355
rect 16451 7287 16507 7321
rect 16451 7253 16462 7287
rect 16496 7253 16507 7287
rect 16451 7219 16507 7253
rect 16451 7185 16462 7219
rect 16496 7185 16507 7219
rect 16451 7151 16507 7185
rect 16451 7117 16462 7151
rect 16496 7117 16507 7151
rect 16451 7083 16507 7117
rect 16451 7049 16462 7083
rect 16496 7049 16507 7083
rect 16451 7015 16507 7049
rect 16451 6981 16462 7015
rect 16496 6981 16507 7015
rect 16451 6969 16507 6981
rect 16537 7967 16593 7979
rect 16537 7933 16548 7967
rect 16582 7933 16593 7967
rect 16537 7899 16593 7933
rect 16537 7865 16548 7899
rect 16582 7865 16593 7899
rect 16537 7831 16593 7865
rect 16537 7797 16548 7831
rect 16582 7797 16593 7831
rect 16537 7763 16593 7797
rect 16537 7729 16548 7763
rect 16582 7729 16593 7763
rect 16537 7695 16593 7729
rect 16537 7661 16548 7695
rect 16582 7661 16593 7695
rect 16537 7627 16593 7661
rect 16537 7593 16548 7627
rect 16582 7593 16593 7627
rect 16537 7559 16593 7593
rect 16537 7525 16548 7559
rect 16582 7525 16593 7559
rect 16537 7491 16593 7525
rect 16537 7457 16548 7491
rect 16582 7457 16593 7491
rect 16537 7423 16593 7457
rect 16537 7389 16548 7423
rect 16582 7389 16593 7423
rect 16537 7355 16593 7389
rect 16537 7321 16548 7355
rect 16582 7321 16593 7355
rect 16537 7287 16593 7321
rect 16537 7253 16548 7287
rect 16582 7253 16593 7287
rect 16537 7219 16593 7253
rect 16537 7185 16548 7219
rect 16582 7185 16593 7219
rect 16537 7151 16593 7185
rect 16537 7117 16548 7151
rect 16582 7117 16593 7151
rect 16537 7083 16593 7117
rect 16537 7049 16548 7083
rect 16582 7049 16593 7083
rect 16537 7015 16593 7049
rect 16537 6981 16548 7015
rect 16582 6981 16593 7015
rect 16537 6969 16593 6981
rect 16623 7967 16679 7979
rect 16623 7933 16634 7967
rect 16668 7933 16679 7967
rect 16623 7899 16679 7933
rect 16623 7865 16634 7899
rect 16668 7865 16679 7899
rect 16623 7831 16679 7865
rect 16623 7797 16634 7831
rect 16668 7797 16679 7831
rect 16623 7763 16679 7797
rect 16623 7729 16634 7763
rect 16668 7729 16679 7763
rect 16623 7695 16679 7729
rect 16623 7661 16634 7695
rect 16668 7661 16679 7695
rect 16623 7627 16679 7661
rect 16623 7593 16634 7627
rect 16668 7593 16679 7627
rect 16623 7559 16679 7593
rect 16623 7525 16634 7559
rect 16668 7525 16679 7559
rect 16623 7491 16679 7525
rect 16623 7457 16634 7491
rect 16668 7457 16679 7491
rect 16623 7423 16679 7457
rect 16623 7389 16634 7423
rect 16668 7389 16679 7423
rect 16623 7355 16679 7389
rect 16623 7321 16634 7355
rect 16668 7321 16679 7355
rect 16623 7287 16679 7321
rect 16623 7253 16634 7287
rect 16668 7253 16679 7287
rect 16623 7219 16679 7253
rect 16623 7185 16634 7219
rect 16668 7185 16679 7219
rect 16623 7151 16679 7185
rect 16623 7117 16634 7151
rect 16668 7117 16679 7151
rect 16623 7083 16679 7117
rect 16623 7049 16634 7083
rect 16668 7049 16679 7083
rect 16623 7015 16679 7049
rect 16623 6981 16634 7015
rect 16668 6981 16679 7015
rect 16623 6969 16679 6981
rect 16709 7967 16765 7979
rect 16709 7933 16720 7967
rect 16754 7933 16765 7967
rect 16709 7899 16765 7933
rect 16709 7865 16720 7899
rect 16754 7865 16765 7899
rect 16709 7831 16765 7865
rect 16709 7797 16720 7831
rect 16754 7797 16765 7831
rect 16709 7763 16765 7797
rect 16709 7729 16720 7763
rect 16754 7729 16765 7763
rect 16709 7695 16765 7729
rect 16709 7661 16720 7695
rect 16754 7661 16765 7695
rect 16709 7627 16765 7661
rect 16709 7593 16720 7627
rect 16754 7593 16765 7627
rect 16709 7559 16765 7593
rect 16709 7525 16720 7559
rect 16754 7525 16765 7559
rect 16709 7491 16765 7525
rect 16709 7457 16720 7491
rect 16754 7457 16765 7491
rect 16709 7423 16765 7457
rect 16709 7389 16720 7423
rect 16754 7389 16765 7423
rect 16709 7355 16765 7389
rect 16709 7321 16720 7355
rect 16754 7321 16765 7355
rect 16709 7287 16765 7321
rect 16709 7253 16720 7287
rect 16754 7253 16765 7287
rect 16709 7219 16765 7253
rect 16709 7185 16720 7219
rect 16754 7185 16765 7219
rect 16709 7151 16765 7185
rect 16709 7117 16720 7151
rect 16754 7117 16765 7151
rect 16709 7083 16765 7117
rect 16709 7049 16720 7083
rect 16754 7049 16765 7083
rect 16709 7015 16765 7049
rect 16709 6981 16720 7015
rect 16754 6981 16765 7015
rect 16709 6969 16765 6981
rect 16795 7967 16851 7979
rect 16795 7933 16806 7967
rect 16840 7933 16851 7967
rect 16795 7899 16851 7933
rect 16795 7865 16806 7899
rect 16840 7865 16851 7899
rect 16795 7831 16851 7865
rect 16795 7797 16806 7831
rect 16840 7797 16851 7831
rect 16795 7763 16851 7797
rect 16795 7729 16806 7763
rect 16840 7729 16851 7763
rect 16795 7695 16851 7729
rect 16795 7661 16806 7695
rect 16840 7661 16851 7695
rect 16795 7627 16851 7661
rect 16795 7593 16806 7627
rect 16840 7593 16851 7627
rect 16795 7559 16851 7593
rect 16795 7525 16806 7559
rect 16840 7525 16851 7559
rect 16795 7491 16851 7525
rect 16795 7457 16806 7491
rect 16840 7457 16851 7491
rect 16795 7423 16851 7457
rect 16795 7389 16806 7423
rect 16840 7389 16851 7423
rect 16795 7355 16851 7389
rect 16795 7321 16806 7355
rect 16840 7321 16851 7355
rect 16795 7287 16851 7321
rect 16795 7253 16806 7287
rect 16840 7253 16851 7287
rect 16795 7219 16851 7253
rect 16795 7185 16806 7219
rect 16840 7185 16851 7219
rect 16795 7151 16851 7185
rect 16795 7117 16806 7151
rect 16840 7117 16851 7151
rect 16795 7083 16851 7117
rect 16795 7049 16806 7083
rect 16840 7049 16851 7083
rect 16795 7015 16851 7049
rect 16795 6981 16806 7015
rect 16840 6981 16851 7015
rect 16795 6969 16851 6981
rect 16881 7967 16937 7979
rect 16881 7933 16892 7967
rect 16926 7933 16937 7967
rect 16881 7899 16937 7933
rect 16881 7865 16892 7899
rect 16926 7865 16937 7899
rect 16881 7831 16937 7865
rect 16881 7797 16892 7831
rect 16926 7797 16937 7831
rect 16881 7763 16937 7797
rect 16881 7729 16892 7763
rect 16926 7729 16937 7763
rect 16881 7695 16937 7729
rect 16881 7661 16892 7695
rect 16926 7661 16937 7695
rect 16881 7627 16937 7661
rect 16881 7593 16892 7627
rect 16926 7593 16937 7627
rect 16881 7559 16937 7593
rect 16881 7525 16892 7559
rect 16926 7525 16937 7559
rect 16881 7491 16937 7525
rect 16881 7457 16892 7491
rect 16926 7457 16937 7491
rect 16881 7423 16937 7457
rect 16881 7389 16892 7423
rect 16926 7389 16937 7423
rect 16881 7355 16937 7389
rect 16881 7321 16892 7355
rect 16926 7321 16937 7355
rect 16881 7287 16937 7321
rect 16881 7253 16892 7287
rect 16926 7253 16937 7287
rect 16881 7219 16937 7253
rect 16881 7185 16892 7219
rect 16926 7185 16937 7219
rect 16881 7151 16937 7185
rect 16881 7117 16892 7151
rect 16926 7117 16937 7151
rect 16881 7083 16937 7117
rect 16881 7049 16892 7083
rect 16926 7049 16937 7083
rect 16881 7015 16937 7049
rect 16881 6981 16892 7015
rect 16926 6981 16937 7015
rect 16881 6969 16937 6981
rect 16967 7967 17023 7979
rect 16967 7933 16978 7967
rect 17012 7933 17023 7967
rect 16967 7899 17023 7933
rect 16967 7865 16978 7899
rect 17012 7865 17023 7899
rect 16967 7831 17023 7865
rect 16967 7797 16978 7831
rect 17012 7797 17023 7831
rect 16967 7763 17023 7797
rect 16967 7729 16978 7763
rect 17012 7729 17023 7763
rect 16967 7695 17023 7729
rect 16967 7661 16978 7695
rect 17012 7661 17023 7695
rect 16967 7627 17023 7661
rect 16967 7593 16978 7627
rect 17012 7593 17023 7627
rect 16967 7559 17023 7593
rect 16967 7525 16978 7559
rect 17012 7525 17023 7559
rect 16967 7491 17023 7525
rect 16967 7457 16978 7491
rect 17012 7457 17023 7491
rect 16967 7423 17023 7457
rect 16967 7389 16978 7423
rect 17012 7389 17023 7423
rect 16967 7355 17023 7389
rect 16967 7321 16978 7355
rect 17012 7321 17023 7355
rect 16967 7287 17023 7321
rect 16967 7253 16978 7287
rect 17012 7253 17023 7287
rect 16967 7219 17023 7253
rect 16967 7185 16978 7219
rect 17012 7185 17023 7219
rect 16967 7151 17023 7185
rect 16967 7117 16978 7151
rect 17012 7117 17023 7151
rect 16967 7083 17023 7117
rect 16967 7049 16978 7083
rect 17012 7049 17023 7083
rect 16967 7015 17023 7049
rect 16967 6981 16978 7015
rect 17012 6981 17023 7015
rect 16967 6969 17023 6981
rect 17053 7967 17109 7979
rect 17053 7933 17064 7967
rect 17098 7933 17109 7967
rect 17053 7899 17109 7933
rect 17053 7865 17064 7899
rect 17098 7865 17109 7899
rect 17053 7831 17109 7865
rect 17053 7797 17064 7831
rect 17098 7797 17109 7831
rect 17053 7763 17109 7797
rect 17053 7729 17064 7763
rect 17098 7729 17109 7763
rect 17053 7695 17109 7729
rect 17053 7661 17064 7695
rect 17098 7661 17109 7695
rect 17053 7627 17109 7661
rect 17053 7593 17064 7627
rect 17098 7593 17109 7627
rect 17053 7559 17109 7593
rect 17053 7525 17064 7559
rect 17098 7525 17109 7559
rect 17053 7491 17109 7525
rect 17053 7457 17064 7491
rect 17098 7457 17109 7491
rect 17053 7423 17109 7457
rect 17053 7389 17064 7423
rect 17098 7389 17109 7423
rect 17053 7355 17109 7389
rect 17053 7321 17064 7355
rect 17098 7321 17109 7355
rect 17053 7287 17109 7321
rect 17053 7253 17064 7287
rect 17098 7253 17109 7287
rect 17053 7219 17109 7253
rect 17053 7185 17064 7219
rect 17098 7185 17109 7219
rect 17053 7151 17109 7185
rect 17053 7117 17064 7151
rect 17098 7117 17109 7151
rect 17053 7083 17109 7117
rect 17053 7049 17064 7083
rect 17098 7049 17109 7083
rect 17053 7015 17109 7049
rect 17053 6981 17064 7015
rect 17098 6981 17109 7015
rect 17053 6969 17109 6981
rect 17139 7967 17195 7979
rect 17139 7933 17150 7967
rect 17184 7933 17195 7967
rect 17139 7899 17195 7933
rect 17139 7865 17150 7899
rect 17184 7865 17195 7899
rect 17139 7831 17195 7865
rect 17139 7797 17150 7831
rect 17184 7797 17195 7831
rect 17139 7763 17195 7797
rect 17139 7729 17150 7763
rect 17184 7729 17195 7763
rect 17139 7695 17195 7729
rect 17139 7661 17150 7695
rect 17184 7661 17195 7695
rect 17139 7627 17195 7661
rect 17139 7593 17150 7627
rect 17184 7593 17195 7627
rect 17139 7559 17195 7593
rect 17139 7525 17150 7559
rect 17184 7525 17195 7559
rect 17139 7491 17195 7525
rect 17139 7457 17150 7491
rect 17184 7457 17195 7491
rect 17139 7423 17195 7457
rect 17139 7389 17150 7423
rect 17184 7389 17195 7423
rect 17139 7355 17195 7389
rect 17139 7321 17150 7355
rect 17184 7321 17195 7355
rect 17139 7287 17195 7321
rect 17139 7253 17150 7287
rect 17184 7253 17195 7287
rect 17139 7219 17195 7253
rect 17139 7185 17150 7219
rect 17184 7185 17195 7219
rect 17139 7151 17195 7185
rect 17139 7117 17150 7151
rect 17184 7117 17195 7151
rect 17139 7083 17195 7117
rect 17139 7049 17150 7083
rect 17184 7049 17195 7083
rect 17139 7015 17195 7049
rect 17139 6981 17150 7015
rect 17184 6981 17195 7015
rect 17139 6969 17195 6981
rect 11774 6846 11830 6858
rect 11774 6812 11785 6846
rect 11819 6812 11830 6846
rect 11774 6778 11830 6812
rect 11774 6744 11785 6778
rect 11819 6744 11830 6778
rect 11774 6710 11830 6744
rect 11774 6676 11785 6710
rect 11819 6676 11830 6710
rect 11774 6642 11830 6676
rect 11774 6608 11785 6642
rect 11819 6608 11830 6642
rect 11774 6574 11830 6608
rect 11774 6540 11785 6574
rect 11819 6540 11830 6574
rect 11774 6506 11830 6540
rect 11774 6472 11785 6506
rect 11819 6472 11830 6506
rect 11774 6438 11830 6472
rect 11774 6404 11785 6438
rect 11819 6404 11830 6438
rect 11774 6370 11830 6404
rect 11774 6336 11785 6370
rect 11819 6336 11830 6370
rect 11774 6302 11830 6336
rect 11774 6268 11785 6302
rect 11819 6268 11830 6302
rect 11774 6234 11830 6268
rect 11774 6200 11785 6234
rect 11819 6200 11830 6234
rect 11774 6166 11830 6200
rect 11774 6132 11785 6166
rect 11819 6132 11830 6166
rect 11774 6098 11830 6132
rect 11774 6064 11785 6098
rect 11819 6064 11830 6098
rect 11774 6030 11830 6064
rect 11774 5996 11785 6030
rect 11819 5996 11830 6030
rect 11774 5962 11830 5996
rect 11774 5928 11785 5962
rect 11819 5928 11830 5962
rect 11774 5894 11830 5928
rect 11774 5860 11785 5894
rect 11819 5860 11830 5894
rect 11774 5848 11830 5860
rect 11860 6846 11916 6858
rect 11860 6812 11871 6846
rect 11905 6812 11916 6846
rect 11860 6778 11916 6812
rect 11860 6744 11871 6778
rect 11905 6744 11916 6778
rect 11860 6710 11916 6744
rect 11860 6676 11871 6710
rect 11905 6676 11916 6710
rect 11860 6642 11916 6676
rect 11860 6608 11871 6642
rect 11905 6608 11916 6642
rect 11860 6574 11916 6608
rect 11860 6540 11871 6574
rect 11905 6540 11916 6574
rect 11860 6506 11916 6540
rect 11860 6472 11871 6506
rect 11905 6472 11916 6506
rect 11860 6438 11916 6472
rect 11860 6404 11871 6438
rect 11905 6404 11916 6438
rect 11860 6370 11916 6404
rect 11860 6336 11871 6370
rect 11905 6336 11916 6370
rect 11860 6302 11916 6336
rect 11860 6268 11871 6302
rect 11905 6268 11916 6302
rect 11860 6234 11916 6268
rect 11860 6200 11871 6234
rect 11905 6200 11916 6234
rect 11860 6166 11916 6200
rect 11860 6132 11871 6166
rect 11905 6132 11916 6166
rect 11860 6098 11916 6132
rect 11860 6064 11871 6098
rect 11905 6064 11916 6098
rect 11860 6030 11916 6064
rect 11860 5996 11871 6030
rect 11905 5996 11916 6030
rect 11860 5962 11916 5996
rect 11860 5928 11871 5962
rect 11905 5928 11916 5962
rect 11860 5894 11916 5928
rect 11860 5860 11871 5894
rect 11905 5860 11916 5894
rect 11860 5848 11916 5860
rect 11946 6846 12002 6858
rect 11946 6812 11957 6846
rect 11991 6812 12002 6846
rect 11946 6778 12002 6812
rect 11946 6744 11957 6778
rect 11991 6744 12002 6778
rect 11946 6710 12002 6744
rect 11946 6676 11957 6710
rect 11991 6676 12002 6710
rect 11946 6642 12002 6676
rect 11946 6608 11957 6642
rect 11991 6608 12002 6642
rect 11946 6574 12002 6608
rect 11946 6540 11957 6574
rect 11991 6540 12002 6574
rect 11946 6506 12002 6540
rect 11946 6472 11957 6506
rect 11991 6472 12002 6506
rect 11946 6438 12002 6472
rect 11946 6404 11957 6438
rect 11991 6404 12002 6438
rect 11946 6370 12002 6404
rect 11946 6336 11957 6370
rect 11991 6336 12002 6370
rect 11946 6302 12002 6336
rect 11946 6268 11957 6302
rect 11991 6268 12002 6302
rect 11946 6234 12002 6268
rect 11946 6200 11957 6234
rect 11991 6200 12002 6234
rect 11946 6166 12002 6200
rect 11946 6132 11957 6166
rect 11991 6132 12002 6166
rect 11946 6098 12002 6132
rect 11946 6064 11957 6098
rect 11991 6064 12002 6098
rect 11946 6030 12002 6064
rect 11946 5996 11957 6030
rect 11991 5996 12002 6030
rect 11946 5962 12002 5996
rect 11946 5928 11957 5962
rect 11991 5928 12002 5962
rect 11946 5894 12002 5928
rect 11946 5860 11957 5894
rect 11991 5860 12002 5894
rect 11946 5848 12002 5860
rect 12032 6846 12088 6858
rect 12032 6812 12043 6846
rect 12077 6812 12088 6846
rect 12032 6778 12088 6812
rect 12032 6744 12043 6778
rect 12077 6744 12088 6778
rect 12032 6710 12088 6744
rect 12032 6676 12043 6710
rect 12077 6676 12088 6710
rect 12032 6642 12088 6676
rect 12032 6608 12043 6642
rect 12077 6608 12088 6642
rect 12032 6574 12088 6608
rect 12032 6540 12043 6574
rect 12077 6540 12088 6574
rect 12032 6506 12088 6540
rect 12032 6472 12043 6506
rect 12077 6472 12088 6506
rect 12032 6438 12088 6472
rect 12032 6404 12043 6438
rect 12077 6404 12088 6438
rect 12032 6370 12088 6404
rect 12032 6336 12043 6370
rect 12077 6336 12088 6370
rect 12032 6302 12088 6336
rect 12032 6268 12043 6302
rect 12077 6268 12088 6302
rect 12032 6234 12088 6268
rect 12032 6200 12043 6234
rect 12077 6200 12088 6234
rect 12032 6166 12088 6200
rect 12032 6132 12043 6166
rect 12077 6132 12088 6166
rect 12032 6098 12088 6132
rect 12032 6064 12043 6098
rect 12077 6064 12088 6098
rect 12032 6030 12088 6064
rect 12032 5996 12043 6030
rect 12077 5996 12088 6030
rect 12032 5962 12088 5996
rect 12032 5928 12043 5962
rect 12077 5928 12088 5962
rect 12032 5894 12088 5928
rect 12032 5860 12043 5894
rect 12077 5860 12088 5894
rect 12032 5848 12088 5860
rect 12118 6846 12174 6858
rect 12118 6812 12129 6846
rect 12163 6812 12174 6846
rect 12118 6778 12174 6812
rect 12118 6744 12129 6778
rect 12163 6744 12174 6778
rect 12118 6710 12174 6744
rect 12118 6676 12129 6710
rect 12163 6676 12174 6710
rect 12118 6642 12174 6676
rect 12118 6608 12129 6642
rect 12163 6608 12174 6642
rect 12118 6574 12174 6608
rect 12118 6540 12129 6574
rect 12163 6540 12174 6574
rect 12118 6506 12174 6540
rect 12118 6472 12129 6506
rect 12163 6472 12174 6506
rect 12118 6438 12174 6472
rect 12118 6404 12129 6438
rect 12163 6404 12174 6438
rect 12118 6370 12174 6404
rect 12118 6336 12129 6370
rect 12163 6336 12174 6370
rect 12118 6302 12174 6336
rect 12118 6268 12129 6302
rect 12163 6268 12174 6302
rect 12118 6234 12174 6268
rect 12118 6200 12129 6234
rect 12163 6200 12174 6234
rect 12118 6166 12174 6200
rect 12118 6132 12129 6166
rect 12163 6132 12174 6166
rect 12118 6098 12174 6132
rect 12118 6064 12129 6098
rect 12163 6064 12174 6098
rect 12118 6030 12174 6064
rect 12118 5996 12129 6030
rect 12163 5996 12174 6030
rect 12118 5962 12174 5996
rect 12118 5928 12129 5962
rect 12163 5928 12174 5962
rect 12118 5894 12174 5928
rect 12118 5860 12129 5894
rect 12163 5860 12174 5894
rect 12118 5848 12174 5860
rect 12340 6846 12396 6858
rect 12340 6812 12351 6846
rect 12385 6812 12396 6846
rect 12340 6778 12396 6812
rect 12340 6744 12351 6778
rect 12385 6744 12396 6778
rect 12340 6710 12396 6744
rect 12340 6676 12351 6710
rect 12385 6676 12396 6710
rect 12340 6642 12396 6676
rect 12340 6608 12351 6642
rect 12385 6608 12396 6642
rect 12340 6574 12396 6608
rect 12340 6540 12351 6574
rect 12385 6540 12396 6574
rect 12340 6506 12396 6540
rect 12340 6472 12351 6506
rect 12385 6472 12396 6506
rect 12340 6438 12396 6472
rect 12340 6404 12351 6438
rect 12385 6404 12396 6438
rect 12340 6370 12396 6404
rect 12340 6336 12351 6370
rect 12385 6336 12396 6370
rect 12340 6302 12396 6336
rect 12340 6268 12351 6302
rect 12385 6268 12396 6302
rect 12340 6234 12396 6268
rect 12340 6200 12351 6234
rect 12385 6200 12396 6234
rect 12340 6166 12396 6200
rect 12340 6132 12351 6166
rect 12385 6132 12396 6166
rect 12340 6098 12396 6132
rect 12340 6064 12351 6098
rect 12385 6064 12396 6098
rect 12340 6030 12396 6064
rect 12340 5996 12351 6030
rect 12385 5996 12396 6030
rect 12340 5962 12396 5996
rect 12340 5928 12351 5962
rect 12385 5928 12396 5962
rect 12340 5894 12396 5928
rect 12340 5860 12351 5894
rect 12385 5860 12396 5894
rect 12340 5848 12396 5860
rect 12426 6846 12482 6858
rect 12426 6812 12437 6846
rect 12471 6812 12482 6846
rect 12426 6778 12482 6812
rect 12426 6744 12437 6778
rect 12471 6744 12482 6778
rect 12426 6710 12482 6744
rect 12426 6676 12437 6710
rect 12471 6676 12482 6710
rect 12426 6642 12482 6676
rect 12426 6608 12437 6642
rect 12471 6608 12482 6642
rect 12426 6574 12482 6608
rect 12426 6540 12437 6574
rect 12471 6540 12482 6574
rect 12426 6506 12482 6540
rect 12426 6472 12437 6506
rect 12471 6472 12482 6506
rect 12426 6438 12482 6472
rect 12426 6404 12437 6438
rect 12471 6404 12482 6438
rect 12426 6370 12482 6404
rect 12426 6336 12437 6370
rect 12471 6336 12482 6370
rect 12426 6302 12482 6336
rect 12426 6268 12437 6302
rect 12471 6268 12482 6302
rect 12426 6234 12482 6268
rect 12426 6200 12437 6234
rect 12471 6200 12482 6234
rect 12426 6166 12482 6200
rect 12426 6132 12437 6166
rect 12471 6132 12482 6166
rect 12426 6098 12482 6132
rect 12426 6064 12437 6098
rect 12471 6064 12482 6098
rect 12426 6030 12482 6064
rect 12426 5996 12437 6030
rect 12471 5996 12482 6030
rect 12426 5962 12482 5996
rect 12426 5928 12437 5962
rect 12471 5928 12482 5962
rect 12426 5894 12482 5928
rect 12426 5860 12437 5894
rect 12471 5860 12482 5894
rect 12426 5848 12482 5860
rect 12512 6846 12568 6858
rect 12512 6812 12523 6846
rect 12557 6812 12568 6846
rect 12512 6778 12568 6812
rect 12512 6744 12523 6778
rect 12557 6744 12568 6778
rect 12512 6710 12568 6744
rect 12512 6676 12523 6710
rect 12557 6676 12568 6710
rect 12512 6642 12568 6676
rect 12512 6608 12523 6642
rect 12557 6608 12568 6642
rect 12512 6574 12568 6608
rect 12512 6540 12523 6574
rect 12557 6540 12568 6574
rect 12512 6506 12568 6540
rect 12512 6472 12523 6506
rect 12557 6472 12568 6506
rect 12512 6438 12568 6472
rect 12512 6404 12523 6438
rect 12557 6404 12568 6438
rect 12512 6370 12568 6404
rect 12512 6336 12523 6370
rect 12557 6336 12568 6370
rect 12512 6302 12568 6336
rect 12512 6268 12523 6302
rect 12557 6268 12568 6302
rect 12512 6234 12568 6268
rect 12512 6200 12523 6234
rect 12557 6200 12568 6234
rect 12512 6166 12568 6200
rect 12512 6132 12523 6166
rect 12557 6132 12568 6166
rect 12512 6098 12568 6132
rect 12512 6064 12523 6098
rect 12557 6064 12568 6098
rect 12512 6030 12568 6064
rect 12512 5996 12523 6030
rect 12557 5996 12568 6030
rect 12512 5962 12568 5996
rect 12512 5928 12523 5962
rect 12557 5928 12568 5962
rect 12512 5894 12568 5928
rect 12512 5860 12523 5894
rect 12557 5860 12568 5894
rect 12512 5848 12568 5860
rect 12598 6846 12654 6858
rect 12598 6812 12609 6846
rect 12643 6812 12654 6846
rect 12598 6778 12654 6812
rect 12598 6744 12609 6778
rect 12643 6744 12654 6778
rect 12598 6710 12654 6744
rect 12598 6676 12609 6710
rect 12643 6676 12654 6710
rect 12598 6642 12654 6676
rect 12598 6608 12609 6642
rect 12643 6608 12654 6642
rect 12598 6574 12654 6608
rect 12598 6540 12609 6574
rect 12643 6540 12654 6574
rect 12598 6506 12654 6540
rect 12598 6472 12609 6506
rect 12643 6472 12654 6506
rect 12598 6438 12654 6472
rect 12598 6404 12609 6438
rect 12643 6404 12654 6438
rect 12598 6370 12654 6404
rect 12598 6336 12609 6370
rect 12643 6336 12654 6370
rect 12598 6302 12654 6336
rect 12598 6268 12609 6302
rect 12643 6268 12654 6302
rect 12598 6234 12654 6268
rect 12598 6200 12609 6234
rect 12643 6200 12654 6234
rect 12598 6166 12654 6200
rect 12598 6132 12609 6166
rect 12643 6132 12654 6166
rect 12598 6098 12654 6132
rect 12598 6064 12609 6098
rect 12643 6064 12654 6098
rect 12598 6030 12654 6064
rect 12598 5996 12609 6030
rect 12643 5996 12654 6030
rect 12598 5962 12654 5996
rect 12598 5928 12609 5962
rect 12643 5928 12654 5962
rect 12598 5894 12654 5928
rect 12598 5860 12609 5894
rect 12643 5860 12654 5894
rect 12598 5848 12654 5860
rect 12684 6846 12740 6858
rect 12684 6812 12695 6846
rect 12729 6812 12740 6846
rect 12684 6778 12740 6812
rect 12684 6744 12695 6778
rect 12729 6744 12740 6778
rect 12684 6710 12740 6744
rect 12684 6676 12695 6710
rect 12729 6676 12740 6710
rect 12684 6642 12740 6676
rect 12684 6608 12695 6642
rect 12729 6608 12740 6642
rect 12684 6574 12740 6608
rect 12684 6540 12695 6574
rect 12729 6540 12740 6574
rect 12684 6506 12740 6540
rect 12684 6472 12695 6506
rect 12729 6472 12740 6506
rect 12684 6438 12740 6472
rect 12684 6404 12695 6438
rect 12729 6404 12740 6438
rect 12684 6370 12740 6404
rect 12684 6336 12695 6370
rect 12729 6336 12740 6370
rect 12684 6302 12740 6336
rect 12684 6268 12695 6302
rect 12729 6268 12740 6302
rect 12684 6234 12740 6268
rect 12684 6200 12695 6234
rect 12729 6200 12740 6234
rect 12684 6166 12740 6200
rect 12684 6132 12695 6166
rect 12729 6132 12740 6166
rect 12684 6098 12740 6132
rect 12684 6064 12695 6098
rect 12729 6064 12740 6098
rect 12684 6030 12740 6064
rect 12684 5996 12695 6030
rect 12729 5996 12740 6030
rect 12684 5962 12740 5996
rect 12684 5928 12695 5962
rect 12729 5928 12740 5962
rect 12684 5894 12740 5928
rect 12684 5860 12695 5894
rect 12729 5860 12740 5894
rect 12684 5848 12740 5860
rect 12906 6846 12962 6858
rect 12906 6812 12917 6846
rect 12951 6812 12962 6846
rect 12906 6778 12962 6812
rect 12906 6744 12917 6778
rect 12951 6744 12962 6778
rect 12906 6710 12962 6744
rect 12906 6676 12917 6710
rect 12951 6676 12962 6710
rect 12906 6642 12962 6676
rect 12906 6608 12917 6642
rect 12951 6608 12962 6642
rect 12906 6574 12962 6608
rect 12906 6540 12917 6574
rect 12951 6540 12962 6574
rect 12906 6506 12962 6540
rect 12906 6472 12917 6506
rect 12951 6472 12962 6506
rect 12906 6438 12962 6472
rect 12906 6404 12917 6438
rect 12951 6404 12962 6438
rect 12906 6370 12962 6404
rect 12906 6336 12917 6370
rect 12951 6336 12962 6370
rect 12906 6302 12962 6336
rect 12906 6268 12917 6302
rect 12951 6268 12962 6302
rect 12906 6234 12962 6268
rect 12906 6200 12917 6234
rect 12951 6200 12962 6234
rect 12906 6166 12962 6200
rect 12906 6132 12917 6166
rect 12951 6132 12962 6166
rect 12906 6098 12962 6132
rect 12906 6064 12917 6098
rect 12951 6064 12962 6098
rect 12906 6030 12962 6064
rect 12906 5996 12917 6030
rect 12951 5996 12962 6030
rect 12906 5962 12962 5996
rect 12906 5928 12917 5962
rect 12951 5928 12962 5962
rect 12906 5894 12962 5928
rect 12906 5860 12917 5894
rect 12951 5860 12962 5894
rect 12906 5848 12962 5860
rect 12992 6846 13048 6858
rect 12992 6812 13003 6846
rect 13037 6812 13048 6846
rect 12992 6778 13048 6812
rect 12992 6744 13003 6778
rect 13037 6744 13048 6778
rect 12992 6710 13048 6744
rect 12992 6676 13003 6710
rect 13037 6676 13048 6710
rect 12992 6642 13048 6676
rect 12992 6608 13003 6642
rect 13037 6608 13048 6642
rect 12992 6574 13048 6608
rect 12992 6540 13003 6574
rect 13037 6540 13048 6574
rect 12992 6506 13048 6540
rect 12992 6472 13003 6506
rect 13037 6472 13048 6506
rect 12992 6438 13048 6472
rect 12992 6404 13003 6438
rect 13037 6404 13048 6438
rect 12992 6370 13048 6404
rect 12992 6336 13003 6370
rect 13037 6336 13048 6370
rect 12992 6302 13048 6336
rect 12992 6268 13003 6302
rect 13037 6268 13048 6302
rect 12992 6234 13048 6268
rect 12992 6200 13003 6234
rect 13037 6200 13048 6234
rect 12992 6166 13048 6200
rect 12992 6132 13003 6166
rect 13037 6132 13048 6166
rect 12992 6098 13048 6132
rect 12992 6064 13003 6098
rect 13037 6064 13048 6098
rect 12992 6030 13048 6064
rect 12992 5996 13003 6030
rect 13037 5996 13048 6030
rect 12992 5962 13048 5996
rect 12992 5928 13003 5962
rect 13037 5928 13048 5962
rect 12992 5894 13048 5928
rect 12992 5860 13003 5894
rect 13037 5860 13048 5894
rect 12992 5848 13048 5860
rect 13078 6846 13134 6858
rect 13078 6812 13089 6846
rect 13123 6812 13134 6846
rect 13078 6778 13134 6812
rect 13078 6744 13089 6778
rect 13123 6744 13134 6778
rect 13078 6710 13134 6744
rect 13078 6676 13089 6710
rect 13123 6676 13134 6710
rect 13078 6642 13134 6676
rect 13078 6608 13089 6642
rect 13123 6608 13134 6642
rect 13078 6574 13134 6608
rect 13078 6540 13089 6574
rect 13123 6540 13134 6574
rect 13078 6506 13134 6540
rect 13078 6472 13089 6506
rect 13123 6472 13134 6506
rect 13078 6438 13134 6472
rect 13078 6404 13089 6438
rect 13123 6404 13134 6438
rect 13078 6370 13134 6404
rect 13078 6336 13089 6370
rect 13123 6336 13134 6370
rect 13078 6302 13134 6336
rect 13078 6268 13089 6302
rect 13123 6268 13134 6302
rect 13078 6234 13134 6268
rect 13078 6200 13089 6234
rect 13123 6200 13134 6234
rect 13078 6166 13134 6200
rect 13078 6132 13089 6166
rect 13123 6132 13134 6166
rect 13078 6098 13134 6132
rect 13078 6064 13089 6098
rect 13123 6064 13134 6098
rect 13078 6030 13134 6064
rect 13078 5996 13089 6030
rect 13123 5996 13134 6030
rect 13078 5962 13134 5996
rect 13078 5928 13089 5962
rect 13123 5928 13134 5962
rect 13078 5894 13134 5928
rect 13078 5860 13089 5894
rect 13123 5860 13134 5894
rect 13078 5848 13134 5860
rect 13164 6846 13220 6858
rect 13164 6812 13175 6846
rect 13209 6812 13220 6846
rect 13164 6778 13220 6812
rect 13164 6744 13175 6778
rect 13209 6744 13220 6778
rect 13164 6710 13220 6744
rect 13164 6676 13175 6710
rect 13209 6676 13220 6710
rect 13164 6642 13220 6676
rect 13164 6608 13175 6642
rect 13209 6608 13220 6642
rect 13164 6574 13220 6608
rect 13164 6540 13175 6574
rect 13209 6540 13220 6574
rect 13164 6506 13220 6540
rect 13164 6472 13175 6506
rect 13209 6472 13220 6506
rect 13164 6438 13220 6472
rect 13164 6404 13175 6438
rect 13209 6404 13220 6438
rect 13164 6370 13220 6404
rect 13164 6336 13175 6370
rect 13209 6336 13220 6370
rect 13164 6302 13220 6336
rect 13164 6268 13175 6302
rect 13209 6268 13220 6302
rect 13164 6234 13220 6268
rect 13164 6200 13175 6234
rect 13209 6200 13220 6234
rect 13164 6166 13220 6200
rect 13164 6132 13175 6166
rect 13209 6132 13220 6166
rect 13164 6098 13220 6132
rect 13164 6064 13175 6098
rect 13209 6064 13220 6098
rect 13164 6030 13220 6064
rect 13164 5996 13175 6030
rect 13209 5996 13220 6030
rect 13164 5962 13220 5996
rect 13164 5928 13175 5962
rect 13209 5928 13220 5962
rect 13164 5894 13220 5928
rect 13164 5860 13175 5894
rect 13209 5860 13220 5894
rect 13164 5848 13220 5860
rect 13250 6846 13306 6858
rect 13250 6812 13261 6846
rect 13295 6812 13306 6846
rect 13250 6778 13306 6812
rect 13250 6744 13261 6778
rect 13295 6744 13306 6778
rect 13250 6710 13306 6744
rect 13250 6676 13261 6710
rect 13295 6676 13306 6710
rect 13250 6642 13306 6676
rect 13250 6608 13261 6642
rect 13295 6608 13306 6642
rect 13250 6574 13306 6608
rect 13250 6540 13261 6574
rect 13295 6540 13306 6574
rect 13250 6506 13306 6540
rect 13250 6472 13261 6506
rect 13295 6472 13306 6506
rect 13250 6438 13306 6472
rect 13250 6404 13261 6438
rect 13295 6404 13306 6438
rect 13250 6370 13306 6404
rect 13250 6336 13261 6370
rect 13295 6336 13306 6370
rect 13250 6302 13306 6336
rect 13250 6268 13261 6302
rect 13295 6268 13306 6302
rect 13250 6234 13306 6268
rect 13250 6200 13261 6234
rect 13295 6200 13306 6234
rect 13250 6166 13306 6200
rect 13250 6132 13261 6166
rect 13295 6132 13306 6166
rect 13250 6098 13306 6132
rect 13250 6064 13261 6098
rect 13295 6064 13306 6098
rect 13250 6030 13306 6064
rect 13250 5996 13261 6030
rect 13295 5996 13306 6030
rect 13250 5962 13306 5996
rect 13250 5928 13261 5962
rect 13295 5928 13306 5962
rect 13250 5894 13306 5928
rect 13250 5860 13261 5894
rect 13295 5860 13306 5894
rect 13250 5848 13306 5860
rect 13472 6846 13528 6858
rect 13472 6812 13483 6846
rect 13517 6812 13528 6846
rect 13472 6778 13528 6812
rect 13472 6744 13483 6778
rect 13517 6744 13528 6778
rect 13472 6710 13528 6744
rect 13472 6676 13483 6710
rect 13517 6676 13528 6710
rect 13472 6642 13528 6676
rect 13472 6608 13483 6642
rect 13517 6608 13528 6642
rect 13472 6574 13528 6608
rect 13472 6540 13483 6574
rect 13517 6540 13528 6574
rect 13472 6506 13528 6540
rect 13472 6472 13483 6506
rect 13517 6472 13528 6506
rect 13472 6438 13528 6472
rect 13472 6404 13483 6438
rect 13517 6404 13528 6438
rect 13472 6370 13528 6404
rect 13472 6336 13483 6370
rect 13517 6336 13528 6370
rect 13472 6302 13528 6336
rect 13472 6268 13483 6302
rect 13517 6268 13528 6302
rect 13472 6234 13528 6268
rect 13472 6200 13483 6234
rect 13517 6200 13528 6234
rect 13472 6166 13528 6200
rect 13472 6132 13483 6166
rect 13517 6132 13528 6166
rect 13472 6098 13528 6132
rect 13472 6064 13483 6098
rect 13517 6064 13528 6098
rect 13472 6030 13528 6064
rect 13472 5996 13483 6030
rect 13517 5996 13528 6030
rect 13472 5962 13528 5996
rect 13472 5928 13483 5962
rect 13517 5928 13528 5962
rect 13472 5894 13528 5928
rect 13472 5860 13483 5894
rect 13517 5860 13528 5894
rect 13472 5848 13528 5860
rect 13558 6846 13614 6858
rect 13558 6812 13569 6846
rect 13603 6812 13614 6846
rect 13558 6778 13614 6812
rect 13558 6744 13569 6778
rect 13603 6744 13614 6778
rect 13558 6710 13614 6744
rect 13558 6676 13569 6710
rect 13603 6676 13614 6710
rect 13558 6642 13614 6676
rect 13558 6608 13569 6642
rect 13603 6608 13614 6642
rect 13558 6574 13614 6608
rect 13558 6540 13569 6574
rect 13603 6540 13614 6574
rect 13558 6506 13614 6540
rect 13558 6472 13569 6506
rect 13603 6472 13614 6506
rect 13558 6438 13614 6472
rect 13558 6404 13569 6438
rect 13603 6404 13614 6438
rect 13558 6370 13614 6404
rect 13558 6336 13569 6370
rect 13603 6336 13614 6370
rect 13558 6302 13614 6336
rect 13558 6268 13569 6302
rect 13603 6268 13614 6302
rect 13558 6234 13614 6268
rect 13558 6200 13569 6234
rect 13603 6200 13614 6234
rect 13558 6166 13614 6200
rect 13558 6132 13569 6166
rect 13603 6132 13614 6166
rect 13558 6098 13614 6132
rect 13558 6064 13569 6098
rect 13603 6064 13614 6098
rect 13558 6030 13614 6064
rect 13558 5996 13569 6030
rect 13603 5996 13614 6030
rect 13558 5962 13614 5996
rect 13558 5928 13569 5962
rect 13603 5928 13614 5962
rect 13558 5894 13614 5928
rect 13558 5860 13569 5894
rect 13603 5860 13614 5894
rect 13558 5848 13614 5860
rect 13644 6846 13700 6858
rect 13644 6812 13655 6846
rect 13689 6812 13700 6846
rect 13644 6778 13700 6812
rect 13644 6744 13655 6778
rect 13689 6744 13700 6778
rect 13644 6710 13700 6744
rect 13644 6676 13655 6710
rect 13689 6676 13700 6710
rect 13644 6642 13700 6676
rect 13644 6608 13655 6642
rect 13689 6608 13700 6642
rect 13644 6574 13700 6608
rect 13644 6540 13655 6574
rect 13689 6540 13700 6574
rect 13644 6506 13700 6540
rect 13644 6472 13655 6506
rect 13689 6472 13700 6506
rect 13644 6438 13700 6472
rect 13644 6404 13655 6438
rect 13689 6404 13700 6438
rect 13644 6370 13700 6404
rect 13644 6336 13655 6370
rect 13689 6336 13700 6370
rect 13644 6302 13700 6336
rect 13644 6268 13655 6302
rect 13689 6268 13700 6302
rect 13644 6234 13700 6268
rect 13644 6200 13655 6234
rect 13689 6200 13700 6234
rect 13644 6166 13700 6200
rect 13644 6132 13655 6166
rect 13689 6132 13700 6166
rect 13644 6098 13700 6132
rect 13644 6064 13655 6098
rect 13689 6064 13700 6098
rect 13644 6030 13700 6064
rect 13644 5996 13655 6030
rect 13689 5996 13700 6030
rect 13644 5962 13700 5996
rect 13644 5928 13655 5962
rect 13689 5928 13700 5962
rect 13644 5894 13700 5928
rect 13644 5860 13655 5894
rect 13689 5860 13700 5894
rect 13644 5848 13700 5860
rect 13730 6846 13786 6858
rect 13730 6812 13741 6846
rect 13775 6812 13786 6846
rect 13730 6778 13786 6812
rect 13730 6744 13741 6778
rect 13775 6744 13786 6778
rect 13730 6710 13786 6744
rect 13730 6676 13741 6710
rect 13775 6676 13786 6710
rect 13730 6642 13786 6676
rect 13730 6608 13741 6642
rect 13775 6608 13786 6642
rect 13730 6574 13786 6608
rect 13730 6540 13741 6574
rect 13775 6540 13786 6574
rect 13730 6506 13786 6540
rect 13730 6472 13741 6506
rect 13775 6472 13786 6506
rect 13730 6438 13786 6472
rect 13730 6404 13741 6438
rect 13775 6404 13786 6438
rect 13730 6370 13786 6404
rect 13730 6336 13741 6370
rect 13775 6336 13786 6370
rect 13730 6302 13786 6336
rect 13730 6268 13741 6302
rect 13775 6268 13786 6302
rect 13730 6234 13786 6268
rect 13730 6200 13741 6234
rect 13775 6200 13786 6234
rect 13730 6166 13786 6200
rect 13730 6132 13741 6166
rect 13775 6132 13786 6166
rect 13730 6098 13786 6132
rect 13730 6064 13741 6098
rect 13775 6064 13786 6098
rect 13730 6030 13786 6064
rect 13730 5996 13741 6030
rect 13775 5996 13786 6030
rect 13730 5962 13786 5996
rect 13730 5928 13741 5962
rect 13775 5928 13786 5962
rect 13730 5894 13786 5928
rect 13730 5860 13741 5894
rect 13775 5860 13786 5894
rect 13730 5848 13786 5860
rect 13816 6846 13872 6858
rect 13816 6812 13827 6846
rect 13861 6812 13872 6846
rect 13816 6778 13872 6812
rect 13816 6744 13827 6778
rect 13861 6744 13872 6778
rect 13816 6710 13872 6744
rect 13816 6676 13827 6710
rect 13861 6676 13872 6710
rect 13816 6642 13872 6676
rect 13816 6608 13827 6642
rect 13861 6608 13872 6642
rect 13816 6574 13872 6608
rect 13816 6540 13827 6574
rect 13861 6540 13872 6574
rect 13816 6506 13872 6540
rect 13816 6472 13827 6506
rect 13861 6472 13872 6506
rect 13816 6438 13872 6472
rect 13816 6404 13827 6438
rect 13861 6404 13872 6438
rect 13816 6370 13872 6404
rect 13816 6336 13827 6370
rect 13861 6336 13872 6370
rect 13816 6302 13872 6336
rect 13816 6268 13827 6302
rect 13861 6268 13872 6302
rect 13816 6234 13872 6268
rect 13816 6200 13827 6234
rect 13861 6200 13872 6234
rect 13816 6166 13872 6200
rect 13816 6132 13827 6166
rect 13861 6132 13872 6166
rect 13816 6098 13872 6132
rect 13816 6064 13827 6098
rect 13861 6064 13872 6098
rect 13816 6030 13872 6064
rect 13816 5996 13827 6030
rect 13861 5996 13872 6030
rect 13816 5962 13872 5996
rect 13816 5928 13827 5962
rect 13861 5928 13872 5962
rect 13816 5894 13872 5928
rect 13816 5860 13827 5894
rect 13861 5860 13872 5894
rect 13816 5848 13872 5860
rect 14038 6846 14094 6858
rect 14038 6812 14049 6846
rect 14083 6812 14094 6846
rect 14038 6778 14094 6812
rect 14038 6744 14049 6778
rect 14083 6744 14094 6778
rect 14038 6710 14094 6744
rect 14038 6676 14049 6710
rect 14083 6676 14094 6710
rect 14038 6642 14094 6676
rect 14038 6608 14049 6642
rect 14083 6608 14094 6642
rect 14038 6574 14094 6608
rect 14038 6540 14049 6574
rect 14083 6540 14094 6574
rect 14038 6506 14094 6540
rect 14038 6472 14049 6506
rect 14083 6472 14094 6506
rect 14038 6438 14094 6472
rect 14038 6404 14049 6438
rect 14083 6404 14094 6438
rect 14038 6370 14094 6404
rect 14038 6336 14049 6370
rect 14083 6336 14094 6370
rect 14038 6302 14094 6336
rect 14038 6268 14049 6302
rect 14083 6268 14094 6302
rect 14038 6234 14094 6268
rect 14038 6200 14049 6234
rect 14083 6200 14094 6234
rect 14038 6166 14094 6200
rect 14038 6132 14049 6166
rect 14083 6132 14094 6166
rect 14038 6098 14094 6132
rect 14038 6064 14049 6098
rect 14083 6064 14094 6098
rect 14038 6030 14094 6064
rect 14038 5996 14049 6030
rect 14083 5996 14094 6030
rect 14038 5962 14094 5996
rect 14038 5928 14049 5962
rect 14083 5928 14094 5962
rect 14038 5894 14094 5928
rect 14038 5860 14049 5894
rect 14083 5860 14094 5894
rect 14038 5848 14094 5860
rect 14124 6846 14180 6858
rect 14124 6812 14135 6846
rect 14169 6812 14180 6846
rect 14124 6778 14180 6812
rect 14124 6744 14135 6778
rect 14169 6744 14180 6778
rect 14124 6710 14180 6744
rect 14124 6676 14135 6710
rect 14169 6676 14180 6710
rect 14124 6642 14180 6676
rect 14124 6608 14135 6642
rect 14169 6608 14180 6642
rect 14124 6574 14180 6608
rect 14124 6540 14135 6574
rect 14169 6540 14180 6574
rect 14124 6506 14180 6540
rect 14124 6472 14135 6506
rect 14169 6472 14180 6506
rect 14124 6438 14180 6472
rect 14124 6404 14135 6438
rect 14169 6404 14180 6438
rect 14124 6370 14180 6404
rect 14124 6336 14135 6370
rect 14169 6336 14180 6370
rect 14124 6302 14180 6336
rect 14124 6268 14135 6302
rect 14169 6268 14180 6302
rect 14124 6234 14180 6268
rect 14124 6200 14135 6234
rect 14169 6200 14180 6234
rect 14124 6166 14180 6200
rect 14124 6132 14135 6166
rect 14169 6132 14180 6166
rect 14124 6098 14180 6132
rect 14124 6064 14135 6098
rect 14169 6064 14180 6098
rect 14124 6030 14180 6064
rect 14124 5996 14135 6030
rect 14169 5996 14180 6030
rect 14124 5962 14180 5996
rect 14124 5928 14135 5962
rect 14169 5928 14180 5962
rect 14124 5894 14180 5928
rect 14124 5860 14135 5894
rect 14169 5860 14180 5894
rect 14124 5848 14180 5860
rect 14210 6846 14266 6858
rect 14210 6812 14221 6846
rect 14255 6812 14266 6846
rect 14210 6778 14266 6812
rect 14210 6744 14221 6778
rect 14255 6744 14266 6778
rect 14210 6710 14266 6744
rect 14210 6676 14221 6710
rect 14255 6676 14266 6710
rect 14210 6642 14266 6676
rect 14210 6608 14221 6642
rect 14255 6608 14266 6642
rect 14210 6574 14266 6608
rect 14210 6540 14221 6574
rect 14255 6540 14266 6574
rect 14210 6506 14266 6540
rect 14210 6472 14221 6506
rect 14255 6472 14266 6506
rect 14210 6438 14266 6472
rect 14210 6404 14221 6438
rect 14255 6404 14266 6438
rect 14210 6370 14266 6404
rect 14210 6336 14221 6370
rect 14255 6336 14266 6370
rect 14210 6302 14266 6336
rect 14210 6268 14221 6302
rect 14255 6268 14266 6302
rect 14210 6234 14266 6268
rect 14210 6200 14221 6234
rect 14255 6200 14266 6234
rect 14210 6166 14266 6200
rect 14210 6132 14221 6166
rect 14255 6132 14266 6166
rect 14210 6098 14266 6132
rect 14210 6064 14221 6098
rect 14255 6064 14266 6098
rect 14210 6030 14266 6064
rect 14210 5996 14221 6030
rect 14255 5996 14266 6030
rect 14210 5962 14266 5996
rect 14210 5928 14221 5962
rect 14255 5928 14266 5962
rect 14210 5894 14266 5928
rect 14210 5860 14221 5894
rect 14255 5860 14266 5894
rect 14210 5848 14266 5860
rect 14296 6846 14352 6858
rect 14296 6812 14307 6846
rect 14341 6812 14352 6846
rect 14296 6778 14352 6812
rect 14296 6744 14307 6778
rect 14341 6744 14352 6778
rect 14296 6710 14352 6744
rect 14296 6676 14307 6710
rect 14341 6676 14352 6710
rect 14296 6642 14352 6676
rect 14296 6608 14307 6642
rect 14341 6608 14352 6642
rect 14296 6574 14352 6608
rect 14296 6540 14307 6574
rect 14341 6540 14352 6574
rect 14296 6506 14352 6540
rect 14296 6472 14307 6506
rect 14341 6472 14352 6506
rect 14296 6438 14352 6472
rect 14296 6404 14307 6438
rect 14341 6404 14352 6438
rect 14296 6370 14352 6404
rect 14296 6336 14307 6370
rect 14341 6336 14352 6370
rect 14296 6302 14352 6336
rect 14296 6268 14307 6302
rect 14341 6268 14352 6302
rect 14296 6234 14352 6268
rect 14296 6200 14307 6234
rect 14341 6200 14352 6234
rect 14296 6166 14352 6200
rect 14296 6132 14307 6166
rect 14341 6132 14352 6166
rect 14296 6098 14352 6132
rect 14296 6064 14307 6098
rect 14341 6064 14352 6098
rect 14296 6030 14352 6064
rect 14296 5996 14307 6030
rect 14341 5996 14352 6030
rect 14296 5962 14352 5996
rect 14296 5928 14307 5962
rect 14341 5928 14352 5962
rect 14296 5894 14352 5928
rect 14296 5860 14307 5894
rect 14341 5860 14352 5894
rect 14296 5848 14352 5860
rect 14382 6846 14438 6858
rect 14382 6812 14393 6846
rect 14427 6812 14438 6846
rect 14382 6778 14438 6812
rect 14382 6744 14393 6778
rect 14427 6744 14438 6778
rect 14382 6710 14438 6744
rect 14382 6676 14393 6710
rect 14427 6676 14438 6710
rect 14382 6642 14438 6676
rect 14382 6608 14393 6642
rect 14427 6608 14438 6642
rect 14382 6574 14438 6608
rect 14382 6540 14393 6574
rect 14427 6540 14438 6574
rect 14382 6506 14438 6540
rect 14382 6472 14393 6506
rect 14427 6472 14438 6506
rect 14382 6438 14438 6472
rect 14382 6404 14393 6438
rect 14427 6404 14438 6438
rect 14382 6370 14438 6404
rect 14382 6336 14393 6370
rect 14427 6336 14438 6370
rect 14382 6302 14438 6336
rect 14382 6268 14393 6302
rect 14427 6268 14438 6302
rect 14382 6234 14438 6268
rect 14382 6200 14393 6234
rect 14427 6200 14438 6234
rect 14382 6166 14438 6200
rect 14382 6132 14393 6166
rect 14427 6132 14438 6166
rect 14382 6098 14438 6132
rect 14382 6064 14393 6098
rect 14427 6064 14438 6098
rect 14382 6030 14438 6064
rect 14382 5996 14393 6030
rect 14427 5996 14438 6030
rect 14382 5962 14438 5996
rect 14382 5928 14393 5962
rect 14427 5928 14438 5962
rect 14382 5894 14438 5928
rect 14382 5860 14393 5894
rect 14427 5860 14438 5894
rect 14382 5848 14438 5860
rect 14604 6846 14660 6858
rect 14604 6812 14615 6846
rect 14649 6812 14660 6846
rect 14604 6778 14660 6812
rect 14604 6744 14615 6778
rect 14649 6744 14660 6778
rect 14604 6710 14660 6744
rect 14604 6676 14615 6710
rect 14649 6676 14660 6710
rect 14604 6642 14660 6676
rect 14604 6608 14615 6642
rect 14649 6608 14660 6642
rect 14604 6574 14660 6608
rect 14604 6540 14615 6574
rect 14649 6540 14660 6574
rect 14604 6506 14660 6540
rect 14604 6472 14615 6506
rect 14649 6472 14660 6506
rect 14604 6438 14660 6472
rect 14604 6404 14615 6438
rect 14649 6404 14660 6438
rect 14604 6370 14660 6404
rect 14604 6336 14615 6370
rect 14649 6336 14660 6370
rect 14604 6302 14660 6336
rect 14604 6268 14615 6302
rect 14649 6268 14660 6302
rect 14604 6234 14660 6268
rect 14604 6200 14615 6234
rect 14649 6200 14660 6234
rect 14604 6166 14660 6200
rect 14604 6132 14615 6166
rect 14649 6132 14660 6166
rect 14604 6098 14660 6132
rect 14604 6064 14615 6098
rect 14649 6064 14660 6098
rect 14604 6030 14660 6064
rect 14604 5996 14615 6030
rect 14649 5996 14660 6030
rect 14604 5962 14660 5996
rect 14604 5928 14615 5962
rect 14649 5928 14660 5962
rect 14604 5894 14660 5928
rect 14604 5860 14615 5894
rect 14649 5860 14660 5894
rect 14604 5848 14660 5860
rect 14690 6846 14746 6858
rect 14690 6812 14701 6846
rect 14735 6812 14746 6846
rect 14690 6778 14746 6812
rect 14690 6744 14701 6778
rect 14735 6744 14746 6778
rect 14690 6710 14746 6744
rect 14690 6676 14701 6710
rect 14735 6676 14746 6710
rect 14690 6642 14746 6676
rect 14690 6608 14701 6642
rect 14735 6608 14746 6642
rect 14690 6574 14746 6608
rect 14690 6540 14701 6574
rect 14735 6540 14746 6574
rect 14690 6506 14746 6540
rect 14690 6472 14701 6506
rect 14735 6472 14746 6506
rect 14690 6438 14746 6472
rect 14690 6404 14701 6438
rect 14735 6404 14746 6438
rect 14690 6370 14746 6404
rect 14690 6336 14701 6370
rect 14735 6336 14746 6370
rect 14690 6302 14746 6336
rect 14690 6268 14701 6302
rect 14735 6268 14746 6302
rect 14690 6234 14746 6268
rect 14690 6200 14701 6234
rect 14735 6200 14746 6234
rect 14690 6166 14746 6200
rect 14690 6132 14701 6166
rect 14735 6132 14746 6166
rect 14690 6098 14746 6132
rect 14690 6064 14701 6098
rect 14735 6064 14746 6098
rect 14690 6030 14746 6064
rect 14690 5996 14701 6030
rect 14735 5996 14746 6030
rect 14690 5962 14746 5996
rect 14690 5928 14701 5962
rect 14735 5928 14746 5962
rect 14690 5894 14746 5928
rect 14690 5860 14701 5894
rect 14735 5860 14746 5894
rect 14690 5848 14746 5860
rect 14776 6846 14832 6858
rect 14776 6812 14787 6846
rect 14821 6812 14832 6846
rect 14776 6778 14832 6812
rect 14776 6744 14787 6778
rect 14821 6744 14832 6778
rect 14776 6710 14832 6744
rect 14776 6676 14787 6710
rect 14821 6676 14832 6710
rect 14776 6642 14832 6676
rect 14776 6608 14787 6642
rect 14821 6608 14832 6642
rect 14776 6574 14832 6608
rect 14776 6540 14787 6574
rect 14821 6540 14832 6574
rect 14776 6506 14832 6540
rect 14776 6472 14787 6506
rect 14821 6472 14832 6506
rect 14776 6438 14832 6472
rect 14776 6404 14787 6438
rect 14821 6404 14832 6438
rect 14776 6370 14832 6404
rect 14776 6336 14787 6370
rect 14821 6336 14832 6370
rect 14776 6302 14832 6336
rect 14776 6268 14787 6302
rect 14821 6268 14832 6302
rect 14776 6234 14832 6268
rect 14776 6200 14787 6234
rect 14821 6200 14832 6234
rect 14776 6166 14832 6200
rect 14776 6132 14787 6166
rect 14821 6132 14832 6166
rect 14776 6098 14832 6132
rect 14776 6064 14787 6098
rect 14821 6064 14832 6098
rect 14776 6030 14832 6064
rect 14776 5996 14787 6030
rect 14821 5996 14832 6030
rect 14776 5962 14832 5996
rect 14776 5928 14787 5962
rect 14821 5928 14832 5962
rect 14776 5894 14832 5928
rect 14776 5860 14787 5894
rect 14821 5860 14832 5894
rect 14776 5848 14832 5860
rect 14862 6846 14918 6858
rect 14862 6812 14873 6846
rect 14907 6812 14918 6846
rect 14862 6778 14918 6812
rect 14862 6744 14873 6778
rect 14907 6744 14918 6778
rect 14862 6710 14918 6744
rect 14862 6676 14873 6710
rect 14907 6676 14918 6710
rect 14862 6642 14918 6676
rect 14862 6608 14873 6642
rect 14907 6608 14918 6642
rect 14862 6574 14918 6608
rect 14862 6540 14873 6574
rect 14907 6540 14918 6574
rect 14862 6506 14918 6540
rect 14862 6472 14873 6506
rect 14907 6472 14918 6506
rect 14862 6438 14918 6472
rect 14862 6404 14873 6438
rect 14907 6404 14918 6438
rect 14862 6370 14918 6404
rect 14862 6336 14873 6370
rect 14907 6336 14918 6370
rect 14862 6302 14918 6336
rect 14862 6268 14873 6302
rect 14907 6268 14918 6302
rect 14862 6234 14918 6268
rect 14862 6200 14873 6234
rect 14907 6200 14918 6234
rect 14862 6166 14918 6200
rect 14862 6132 14873 6166
rect 14907 6132 14918 6166
rect 14862 6098 14918 6132
rect 14862 6064 14873 6098
rect 14907 6064 14918 6098
rect 14862 6030 14918 6064
rect 14862 5996 14873 6030
rect 14907 5996 14918 6030
rect 14862 5962 14918 5996
rect 14862 5928 14873 5962
rect 14907 5928 14918 5962
rect 14862 5894 14918 5928
rect 14862 5860 14873 5894
rect 14907 5860 14918 5894
rect 14862 5848 14918 5860
rect 14948 6846 15004 6858
rect 14948 6812 14959 6846
rect 14993 6812 15004 6846
rect 14948 6778 15004 6812
rect 14948 6744 14959 6778
rect 14993 6744 15004 6778
rect 14948 6710 15004 6744
rect 14948 6676 14959 6710
rect 14993 6676 15004 6710
rect 14948 6642 15004 6676
rect 14948 6608 14959 6642
rect 14993 6608 15004 6642
rect 14948 6574 15004 6608
rect 14948 6540 14959 6574
rect 14993 6540 15004 6574
rect 14948 6506 15004 6540
rect 14948 6472 14959 6506
rect 14993 6472 15004 6506
rect 14948 6438 15004 6472
rect 14948 6404 14959 6438
rect 14993 6404 15004 6438
rect 14948 6370 15004 6404
rect 14948 6336 14959 6370
rect 14993 6336 15004 6370
rect 14948 6302 15004 6336
rect 14948 6268 14959 6302
rect 14993 6268 15004 6302
rect 14948 6234 15004 6268
rect 14948 6200 14959 6234
rect 14993 6200 15004 6234
rect 14948 6166 15004 6200
rect 14948 6132 14959 6166
rect 14993 6132 15004 6166
rect 14948 6098 15004 6132
rect 14948 6064 14959 6098
rect 14993 6064 15004 6098
rect 14948 6030 15004 6064
rect 14948 5996 14959 6030
rect 14993 5996 15004 6030
rect 14948 5962 15004 5996
rect 14948 5928 14959 5962
rect 14993 5928 15004 5962
rect 14948 5894 15004 5928
rect 14948 5860 14959 5894
rect 14993 5860 15004 5894
rect 14948 5848 15004 5860
rect 15170 6846 15226 6858
rect 15170 6812 15181 6846
rect 15215 6812 15226 6846
rect 15170 6778 15226 6812
rect 15170 6744 15181 6778
rect 15215 6744 15226 6778
rect 15170 6710 15226 6744
rect 15170 6676 15181 6710
rect 15215 6676 15226 6710
rect 15170 6642 15226 6676
rect 15170 6608 15181 6642
rect 15215 6608 15226 6642
rect 15170 6574 15226 6608
rect 15170 6540 15181 6574
rect 15215 6540 15226 6574
rect 15170 6506 15226 6540
rect 15170 6472 15181 6506
rect 15215 6472 15226 6506
rect 15170 6438 15226 6472
rect 15170 6404 15181 6438
rect 15215 6404 15226 6438
rect 15170 6370 15226 6404
rect 15170 6336 15181 6370
rect 15215 6336 15226 6370
rect 15170 6302 15226 6336
rect 15170 6268 15181 6302
rect 15215 6268 15226 6302
rect 15170 6234 15226 6268
rect 15170 6200 15181 6234
rect 15215 6200 15226 6234
rect 15170 6166 15226 6200
rect 15170 6132 15181 6166
rect 15215 6132 15226 6166
rect 15170 6098 15226 6132
rect 15170 6064 15181 6098
rect 15215 6064 15226 6098
rect 15170 6030 15226 6064
rect 15170 5996 15181 6030
rect 15215 5996 15226 6030
rect 15170 5962 15226 5996
rect 15170 5928 15181 5962
rect 15215 5928 15226 5962
rect 15170 5894 15226 5928
rect 15170 5860 15181 5894
rect 15215 5860 15226 5894
rect 15170 5848 15226 5860
rect 15256 6846 15312 6858
rect 15256 6812 15267 6846
rect 15301 6812 15312 6846
rect 15256 6778 15312 6812
rect 15256 6744 15267 6778
rect 15301 6744 15312 6778
rect 15256 6710 15312 6744
rect 15256 6676 15267 6710
rect 15301 6676 15312 6710
rect 15256 6642 15312 6676
rect 15256 6608 15267 6642
rect 15301 6608 15312 6642
rect 15256 6574 15312 6608
rect 15256 6540 15267 6574
rect 15301 6540 15312 6574
rect 15256 6506 15312 6540
rect 15256 6472 15267 6506
rect 15301 6472 15312 6506
rect 15256 6438 15312 6472
rect 15256 6404 15267 6438
rect 15301 6404 15312 6438
rect 15256 6370 15312 6404
rect 15256 6336 15267 6370
rect 15301 6336 15312 6370
rect 15256 6302 15312 6336
rect 15256 6268 15267 6302
rect 15301 6268 15312 6302
rect 15256 6234 15312 6268
rect 15256 6200 15267 6234
rect 15301 6200 15312 6234
rect 15256 6166 15312 6200
rect 15256 6132 15267 6166
rect 15301 6132 15312 6166
rect 15256 6098 15312 6132
rect 15256 6064 15267 6098
rect 15301 6064 15312 6098
rect 15256 6030 15312 6064
rect 15256 5996 15267 6030
rect 15301 5996 15312 6030
rect 15256 5962 15312 5996
rect 15256 5928 15267 5962
rect 15301 5928 15312 5962
rect 15256 5894 15312 5928
rect 15256 5860 15267 5894
rect 15301 5860 15312 5894
rect 15256 5848 15312 5860
rect 15342 6846 15398 6858
rect 15342 6812 15353 6846
rect 15387 6812 15398 6846
rect 15342 6778 15398 6812
rect 15342 6744 15353 6778
rect 15387 6744 15398 6778
rect 15342 6710 15398 6744
rect 15342 6676 15353 6710
rect 15387 6676 15398 6710
rect 15342 6642 15398 6676
rect 15342 6608 15353 6642
rect 15387 6608 15398 6642
rect 15342 6574 15398 6608
rect 15342 6540 15353 6574
rect 15387 6540 15398 6574
rect 15342 6506 15398 6540
rect 15342 6472 15353 6506
rect 15387 6472 15398 6506
rect 15342 6438 15398 6472
rect 15342 6404 15353 6438
rect 15387 6404 15398 6438
rect 15342 6370 15398 6404
rect 15342 6336 15353 6370
rect 15387 6336 15398 6370
rect 15342 6302 15398 6336
rect 15342 6268 15353 6302
rect 15387 6268 15398 6302
rect 15342 6234 15398 6268
rect 15342 6200 15353 6234
rect 15387 6200 15398 6234
rect 15342 6166 15398 6200
rect 15342 6132 15353 6166
rect 15387 6132 15398 6166
rect 15342 6098 15398 6132
rect 15342 6064 15353 6098
rect 15387 6064 15398 6098
rect 15342 6030 15398 6064
rect 15342 5996 15353 6030
rect 15387 5996 15398 6030
rect 15342 5962 15398 5996
rect 15342 5928 15353 5962
rect 15387 5928 15398 5962
rect 15342 5894 15398 5928
rect 15342 5860 15353 5894
rect 15387 5860 15398 5894
rect 15342 5848 15398 5860
rect 15428 6846 15484 6858
rect 15428 6812 15439 6846
rect 15473 6812 15484 6846
rect 15428 6778 15484 6812
rect 15428 6744 15439 6778
rect 15473 6744 15484 6778
rect 15428 6710 15484 6744
rect 15428 6676 15439 6710
rect 15473 6676 15484 6710
rect 15428 6642 15484 6676
rect 15428 6608 15439 6642
rect 15473 6608 15484 6642
rect 15428 6574 15484 6608
rect 15428 6540 15439 6574
rect 15473 6540 15484 6574
rect 15428 6506 15484 6540
rect 15428 6472 15439 6506
rect 15473 6472 15484 6506
rect 15428 6438 15484 6472
rect 15428 6404 15439 6438
rect 15473 6404 15484 6438
rect 15428 6370 15484 6404
rect 15428 6336 15439 6370
rect 15473 6336 15484 6370
rect 15428 6302 15484 6336
rect 15428 6268 15439 6302
rect 15473 6268 15484 6302
rect 15428 6234 15484 6268
rect 15428 6200 15439 6234
rect 15473 6200 15484 6234
rect 15428 6166 15484 6200
rect 15428 6132 15439 6166
rect 15473 6132 15484 6166
rect 15428 6098 15484 6132
rect 15428 6064 15439 6098
rect 15473 6064 15484 6098
rect 15428 6030 15484 6064
rect 15428 5996 15439 6030
rect 15473 5996 15484 6030
rect 15428 5962 15484 5996
rect 15428 5928 15439 5962
rect 15473 5928 15484 5962
rect 15428 5894 15484 5928
rect 15428 5860 15439 5894
rect 15473 5860 15484 5894
rect 15428 5848 15484 5860
rect 15514 6846 15570 6858
rect 15514 6812 15525 6846
rect 15559 6812 15570 6846
rect 15514 6778 15570 6812
rect 15514 6744 15525 6778
rect 15559 6744 15570 6778
rect 15514 6710 15570 6744
rect 15514 6676 15525 6710
rect 15559 6676 15570 6710
rect 15514 6642 15570 6676
rect 15514 6608 15525 6642
rect 15559 6608 15570 6642
rect 15514 6574 15570 6608
rect 15514 6540 15525 6574
rect 15559 6540 15570 6574
rect 15514 6506 15570 6540
rect 15514 6472 15525 6506
rect 15559 6472 15570 6506
rect 15514 6438 15570 6472
rect 15514 6404 15525 6438
rect 15559 6404 15570 6438
rect 15514 6370 15570 6404
rect 15514 6336 15525 6370
rect 15559 6336 15570 6370
rect 15514 6302 15570 6336
rect 15514 6268 15525 6302
rect 15559 6268 15570 6302
rect 15514 6234 15570 6268
rect 15514 6200 15525 6234
rect 15559 6200 15570 6234
rect 15514 6166 15570 6200
rect 15514 6132 15525 6166
rect 15559 6132 15570 6166
rect 15514 6098 15570 6132
rect 15514 6064 15525 6098
rect 15559 6064 15570 6098
rect 15514 6030 15570 6064
rect 15514 5996 15525 6030
rect 15559 5996 15570 6030
rect 15514 5962 15570 5996
rect 15514 5928 15525 5962
rect 15559 5928 15570 5962
rect 15514 5894 15570 5928
rect 15514 5860 15525 5894
rect 15559 5860 15570 5894
rect 15514 5848 15570 5860
rect 16107 6179 16163 6191
rect 16107 6145 16118 6179
rect 16152 6145 16163 6179
rect 16107 6111 16163 6145
rect 16107 6077 16118 6111
rect 16152 6077 16163 6111
rect 16107 6043 16163 6077
rect 16107 6009 16118 6043
rect 16152 6009 16163 6043
rect 16107 5975 16163 6009
rect 16107 5941 16118 5975
rect 16152 5941 16163 5975
rect 16107 5907 16163 5941
rect 16107 5873 16118 5907
rect 16152 5873 16163 5907
rect 16107 5839 16163 5873
rect 16107 5805 16118 5839
rect 16152 5805 16163 5839
rect 16107 5771 16163 5805
rect 16107 5737 16118 5771
rect 16152 5737 16163 5771
rect 16107 5703 16163 5737
rect 16107 5669 16118 5703
rect 16152 5669 16163 5703
rect 16107 5635 16163 5669
rect 16107 5601 16118 5635
rect 16152 5601 16163 5635
rect 16107 5567 16163 5601
rect 16107 5533 16118 5567
rect 16152 5533 16163 5567
rect 16107 5499 16163 5533
rect 16107 5465 16118 5499
rect 16152 5465 16163 5499
rect 16107 5431 16163 5465
rect 16107 5397 16118 5431
rect 16152 5397 16163 5431
rect 16107 5363 16163 5397
rect 16107 5329 16118 5363
rect 16152 5329 16163 5363
rect 16107 5295 16163 5329
rect 16107 5261 16118 5295
rect 16152 5261 16163 5295
rect 16107 5227 16163 5261
rect 16107 5193 16118 5227
rect 16152 5193 16163 5227
rect 16107 5181 16163 5193
rect 16193 6179 16249 6191
rect 16193 6145 16204 6179
rect 16238 6145 16249 6179
rect 16193 6111 16249 6145
rect 16193 6077 16204 6111
rect 16238 6077 16249 6111
rect 16193 6043 16249 6077
rect 16193 6009 16204 6043
rect 16238 6009 16249 6043
rect 16193 5975 16249 6009
rect 16193 5941 16204 5975
rect 16238 5941 16249 5975
rect 16193 5907 16249 5941
rect 16193 5873 16204 5907
rect 16238 5873 16249 5907
rect 16193 5839 16249 5873
rect 16193 5805 16204 5839
rect 16238 5805 16249 5839
rect 16193 5771 16249 5805
rect 16193 5737 16204 5771
rect 16238 5737 16249 5771
rect 16193 5703 16249 5737
rect 16193 5669 16204 5703
rect 16238 5669 16249 5703
rect 16193 5635 16249 5669
rect 16193 5601 16204 5635
rect 16238 5601 16249 5635
rect 16193 5567 16249 5601
rect 16193 5533 16204 5567
rect 16238 5533 16249 5567
rect 16193 5499 16249 5533
rect 16193 5465 16204 5499
rect 16238 5465 16249 5499
rect 16193 5431 16249 5465
rect 16193 5397 16204 5431
rect 16238 5397 16249 5431
rect 16193 5363 16249 5397
rect 16193 5329 16204 5363
rect 16238 5329 16249 5363
rect 16193 5295 16249 5329
rect 16193 5261 16204 5295
rect 16238 5261 16249 5295
rect 16193 5227 16249 5261
rect 16193 5193 16204 5227
rect 16238 5193 16249 5227
rect 16193 5181 16249 5193
rect 16279 6179 16335 6191
rect 16279 6145 16290 6179
rect 16324 6145 16335 6179
rect 16279 6111 16335 6145
rect 16279 6077 16290 6111
rect 16324 6077 16335 6111
rect 16279 6043 16335 6077
rect 16279 6009 16290 6043
rect 16324 6009 16335 6043
rect 16279 5975 16335 6009
rect 16279 5941 16290 5975
rect 16324 5941 16335 5975
rect 16279 5907 16335 5941
rect 16279 5873 16290 5907
rect 16324 5873 16335 5907
rect 16279 5839 16335 5873
rect 16279 5805 16290 5839
rect 16324 5805 16335 5839
rect 16279 5771 16335 5805
rect 16279 5737 16290 5771
rect 16324 5737 16335 5771
rect 16279 5703 16335 5737
rect 16279 5669 16290 5703
rect 16324 5669 16335 5703
rect 16279 5635 16335 5669
rect 16279 5601 16290 5635
rect 16324 5601 16335 5635
rect 16279 5567 16335 5601
rect 16279 5533 16290 5567
rect 16324 5533 16335 5567
rect 16279 5499 16335 5533
rect 16279 5465 16290 5499
rect 16324 5465 16335 5499
rect 16279 5431 16335 5465
rect 16279 5397 16290 5431
rect 16324 5397 16335 5431
rect 16279 5363 16335 5397
rect 16279 5329 16290 5363
rect 16324 5329 16335 5363
rect 16279 5295 16335 5329
rect 16279 5261 16290 5295
rect 16324 5261 16335 5295
rect 16279 5227 16335 5261
rect 16279 5193 16290 5227
rect 16324 5193 16335 5227
rect 16279 5181 16335 5193
rect 16365 6179 16421 6191
rect 16365 6145 16376 6179
rect 16410 6145 16421 6179
rect 16365 6111 16421 6145
rect 16365 6077 16376 6111
rect 16410 6077 16421 6111
rect 16365 6043 16421 6077
rect 16365 6009 16376 6043
rect 16410 6009 16421 6043
rect 16365 5975 16421 6009
rect 16365 5941 16376 5975
rect 16410 5941 16421 5975
rect 16365 5907 16421 5941
rect 16365 5873 16376 5907
rect 16410 5873 16421 5907
rect 16365 5839 16421 5873
rect 16365 5805 16376 5839
rect 16410 5805 16421 5839
rect 16365 5771 16421 5805
rect 16365 5737 16376 5771
rect 16410 5737 16421 5771
rect 16365 5703 16421 5737
rect 16365 5669 16376 5703
rect 16410 5669 16421 5703
rect 16365 5635 16421 5669
rect 16365 5601 16376 5635
rect 16410 5601 16421 5635
rect 16365 5567 16421 5601
rect 16365 5533 16376 5567
rect 16410 5533 16421 5567
rect 16365 5499 16421 5533
rect 16365 5465 16376 5499
rect 16410 5465 16421 5499
rect 16365 5431 16421 5465
rect 16365 5397 16376 5431
rect 16410 5397 16421 5431
rect 16365 5363 16421 5397
rect 16365 5329 16376 5363
rect 16410 5329 16421 5363
rect 16365 5295 16421 5329
rect 16365 5261 16376 5295
rect 16410 5261 16421 5295
rect 16365 5227 16421 5261
rect 16365 5193 16376 5227
rect 16410 5193 16421 5227
rect 16365 5181 16421 5193
rect 16451 6179 16507 6191
rect 16451 6145 16462 6179
rect 16496 6145 16507 6179
rect 16451 6111 16507 6145
rect 16451 6077 16462 6111
rect 16496 6077 16507 6111
rect 16451 6043 16507 6077
rect 16451 6009 16462 6043
rect 16496 6009 16507 6043
rect 16451 5975 16507 6009
rect 16451 5941 16462 5975
rect 16496 5941 16507 5975
rect 16451 5907 16507 5941
rect 16451 5873 16462 5907
rect 16496 5873 16507 5907
rect 16451 5839 16507 5873
rect 16451 5805 16462 5839
rect 16496 5805 16507 5839
rect 16451 5771 16507 5805
rect 16451 5737 16462 5771
rect 16496 5737 16507 5771
rect 16451 5703 16507 5737
rect 16451 5669 16462 5703
rect 16496 5669 16507 5703
rect 16451 5635 16507 5669
rect 16451 5601 16462 5635
rect 16496 5601 16507 5635
rect 16451 5567 16507 5601
rect 16451 5533 16462 5567
rect 16496 5533 16507 5567
rect 16451 5499 16507 5533
rect 16451 5465 16462 5499
rect 16496 5465 16507 5499
rect 16451 5431 16507 5465
rect 16451 5397 16462 5431
rect 16496 5397 16507 5431
rect 16451 5363 16507 5397
rect 16451 5329 16462 5363
rect 16496 5329 16507 5363
rect 16451 5295 16507 5329
rect 16451 5261 16462 5295
rect 16496 5261 16507 5295
rect 16451 5227 16507 5261
rect 16451 5193 16462 5227
rect 16496 5193 16507 5227
rect 16451 5181 16507 5193
rect 16537 6179 16593 6191
rect 16537 6145 16548 6179
rect 16582 6145 16593 6179
rect 16537 6111 16593 6145
rect 16537 6077 16548 6111
rect 16582 6077 16593 6111
rect 16537 6043 16593 6077
rect 16537 6009 16548 6043
rect 16582 6009 16593 6043
rect 16537 5975 16593 6009
rect 16537 5941 16548 5975
rect 16582 5941 16593 5975
rect 16537 5907 16593 5941
rect 16537 5873 16548 5907
rect 16582 5873 16593 5907
rect 16537 5839 16593 5873
rect 16537 5805 16548 5839
rect 16582 5805 16593 5839
rect 16537 5771 16593 5805
rect 16537 5737 16548 5771
rect 16582 5737 16593 5771
rect 16537 5703 16593 5737
rect 16537 5669 16548 5703
rect 16582 5669 16593 5703
rect 16537 5635 16593 5669
rect 16537 5601 16548 5635
rect 16582 5601 16593 5635
rect 16537 5567 16593 5601
rect 16537 5533 16548 5567
rect 16582 5533 16593 5567
rect 16537 5499 16593 5533
rect 16537 5465 16548 5499
rect 16582 5465 16593 5499
rect 16537 5431 16593 5465
rect 16537 5397 16548 5431
rect 16582 5397 16593 5431
rect 16537 5363 16593 5397
rect 16537 5329 16548 5363
rect 16582 5329 16593 5363
rect 16537 5295 16593 5329
rect 16537 5261 16548 5295
rect 16582 5261 16593 5295
rect 16537 5227 16593 5261
rect 16537 5193 16548 5227
rect 16582 5193 16593 5227
rect 16537 5181 16593 5193
rect 16623 6179 16679 6191
rect 16623 6145 16634 6179
rect 16668 6145 16679 6179
rect 16623 6111 16679 6145
rect 16623 6077 16634 6111
rect 16668 6077 16679 6111
rect 16623 6043 16679 6077
rect 16623 6009 16634 6043
rect 16668 6009 16679 6043
rect 16623 5975 16679 6009
rect 16623 5941 16634 5975
rect 16668 5941 16679 5975
rect 16623 5907 16679 5941
rect 16623 5873 16634 5907
rect 16668 5873 16679 5907
rect 16623 5839 16679 5873
rect 16623 5805 16634 5839
rect 16668 5805 16679 5839
rect 16623 5771 16679 5805
rect 16623 5737 16634 5771
rect 16668 5737 16679 5771
rect 16623 5703 16679 5737
rect 16623 5669 16634 5703
rect 16668 5669 16679 5703
rect 16623 5635 16679 5669
rect 16623 5601 16634 5635
rect 16668 5601 16679 5635
rect 16623 5567 16679 5601
rect 16623 5533 16634 5567
rect 16668 5533 16679 5567
rect 16623 5499 16679 5533
rect 16623 5465 16634 5499
rect 16668 5465 16679 5499
rect 16623 5431 16679 5465
rect 16623 5397 16634 5431
rect 16668 5397 16679 5431
rect 16623 5363 16679 5397
rect 16623 5329 16634 5363
rect 16668 5329 16679 5363
rect 16623 5295 16679 5329
rect 16623 5261 16634 5295
rect 16668 5261 16679 5295
rect 16623 5227 16679 5261
rect 16623 5193 16634 5227
rect 16668 5193 16679 5227
rect 16623 5181 16679 5193
rect 16709 6179 16765 6191
rect 16709 6145 16720 6179
rect 16754 6145 16765 6179
rect 16709 6111 16765 6145
rect 16709 6077 16720 6111
rect 16754 6077 16765 6111
rect 16709 6043 16765 6077
rect 16709 6009 16720 6043
rect 16754 6009 16765 6043
rect 16709 5975 16765 6009
rect 16709 5941 16720 5975
rect 16754 5941 16765 5975
rect 16709 5907 16765 5941
rect 16709 5873 16720 5907
rect 16754 5873 16765 5907
rect 16709 5839 16765 5873
rect 16709 5805 16720 5839
rect 16754 5805 16765 5839
rect 16709 5771 16765 5805
rect 16709 5737 16720 5771
rect 16754 5737 16765 5771
rect 16709 5703 16765 5737
rect 16709 5669 16720 5703
rect 16754 5669 16765 5703
rect 16709 5635 16765 5669
rect 16709 5601 16720 5635
rect 16754 5601 16765 5635
rect 16709 5567 16765 5601
rect 16709 5533 16720 5567
rect 16754 5533 16765 5567
rect 16709 5499 16765 5533
rect 16709 5465 16720 5499
rect 16754 5465 16765 5499
rect 16709 5431 16765 5465
rect 16709 5397 16720 5431
rect 16754 5397 16765 5431
rect 16709 5363 16765 5397
rect 16709 5329 16720 5363
rect 16754 5329 16765 5363
rect 16709 5295 16765 5329
rect 16709 5261 16720 5295
rect 16754 5261 16765 5295
rect 16709 5227 16765 5261
rect 16709 5193 16720 5227
rect 16754 5193 16765 5227
rect 16709 5181 16765 5193
rect 16795 6179 16851 6191
rect 16795 6145 16806 6179
rect 16840 6145 16851 6179
rect 16795 6111 16851 6145
rect 16795 6077 16806 6111
rect 16840 6077 16851 6111
rect 16795 6043 16851 6077
rect 16795 6009 16806 6043
rect 16840 6009 16851 6043
rect 16795 5975 16851 6009
rect 16795 5941 16806 5975
rect 16840 5941 16851 5975
rect 16795 5907 16851 5941
rect 16795 5873 16806 5907
rect 16840 5873 16851 5907
rect 16795 5839 16851 5873
rect 16795 5805 16806 5839
rect 16840 5805 16851 5839
rect 16795 5771 16851 5805
rect 16795 5737 16806 5771
rect 16840 5737 16851 5771
rect 16795 5703 16851 5737
rect 16795 5669 16806 5703
rect 16840 5669 16851 5703
rect 16795 5635 16851 5669
rect 16795 5601 16806 5635
rect 16840 5601 16851 5635
rect 16795 5567 16851 5601
rect 16795 5533 16806 5567
rect 16840 5533 16851 5567
rect 16795 5499 16851 5533
rect 16795 5465 16806 5499
rect 16840 5465 16851 5499
rect 16795 5431 16851 5465
rect 16795 5397 16806 5431
rect 16840 5397 16851 5431
rect 16795 5363 16851 5397
rect 16795 5329 16806 5363
rect 16840 5329 16851 5363
rect 16795 5295 16851 5329
rect 16795 5261 16806 5295
rect 16840 5261 16851 5295
rect 16795 5227 16851 5261
rect 16795 5193 16806 5227
rect 16840 5193 16851 5227
rect 16795 5181 16851 5193
rect 16881 6179 16937 6191
rect 16881 6145 16892 6179
rect 16926 6145 16937 6179
rect 16881 6111 16937 6145
rect 16881 6077 16892 6111
rect 16926 6077 16937 6111
rect 16881 6043 16937 6077
rect 16881 6009 16892 6043
rect 16926 6009 16937 6043
rect 16881 5975 16937 6009
rect 16881 5941 16892 5975
rect 16926 5941 16937 5975
rect 16881 5907 16937 5941
rect 16881 5873 16892 5907
rect 16926 5873 16937 5907
rect 16881 5839 16937 5873
rect 16881 5805 16892 5839
rect 16926 5805 16937 5839
rect 16881 5771 16937 5805
rect 16881 5737 16892 5771
rect 16926 5737 16937 5771
rect 16881 5703 16937 5737
rect 16881 5669 16892 5703
rect 16926 5669 16937 5703
rect 16881 5635 16937 5669
rect 16881 5601 16892 5635
rect 16926 5601 16937 5635
rect 16881 5567 16937 5601
rect 16881 5533 16892 5567
rect 16926 5533 16937 5567
rect 16881 5499 16937 5533
rect 16881 5465 16892 5499
rect 16926 5465 16937 5499
rect 16881 5431 16937 5465
rect 16881 5397 16892 5431
rect 16926 5397 16937 5431
rect 16881 5363 16937 5397
rect 16881 5329 16892 5363
rect 16926 5329 16937 5363
rect 16881 5295 16937 5329
rect 16881 5261 16892 5295
rect 16926 5261 16937 5295
rect 16881 5227 16937 5261
rect 16881 5193 16892 5227
rect 16926 5193 16937 5227
rect 16881 5181 16937 5193
rect 16967 6179 17023 6191
rect 16967 6145 16978 6179
rect 17012 6145 17023 6179
rect 16967 6111 17023 6145
rect 16967 6077 16978 6111
rect 17012 6077 17023 6111
rect 16967 6043 17023 6077
rect 16967 6009 16978 6043
rect 17012 6009 17023 6043
rect 16967 5975 17023 6009
rect 16967 5941 16978 5975
rect 17012 5941 17023 5975
rect 16967 5907 17023 5941
rect 16967 5873 16978 5907
rect 17012 5873 17023 5907
rect 16967 5839 17023 5873
rect 16967 5805 16978 5839
rect 17012 5805 17023 5839
rect 16967 5771 17023 5805
rect 16967 5737 16978 5771
rect 17012 5737 17023 5771
rect 16967 5703 17023 5737
rect 16967 5669 16978 5703
rect 17012 5669 17023 5703
rect 16967 5635 17023 5669
rect 16967 5601 16978 5635
rect 17012 5601 17023 5635
rect 16967 5567 17023 5601
rect 16967 5533 16978 5567
rect 17012 5533 17023 5567
rect 16967 5499 17023 5533
rect 16967 5465 16978 5499
rect 17012 5465 17023 5499
rect 16967 5431 17023 5465
rect 16967 5397 16978 5431
rect 17012 5397 17023 5431
rect 16967 5363 17023 5397
rect 16967 5329 16978 5363
rect 17012 5329 17023 5363
rect 16967 5295 17023 5329
rect 16967 5261 16978 5295
rect 17012 5261 17023 5295
rect 16967 5227 17023 5261
rect 16967 5193 16978 5227
rect 17012 5193 17023 5227
rect 16967 5181 17023 5193
rect 17053 6179 17109 6191
rect 17053 6145 17064 6179
rect 17098 6145 17109 6179
rect 17053 6111 17109 6145
rect 17053 6077 17064 6111
rect 17098 6077 17109 6111
rect 17053 6043 17109 6077
rect 17053 6009 17064 6043
rect 17098 6009 17109 6043
rect 17053 5975 17109 6009
rect 17053 5941 17064 5975
rect 17098 5941 17109 5975
rect 17053 5907 17109 5941
rect 17053 5873 17064 5907
rect 17098 5873 17109 5907
rect 17053 5839 17109 5873
rect 17053 5805 17064 5839
rect 17098 5805 17109 5839
rect 17053 5771 17109 5805
rect 17053 5737 17064 5771
rect 17098 5737 17109 5771
rect 17053 5703 17109 5737
rect 17053 5669 17064 5703
rect 17098 5669 17109 5703
rect 17053 5635 17109 5669
rect 17053 5601 17064 5635
rect 17098 5601 17109 5635
rect 17053 5567 17109 5601
rect 17053 5533 17064 5567
rect 17098 5533 17109 5567
rect 17053 5499 17109 5533
rect 17053 5465 17064 5499
rect 17098 5465 17109 5499
rect 17053 5431 17109 5465
rect 17053 5397 17064 5431
rect 17098 5397 17109 5431
rect 17053 5363 17109 5397
rect 17053 5329 17064 5363
rect 17098 5329 17109 5363
rect 17053 5295 17109 5329
rect 17053 5261 17064 5295
rect 17098 5261 17109 5295
rect 17053 5227 17109 5261
rect 17053 5193 17064 5227
rect 17098 5193 17109 5227
rect 17053 5181 17109 5193
rect 17139 6179 17195 6191
rect 17139 6145 17150 6179
rect 17184 6145 17195 6179
rect 17139 6111 17195 6145
rect 17139 6077 17150 6111
rect 17184 6077 17195 6111
rect 17139 6043 17195 6077
rect 17139 6009 17150 6043
rect 17184 6009 17195 6043
rect 17139 5975 17195 6009
rect 17139 5941 17150 5975
rect 17184 5941 17195 5975
rect 17139 5907 17195 5941
rect 17139 5873 17150 5907
rect 17184 5873 17195 5907
rect 17139 5839 17195 5873
rect 17139 5805 17150 5839
rect 17184 5805 17195 5839
rect 17139 5771 17195 5805
rect 17139 5737 17150 5771
rect 17184 5737 17195 5771
rect 17139 5703 17195 5737
rect 17139 5669 17150 5703
rect 17184 5669 17195 5703
rect 17139 5635 17195 5669
rect 17139 5601 17150 5635
rect 17184 5601 17195 5635
rect 17139 5567 17195 5601
rect 17139 5533 17150 5567
rect 17184 5533 17195 5567
rect 17139 5499 17195 5533
rect 17139 5465 17150 5499
rect 17184 5465 17195 5499
rect 17139 5431 17195 5465
rect 17139 5397 17150 5431
rect 17184 5397 17195 5431
rect 17139 5363 17195 5397
rect 17139 5329 17150 5363
rect 17184 5329 17195 5363
rect 17139 5295 17195 5329
rect 17139 5261 17150 5295
rect 17184 5261 17195 5295
rect 17139 5227 17195 5261
rect 17139 5193 17150 5227
rect 17184 5193 17195 5227
rect 17139 5181 17195 5193
<< pdiff >>
rect 17614 7908 17667 7957
rect 17614 7874 17622 7908
rect 17656 7874 17667 7908
rect 17614 7836 17667 7874
rect 17614 7802 17622 7836
rect 17656 7802 17667 7836
rect 17614 7764 17667 7802
rect 17614 7730 17622 7764
rect 17656 7730 17667 7764
rect 17614 7692 17667 7730
rect 17614 7658 17622 7692
rect 17656 7658 17667 7692
rect 17614 7620 17667 7658
rect 17614 7586 17622 7620
rect 17656 7586 17667 7620
rect 17614 7548 17667 7586
rect 17614 7514 17622 7548
rect 17656 7514 17667 7548
rect 17614 7476 17667 7514
rect 17614 7442 17622 7476
rect 17656 7442 17667 7476
rect 17614 7404 17667 7442
rect 17614 7370 17622 7404
rect 17656 7370 17667 7404
rect 17614 7332 17667 7370
rect 17614 7298 17622 7332
rect 17656 7298 17667 7332
rect 17614 7260 17667 7298
rect 17614 7226 17622 7260
rect 17656 7226 17667 7260
rect 17614 7188 17667 7226
rect 17614 7154 17622 7188
rect 17656 7154 17667 7188
rect 17614 7116 17667 7154
rect 17614 7082 17622 7116
rect 17656 7082 17667 7116
rect 17614 7044 17667 7082
rect 17614 7010 17622 7044
rect 17656 7010 17667 7044
rect 17614 6957 17667 7010
rect 17697 7908 17753 7957
rect 17697 7874 17708 7908
rect 17742 7874 17753 7908
rect 17697 7836 17753 7874
rect 17697 7802 17708 7836
rect 17742 7802 17753 7836
rect 17697 7764 17753 7802
rect 17697 7730 17708 7764
rect 17742 7730 17753 7764
rect 17697 7692 17753 7730
rect 17697 7658 17708 7692
rect 17742 7658 17753 7692
rect 17697 7620 17753 7658
rect 17697 7586 17708 7620
rect 17742 7586 17753 7620
rect 17697 7548 17753 7586
rect 17697 7514 17708 7548
rect 17742 7514 17753 7548
rect 17697 7476 17753 7514
rect 17697 7442 17708 7476
rect 17742 7442 17753 7476
rect 17697 7404 17753 7442
rect 17697 7370 17708 7404
rect 17742 7370 17753 7404
rect 17697 7332 17753 7370
rect 17697 7298 17708 7332
rect 17742 7298 17753 7332
rect 17697 7260 17753 7298
rect 17697 7226 17708 7260
rect 17742 7226 17753 7260
rect 17697 7188 17753 7226
rect 17697 7154 17708 7188
rect 17742 7154 17753 7188
rect 17697 7116 17753 7154
rect 17697 7082 17708 7116
rect 17742 7082 17753 7116
rect 17697 7044 17753 7082
rect 17697 7010 17708 7044
rect 17742 7010 17753 7044
rect 17697 6957 17753 7010
rect 17783 7908 17839 7957
rect 17783 7874 17794 7908
rect 17828 7874 17839 7908
rect 17783 7836 17839 7874
rect 17783 7802 17794 7836
rect 17828 7802 17839 7836
rect 17783 7764 17839 7802
rect 17783 7730 17794 7764
rect 17828 7730 17839 7764
rect 17783 7692 17839 7730
rect 17783 7658 17794 7692
rect 17828 7658 17839 7692
rect 17783 7620 17839 7658
rect 17783 7586 17794 7620
rect 17828 7586 17839 7620
rect 17783 7548 17839 7586
rect 17783 7514 17794 7548
rect 17828 7514 17839 7548
rect 17783 7476 17839 7514
rect 17783 7442 17794 7476
rect 17828 7442 17839 7476
rect 17783 7404 17839 7442
rect 17783 7370 17794 7404
rect 17828 7370 17839 7404
rect 17783 7332 17839 7370
rect 17783 7298 17794 7332
rect 17828 7298 17839 7332
rect 17783 7260 17839 7298
rect 17783 7226 17794 7260
rect 17828 7226 17839 7260
rect 17783 7188 17839 7226
rect 17783 7154 17794 7188
rect 17828 7154 17839 7188
rect 17783 7116 17839 7154
rect 17783 7082 17794 7116
rect 17828 7082 17839 7116
rect 17783 7044 17839 7082
rect 17783 7010 17794 7044
rect 17828 7010 17839 7044
rect 17783 6957 17839 7010
rect 17869 7908 17925 7957
rect 17869 7874 17880 7908
rect 17914 7874 17925 7908
rect 17869 7836 17925 7874
rect 17869 7802 17880 7836
rect 17914 7802 17925 7836
rect 17869 7764 17925 7802
rect 17869 7730 17880 7764
rect 17914 7730 17925 7764
rect 17869 7692 17925 7730
rect 17869 7658 17880 7692
rect 17914 7658 17925 7692
rect 17869 7620 17925 7658
rect 17869 7586 17880 7620
rect 17914 7586 17925 7620
rect 17869 7548 17925 7586
rect 17869 7514 17880 7548
rect 17914 7514 17925 7548
rect 17869 7476 17925 7514
rect 17869 7442 17880 7476
rect 17914 7442 17925 7476
rect 17869 7404 17925 7442
rect 17869 7370 17880 7404
rect 17914 7370 17925 7404
rect 17869 7332 17925 7370
rect 17869 7298 17880 7332
rect 17914 7298 17925 7332
rect 17869 7260 17925 7298
rect 17869 7226 17880 7260
rect 17914 7226 17925 7260
rect 17869 7188 17925 7226
rect 17869 7154 17880 7188
rect 17914 7154 17925 7188
rect 17869 7116 17925 7154
rect 17869 7082 17880 7116
rect 17914 7082 17925 7116
rect 17869 7044 17925 7082
rect 17869 7010 17880 7044
rect 17914 7010 17925 7044
rect 17869 6957 17925 7010
rect 17955 7908 18011 7957
rect 17955 7874 17966 7908
rect 18000 7874 18011 7908
rect 17955 7836 18011 7874
rect 17955 7802 17966 7836
rect 18000 7802 18011 7836
rect 17955 7764 18011 7802
rect 17955 7730 17966 7764
rect 18000 7730 18011 7764
rect 17955 7692 18011 7730
rect 17955 7658 17966 7692
rect 18000 7658 18011 7692
rect 17955 7620 18011 7658
rect 17955 7586 17966 7620
rect 18000 7586 18011 7620
rect 17955 7548 18011 7586
rect 17955 7514 17966 7548
rect 18000 7514 18011 7548
rect 17955 7476 18011 7514
rect 17955 7442 17966 7476
rect 18000 7442 18011 7476
rect 17955 7404 18011 7442
rect 17955 7370 17966 7404
rect 18000 7370 18011 7404
rect 17955 7332 18011 7370
rect 17955 7298 17966 7332
rect 18000 7298 18011 7332
rect 17955 7260 18011 7298
rect 17955 7226 17966 7260
rect 18000 7226 18011 7260
rect 17955 7188 18011 7226
rect 17955 7154 17966 7188
rect 18000 7154 18011 7188
rect 17955 7116 18011 7154
rect 17955 7082 17966 7116
rect 18000 7082 18011 7116
rect 17955 7044 18011 7082
rect 17955 7010 17966 7044
rect 18000 7010 18011 7044
rect 17955 6957 18011 7010
rect 18041 7908 18097 7957
rect 18041 7874 18052 7908
rect 18086 7874 18097 7908
rect 18041 7836 18097 7874
rect 18041 7802 18052 7836
rect 18086 7802 18097 7836
rect 18041 7764 18097 7802
rect 18041 7730 18052 7764
rect 18086 7730 18097 7764
rect 18041 7692 18097 7730
rect 18041 7658 18052 7692
rect 18086 7658 18097 7692
rect 18041 7620 18097 7658
rect 18041 7586 18052 7620
rect 18086 7586 18097 7620
rect 18041 7548 18097 7586
rect 18041 7514 18052 7548
rect 18086 7514 18097 7548
rect 18041 7476 18097 7514
rect 18041 7442 18052 7476
rect 18086 7442 18097 7476
rect 18041 7404 18097 7442
rect 18041 7370 18052 7404
rect 18086 7370 18097 7404
rect 18041 7332 18097 7370
rect 18041 7298 18052 7332
rect 18086 7298 18097 7332
rect 18041 7260 18097 7298
rect 18041 7226 18052 7260
rect 18086 7226 18097 7260
rect 18041 7188 18097 7226
rect 18041 7154 18052 7188
rect 18086 7154 18097 7188
rect 18041 7116 18097 7154
rect 18041 7082 18052 7116
rect 18086 7082 18097 7116
rect 18041 7044 18097 7082
rect 18041 7010 18052 7044
rect 18086 7010 18097 7044
rect 18041 6957 18097 7010
rect 18127 7908 18183 7957
rect 18127 7874 18138 7908
rect 18172 7874 18183 7908
rect 18127 7836 18183 7874
rect 18127 7802 18138 7836
rect 18172 7802 18183 7836
rect 18127 7764 18183 7802
rect 18127 7730 18138 7764
rect 18172 7730 18183 7764
rect 18127 7692 18183 7730
rect 18127 7658 18138 7692
rect 18172 7658 18183 7692
rect 18127 7620 18183 7658
rect 18127 7586 18138 7620
rect 18172 7586 18183 7620
rect 18127 7548 18183 7586
rect 18127 7514 18138 7548
rect 18172 7514 18183 7548
rect 18127 7476 18183 7514
rect 18127 7442 18138 7476
rect 18172 7442 18183 7476
rect 18127 7404 18183 7442
rect 18127 7370 18138 7404
rect 18172 7370 18183 7404
rect 18127 7332 18183 7370
rect 18127 7298 18138 7332
rect 18172 7298 18183 7332
rect 18127 7260 18183 7298
rect 18127 7226 18138 7260
rect 18172 7226 18183 7260
rect 18127 7188 18183 7226
rect 18127 7154 18138 7188
rect 18172 7154 18183 7188
rect 18127 7116 18183 7154
rect 18127 7082 18138 7116
rect 18172 7082 18183 7116
rect 18127 7044 18183 7082
rect 18127 7010 18138 7044
rect 18172 7010 18183 7044
rect 18127 6957 18183 7010
rect 18213 7908 18269 7957
rect 18213 7874 18224 7908
rect 18258 7874 18269 7908
rect 18213 7836 18269 7874
rect 18213 7802 18224 7836
rect 18258 7802 18269 7836
rect 18213 7764 18269 7802
rect 18213 7730 18224 7764
rect 18258 7730 18269 7764
rect 18213 7692 18269 7730
rect 18213 7658 18224 7692
rect 18258 7658 18269 7692
rect 18213 7620 18269 7658
rect 18213 7586 18224 7620
rect 18258 7586 18269 7620
rect 18213 7548 18269 7586
rect 18213 7514 18224 7548
rect 18258 7514 18269 7548
rect 18213 7476 18269 7514
rect 18213 7442 18224 7476
rect 18258 7442 18269 7476
rect 18213 7404 18269 7442
rect 18213 7370 18224 7404
rect 18258 7370 18269 7404
rect 18213 7332 18269 7370
rect 18213 7298 18224 7332
rect 18258 7298 18269 7332
rect 18213 7260 18269 7298
rect 18213 7226 18224 7260
rect 18258 7226 18269 7260
rect 18213 7188 18269 7226
rect 18213 7154 18224 7188
rect 18258 7154 18269 7188
rect 18213 7116 18269 7154
rect 18213 7082 18224 7116
rect 18258 7082 18269 7116
rect 18213 7044 18269 7082
rect 18213 7010 18224 7044
rect 18258 7010 18269 7044
rect 18213 6957 18269 7010
rect 18299 7908 18355 7957
rect 18299 7874 18310 7908
rect 18344 7874 18355 7908
rect 18299 7836 18355 7874
rect 18299 7802 18310 7836
rect 18344 7802 18355 7836
rect 18299 7764 18355 7802
rect 18299 7730 18310 7764
rect 18344 7730 18355 7764
rect 18299 7692 18355 7730
rect 18299 7658 18310 7692
rect 18344 7658 18355 7692
rect 18299 7620 18355 7658
rect 18299 7586 18310 7620
rect 18344 7586 18355 7620
rect 18299 7548 18355 7586
rect 18299 7514 18310 7548
rect 18344 7514 18355 7548
rect 18299 7476 18355 7514
rect 18299 7442 18310 7476
rect 18344 7442 18355 7476
rect 18299 7404 18355 7442
rect 18299 7370 18310 7404
rect 18344 7370 18355 7404
rect 18299 7332 18355 7370
rect 18299 7298 18310 7332
rect 18344 7298 18355 7332
rect 18299 7260 18355 7298
rect 18299 7226 18310 7260
rect 18344 7226 18355 7260
rect 18299 7188 18355 7226
rect 18299 7154 18310 7188
rect 18344 7154 18355 7188
rect 18299 7116 18355 7154
rect 18299 7082 18310 7116
rect 18344 7082 18355 7116
rect 18299 7044 18355 7082
rect 18299 7010 18310 7044
rect 18344 7010 18355 7044
rect 18299 6957 18355 7010
rect 18385 7908 18441 7957
rect 18385 7874 18396 7908
rect 18430 7874 18441 7908
rect 18385 7836 18441 7874
rect 18385 7802 18396 7836
rect 18430 7802 18441 7836
rect 18385 7764 18441 7802
rect 18385 7730 18396 7764
rect 18430 7730 18441 7764
rect 18385 7692 18441 7730
rect 18385 7658 18396 7692
rect 18430 7658 18441 7692
rect 18385 7620 18441 7658
rect 18385 7586 18396 7620
rect 18430 7586 18441 7620
rect 18385 7548 18441 7586
rect 18385 7514 18396 7548
rect 18430 7514 18441 7548
rect 18385 7476 18441 7514
rect 18385 7442 18396 7476
rect 18430 7442 18441 7476
rect 18385 7404 18441 7442
rect 18385 7370 18396 7404
rect 18430 7370 18441 7404
rect 18385 7332 18441 7370
rect 18385 7298 18396 7332
rect 18430 7298 18441 7332
rect 18385 7260 18441 7298
rect 18385 7226 18396 7260
rect 18430 7226 18441 7260
rect 18385 7188 18441 7226
rect 18385 7154 18396 7188
rect 18430 7154 18441 7188
rect 18385 7116 18441 7154
rect 18385 7082 18396 7116
rect 18430 7082 18441 7116
rect 18385 7044 18441 7082
rect 18385 7010 18396 7044
rect 18430 7010 18441 7044
rect 18385 6957 18441 7010
rect 18471 7908 18527 7957
rect 18471 7874 18482 7908
rect 18516 7874 18527 7908
rect 18471 7836 18527 7874
rect 18471 7802 18482 7836
rect 18516 7802 18527 7836
rect 18471 7764 18527 7802
rect 18471 7730 18482 7764
rect 18516 7730 18527 7764
rect 18471 7692 18527 7730
rect 18471 7658 18482 7692
rect 18516 7658 18527 7692
rect 18471 7620 18527 7658
rect 18471 7586 18482 7620
rect 18516 7586 18527 7620
rect 18471 7548 18527 7586
rect 18471 7514 18482 7548
rect 18516 7514 18527 7548
rect 18471 7476 18527 7514
rect 18471 7442 18482 7476
rect 18516 7442 18527 7476
rect 18471 7404 18527 7442
rect 18471 7370 18482 7404
rect 18516 7370 18527 7404
rect 18471 7332 18527 7370
rect 18471 7298 18482 7332
rect 18516 7298 18527 7332
rect 18471 7260 18527 7298
rect 18471 7226 18482 7260
rect 18516 7226 18527 7260
rect 18471 7188 18527 7226
rect 18471 7154 18482 7188
rect 18516 7154 18527 7188
rect 18471 7116 18527 7154
rect 18471 7082 18482 7116
rect 18516 7082 18527 7116
rect 18471 7044 18527 7082
rect 18471 7010 18482 7044
rect 18516 7010 18527 7044
rect 18471 6957 18527 7010
rect 18557 7908 18613 7957
rect 18557 7874 18568 7908
rect 18602 7874 18613 7908
rect 18557 7836 18613 7874
rect 18557 7802 18568 7836
rect 18602 7802 18613 7836
rect 18557 7764 18613 7802
rect 18557 7730 18568 7764
rect 18602 7730 18613 7764
rect 18557 7692 18613 7730
rect 18557 7658 18568 7692
rect 18602 7658 18613 7692
rect 18557 7620 18613 7658
rect 18557 7586 18568 7620
rect 18602 7586 18613 7620
rect 18557 7548 18613 7586
rect 18557 7514 18568 7548
rect 18602 7514 18613 7548
rect 18557 7476 18613 7514
rect 18557 7442 18568 7476
rect 18602 7442 18613 7476
rect 18557 7404 18613 7442
rect 18557 7370 18568 7404
rect 18602 7370 18613 7404
rect 18557 7332 18613 7370
rect 18557 7298 18568 7332
rect 18602 7298 18613 7332
rect 18557 7260 18613 7298
rect 18557 7226 18568 7260
rect 18602 7226 18613 7260
rect 18557 7188 18613 7226
rect 18557 7154 18568 7188
rect 18602 7154 18613 7188
rect 18557 7116 18613 7154
rect 18557 7082 18568 7116
rect 18602 7082 18613 7116
rect 18557 7044 18613 7082
rect 18557 7010 18568 7044
rect 18602 7010 18613 7044
rect 18557 6957 18613 7010
rect 18643 7908 18699 7957
rect 18643 7874 18654 7908
rect 18688 7874 18699 7908
rect 18643 7836 18699 7874
rect 18643 7802 18654 7836
rect 18688 7802 18699 7836
rect 18643 7764 18699 7802
rect 18643 7730 18654 7764
rect 18688 7730 18699 7764
rect 18643 7692 18699 7730
rect 18643 7658 18654 7692
rect 18688 7658 18699 7692
rect 18643 7620 18699 7658
rect 18643 7586 18654 7620
rect 18688 7586 18699 7620
rect 18643 7548 18699 7586
rect 18643 7514 18654 7548
rect 18688 7514 18699 7548
rect 18643 7476 18699 7514
rect 18643 7442 18654 7476
rect 18688 7442 18699 7476
rect 18643 7404 18699 7442
rect 18643 7370 18654 7404
rect 18688 7370 18699 7404
rect 18643 7332 18699 7370
rect 18643 7298 18654 7332
rect 18688 7298 18699 7332
rect 18643 7260 18699 7298
rect 18643 7226 18654 7260
rect 18688 7226 18699 7260
rect 18643 7188 18699 7226
rect 18643 7154 18654 7188
rect 18688 7154 18699 7188
rect 18643 7116 18699 7154
rect 18643 7082 18654 7116
rect 18688 7082 18699 7116
rect 18643 7044 18699 7082
rect 18643 7010 18654 7044
rect 18688 7010 18699 7044
rect 18643 6957 18699 7010
rect 18729 7908 18785 7957
rect 18729 7874 18740 7908
rect 18774 7874 18785 7908
rect 18729 7836 18785 7874
rect 18729 7802 18740 7836
rect 18774 7802 18785 7836
rect 18729 7764 18785 7802
rect 18729 7730 18740 7764
rect 18774 7730 18785 7764
rect 18729 7692 18785 7730
rect 18729 7658 18740 7692
rect 18774 7658 18785 7692
rect 18729 7620 18785 7658
rect 18729 7586 18740 7620
rect 18774 7586 18785 7620
rect 18729 7548 18785 7586
rect 18729 7514 18740 7548
rect 18774 7514 18785 7548
rect 18729 7476 18785 7514
rect 18729 7442 18740 7476
rect 18774 7442 18785 7476
rect 18729 7404 18785 7442
rect 18729 7370 18740 7404
rect 18774 7370 18785 7404
rect 18729 7332 18785 7370
rect 18729 7298 18740 7332
rect 18774 7298 18785 7332
rect 18729 7260 18785 7298
rect 18729 7226 18740 7260
rect 18774 7226 18785 7260
rect 18729 7188 18785 7226
rect 18729 7154 18740 7188
rect 18774 7154 18785 7188
rect 18729 7116 18785 7154
rect 18729 7082 18740 7116
rect 18774 7082 18785 7116
rect 18729 7044 18785 7082
rect 18729 7010 18740 7044
rect 18774 7010 18785 7044
rect 18729 6957 18785 7010
rect 18815 7908 18871 7957
rect 18815 7874 18826 7908
rect 18860 7874 18871 7908
rect 18815 7836 18871 7874
rect 18815 7802 18826 7836
rect 18860 7802 18871 7836
rect 18815 7764 18871 7802
rect 18815 7730 18826 7764
rect 18860 7730 18871 7764
rect 18815 7692 18871 7730
rect 18815 7658 18826 7692
rect 18860 7658 18871 7692
rect 18815 7620 18871 7658
rect 18815 7586 18826 7620
rect 18860 7586 18871 7620
rect 18815 7548 18871 7586
rect 18815 7514 18826 7548
rect 18860 7514 18871 7548
rect 18815 7476 18871 7514
rect 18815 7442 18826 7476
rect 18860 7442 18871 7476
rect 18815 7404 18871 7442
rect 18815 7370 18826 7404
rect 18860 7370 18871 7404
rect 18815 7332 18871 7370
rect 18815 7298 18826 7332
rect 18860 7298 18871 7332
rect 18815 7260 18871 7298
rect 18815 7226 18826 7260
rect 18860 7226 18871 7260
rect 18815 7188 18871 7226
rect 18815 7154 18826 7188
rect 18860 7154 18871 7188
rect 18815 7116 18871 7154
rect 18815 7082 18826 7116
rect 18860 7082 18871 7116
rect 18815 7044 18871 7082
rect 18815 7010 18826 7044
rect 18860 7010 18871 7044
rect 18815 6957 18871 7010
rect 18901 7908 18957 7957
rect 18901 7874 18912 7908
rect 18946 7874 18957 7908
rect 18901 7836 18957 7874
rect 18901 7802 18912 7836
rect 18946 7802 18957 7836
rect 18901 7764 18957 7802
rect 18901 7730 18912 7764
rect 18946 7730 18957 7764
rect 18901 7692 18957 7730
rect 18901 7658 18912 7692
rect 18946 7658 18957 7692
rect 18901 7620 18957 7658
rect 18901 7586 18912 7620
rect 18946 7586 18957 7620
rect 18901 7548 18957 7586
rect 18901 7514 18912 7548
rect 18946 7514 18957 7548
rect 18901 7476 18957 7514
rect 18901 7442 18912 7476
rect 18946 7442 18957 7476
rect 18901 7404 18957 7442
rect 18901 7370 18912 7404
rect 18946 7370 18957 7404
rect 18901 7332 18957 7370
rect 18901 7298 18912 7332
rect 18946 7298 18957 7332
rect 18901 7260 18957 7298
rect 18901 7226 18912 7260
rect 18946 7226 18957 7260
rect 18901 7188 18957 7226
rect 18901 7154 18912 7188
rect 18946 7154 18957 7188
rect 18901 7116 18957 7154
rect 18901 7082 18912 7116
rect 18946 7082 18957 7116
rect 18901 7044 18957 7082
rect 18901 7010 18912 7044
rect 18946 7010 18957 7044
rect 18901 6957 18957 7010
rect 18987 7908 19043 7957
rect 18987 7874 18998 7908
rect 19032 7874 19043 7908
rect 18987 7836 19043 7874
rect 18987 7802 18998 7836
rect 19032 7802 19043 7836
rect 18987 7764 19043 7802
rect 18987 7730 18998 7764
rect 19032 7730 19043 7764
rect 18987 7692 19043 7730
rect 18987 7658 18998 7692
rect 19032 7658 19043 7692
rect 18987 7620 19043 7658
rect 18987 7586 18998 7620
rect 19032 7586 19043 7620
rect 18987 7548 19043 7586
rect 18987 7514 18998 7548
rect 19032 7514 19043 7548
rect 18987 7476 19043 7514
rect 18987 7442 18998 7476
rect 19032 7442 19043 7476
rect 18987 7404 19043 7442
rect 18987 7370 18998 7404
rect 19032 7370 19043 7404
rect 18987 7332 19043 7370
rect 18987 7298 18998 7332
rect 19032 7298 19043 7332
rect 18987 7260 19043 7298
rect 18987 7226 18998 7260
rect 19032 7226 19043 7260
rect 18987 7188 19043 7226
rect 18987 7154 18998 7188
rect 19032 7154 19043 7188
rect 18987 7116 19043 7154
rect 18987 7082 18998 7116
rect 19032 7082 19043 7116
rect 18987 7044 19043 7082
rect 18987 7010 18998 7044
rect 19032 7010 19043 7044
rect 18987 6957 19043 7010
rect 19073 7908 19129 7957
rect 19073 7874 19084 7908
rect 19118 7874 19129 7908
rect 19073 7836 19129 7874
rect 19073 7802 19084 7836
rect 19118 7802 19129 7836
rect 19073 7764 19129 7802
rect 19073 7730 19084 7764
rect 19118 7730 19129 7764
rect 19073 7692 19129 7730
rect 19073 7658 19084 7692
rect 19118 7658 19129 7692
rect 19073 7620 19129 7658
rect 19073 7586 19084 7620
rect 19118 7586 19129 7620
rect 19073 7548 19129 7586
rect 19073 7514 19084 7548
rect 19118 7514 19129 7548
rect 19073 7476 19129 7514
rect 19073 7442 19084 7476
rect 19118 7442 19129 7476
rect 19073 7404 19129 7442
rect 19073 7370 19084 7404
rect 19118 7370 19129 7404
rect 19073 7332 19129 7370
rect 19073 7298 19084 7332
rect 19118 7298 19129 7332
rect 19073 7260 19129 7298
rect 19073 7226 19084 7260
rect 19118 7226 19129 7260
rect 19073 7188 19129 7226
rect 19073 7154 19084 7188
rect 19118 7154 19129 7188
rect 19073 7116 19129 7154
rect 19073 7082 19084 7116
rect 19118 7082 19129 7116
rect 19073 7044 19129 7082
rect 19073 7010 19084 7044
rect 19118 7010 19129 7044
rect 19073 6957 19129 7010
rect 19159 7908 19215 7957
rect 19159 7874 19170 7908
rect 19204 7874 19215 7908
rect 19159 7836 19215 7874
rect 19159 7802 19170 7836
rect 19204 7802 19215 7836
rect 19159 7764 19215 7802
rect 19159 7730 19170 7764
rect 19204 7730 19215 7764
rect 19159 7692 19215 7730
rect 19159 7658 19170 7692
rect 19204 7658 19215 7692
rect 19159 7620 19215 7658
rect 19159 7586 19170 7620
rect 19204 7586 19215 7620
rect 19159 7548 19215 7586
rect 19159 7514 19170 7548
rect 19204 7514 19215 7548
rect 19159 7476 19215 7514
rect 19159 7442 19170 7476
rect 19204 7442 19215 7476
rect 19159 7404 19215 7442
rect 19159 7370 19170 7404
rect 19204 7370 19215 7404
rect 19159 7332 19215 7370
rect 19159 7298 19170 7332
rect 19204 7298 19215 7332
rect 19159 7260 19215 7298
rect 19159 7226 19170 7260
rect 19204 7226 19215 7260
rect 19159 7188 19215 7226
rect 19159 7154 19170 7188
rect 19204 7154 19215 7188
rect 19159 7116 19215 7154
rect 19159 7082 19170 7116
rect 19204 7082 19215 7116
rect 19159 7044 19215 7082
rect 19159 7010 19170 7044
rect 19204 7010 19215 7044
rect 19159 6957 19215 7010
rect 19245 7908 19301 7957
rect 19245 7874 19256 7908
rect 19290 7874 19301 7908
rect 19245 7836 19301 7874
rect 19245 7802 19256 7836
rect 19290 7802 19301 7836
rect 19245 7764 19301 7802
rect 19245 7730 19256 7764
rect 19290 7730 19301 7764
rect 19245 7692 19301 7730
rect 19245 7658 19256 7692
rect 19290 7658 19301 7692
rect 19245 7620 19301 7658
rect 19245 7586 19256 7620
rect 19290 7586 19301 7620
rect 19245 7548 19301 7586
rect 19245 7514 19256 7548
rect 19290 7514 19301 7548
rect 19245 7476 19301 7514
rect 19245 7442 19256 7476
rect 19290 7442 19301 7476
rect 19245 7404 19301 7442
rect 19245 7370 19256 7404
rect 19290 7370 19301 7404
rect 19245 7332 19301 7370
rect 19245 7298 19256 7332
rect 19290 7298 19301 7332
rect 19245 7260 19301 7298
rect 19245 7226 19256 7260
rect 19290 7226 19301 7260
rect 19245 7188 19301 7226
rect 19245 7154 19256 7188
rect 19290 7154 19301 7188
rect 19245 7116 19301 7154
rect 19245 7082 19256 7116
rect 19290 7082 19301 7116
rect 19245 7044 19301 7082
rect 19245 7010 19256 7044
rect 19290 7010 19301 7044
rect 19245 6957 19301 7010
rect 19331 7908 19387 7957
rect 19331 7874 19342 7908
rect 19376 7874 19387 7908
rect 19331 7836 19387 7874
rect 19331 7802 19342 7836
rect 19376 7802 19387 7836
rect 19331 7764 19387 7802
rect 19331 7730 19342 7764
rect 19376 7730 19387 7764
rect 19331 7692 19387 7730
rect 19331 7658 19342 7692
rect 19376 7658 19387 7692
rect 19331 7620 19387 7658
rect 19331 7586 19342 7620
rect 19376 7586 19387 7620
rect 19331 7548 19387 7586
rect 19331 7514 19342 7548
rect 19376 7514 19387 7548
rect 19331 7476 19387 7514
rect 19331 7442 19342 7476
rect 19376 7442 19387 7476
rect 19331 7404 19387 7442
rect 19331 7370 19342 7404
rect 19376 7370 19387 7404
rect 19331 7332 19387 7370
rect 19331 7298 19342 7332
rect 19376 7298 19387 7332
rect 19331 7260 19387 7298
rect 19331 7226 19342 7260
rect 19376 7226 19387 7260
rect 19331 7188 19387 7226
rect 19331 7154 19342 7188
rect 19376 7154 19387 7188
rect 19331 7116 19387 7154
rect 19331 7082 19342 7116
rect 19376 7082 19387 7116
rect 19331 7044 19387 7082
rect 19331 7010 19342 7044
rect 19376 7010 19387 7044
rect 19331 6957 19387 7010
rect 19417 7908 19473 7957
rect 19417 7874 19428 7908
rect 19462 7874 19473 7908
rect 19417 7836 19473 7874
rect 19417 7802 19428 7836
rect 19462 7802 19473 7836
rect 19417 7764 19473 7802
rect 19417 7730 19428 7764
rect 19462 7730 19473 7764
rect 19417 7692 19473 7730
rect 19417 7658 19428 7692
rect 19462 7658 19473 7692
rect 19417 7620 19473 7658
rect 19417 7586 19428 7620
rect 19462 7586 19473 7620
rect 19417 7548 19473 7586
rect 19417 7514 19428 7548
rect 19462 7514 19473 7548
rect 19417 7476 19473 7514
rect 19417 7442 19428 7476
rect 19462 7442 19473 7476
rect 19417 7404 19473 7442
rect 19417 7370 19428 7404
rect 19462 7370 19473 7404
rect 19417 7332 19473 7370
rect 19417 7298 19428 7332
rect 19462 7298 19473 7332
rect 19417 7260 19473 7298
rect 19417 7226 19428 7260
rect 19462 7226 19473 7260
rect 19417 7188 19473 7226
rect 19417 7154 19428 7188
rect 19462 7154 19473 7188
rect 19417 7116 19473 7154
rect 19417 7082 19428 7116
rect 19462 7082 19473 7116
rect 19417 7044 19473 7082
rect 19417 7010 19428 7044
rect 19462 7010 19473 7044
rect 19417 6957 19473 7010
rect 19503 7908 19559 7957
rect 19503 7874 19514 7908
rect 19548 7874 19559 7908
rect 19503 7836 19559 7874
rect 19503 7802 19514 7836
rect 19548 7802 19559 7836
rect 19503 7764 19559 7802
rect 19503 7730 19514 7764
rect 19548 7730 19559 7764
rect 19503 7692 19559 7730
rect 19503 7658 19514 7692
rect 19548 7658 19559 7692
rect 19503 7620 19559 7658
rect 19503 7586 19514 7620
rect 19548 7586 19559 7620
rect 19503 7548 19559 7586
rect 19503 7514 19514 7548
rect 19548 7514 19559 7548
rect 19503 7476 19559 7514
rect 19503 7442 19514 7476
rect 19548 7442 19559 7476
rect 19503 7404 19559 7442
rect 19503 7370 19514 7404
rect 19548 7370 19559 7404
rect 19503 7332 19559 7370
rect 19503 7298 19514 7332
rect 19548 7298 19559 7332
rect 19503 7260 19559 7298
rect 19503 7226 19514 7260
rect 19548 7226 19559 7260
rect 19503 7188 19559 7226
rect 19503 7154 19514 7188
rect 19548 7154 19559 7188
rect 19503 7116 19559 7154
rect 19503 7082 19514 7116
rect 19548 7082 19559 7116
rect 19503 7044 19559 7082
rect 19503 7010 19514 7044
rect 19548 7010 19559 7044
rect 19503 6957 19559 7010
rect 19589 7908 19645 7957
rect 19589 7874 19600 7908
rect 19634 7874 19645 7908
rect 19589 7836 19645 7874
rect 19589 7802 19600 7836
rect 19634 7802 19645 7836
rect 19589 7764 19645 7802
rect 19589 7730 19600 7764
rect 19634 7730 19645 7764
rect 19589 7692 19645 7730
rect 19589 7658 19600 7692
rect 19634 7658 19645 7692
rect 19589 7620 19645 7658
rect 19589 7586 19600 7620
rect 19634 7586 19645 7620
rect 19589 7548 19645 7586
rect 19589 7514 19600 7548
rect 19634 7514 19645 7548
rect 19589 7476 19645 7514
rect 19589 7442 19600 7476
rect 19634 7442 19645 7476
rect 19589 7404 19645 7442
rect 19589 7370 19600 7404
rect 19634 7370 19645 7404
rect 19589 7332 19645 7370
rect 19589 7298 19600 7332
rect 19634 7298 19645 7332
rect 19589 7260 19645 7298
rect 19589 7226 19600 7260
rect 19634 7226 19645 7260
rect 19589 7188 19645 7226
rect 19589 7154 19600 7188
rect 19634 7154 19645 7188
rect 19589 7116 19645 7154
rect 19589 7082 19600 7116
rect 19634 7082 19645 7116
rect 19589 7044 19645 7082
rect 19589 7010 19600 7044
rect 19634 7010 19645 7044
rect 19589 6957 19645 7010
rect 19675 7908 19731 7957
rect 19675 7874 19686 7908
rect 19720 7874 19731 7908
rect 19675 7836 19731 7874
rect 19675 7802 19686 7836
rect 19720 7802 19731 7836
rect 19675 7764 19731 7802
rect 19675 7730 19686 7764
rect 19720 7730 19731 7764
rect 19675 7692 19731 7730
rect 19675 7658 19686 7692
rect 19720 7658 19731 7692
rect 19675 7620 19731 7658
rect 19675 7586 19686 7620
rect 19720 7586 19731 7620
rect 19675 7548 19731 7586
rect 19675 7514 19686 7548
rect 19720 7514 19731 7548
rect 19675 7476 19731 7514
rect 19675 7442 19686 7476
rect 19720 7442 19731 7476
rect 19675 7404 19731 7442
rect 19675 7370 19686 7404
rect 19720 7370 19731 7404
rect 19675 7332 19731 7370
rect 19675 7298 19686 7332
rect 19720 7298 19731 7332
rect 19675 7260 19731 7298
rect 19675 7226 19686 7260
rect 19720 7226 19731 7260
rect 19675 7188 19731 7226
rect 19675 7154 19686 7188
rect 19720 7154 19731 7188
rect 19675 7116 19731 7154
rect 19675 7082 19686 7116
rect 19720 7082 19731 7116
rect 19675 7044 19731 7082
rect 19675 7010 19686 7044
rect 19720 7010 19731 7044
rect 19675 6957 19731 7010
rect 19761 7908 19817 7957
rect 19761 7874 19772 7908
rect 19806 7874 19817 7908
rect 19761 7836 19817 7874
rect 19761 7802 19772 7836
rect 19806 7802 19817 7836
rect 19761 7764 19817 7802
rect 19761 7730 19772 7764
rect 19806 7730 19817 7764
rect 19761 7692 19817 7730
rect 19761 7658 19772 7692
rect 19806 7658 19817 7692
rect 19761 7620 19817 7658
rect 19761 7586 19772 7620
rect 19806 7586 19817 7620
rect 19761 7548 19817 7586
rect 19761 7514 19772 7548
rect 19806 7514 19817 7548
rect 19761 7476 19817 7514
rect 19761 7442 19772 7476
rect 19806 7442 19817 7476
rect 19761 7404 19817 7442
rect 19761 7370 19772 7404
rect 19806 7370 19817 7404
rect 19761 7332 19817 7370
rect 19761 7298 19772 7332
rect 19806 7298 19817 7332
rect 19761 7260 19817 7298
rect 19761 7226 19772 7260
rect 19806 7226 19817 7260
rect 19761 7188 19817 7226
rect 19761 7154 19772 7188
rect 19806 7154 19817 7188
rect 19761 7116 19817 7154
rect 19761 7082 19772 7116
rect 19806 7082 19817 7116
rect 19761 7044 19817 7082
rect 19761 7010 19772 7044
rect 19806 7010 19817 7044
rect 19761 6957 19817 7010
rect 19847 7908 19903 7957
rect 19847 7874 19858 7908
rect 19892 7874 19903 7908
rect 19847 7836 19903 7874
rect 19847 7802 19858 7836
rect 19892 7802 19903 7836
rect 19847 7764 19903 7802
rect 19847 7730 19858 7764
rect 19892 7730 19903 7764
rect 19847 7692 19903 7730
rect 19847 7658 19858 7692
rect 19892 7658 19903 7692
rect 19847 7620 19903 7658
rect 19847 7586 19858 7620
rect 19892 7586 19903 7620
rect 19847 7548 19903 7586
rect 19847 7514 19858 7548
rect 19892 7514 19903 7548
rect 19847 7476 19903 7514
rect 19847 7442 19858 7476
rect 19892 7442 19903 7476
rect 19847 7404 19903 7442
rect 19847 7370 19858 7404
rect 19892 7370 19903 7404
rect 19847 7332 19903 7370
rect 19847 7298 19858 7332
rect 19892 7298 19903 7332
rect 19847 7260 19903 7298
rect 19847 7226 19858 7260
rect 19892 7226 19903 7260
rect 19847 7188 19903 7226
rect 19847 7154 19858 7188
rect 19892 7154 19903 7188
rect 19847 7116 19903 7154
rect 19847 7082 19858 7116
rect 19892 7082 19903 7116
rect 19847 7044 19903 7082
rect 19847 7010 19858 7044
rect 19892 7010 19903 7044
rect 19847 6957 19903 7010
rect 19933 7908 19989 7957
rect 19933 7874 19944 7908
rect 19978 7874 19989 7908
rect 19933 7836 19989 7874
rect 19933 7802 19944 7836
rect 19978 7802 19989 7836
rect 19933 7764 19989 7802
rect 19933 7730 19944 7764
rect 19978 7730 19989 7764
rect 19933 7692 19989 7730
rect 19933 7658 19944 7692
rect 19978 7658 19989 7692
rect 19933 7620 19989 7658
rect 19933 7586 19944 7620
rect 19978 7586 19989 7620
rect 19933 7548 19989 7586
rect 19933 7514 19944 7548
rect 19978 7514 19989 7548
rect 19933 7476 19989 7514
rect 19933 7442 19944 7476
rect 19978 7442 19989 7476
rect 19933 7404 19989 7442
rect 19933 7370 19944 7404
rect 19978 7370 19989 7404
rect 19933 7332 19989 7370
rect 19933 7298 19944 7332
rect 19978 7298 19989 7332
rect 19933 7260 19989 7298
rect 19933 7226 19944 7260
rect 19978 7226 19989 7260
rect 19933 7188 19989 7226
rect 19933 7154 19944 7188
rect 19978 7154 19989 7188
rect 19933 7116 19989 7154
rect 19933 7082 19944 7116
rect 19978 7082 19989 7116
rect 19933 7044 19989 7082
rect 19933 7010 19944 7044
rect 19978 7010 19989 7044
rect 19933 6957 19989 7010
rect 20019 7908 20072 7957
rect 20019 7874 20030 7908
rect 20064 7874 20072 7908
rect 20019 7836 20072 7874
rect 20019 7802 20030 7836
rect 20064 7802 20072 7836
rect 20019 7764 20072 7802
rect 20019 7730 20030 7764
rect 20064 7730 20072 7764
rect 20019 7692 20072 7730
rect 20019 7658 20030 7692
rect 20064 7658 20072 7692
rect 20019 7620 20072 7658
rect 20019 7586 20030 7620
rect 20064 7586 20072 7620
rect 20019 7548 20072 7586
rect 20019 7514 20030 7548
rect 20064 7514 20072 7548
rect 20019 7476 20072 7514
rect 20019 7442 20030 7476
rect 20064 7442 20072 7476
rect 20019 7404 20072 7442
rect 20019 7370 20030 7404
rect 20064 7370 20072 7404
rect 20019 7332 20072 7370
rect 20019 7298 20030 7332
rect 20064 7298 20072 7332
rect 20019 7260 20072 7298
rect 20019 7226 20030 7260
rect 20064 7226 20072 7260
rect 20019 7188 20072 7226
rect 20019 7154 20030 7188
rect 20064 7154 20072 7188
rect 20019 7116 20072 7154
rect 20019 7082 20030 7116
rect 20064 7082 20072 7116
rect 20019 7044 20072 7082
rect 20019 7010 20030 7044
rect 20064 7010 20072 7044
rect 20019 6957 20072 7010
rect 17596 6180 17649 6233
rect 17596 6146 17604 6180
rect 17638 6146 17649 6180
rect 17596 6108 17649 6146
rect 17596 6074 17604 6108
rect 17638 6074 17649 6108
rect 17596 6036 17649 6074
rect 17596 6002 17604 6036
rect 17638 6002 17649 6036
rect 17596 5964 17649 6002
rect 17596 5930 17604 5964
rect 17638 5930 17649 5964
rect 17596 5892 17649 5930
rect 17596 5858 17604 5892
rect 17638 5858 17649 5892
rect 17596 5820 17649 5858
rect 17596 5786 17604 5820
rect 17638 5786 17649 5820
rect 17596 5748 17649 5786
rect 17596 5714 17604 5748
rect 17638 5714 17649 5748
rect 17596 5676 17649 5714
rect 17596 5642 17604 5676
rect 17638 5642 17649 5676
rect 17596 5604 17649 5642
rect 17596 5570 17604 5604
rect 17638 5570 17649 5604
rect 17596 5532 17649 5570
rect 17596 5498 17604 5532
rect 17638 5498 17649 5532
rect 17596 5460 17649 5498
rect 17596 5426 17604 5460
rect 17638 5426 17649 5460
rect 17596 5388 17649 5426
rect 17596 5354 17604 5388
rect 17638 5354 17649 5388
rect 17596 5316 17649 5354
rect 17596 5282 17604 5316
rect 17638 5282 17649 5316
rect 17596 5233 17649 5282
rect 17679 6180 17735 6233
rect 17679 6146 17690 6180
rect 17724 6146 17735 6180
rect 17679 6108 17735 6146
rect 17679 6074 17690 6108
rect 17724 6074 17735 6108
rect 17679 6036 17735 6074
rect 17679 6002 17690 6036
rect 17724 6002 17735 6036
rect 17679 5964 17735 6002
rect 17679 5930 17690 5964
rect 17724 5930 17735 5964
rect 17679 5892 17735 5930
rect 17679 5858 17690 5892
rect 17724 5858 17735 5892
rect 17679 5820 17735 5858
rect 17679 5786 17690 5820
rect 17724 5786 17735 5820
rect 17679 5748 17735 5786
rect 17679 5714 17690 5748
rect 17724 5714 17735 5748
rect 17679 5676 17735 5714
rect 17679 5642 17690 5676
rect 17724 5642 17735 5676
rect 17679 5604 17735 5642
rect 17679 5570 17690 5604
rect 17724 5570 17735 5604
rect 17679 5532 17735 5570
rect 17679 5498 17690 5532
rect 17724 5498 17735 5532
rect 17679 5460 17735 5498
rect 17679 5426 17690 5460
rect 17724 5426 17735 5460
rect 17679 5388 17735 5426
rect 17679 5354 17690 5388
rect 17724 5354 17735 5388
rect 17679 5316 17735 5354
rect 17679 5282 17690 5316
rect 17724 5282 17735 5316
rect 17679 5233 17735 5282
rect 17765 6180 17821 6233
rect 17765 6146 17776 6180
rect 17810 6146 17821 6180
rect 17765 6108 17821 6146
rect 17765 6074 17776 6108
rect 17810 6074 17821 6108
rect 17765 6036 17821 6074
rect 17765 6002 17776 6036
rect 17810 6002 17821 6036
rect 17765 5964 17821 6002
rect 17765 5930 17776 5964
rect 17810 5930 17821 5964
rect 17765 5892 17821 5930
rect 17765 5858 17776 5892
rect 17810 5858 17821 5892
rect 17765 5820 17821 5858
rect 17765 5786 17776 5820
rect 17810 5786 17821 5820
rect 17765 5748 17821 5786
rect 17765 5714 17776 5748
rect 17810 5714 17821 5748
rect 17765 5676 17821 5714
rect 17765 5642 17776 5676
rect 17810 5642 17821 5676
rect 17765 5604 17821 5642
rect 17765 5570 17776 5604
rect 17810 5570 17821 5604
rect 17765 5532 17821 5570
rect 17765 5498 17776 5532
rect 17810 5498 17821 5532
rect 17765 5460 17821 5498
rect 17765 5426 17776 5460
rect 17810 5426 17821 5460
rect 17765 5388 17821 5426
rect 17765 5354 17776 5388
rect 17810 5354 17821 5388
rect 17765 5316 17821 5354
rect 17765 5282 17776 5316
rect 17810 5282 17821 5316
rect 17765 5233 17821 5282
rect 17851 6180 17907 6233
rect 17851 6146 17862 6180
rect 17896 6146 17907 6180
rect 17851 6108 17907 6146
rect 17851 6074 17862 6108
rect 17896 6074 17907 6108
rect 17851 6036 17907 6074
rect 17851 6002 17862 6036
rect 17896 6002 17907 6036
rect 17851 5964 17907 6002
rect 17851 5930 17862 5964
rect 17896 5930 17907 5964
rect 17851 5892 17907 5930
rect 17851 5858 17862 5892
rect 17896 5858 17907 5892
rect 17851 5820 17907 5858
rect 17851 5786 17862 5820
rect 17896 5786 17907 5820
rect 17851 5748 17907 5786
rect 17851 5714 17862 5748
rect 17896 5714 17907 5748
rect 17851 5676 17907 5714
rect 17851 5642 17862 5676
rect 17896 5642 17907 5676
rect 17851 5604 17907 5642
rect 17851 5570 17862 5604
rect 17896 5570 17907 5604
rect 17851 5532 17907 5570
rect 17851 5498 17862 5532
rect 17896 5498 17907 5532
rect 17851 5460 17907 5498
rect 17851 5426 17862 5460
rect 17896 5426 17907 5460
rect 17851 5388 17907 5426
rect 17851 5354 17862 5388
rect 17896 5354 17907 5388
rect 17851 5316 17907 5354
rect 17851 5282 17862 5316
rect 17896 5282 17907 5316
rect 17851 5233 17907 5282
rect 17937 6180 17993 6233
rect 17937 6146 17948 6180
rect 17982 6146 17993 6180
rect 17937 6108 17993 6146
rect 17937 6074 17948 6108
rect 17982 6074 17993 6108
rect 17937 6036 17993 6074
rect 17937 6002 17948 6036
rect 17982 6002 17993 6036
rect 17937 5964 17993 6002
rect 17937 5930 17948 5964
rect 17982 5930 17993 5964
rect 17937 5892 17993 5930
rect 17937 5858 17948 5892
rect 17982 5858 17993 5892
rect 17937 5820 17993 5858
rect 17937 5786 17948 5820
rect 17982 5786 17993 5820
rect 17937 5748 17993 5786
rect 17937 5714 17948 5748
rect 17982 5714 17993 5748
rect 17937 5676 17993 5714
rect 17937 5642 17948 5676
rect 17982 5642 17993 5676
rect 17937 5604 17993 5642
rect 17937 5570 17948 5604
rect 17982 5570 17993 5604
rect 17937 5532 17993 5570
rect 17937 5498 17948 5532
rect 17982 5498 17993 5532
rect 17937 5460 17993 5498
rect 17937 5426 17948 5460
rect 17982 5426 17993 5460
rect 17937 5388 17993 5426
rect 17937 5354 17948 5388
rect 17982 5354 17993 5388
rect 17937 5316 17993 5354
rect 17937 5282 17948 5316
rect 17982 5282 17993 5316
rect 17937 5233 17993 5282
rect 18023 6180 18079 6233
rect 18023 6146 18034 6180
rect 18068 6146 18079 6180
rect 18023 6108 18079 6146
rect 18023 6074 18034 6108
rect 18068 6074 18079 6108
rect 18023 6036 18079 6074
rect 18023 6002 18034 6036
rect 18068 6002 18079 6036
rect 18023 5964 18079 6002
rect 18023 5930 18034 5964
rect 18068 5930 18079 5964
rect 18023 5892 18079 5930
rect 18023 5858 18034 5892
rect 18068 5858 18079 5892
rect 18023 5820 18079 5858
rect 18023 5786 18034 5820
rect 18068 5786 18079 5820
rect 18023 5748 18079 5786
rect 18023 5714 18034 5748
rect 18068 5714 18079 5748
rect 18023 5676 18079 5714
rect 18023 5642 18034 5676
rect 18068 5642 18079 5676
rect 18023 5604 18079 5642
rect 18023 5570 18034 5604
rect 18068 5570 18079 5604
rect 18023 5532 18079 5570
rect 18023 5498 18034 5532
rect 18068 5498 18079 5532
rect 18023 5460 18079 5498
rect 18023 5426 18034 5460
rect 18068 5426 18079 5460
rect 18023 5388 18079 5426
rect 18023 5354 18034 5388
rect 18068 5354 18079 5388
rect 18023 5316 18079 5354
rect 18023 5282 18034 5316
rect 18068 5282 18079 5316
rect 18023 5233 18079 5282
rect 18109 6180 18165 6233
rect 18109 6146 18120 6180
rect 18154 6146 18165 6180
rect 18109 6108 18165 6146
rect 18109 6074 18120 6108
rect 18154 6074 18165 6108
rect 18109 6036 18165 6074
rect 18109 6002 18120 6036
rect 18154 6002 18165 6036
rect 18109 5964 18165 6002
rect 18109 5930 18120 5964
rect 18154 5930 18165 5964
rect 18109 5892 18165 5930
rect 18109 5858 18120 5892
rect 18154 5858 18165 5892
rect 18109 5820 18165 5858
rect 18109 5786 18120 5820
rect 18154 5786 18165 5820
rect 18109 5748 18165 5786
rect 18109 5714 18120 5748
rect 18154 5714 18165 5748
rect 18109 5676 18165 5714
rect 18109 5642 18120 5676
rect 18154 5642 18165 5676
rect 18109 5604 18165 5642
rect 18109 5570 18120 5604
rect 18154 5570 18165 5604
rect 18109 5532 18165 5570
rect 18109 5498 18120 5532
rect 18154 5498 18165 5532
rect 18109 5460 18165 5498
rect 18109 5426 18120 5460
rect 18154 5426 18165 5460
rect 18109 5388 18165 5426
rect 18109 5354 18120 5388
rect 18154 5354 18165 5388
rect 18109 5316 18165 5354
rect 18109 5282 18120 5316
rect 18154 5282 18165 5316
rect 18109 5233 18165 5282
rect 18195 6180 18251 6233
rect 18195 6146 18206 6180
rect 18240 6146 18251 6180
rect 18195 6108 18251 6146
rect 18195 6074 18206 6108
rect 18240 6074 18251 6108
rect 18195 6036 18251 6074
rect 18195 6002 18206 6036
rect 18240 6002 18251 6036
rect 18195 5964 18251 6002
rect 18195 5930 18206 5964
rect 18240 5930 18251 5964
rect 18195 5892 18251 5930
rect 18195 5858 18206 5892
rect 18240 5858 18251 5892
rect 18195 5820 18251 5858
rect 18195 5786 18206 5820
rect 18240 5786 18251 5820
rect 18195 5748 18251 5786
rect 18195 5714 18206 5748
rect 18240 5714 18251 5748
rect 18195 5676 18251 5714
rect 18195 5642 18206 5676
rect 18240 5642 18251 5676
rect 18195 5604 18251 5642
rect 18195 5570 18206 5604
rect 18240 5570 18251 5604
rect 18195 5532 18251 5570
rect 18195 5498 18206 5532
rect 18240 5498 18251 5532
rect 18195 5460 18251 5498
rect 18195 5426 18206 5460
rect 18240 5426 18251 5460
rect 18195 5388 18251 5426
rect 18195 5354 18206 5388
rect 18240 5354 18251 5388
rect 18195 5316 18251 5354
rect 18195 5282 18206 5316
rect 18240 5282 18251 5316
rect 18195 5233 18251 5282
rect 18281 6180 18337 6233
rect 18281 6146 18292 6180
rect 18326 6146 18337 6180
rect 18281 6108 18337 6146
rect 18281 6074 18292 6108
rect 18326 6074 18337 6108
rect 18281 6036 18337 6074
rect 18281 6002 18292 6036
rect 18326 6002 18337 6036
rect 18281 5964 18337 6002
rect 18281 5930 18292 5964
rect 18326 5930 18337 5964
rect 18281 5892 18337 5930
rect 18281 5858 18292 5892
rect 18326 5858 18337 5892
rect 18281 5820 18337 5858
rect 18281 5786 18292 5820
rect 18326 5786 18337 5820
rect 18281 5748 18337 5786
rect 18281 5714 18292 5748
rect 18326 5714 18337 5748
rect 18281 5676 18337 5714
rect 18281 5642 18292 5676
rect 18326 5642 18337 5676
rect 18281 5604 18337 5642
rect 18281 5570 18292 5604
rect 18326 5570 18337 5604
rect 18281 5532 18337 5570
rect 18281 5498 18292 5532
rect 18326 5498 18337 5532
rect 18281 5460 18337 5498
rect 18281 5426 18292 5460
rect 18326 5426 18337 5460
rect 18281 5388 18337 5426
rect 18281 5354 18292 5388
rect 18326 5354 18337 5388
rect 18281 5316 18337 5354
rect 18281 5282 18292 5316
rect 18326 5282 18337 5316
rect 18281 5233 18337 5282
rect 18367 6180 18423 6233
rect 18367 6146 18378 6180
rect 18412 6146 18423 6180
rect 18367 6108 18423 6146
rect 18367 6074 18378 6108
rect 18412 6074 18423 6108
rect 18367 6036 18423 6074
rect 18367 6002 18378 6036
rect 18412 6002 18423 6036
rect 18367 5964 18423 6002
rect 18367 5930 18378 5964
rect 18412 5930 18423 5964
rect 18367 5892 18423 5930
rect 18367 5858 18378 5892
rect 18412 5858 18423 5892
rect 18367 5820 18423 5858
rect 18367 5786 18378 5820
rect 18412 5786 18423 5820
rect 18367 5748 18423 5786
rect 18367 5714 18378 5748
rect 18412 5714 18423 5748
rect 18367 5676 18423 5714
rect 18367 5642 18378 5676
rect 18412 5642 18423 5676
rect 18367 5604 18423 5642
rect 18367 5570 18378 5604
rect 18412 5570 18423 5604
rect 18367 5532 18423 5570
rect 18367 5498 18378 5532
rect 18412 5498 18423 5532
rect 18367 5460 18423 5498
rect 18367 5426 18378 5460
rect 18412 5426 18423 5460
rect 18367 5388 18423 5426
rect 18367 5354 18378 5388
rect 18412 5354 18423 5388
rect 18367 5316 18423 5354
rect 18367 5282 18378 5316
rect 18412 5282 18423 5316
rect 18367 5233 18423 5282
rect 18453 6180 18509 6233
rect 18453 6146 18464 6180
rect 18498 6146 18509 6180
rect 18453 6108 18509 6146
rect 18453 6074 18464 6108
rect 18498 6074 18509 6108
rect 18453 6036 18509 6074
rect 18453 6002 18464 6036
rect 18498 6002 18509 6036
rect 18453 5964 18509 6002
rect 18453 5930 18464 5964
rect 18498 5930 18509 5964
rect 18453 5892 18509 5930
rect 18453 5858 18464 5892
rect 18498 5858 18509 5892
rect 18453 5820 18509 5858
rect 18453 5786 18464 5820
rect 18498 5786 18509 5820
rect 18453 5748 18509 5786
rect 18453 5714 18464 5748
rect 18498 5714 18509 5748
rect 18453 5676 18509 5714
rect 18453 5642 18464 5676
rect 18498 5642 18509 5676
rect 18453 5604 18509 5642
rect 18453 5570 18464 5604
rect 18498 5570 18509 5604
rect 18453 5532 18509 5570
rect 18453 5498 18464 5532
rect 18498 5498 18509 5532
rect 18453 5460 18509 5498
rect 18453 5426 18464 5460
rect 18498 5426 18509 5460
rect 18453 5388 18509 5426
rect 18453 5354 18464 5388
rect 18498 5354 18509 5388
rect 18453 5316 18509 5354
rect 18453 5282 18464 5316
rect 18498 5282 18509 5316
rect 18453 5233 18509 5282
rect 18539 6180 18595 6233
rect 18539 6146 18550 6180
rect 18584 6146 18595 6180
rect 18539 6108 18595 6146
rect 18539 6074 18550 6108
rect 18584 6074 18595 6108
rect 18539 6036 18595 6074
rect 18539 6002 18550 6036
rect 18584 6002 18595 6036
rect 18539 5964 18595 6002
rect 18539 5930 18550 5964
rect 18584 5930 18595 5964
rect 18539 5892 18595 5930
rect 18539 5858 18550 5892
rect 18584 5858 18595 5892
rect 18539 5820 18595 5858
rect 18539 5786 18550 5820
rect 18584 5786 18595 5820
rect 18539 5748 18595 5786
rect 18539 5714 18550 5748
rect 18584 5714 18595 5748
rect 18539 5676 18595 5714
rect 18539 5642 18550 5676
rect 18584 5642 18595 5676
rect 18539 5604 18595 5642
rect 18539 5570 18550 5604
rect 18584 5570 18595 5604
rect 18539 5532 18595 5570
rect 18539 5498 18550 5532
rect 18584 5498 18595 5532
rect 18539 5460 18595 5498
rect 18539 5426 18550 5460
rect 18584 5426 18595 5460
rect 18539 5388 18595 5426
rect 18539 5354 18550 5388
rect 18584 5354 18595 5388
rect 18539 5316 18595 5354
rect 18539 5282 18550 5316
rect 18584 5282 18595 5316
rect 18539 5233 18595 5282
rect 18625 6180 18681 6233
rect 18625 6146 18636 6180
rect 18670 6146 18681 6180
rect 18625 6108 18681 6146
rect 18625 6074 18636 6108
rect 18670 6074 18681 6108
rect 18625 6036 18681 6074
rect 18625 6002 18636 6036
rect 18670 6002 18681 6036
rect 18625 5964 18681 6002
rect 18625 5930 18636 5964
rect 18670 5930 18681 5964
rect 18625 5892 18681 5930
rect 18625 5858 18636 5892
rect 18670 5858 18681 5892
rect 18625 5820 18681 5858
rect 18625 5786 18636 5820
rect 18670 5786 18681 5820
rect 18625 5748 18681 5786
rect 18625 5714 18636 5748
rect 18670 5714 18681 5748
rect 18625 5676 18681 5714
rect 18625 5642 18636 5676
rect 18670 5642 18681 5676
rect 18625 5604 18681 5642
rect 18625 5570 18636 5604
rect 18670 5570 18681 5604
rect 18625 5532 18681 5570
rect 18625 5498 18636 5532
rect 18670 5498 18681 5532
rect 18625 5460 18681 5498
rect 18625 5426 18636 5460
rect 18670 5426 18681 5460
rect 18625 5388 18681 5426
rect 18625 5354 18636 5388
rect 18670 5354 18681 5388
rect 18625 5316 18681 5354
rect 18625 5282 18636 5316
rect 18670 5282 18681 5316
rect 18625 5233 18681 5282
rect 18711 6180 18767 6233
rect 18711 6146 18722 6180
rect 18756 6146 18767 6180
rect 18711 6108 18767 6146
rect 18711 6074 18722 6108
rect 18756 6074 18767 6108
rect 18711 6036 18767 6074
rect 18711 6002 18722 6036
rect 18756 6002 18767 6036
rect 18711 5964 18767 6002
rect 18711 5930 18722 5964
rect 18756 5930 18767 5964
rect 18711 5892 18767 5930
rect 18711 5858 18722 5892
rect 18756 5858 18767 5892
rect 18711 5820 18767 5858
rect 18711 5786 18722 5820
rect 18756 5786 18767 5820
rect 18711 5748 18767 5786
rect 18711 5714 18722 5748
rect 18756 5714 18767 5748
rect 18711 5676 18767 5714
rect 18711 5642 18722 5676
rect 18756 5642 18767 5676
rect 18711 5604 18767 5642
rect 18711 5570 18722 5604
rect 18756 5570 18767 5604
rect 18711 5532 18767 5570
rect 18711 5498 18722 5532
rect 18756 5498 18767 5532
rect 18711 5460 18767 5498
rect 18711 5426 18722 5460
rect 18756 5426 18767 5460
rect 18711 5388 18767 5426
rect 18711 5354 18722 5388
rect 18756 5354 18767 5388
rect 18711 5316 18767 5354
rect 18711 5282 18722 5316
rect 18756 5282 18767 5316
rect 18711 5233 18767 5282
rect 18797 6180 18853 6233
rect 18797 6146 18808 6180
rect 18842 6146 18853 6180
rect 18797 6108 18853 6146
rect 18797 6074 18808 6108
rect 18842 6074 18853 6108
rect 18797 6036 18853 6074
rect 18797 6002 18808 6036
rect 18842 6002 18853 6036
rect 18797 5964 18853 6002
rect 18797 5930 18808 5964
rect 18842 5930 18853 5964
rect 18797 5892 18853 5930
rect 18797 5858 18808 5892
rect 18842 5858 18853 5892
rect 18797 5820 18853 5858
rect 18797 5786 18808 5820
rect 18842 5786 18853 5820
rect 18797 5748 18853 5786
rect 18797 5714 18808 5748
rect 18842 5714 18853 5748
rect 18797 5676 18853 5714
rect 18797 5642 18808 5676
rect 18842 5642 18853 5676
rect 18797 5604 18853 5642
rect 18797 5570 18808 5604
rect 18842 5570 18853 5604
rect 18797 5532 18853 5570
rect 18797 5498 18808 5532
rect 18842 5498 18853 5532
rect 18797 5460 18853 5498
rect 18797 5426 18808 5460
rect 18842 5426 18853 5460
rect 18797 5388 18853 5426
rect 18797 5354 18808 5388
rect 18842 5354 18853 5388
rect 18797 5316 18853 5354
rect 18797 5282 18808 5316
rect 18842 5282 18853 5316
rect 18797 5233 18853 5282
rect 18883 6180 18939 6233
rect 18883 6146 18894 6180
rect 18928 6146 18939 6180
rect 18883 6108 18939 6146
rect 18883 6074 18894 6108
rect 18928 6074 18939 6108
rect 18883 6036 18939 6074
rect 18883 6002 18894 6036
rect 18928 6002 18939 6036
rect 18883 5964 18939 6002
rect 18883 5930 18894 5964
rect 18928 5930 18939 5964
rect 18883 5892 18939 5930
rect 18883 5858 18894 5892
rect 18928 5858 18939 5892
rect 18883 5820 18939 5858
rect 18883 5786 18894 5820
rect 18928 5786 18939 5820
rect 18883 5748 18939 5786
rect 18883 5714 18894 5748
rect 18928 5714 18939 5748
rect 18883 5676 18939 5714
rect 18883 5642 18894 5676
rect 18928 5642 18939 5676
rect 18883 5604 18939 5642
rect 18883 5570 18894 5604
rect 18928 5570 18939 5604
rect 18883 5532 18939 5570
rect 18883 5498 18894 5532
rect 18928 5498 18939 5532
rect 18883 5460 18939 5498
rect 18883 5426 18894 5460
rect 18928 5426 18939 5460
rect 18883 5388 18939 5426
rect 18883 5354 18894 5388
rect 18928 5354 18939 5388
rect 18883 5316 18939 5354
rect 18883 5282 18894 5316
rect 18928 5282 18939 5316
rect 18883 5233 18939 5282
rect 18969 6180 19025 6233
rect 18969 6146 18980 6180
rect 19014 6146 19025 6180
rect 18969 6108 19025 6146
rect 18969 6074 18980 6108
rect 19014 6074 19025 6108
rect 18969 6036 19025 6074
rect 18969 6002 18980 6036
rect 19014 6002 19025 6036
rect 18969 5964 19025 6002
rect 18969 5930 18980 5964
rect 19014 5930 19025 5964
rect 18969 5892 19025 5930
rect 18969 5858 18980 5892
rect 19014 5858 19025 5892
rect 18969 5820 19025 5858
rect 18969 5786 18980 5820
rect 19014 5786 19025 5820
rect 18969 5748 19025 5786
rect 18969 5714 18980 5748
rect 19014 5714 19025 5748
rect 18969 5676 19025 5714
rect 18969 5642 18980 5676
rect 19014 5642 19025 5676
rect 18969 5604 19025 5642
rect 18969 5570 18980 5604
rect 19014 5570 19025 5604
rect 18969 5532 19025 5570
rect 18969 5498 18980 5532
rect 19014 5498 19025 5532
rect 18969 5460 19025 5498
rect 18969 5426 18980 5460
rect 19014 5426 19025 5460
rect 18969 5388 19025 5426
rect 18969 5354 18980 5388
rect 19014 5354 19025 5388
rect 18969 5316 19025 5354
rect 18969 5282 18980 5316
rect 19014 5282 19025 5316
rect 18969 5233 19025 5282
rect 19055 6180 19111 6233
rect 19055 6146 19066 6180
rect 19100 6146 19111 6180
rect 19055 6108 19111 6146
rect 19055 6074 19066 6108
rect 19100 6074 19111 6108
rect 19055 6036 19111 6074
rect 19055 6002 19066 6036
rect 19100 6002 19111 6036
rect 19055 5964 19111 6002
rect 19055 5930 19066 5964
rect 19100 5930 19111 5964
rect 19055 5892 19111 5930
rect 19055 5858 19066 5892
rect 19100 5858 19111 5892
rect 19055 5820 19111 5858
rect 19055 5786 19066 5820
rect 19100 5786 19111 5820
rect 19055 5748 19111 5786
rect 19055 5714 19066 5748
rect 19100 5714 19111 5748
rect 19055 5676 19111 5714
rect 19055 5642 19066 5676
rect 19100 5642 19111 5676
rect 19055 5604 19111 5642
rect 19055 5570 19066 5604
rect 19100 5570 19111 5604
rect 19055 5532 19111 5570
rect 19055 5498 19066 5532
rect 19100 5498 19111 5532
rect 19055 5460 19111 5498
rect 19055 5426 19066 5460
rect 19100 5426 19111 5460
rect 19055 5388 19111 5426
rect 19055 5354 19066 5388
rect 19100 5354 19111 5388
rect 19055 5316 19111 5354
rect 19055 5282 19066 5316
rect 19100 5282 19111 5316
rect 19055 5233 19111 5282
rect 19141 6180 19197 6233
rect 19141 6146 19152 6180
rect 19186 6146 19197 6180
rect 19141 6108 19197 6146
rect 19141 6074 19152 6108
rect 19186 6074 19197 6108
rect 19141 6036 19197 6074
rect 19141 6002 19152 6036
rect 19186 6002 19197 6036
rect 19141 5964 19197 6002
rect 19141 5930 19152 5964
rect 19186 5930 19197 5964
rect 19141 5892 19197 5930
rect 19141 5858 19152 5892
rect 19186 5858 19197 5892
rect 19141 5820 19197 5858
rect 19141 5786 19152 5820
rect 19186 5786 19197 5820
rect 19141 5748 19197 5786
rect 19141 5714 19152 5748
rect 19186 5714 19197 5748
rect 19141 5676 19197 5714
rect 19141 5642 19152 5676
rect 19186 5642 19197 5676
rect 19141 5604 19197 5642
rect 19141 5570 19152 5604
rect 19186 5570 19197 5604
rect 19141 5532 19197 5570
rect 19141 5498 19152 5532
rect 19186 5498 19197 5532
rect 19141 5460 19197 5498
rect 19141 5426 19152 5460
rect 19186 5426 19197 5460
rect 19141 5388 19197 5426
rect 19141 5354 19152 5388
rect 19186 5354 19197 5388
rect 19141 5316 19197 5354
rect 19141 5282 19152 5316
rect 19186 5282 19197 5316
rect 19141 5233 19197 5282
rect 19227 6180 19283 6233
rect 19227 6146 19238 6180
rect 19272 6146 19283 6180
rect 19227 6108 19283 6146
rect 19227 6074 19238 6108
rect 19272 6074 19283 6108
rect 19227 6036 19283 6074
rect 19227 6002 19238 6036
rect 19272 6002 19283 6036
rect 19227 5964 19283 6002
rect 19227 5930 19238 5964
rect 19272 5930 19283 5964
rect 19227 5892 19283 5930
rect 19227 5858 19238 5892
rect 19272 5858 19283 5892
rect 19227 5820 19283 5858
rect 19227 5786 19238 5820
rect 19272 5786 19283 5820
rect 19227 5748 19283 5786
rect 19227 5714 19238 5748
rect 19272 5714 19283 5748
rect 19227 5676 19283 5714
rect 19227 5642 19238 5676
rect 19272 5642 19283 5676
rect 19227 5604 19283 5642
rect 19227 5570 19238 5604
rect 19272 5570 19283 5604
rect 19227 5532 19283 5570
rect 19227 5498 19238 5532
rect 19272 5498 19283 5532
rect 19227 5460 19283 5498
rect 19227 5426 19238 5460
rect 19272 5426 19283 5460
rect 19227 5388 19283 5426
rect 19227 5354 19238 5388
rect 19272 5354 19283 5388
rect 19227 5316 19283 5354
rect 19227 5282 19238 5316
rect 19272 5282 19283 5316
rect 19227 5233 19283 5282
rect 19313 6180 19369 6233
rect 19313 6146 19324 6180
rect 19358 6146 19369 6180
rect 19313 6108 19369 6146
rect 19313 6074 19324 6108
rect 19358 6074 19369 6108
rect 19313 6036 19369 6074
rect 19313 6002 19324 6036
rect 19358 6002 19369 6036
rect 19313 5964 19369 6002
rect 19313 5930 19324 5964
rect 19358 5930 19369 5964
rect 19313 5892 19369 5930
rect 19313 5858 19324 5892
rect 19358 5858 19369 5892
rect 19313 5820 19369 5858
rect 19313 5786 19324 5820
rect 19358 5786 19369 5820
rect 19313 5748 19369 5786
rect 19313 5714 19324 5748
rect 19358 5714 19369 5748
rect 19313 5676 19369 5714
rect 19313 5642 19324 5676
rect 19358 5642 19369 5676
rect 19313 5604 19369 5642
rect 19313 5570 19324 5604
rect 19358 5570 19369 5604
rect 19313 5532 19369 5570
rect 19313 5498 19324 5532
rect 19358 5498 19369 5532
rect 19313 5460 19369 5498
rect 19313 5426 19324 5460
rect 19358 5426 19369 5460
rect 19313 5388 19369 5426
rect 19313 5354 19324 5388
rect 19358 5354 19369 5388
rect 19313 5316 19369 5354
rect 19313 5282 19324 5316
rect 19358 5282 19369 5316
rect 19313 5233 19369 5282
rect 19399 6180 19455 6233
rect 19399 6146 19410 6180
rect 19444 6146 19455 6180
rect 19399 6108 19455 6146
rect 19399 6074 19410 6108
rect 19444 6074 19455 6108
rect 19399 6036 19455 6074
rect 19399 6002 19410 6036
rect 19444 6002 19455 6036
rect 19399 5964 19455 6002
rect 19399 5930 19410 5964
rect 19444 5930 19455 5964
rect 19399 5892 19455 5930
rect 19399 5858 19410 5892
rect 19444 5858 19455 5892
rect 19399 5820 19455 5858
rect 19399 5786 19410 5820
rect 19444 5786 19455 5820
rect 19399 5748 19455 5786
rect 19399 5714 19410 5748
rect 19444 5714 19455 5748
rect 19399 5676 19455 5714
rect 19399 5642 19410 5676
rect 19444 5642 19455 5676
rect 19399 5604 19455 5642
rect 19399 5570 19410 5604
rect 19444 5570 19455 5604
rect 19399 5532 19455 5570
rect 19399 5498 19410 5532
rect 19444 5498 19455 5532
rect 19399 5460 19455 5498
rect 19399 5426 19410 5460
rect 19444 5426 19455 5460
rect 19399 5388 19455 5426
rect 19399 5354 19410 5388
rect 19444 5354 19455 5388
rect 19399 5316 19455 5354
rect 19399 5282 19410 5316
rect 19444 5282 19455 5316
rect 19399 5233 19455 5282
rect 19485 6180 19541 6233
rect 19485 6146 19496 6180
rect 19530 6146 19541 6180
rect 19485 6108 19541 6146
rect 19485 6074 19496 6108
rect 19530 6074 19541 6108
rect 19485 6036 19541 6074
rect 19485 6002 19496 6036
rect 19530 6002 19541 6036
rect 19485 5964 19541 6002
rect 19485 5930 19496 5964
rect 19530 5930 19541 5964
rect 19485 5892 19541 5930
rect 19485 5858 19496 5892
rect 19530 5858 19541 5892
rect 19485 5820 19541 5858
rect 19485 5786 19496 5820
rect 19530 5786 19541 5820
rect 19485 5748 19541 5786
rect 19485 5714 19496 5748
rect 19530 5714 19541 5748
rect 19485 5676 19541 5714
rect 19485 5642 19496 5676
rect 19530 5642 19541 5676
rect 19485 5604 19541 5642
rect 19485 5570 19496 5604
rect 19530 5570 19541 5604
rect 19485 5532 19541 5570
rect 19485 5498 19496 5532
rect 19530 5498 19541 5532
rect 19485 5460 19541 5498
rect 19485 5426 19496 5460
rect 19530 5426 19541 5460
rect 19485 5388 19541 5426
rect 19485 5354 19496 5388
rect 19530 5354 19541 5388
rect 19485 5316 19541 5354
rect 19485 5282 19496 5316
rect 19530 5282 19541 5316
rect 19485 5233 19541 5282
rect 19571 6180 19627 6233
rect 19571 6146 19582 6180
rect 19616 6146 19627 6180
rect 19571 6108 19627 6146
rect 19571 6074 19582 6108
rect 19616 6074 19627 6108
rect 19571 6036 19627 6074
rect 19571 6002 19582 6036
rect 19616 6002 19627 6036
rect 19571 5964 19627 6002
rect 19571 5930 19582 5964
rect 19616 5930 19627 5964
rect 19571 5892 19627 5930
rect 19571 5858 19582 5892
rect 19616 5858 19627 5892
rect 19571 5820 19627 5858
rect 19571 5786 19582 5820
rect 19616 5786 19627 5820
rect 19571 5748 19627 5786
rect 19571 5714 19582 5748
rect 19616 5714 19627 5748
rect 19571 5676 19627 5714
rect 19571 5642 19582 5676
rect 19616 5642 19627 5676
rect 19571 5604 19627 5642
rect 19571 5570 19582 5604
rect 19616 5570 19627 5604
rect 19571 5532 19627 5570
rect 19571 5498 19582 5532
rect 19616 5498 19627 5532
rect 19571 5460 19627 5498
rect 19571 5426 19582 5460
rect 19616 5426 19627 5460
rect 19571 5388 19627 5426
rect 19571 5354 19582 5388
rect 19616 5354 19627 5388
rect 19571 5316 19627 5354
rect 19571 5282 19582 5316
rect 19616 5282 19627 5316
rect 19571 5233 19627 5282
rect 19657 6180 19713 6233
rect 19657 6146 19668 6180
rect 19702 6146 19713 6180
rect 19657 6108 19713 6146
rect 19657 6074 19668 6108
rect 19702 6074 19713 6108
rect 19657 6036 19713 6074
rect 19657 6002 19668 6036
rect 19702 6002 19713 6036
rect 19657 5964 19713 6002
rect 19657 5930 19668 5964
rect 19702 5930 19713 5964
rect 19657 5892 19713 5930
rect 19657 5858 19668 5892
rect 19702 5858 19713 5892
rect 19657 5820 19713 5858
rect 19657 5786 19668 5820
rect 19702 5786 19713 5820
rect 19657 5748 19713 5786
rect 19657 5714 19668 5748
rect 19702 5714 19713 5748
rect 19657 5676 19713 5714
rect 19657 5642 19668 5676
rect 19702 5642 19713 5676
rect 19657 5604 19713 5642
rect 19657 5570 19668 5604
rect 19702 5570 19713 5604
rect 19657 5532 19713 5570
rect 19657 5498 19668 5532
rect 19702 5498 19713 5532
rect 19657 5460 19713 5498
rect 19657 5426 19668 5460
rect 19702 5426 19713 5460
rect 19657 5388 19713 5426
rect 19657 5354 19668 5388
rect 19702 5354 19713 5388
rect 19657 5316 19713 5354
rect 19657 5282 19668 5316
rect 19702 5282 19713 5316
rect 19657 5233 19713 5282
rect 19743 6180 19799 6233
rect 19743 6146 19754 6180
rect 19788 6146 19799 6180
rect 19743 6108 19799 6146
rect 19743 6074 19754 6108
rect 19788 6074 19799 6108
rect 19743 6036 19799 6074
rect 19743 6002 19754 6036
rect 19788 6002 19799 6036
rect 19743 5964 19799 6002
rect 19743 5930 19754 5964
rect 19788 5930 19799 5964
rect 19743 5892 19799 5930
rect 19743 5858 19754 5892
rect 19788 5858 19799 5892
rect 19743 5820 19799 5858
rect 19743 5786 19754 5820
rect 19788 5786 19799 5820
rect 19743 5748 19799 5786
rect 19743 5714 19754 5748
rect 19788 5714 19799 5748
rect 19743 5676 19799 5714
rect 19743 5642 19754 5676
rect 19788 5642 19799 5676
rect 19743 5604 19799 5642
rect 19743 5570 19754 5604
rect 19788 5570 19799 5604
rect 19743 5532 19799 5570
rect 19743 5498 19754 5532
rect 19788 5498 19799 5532
rect 19743 5460 19799 5498
rect 19743 5426 19754 5460
rect 19788 5426 19799 5460
rect 19743 5388 19799 5426
rect 19743 5354 19754 5388
rect 19788 5354 19799 5388
rect 19743 5316 19799 5354
rect 19743 5282 19754 5316
rect 19788 5282 19799 5316
rect 19743 5233 19799 5282
rect 19829 6180 19885 6233
rect 19829 6146 19840 6180
rect 19874 6146 19885 6180
rect 19829 6108 19885 6146
rect 19829 6074 19840 6108
rect 19874 6074 19885 6108
rect 19829 6036 19885 6074
rect 19829 6002 19840 6036
rect 19874 6002 19885 6036
rect 19829 5964 19885 6002
rect 19829 5930 19840 5964
rect 19874 5930 19885 5964
rect 19829 5892 19885 5930
rect 19829 5858 19840 5892
rect 19874 5858 19885 5892
rect 19829 5820 19885 5858
rect 19829 5786 19840 5820
rect 19874 5786 19885 5820
rect 19829 5748 19885 5786
rect 19829 5714 19840 5748
rect 19874 5714 19885 5748
rect 19829 5676 19885 5714
rect 19829 5642 19840 5676
rect 19874 5642 19885 5676
rect 19829 5604 19885 5642
rect 19829 5570 19840 5604
rect 19874 5570 19885 5604
rect 19829 5532 19885 5570
rect 19829 5498 19840 5532
rect 19874 5498 19885 5532
rect 19829 5460 19885 5498
rect 19829 5426 19840 5460
rect 19874 5426 19885 5460
rect 19829 5388 19885 5426
rect 19829 5354 19840 5388
rect 19874 5354 19885 5388
rect 19829 5316 19885 5354
rect 19829 5282 19840 5316
rect 19874 5282 19885 5316
rect 19829 5233 19885 5282
rect 19915 6180 19971 6233
rect 19915 6146 19926 6180
rect 19960 6146 19971 6180
rect 19915 6108 19971 6146
rect 19915 6074 19926 6108
rect 19960 6074 19971 6108
rect 19915 6036 19971 6074
rect 19915 6002 19926 6036
rect 19960 6002 19971 6036
rect 19915 5964 19971 6002
rect 19915 5930 19926 5964
rect 19960 5930 19971 5964
rect 19915 5892 19971 5930
rect 19915 5858 19926 5892
rect 19960 5858 19971 5892
rect 19915 5820 19971 5858
rect 19915 5786 19926 5820
rect 19960 5786 19971 5820
rect 19915 5748 19971 5786
rect 19915 5714 19926 5748
rect 19960 5714 19971 5748
rect 19915 5676 19971 5714
rect 19915 5642 19926 5676
rect 19960 5642 19971 5676
rect 19915 5604 19971 5642
rect 19915 5570 19926 5604
rect 19960 5570 19971 5604
rect 19915 5532 19971 5570
rect 19915 5498 19926 5532
rect 19960 5498 19971 5532
rect 19915 5460 19971 5498
rect 19915 5426 19926 5460
rect 19960 5426 19971 5460
rect 19915 5388 19971 5426
rect 19915 5354 19926 5388
rect 19960 5354 19971 5388
rect 19915 5316 19971 5354
rect 19915 5282 19926 5316
rect 19960 5282 19971 5316
rect 19915 5233 19971 5282
rect 20001 6180 20054 6233
rect 20001 6146 20012 6180
rect 20046 6146 20054 6180
rect 20001 6108 20054 6146
rect 20001 6074 20012 6108
rect 20046 6074 20054 6108
rect 20001 6036 20054 6074
rect 20001 6002 20012 6036
rect 20046 6002 20054 6036
rect 20001 5964 20054 6002
rect 20001 5930 20012 5964
rect 20046 5930 20054 5964
rect 20001 5892 20054 5930
rect 20001 5858 20012 5892
rect 20046 5858 20054 5892
rect 20001 5820 20054 5858
rect 20001 5786 20012 5820
rect 20046 5786 20054 5820
rect 20001 5748 20054 5786
rect 20001 5714 20012 5748
rect 20046 5714 20054 5748
rect 20001 5676 20054 5714
rect 20001 5642 20012 5676
rect 20046 5642 20054 5676
rect 20001 5604 20054 5642
rect 20001 5570 20012 5604
rect 20046 5570 20054 5604
rect 20001 5532 20054 5570
rect 20001 5498 20012 5532
rect 20046 5498 20054 5532
rect 20001 5460 20054 5498
rect 20001 5426 20012 5460
rect 20046 5426 20054 5460
rect 20001 5388 20054 5426
rect 20001 5354 20012 5388
rect 20046 5354 20054 5388
rect 20001 5316 20054 5354
rect 20001 5282 20012 5316
rect 20046 5282 20054 5316
rect 20001 5233 20054 5282
<< ndiffc >>
rect 16118 7933 16152 7967
rect 16118 7865 16152 7899
rect 16118 7797 16152 7831
rect 16118 7729 16152 7763
rect 16118 7661 16152 7695
rect 16118 7593 16152 7627
rect 16118 7525 16152 7559
rect 16118 7457 16152 7491
rect 16118 7389 16152 7423
rect 16118 7321 16152 7355
rect 16118 7253 16152 7287
rect 16118 7185 16152 7219
rect 16118 7117 16152 7151
rect 16118 7049 16152 7083
rect 16118 6981 16152 7015
rect 16204 7933 16238 7967
rect 16204 7865 16238 7899
rect 16204 7797 16238 7831
rect 16204 7729 16238 7763
rect 16204 7661 16238 7695
rect 16204 7593 16238 7627
rect 16204 7525 16238 7559
rect 16204 7457 16238 7491
rect 16204 7389 16238 7423
rect 16204 7321 16238 7355
rect 16204 7253 16238 7287
rect 16204 7185 16238 7219
rect 16204 7117 16238 7151
rect 16204 7049 16238 7083
rect 16204 6981 16238 7015
rect 16290 7933 16324 7967
rect 16290 7865 16324 7899
rect 16290 7797 16324 7831
rect 16290 7729 16324 7763
rect 16290 7661 16324 7695
rect 16290 7593 16324 7627
rect 16290 7525 16324 7559
rect 16290 7457 16324 7491
rect 16290 7389 16324 7423
rect 16290 7321 16324 7355
rect 16290 7253 16324 7287
rect 16290 7185 16324 7219
rect 16290 7117 16324 7151
rect 16290 7049 16324 7083
rect 16290 6981 16324 7015
rect 16376 7933 16410 7967
rect 16376 7865 16410 7899
rect 16376 7797 16410 7831
rect 16376 7729 16410 7763
rect 16376 7661 16410 7695
rect 16376 7593 16410 7627
rect 16376 7525 16410 7559
rect 16376 7457 16410 7491
rect 16376 7389 16410 7423
rect 16376 7321 16410 7355
rect 16376 7253 16410 7287
rect 16376 7185 16410 7219
rect 16376 7117 16410 7151
rect 16376 7049 16410 7083
rect 16376 6981 16410 7015
rect 16462 7933 16496 7967
rect 16462 7865 16496 7899
rect 16462 7797 16496 7831
rect 16462 7729 16496 7763
rect 16462 7661 16496 7695
rect 16462 7593 16496 7627
rect 16462 7525 16496 7559
rect 16462 7457 16496 7491
rect 16462 7389 16496 7423
rect 16462 7321 16496 7355
rect 16462 7253 16496 7287
rect 16462 7185 16496 7219
rect 16462 7117 16496 7151
rect 16462 7049 16496 7083
rect 16462 6981 16496 7015
rect 16548 7933 16582 7967
rect 16548 7865 16582 7899
rect 16548 7797 16582 7831
rect 16548 7729 16582 7763
rect 16548 7661 16582 7695
rect 16548 7593 16582 7627
rect 16548 7525 16582 7559
rect 16548 7457 16582 7491
rect 16548 7389 16582 7423
rect 16548 7321 16582 7355
rect 16548 7253 16582 7287
rect 16548 7185 16582 7219
rect 16548 7117 16582 7151
rect 16548 7049 16582 7083
rect 16548 6981 16582 7015
rect 16634 7933 16668 7967
rect 16634 7865 16668 7899
rect 16634 7797 16668 7831
rect 16634 7729 16668 7763
rect 16634 7661 16668 7695
rect 16634 7593 16668 7627
rect 16634 7525 16668 7559
rect 16634 7457 16668 7491
rect 16634 7389 16668 7423
rect 16634 7321 16668 7355
rect 16634 7253 16668 7287
rect 16634 7185 16668 7219
rect 16634 7117 16668 7151
rect 16634 7049 16668 7083
rect 16634 6981 16668 7015
rect 16720 7933 16754 7967
rect 16720 7865 16754 7899
rect 16720 7797 16754 7831
rect 16720 7729 16754 7763
rect 16720 7661 16754 7695
rect 16720 7593 16754 7627
rect 16720 7525 16754 7559
rect 16720 7457 16754 7491
rect 16720 7389 16754 7423
rect 16720 7321 16754 7355
rect 16720 7253 16754 7287
rect 16720 7185 16754 7219
rect 16720 7117 16754 7151
rect 16720 7049 16754 7083
rect 16720 6981 16754 7015
rect 16806 7933 16840 7967
rect 16806 7865 16840 7899
rect 16806 7797 16840 7831
rect 16806 7729 16840 7763
rect 16806 7661 16840 7695
rect 16806 7593 16840 7627
rect 16806 7525 16840 7559
rect 16806 7457 16840 7491
rect 16806 7389 16840 7423
rect 16806 7321 16840 7355
rect 16806 7253 16840 7287
rect 16806 7185 16840 7219
rect 16806 7117 16840 7151
rect 16806 7049 16840 7083
rect 16806 6981 16840 7015
rect 16892 7933 16926 7967
rect 16892 7865 16926 7899
rect 16892 7797 16926 7831
rect 16892 7729 16926 7763
rect 16892 7661 16926 7695
rect 16892 7593 16926 7627
rect 16892 7525 16926 7559
rect 16892 7457 16926 7491
rect 16892 7389 16926 7423
rect 16892 7321 16926 7355
rect 16892 7253 16926 7287
rect 16892 7185 16926 7219
rect 16892 7117 16926 7151
rect 16892 7049 16926 7083
rect 16892 6981 16926 7015
rect 16978 7933 17012 7967
rect 16978 7865 17012 7899
rect 16978 7797 17012 7831
rect 16978 7729 17012 7763
rect 16978 7661 17012 7695
rect 16978 7593 17012 7627
rect 16978 7525 17012 7559
rect 16978 7457 17012 7491
rect 16978 7389 17012 7423
rect 16978 7321 17012 7355
rect 16978 7253 17012 7287
rect 16978 7185 17012 7219
rect 16978 7117 17012 7151
rect 16978 7049 17012 7083
rect 16978 6981 17012 7015
rect 17064 7933 17098 7967
rect 17064 7865 17098 7899
rect 17064 7797 17098 7831
rect 17064 7729 17098 7763
rect 17064 7661 17098 7695
rect 17064 7593 17098 7627
rect 17064 7525 17098 7559
rect 17064 7457 17098 7491
rect 17064 7389 17098 7423
rect 17064 7321 17098 7355
rect 17064 7253 17098 7287
rect 17064 7185 17098 7219
rect 17064 7117 17098 7151
rect 17064 7049 17098 7083
rect 17064 6981 17098 7015
rect 17150 7933 17184 7967
rect 17150 7865 17184 7899
rect 17150 7797 17184 7831
rect 17150 7729 17184 7763
rect 17150 7661 17184 7695
rect 17150 7593 17184 7627
rect 17150 7525 17184 7559
rect 17150 7457 17184 7491
rect 17150 7389 17184 7423
rect 17150 7321 17184 7355
rect 17150 7253 17184 7287
rect 17150 7185 17184 7219
rect 17150 7117 17184 7151
rect 17150 7049 17184 7083
rect 17150 6981 17184 7015
rect 11785 6812 11819 6846
rect 11785 6744 11819 6778
rect 11785 6676 11819 6710
rect 11785 6608 11819 6642
rect 11785 6540 11819 6574
rect 11785 6472 11819 6506
rect 11785 6404 11819 6438
rect 11785 6336 11819 6370
rect 11785 6268 11819 6302
rect 11785 6200 11819 6234
rect 11785 6132 11819 6166
rect 11785 6064 11819 6098
rect 11785 5996 11819 6030
rect 11785 5928 11819 5962
rect 11785 5860 11819 5894
rect 11871 6812 11905 6846
rect 11871 6744 11905 6778
rect 11871 6676 11905 6710
rect 11871 6608 11905 6642
rect 11871 6540 11905 6574
rect 11871 6472 11905 6506
rect 11871 6404 11905 6438
rect 11871 6336 11905 6370
rect 11871 6268 11905 6302
rect 11871 6200 11905 6234
rect 11871 6132 11905 6166
rect 11871 6064 11905 6098
rect 11871 5996 11905 6030
rect 11871 5928 11905 5962
rect 11871 5860 11905 5894
rect 11957 6812 11991 6846
rect 11957 6744 11991 6778
rect 11957 6676 11991 6710
rect 11957 6608 11991 6642
rect 11957 6540 11991 6574
rect 11957 6472 11991 6506
rect 11957 6404 11991 6438
rect 11957 6336 11991 6370
rect 11957 6268 11991 6302
rect 11957 6200 11991 6234
rect 11957 6132 11991 6166
rect 11957 6064 11991 6098
rect 11957 5996 11991 6030
rect 11957 5928 11991 5962
rect 11957 5860 11991 5894
rect 12043 6812 12077 6846
rect 12043 6744 12077 6778
rect 12043 6676 12077 6710
rect 12043 6608 12077 6642
rect 12043 6540 12077 6574
rect 12043 6472 12077 6506
rect 12043 6404 12077 6438
rect 12043 6336 12077 6370
rect 12043 6268 12077 6302
rect 12043 6200 12077 6234
rect 12043 6132 12077 6166
rect 12043 6064 12077 6098
rect 12043 5996 12077 6030
rect 12043 5928 12077 5962
rect 12043 5860 12077 5894
rect 12129 6812 12163 6846
rect 12129 6744 12163 6778
rect 12129 6676 12163 6710
rect 12129 6608 12163 6642
rect 12129 6540 12163 6574
rect 12129 6472 12163 6506
rect 12129 6404 12163 6438
rect 12129 6336 12163 6370
rect 12129 6268 12163 6302
rect 12129 6200 12163 6234
rect 12129 6132 12163 6166
rect 12129 6064 12163 6098
rect 12129 5996 12163 6030
rect 12129 5928 12163 5962
rect 12129 5860 12163 5894
rect 12351 6812 12385 6846
rect 12351 6744 12385 6778
rect 12351 6676 12385 6710
rect 12351 6608 12385 6642
rect 12351 6540 12385 6574
rect 12351 6472 12385 6506
rect 12351 6404 12385 6438
rect 12351 6336 12385 6370
rect 12351 6268 12385 6302
rect 12351 6200 12385 6234
rect 12351 6132 12385 6166
rect 12351 6064 12385 6098
rect 12351 5996 12385 6030
rect 12351 5928 12385 5962
rect 12351 5860 12385 5894
rect 12437 6812 12471 6846
rect 12437 6744 12471 6778
rect 12437 6676 12471 6710
rect 12437 6608 12471 6642
rect 12437 6540 12471 6574
rect 12437 6472 12471 6506
rect 12437 6404 12471 6438
rect 12437 6336 12471 6370
rect 12437 6268 12471 6302
rect 12437 6200 12471 6234
rect 12437 6132 12471 6166
rect 12437 6064 12471 6098
rect 12437 5996 12471 6030
rect 12437 5928 12471 5962
rect 12437 5860 12471 5894
rect 12523 6812 12557 6846
rect 12523 6744 12557 6778
rect 12523 6676 12557 6710
rect 12523 6608 12557 6642
rect 12523 6540 12557 6574
rect 12523 6472 12557 6506
rect 12523 6404 12557 6438
rect 12523 6336 12557 6370
rect 12523 6268 12557 6302
rect 12523 6200 12557 6234
rect 12523 6132 12557 6166
rect 12523 6064 12557 6098
rect 12523 5996 12557 6030
rect 12523 5928 12557 5962
rect 12523 5860 12557 5894
rect 12609 6812 12643 6846
rect 12609 6744 12643 6778
rect 12609 6676 12643 6710
rect 12609 6608 12643 6642
rect 12609 6540 12643 6574
rect 12609 6472 12643 6506
rect 12609 6404 12643 6438
rect 12609 6336 12643 6370
rect 12609 6268 12643 6302
rect 12609 6200 12643 6234
rect 12609 6132 12643 6166
rect 12609 6064 12643 6098
rect 12609 5996 12643 6030
rect 12609 5928 12643 5962
rect 12609 5860 12643 5894
rect 12695 6812 12729 6846
rect 12695 6744 12729 6778
rect 12695 6676 12729 6710
rect 12695 6608 12729 6642
rect 12695 6540 12729 6574
rect 12695 6472 12729 6506
rect 12695 6404 12729 6438
rect 12695 6336 12729 6370
rect 12695 6268 12729 6302
rect 12695 6200 12729 6234
rect 12695 6132 12729 6166
rect 12695 6064 12729 6098
rect 12695 5996 12729 6030
rect 12695 5928 12729 5962
rect 12695 5860 12729 5894
rect 12917 6812 12951 6846
rect 12917 6744 12951 6778
rect 12917 6676 12951 6710
rect 12917 6608 12951 6642
rect 12917 6540 12951 6574
rect 12917 6472 12951 6506
rect 12917 6404 12951 6438
rect 12917 6336 12951 6370
rect 12917 6268 12951 6302
rect 12917 6200 12951 6234
rect 12917 6132 12951 6166
rect 12917 6064 12951 6098
rect 12917 5996 12951 6030
rect 12917 5928 12951 5962
rect 12917 5860 12951 5894
rect 13003 6812 13037 6846
rect 13003 6744 13037 6778
rect 13003 6676 13037 6710
rect 13003 6608 13037 6642
rect 13003 6540 13037 6574
rect 13003 6472 13037 6506
rect 13003 6404 13037 6438
rect 13003 6336 13037 6370
rect 13003 6268 13037 6302
rect 13003 6200 13037 6234
rect 13003 6132 13037 6166
rect 13003 6064 13037 6098
rect 13003 5996 13037 6030
rect 13003 5928 13037 5962
rect 13003 5860 13037 5894
rect 13089 6812 13123 6846
rect 13089 6744 13123 6778
rect 13089 6676 13123 6710
rect 13089 6608 13123 6642
rect 13089 6540 13123 6574
rect 13089 6472 13123 6506
rect 13089 6404 13123 6438
rect 13089 6336 13123 6370
rect 13089 6268 13123 6302
rect 13089 6200 13123 6234
rect 13089 6132 13123 6166
rect 13089 6064 13123 6098
rect 13089 5996 13123 6030
rect 13089 5928 13123 5962
rect 13089 5860 13123 5894
rect 13175 6812 13209 6846
rect 13175 6744 13209 6778
rect 13175 6676 13209 6710
rect 13175 6608 13209 6642
rect 13175 6540 13209 6574
rect 13175 6472 13209 6506
rect 13175 6404 13209 6438
rect 13175 6336 13209 6370
rect 13175 6268 13209 6302
rect 13175 6200 13209 6234
rect 13175 6132 13209 6166
rect 13175 6064 13209 6098
rect 13175 5996 13209 6030
rect 13175 5928 13209 5962
rect 13175 5860 13209 5894
rect 13261 6812 13295 6846
rect 13261 6744 13295 6778
rect 13261 6676 13295 6710
rect 13261 6608 13295 6642
rect 13261 6540 13295 6574
rect 13261 6472 13295 6506
rect 13261 6404 13295 6438
rect 13261 6336 13295 6370
rect 13261 6268 13295 6302
rect 13261 6200 13295 6234
rect 13261 6132 13295 6166
rect 13261 6064 13295 6098
rect 13261 5996 13295 6030
rect 13261 5928 13295 5962
rect 13261 5860 13295 5894
rect 13483 6812 13517 6846
rect 13483 6744 13517 6778
rect 13483 6676 13517 6710
rect 13483 6608 13517 6642
rect 13483 6540 13517 6574
rect 13483 6472 13517 6506
rect 13483 6404 13517 6438
rect 13483 6336 13517 6370
rect 13483 6268 13517 6302
rect 13483 6200 13517 6234
rect 13483 6132 13517 6166
rect 13483 6064 13517 6098
rect 13483 5996 13517 6030
rect 13483 5928 13517 5962
rect 13483 5860 13517 5894
rect 13569 6812 13603 6846
rect 13569 6744 13603 6778
rect 13569 6676 13603 6710
rect 13569 6608 13603 6642
rect 13569 6540 13603 6574
rect 13569 6472 13603 6506
rect 13569 6404 13603 6438
rect 13569 6336 13603 6370
rect 13569 6268 13603 6302
rect 13569 6200 13603 6234
rect 13569 6132 13603 6166
rect 13569 6064 13603 6098
rect 13569 5996 13603 6030
rect 13569 5928 13603 5962
rect 13569 5860 13603 5894
rect 13655 6812 13689 6846
rect 13655 6744 13689 6778
rect 13655 6676 13689 6710
rect 13655 6608 13689 6642
rect 13655 6540 13689 6574
rect 13655 6472 13689 6506
rect 13655 6404 13689 6438
rect 13655 6336 13689 6370
rect 13655 6268 13689 6302
rect 13655 6200 13689 6234
rect 13655 6132 13689 6166
rect 13655 6064 13689 6098
rect 13655 5996 13689 6030
rect 13655 5928 13689 5962
rect 13655 5860 13689 5894
rect 13741 6812 13775 6846
rect 13741 6744 13775 6778
rect 13741 6676 13775 6710
rect 13741 6608 13775 6642
rect 13741 6540 13775 6574
rect 13741 6472 13775 6506
rect 13741 6404 13775 6438
rect 13741 6336 13775 6370
rect 13741 6268 13775 6302
rect 13741 6200 13775 6234
rect 13741 6132 13775 6166
rect 13741 6064 13775 6098
rect 13741 5996 13775 6030
rect 13741 5928 13775 5962
rect 13741 5860 13775 5894
rect 13827 6812 13861 6846
rect 13827 6744 13861 6778
rect 13827 6676 13861 6710
rect 13827 6608 13861 6642
rect 13827 6540 13861 6574
rect 13827 6472 13861 6506
rect 13827 6404 13861 6438
rect 13827 6336 13861 6370
rect 13827 6268 13861 6302
rect 13827 6200 13861 6234
rect 13827 6132 13861 6166
rect 13827 6064 13861 6098
rect 13827 5996 13861 6030
rect 13827 5928 13861 5962
rect 13827 5860 13861 5894
rect 14049 6812 14083 6846
rect 14049 6744 14083 6778
rect 14049 6676 14083 6710
rect 14049 6608 14083 6642
rect 14049 6540 14083 6574
rect 14049 6472 14083 6506
rect 14049 6404 14083 6438
rect 14049 6336 14083 6370
rect 14049 6268 14083 6302
rect 14049 6200 14083 6234
rect 14049 6132 14083 6166
rect 14049 6064 14083 6098
rect 14049 5996 14083 6030
rect 14049 5928 14083 5962
rect 14049 5860 14083 5894
rect 14135 6812 14169 6846
rect 14135 6744 14169 6778
rect 14135 6676 14169 6710
rect 14135 6608 14169 6642
rect 14135 6540 14169 6574
rect 14135 6472 14169 6506
rect 14135 6404 14169 6438
rect 14135 6336 14169 6370
rect 14135 6268 14169 6302
rect 14135 6200 14169 6234
rect 14135 6132 14169 6166
rect 14135 6064 14169 6098
rect 14135 5996 14169 6030
rect 14135 5928 14169 5962
rect 14135 5860 14169 5894
rect 14221 6812 14255 6846
rect 14221 6744 14255 6778
rect 14221 6676 14255 6710
rect 14221 6608 14255 6642
rect 14221 6540 14255 6574
rect 14221 6472 14255 6506
rect 14221 6404 14255 6438
rect 14221 6336 14255 6370
rect 14221 6268 14255 6302
rect 14221 6200 14255 6234
rect 14221 6132 14255 6166
rect 14221 6064 14255 6098
rect 14221 5996 14255 6030
rect 14221 5928 14255 5962
rect 14221 5860 14255 5894
rect 14307 6812 14341 6846
rect 14307 6744 14341 6778
rect 14307 6676 14341 6710
rect 14307 6608 14341 6642
rect 14307 6540 14341 6574
rect 14307 6472 14341 6506
rect 14307 6404 14341 6438
rect 14307 6336 14341 6370
rect 14307 6268 14341 6302
rect 14307 6200 14341 6234
rect 14307 6132 14341 6166
rect 14307 6064 14341 6098
rect 14307 5996 14341 6030
rect 14307 5928 14341 5962
rect 14307 5860 14341 5894
rect 14393 6812 14427 6846
rect 14393 6744 14427 6778
rect 14393 6676 14427 6710
rect 14393 6608 14427 6642
rect 14393 6540 14427 6574
rect 14393 6472 14427 6506
rect 14393 6404 14427 6438
rect 14393 6336 14427 6370
rect 14393 6268 14427 6302
rect 14393 6200 14427 6234
rect 14393 6132 14427 6166
rect 14393 6064 14427 6098
rect 14393 5996 14427 6030
rect 14393 5928 14427 5962
rect 14393 5860 14427 5894
rect 14615 6812 14649 6846
rect 14615 6744 14649 6778
rect 14615 6676 14649 6710
rect 14615 6608 14649 6642
rect 14615 6540 14649 6574
rect 14615 6472 14649 6506
rect 14615 6404 14649 6438
rect 14615 6336 14649 6370
rect 14615 6268 14649 6302
rect 14615 6200 14649 6234
rect 14615 6132 14649 6166
rect 14615 6064 14649 6098
rect 14615 5996 14649 6030
rect 14615 5928 14649 5962
rect 14615 5860 14649 5894
rect 14701 6812 14735 6846
rect 14701 6744 14735 6778
rect 14701 6676 14735 6710
rect 14701 6608 14735 6642
rect 14701 6540 14735 6574
rect 14701 6472 14735 6506
rect 14701 6404 14735 6438
rect 14701 6336 14735 6370
rect 14701 6268 14735 6302
rect 14701 6200 14735 6234
rect 14701 6132 14735 6166
rect 14701 6064 14735 6098
rect 14701 5996 14735 6030
rect 14701 5928 14735 5962
rect 14701 5860 14735 5894
rect 14787 6812 14821 6846
rect 14787 6744 14821 6778
rect 14787 6676 14821 6710
rect 14787 6608 14821 6642
rect 14787 6540 14821 6574
rect 14787 6472 14821 6506
rect 14787 6404 14821 6438
rect 14787 6336 14821 6370
rect 14787 6268 14821 6302
rect 14787 6200 14821 6234
rect 14787 6132 14821 6166
rect 14787 6064 14821 6098
rect 14787 5996 14821 6030
rect 14787 5928 14821 5962
rect 14787 5860 14821 5894
rect 14873 6812 14907 6846
rect 14873 6744 14907 6778
rect 14873 6676 14907 6710
rect 14873 6608 14907 6642
rect 14873 6540 14907 6574
rect 14873 6472 14907 6506
rect 14873 6404 14907 6438
rect 14873 6336 14907 6370
rect 14873 6268 14907 6302
rect 14873 6200 14907 6234
rect 14873 6132 14907 6166
rect 14873 6064 14907 6098
rect 14873 5996 14907 6030
rect 14873 5928 14907 5962
rect 14873 5860 14907 5894
rect 14959 6812 14993 6846
rect 14959 6744 14993 6778
rect 14959 6676 14993 6710
rect 14959 6608 14993 6642
rect 14959 6540 14993 6574
rect 14959 6472 14993 6506
rect 14959 6404 14993 6438
rect 14959 6336 14993 6370
rect 14959 6268 14993 6302
rect 14959 6200 14993 6234
rect 14959 6132 14993 6166
rect 14959 6064 14993 6098
rect 14959 5996 14993 6030
rect 14959 5928 14993 5962
rect 14959 5860 14993 5894
rect 15181 6812 15215 6846
rect 15181 6744 15215 6778
rect 15181 6676 15215 6710
rect 15181 6608 15215 6642
rect 15181 6540 15215 6574
rect 15181 6472 15215 6506
rect 15181 6404 15215 6438
rect 15181 6336 15215 6370
rect 15181 6268 15215 6302
rect 15181 6200 15215 6234
rect 15181 6132 15215 6166
rect 15181 6064 15215 6098
rect 15181 5996 15215 6030
rect 15181 5928 15215 5962
rect 15181 5860 15215 5894
rect 15267 6812 15301 6846
rect 15267 6744 15301 6778
rect 15267 6676 15301 6710
rect 15267 6608 15301 6642
rect 15267 6540 15301 6574
rect 15267 6472 15301 6506
rect 15267 6404 15301 6438
rect 15267 6336 15301 6370
rect 15267 6268 15301 6302
rect 15267 6200 15301 6234
rect 15267 6132 15301 6166
rect 15267 6064 15301 6098
rect 15267 5996 15301 6030
rect 15267 5928 15301 5962
rect 15267 5860 15301 5894
rect 15353 6812 15387 6846
rect 15353 6744 15387 6778
rect 15353 6676 15387 6710
rect 15353 6608 15387 6642
rect 15353 6540 15387 6574
rect 15353 6472 15387 6506
rect 15353 6404 15387 6438
rect 15353 6336 15387 6370
rect 15353 6268 15387 6302
rect 15353 6200 15387 6234
rect 15353 6132 15387 6166
rect 15353 6064 15387 6098
rect 15353 5996 15387 6030
rect 15353 5928 15387 5962
rect 15353 5860 15387 5894
rect 15439 6812 15473 6846
rect 15439 6744 15473 6778
rect 15439 6676 15473 6710
rect 15439 6608 15473 6642
rect 15439 6540 15473 6574
rect 15439 6472 15473 6506
rect 15439 6404 15473 6438
rect 15439 6336 15473 6370
rect 15439 6268 15473 6302
rect 15439 6200 15473 6234
rect 15439 6132 15473 6166
rect 15439 6064 15473 6098
rect 15439 5996 15473 6030
rect 15439 5928 15473 5962
rect 15439 5860 15473 5894
rect 15525 6812 15559 6846
rect 15525 6744 15559 6778
rect 15525 6676 15559 6710
rect 15525 6608 15559 6642
rect 15525 6540 15559 6574
rect 15525 6472 15559 6506
rect 15525 6404 15559 6438
rect 15525 6336 15559 6370
rect 15525 6268 15559 6302
rect 15525 6200 15559 6234
rect 15525 6132 15559 6166
rect 15525 6064 15559 6098
rect 15525 5996 15559 6030
rect 15525 5928 15559 5962
rect 15525 5860 15559 5894
rect 16118 6145 16152 6179
rect 16118 6077 16152 6111
rect 16118 6009 16152 6043
rect 16118 5941 16152 5975
rect 16118 5873 16152 5907
rect 16118 5805 16152 5839
rect 16118 5737 16152 5771
rect 16118 5669 16152 5703
rect 16118 5601 16152 5635
rect 16118 5533 16152 5567
rect 16118 5465 16152 5499
rect 16118 5397 16152 5431
rect 16118 5329 16152 5363
rect 16118 5261 16152 5295
rect 16118 5193 16152 5227
rect 16204 6145 16238 6179
rect 16204 6077 16238 6111
rect 16204 6009 16238 6043
rect 16204 5941 16238 5975
rect 16204 5873 16238 5907
rect 16204 5805 16238 5839
rect 16204 5737 16238 5771
rect 16204 5669 16238 5703
rect 16204 5601 16238 5635
rect 16204 5533 16238 5567
rect 16204 5465 16238 5499
rect 16204 5397 16238 5431
rect 16204 5329 16238 5363
rect 16204 5261 16238 5295
rect 16204 5193 16238 5227
rect 16290 6145 16324 6179
rect 16290 6077 16324 6111
rect 16290 6009 16324 6043
rect 16290 5941 16324 5975
rect 16290 5873 16324 5907
rect 16290 5805 16324 5839
rect 16290 5737 16324 5771
rect 16290 5669 16324 5703
rect 16290 5601 16324 5635
rect 16290 5533 16324 5567
rect 16290 5465 16324 5499
rect 16290 5397 16324 5431
rect 16290 5329 16324 5363
rect 16290 5261 16324 5295
rect 16290 5193 16324 5227
rect 16376 6145 16410 6179
rect 16376 6077 16410 6111
rect 16376 6009 16410 6043
rect 16376 5941 16410 5975
rect 16376 5873 16410 5907
rect 16376 5805 16410 5839
rect 16376 5737 16410 5771
rect 16376 5669 16410 5703
rect 16376 5601 16410 5635
rect 16376 5533 16410 5567
rect 16376 5465 16410 5499
rect 16376 5397 16410 5431
rect 16376 5329 16410 5363
rect 16376 5261 16410 5295
rect 16376 5193 16410 5227
rect 16462 6145 16496 6179
rect 16462 6077 16496 6111
rect 16462 6009 16496 6043
rect 16462 5941 16496 5975
rect 16462 5873 16496 5907
rect 16462 5805 16496 5839
rect 16462 5737 16496 5771
rect 16462 5669 16496 5703
rect 16462 5601 16496 5635
rect 16462 5533 16496 5567
rect 16462 5465 16496 5499
rect 16462 5397 16496 5431
rect 16462 5329 16496 5363
rect 16462 5261 16496 5295
rect 16462 5193 16496 5227
rect 16548 6145 16582 6179
rect 16548 6077 16582 6111
rect 16548 6009 16582 6043
rect 16548 5941 16582 5975
rect 16548 5873 16582 5907
rect 16548 5805 16582 5839
rect 16548 5737 16582 5771
rect 16548 5669 16582 5703
rect 16548 5601 16582 5635
rect 16548 5533 16582 5567
rect 16548 5465 16582 5499
rect 16548 5397 16582 5431
rect 16548 5329 16582 5363
rect 16548 5261 16582 5295
rect 16548 5193 16582 5227
rect 16634 6145 16668 6179
rect 16634 6077 16668 6111
rect 16634 6009 16668 6043
rect 16634 5941 16668 5975
rect 16634 5873 16668 5907
rect 16634 5805 16668 5839
rect 16634 5737 16668 5771
rect 16634 5669 16668 5703
rect 16634 5601 16668 5635
rect 16634 5533 16668 5567
rect 16634 5465 16668 5499
rect 16634 5397 16668 5431
rect 16634 5329 16668 5363
rect 16634 5261 16668 5295
rect 16634 5193 16668 5227
rect 16720 6145 16754 6179
rect 16720 6077 16754 6111
rect 16720 6009 16754 6043
rect 16720 5941 16754 5975
rect 16720 5873 16754 5907
rect 16720 5805 16754 5839
rect 16720 5737 16754 5771
rect 16720 5669 16754 5703
rect 16720 5601 16754 5635
rect 16720 5533 16754 5567
rect 16720 5465 16754 5499
rect 16720 5397 16754 5431
rect 16720 5329 16754 5363
rect 16720 5261 16754 5295
rect 16720 5193 16754 5227
rect 16806 6145 16840 6179
rect 16806 6077 16840 6111
rect 16806 6009 16840 6043
rect 16806 5941 16840 5975
rect 16806 5873 16840 5907
rect 16806 5805 16840 5839
rect 16806 5737 16840 5771
rect 16806 5669 16840 5703
rect 16806 5601 16840 5635
rect 16806 5533 16840 5567
rect 16806 5465 16840 5499
rect 16806 5397 16840 5431
rect 16806 5329 16840 5363
rect 16806 5261 16840 5295
rect 16806 5193 16840 5227
rect 16892 6145 16926 6179
rect 16892 6077 16926 6111
rect 16892 6009 16926 6043
rect 16892 5941 16926 5975
rect 16892 5873 16926 5907
rect 16892 5805 16926 5839
rect 16892 5737 16926 5771
rect 16892 5669 16926 5703
rect 16892 5601 16926 5635
rect 16892 5533 16926 5567
rect 16892 5465 16926 5499
rect 16892 5397 16926 5431
rect 16892 5329 16926 5363
rect 16892 5261 16926 5295
rect 16892 5193 16926 5227
rect 16978 6145 17012 6179
rect 16978 6077 17012 6111
rect 16978 6009 17012 6043
rect 16978 5941 17012 5975
rect 16978 5873 17012 5907
rect 16978 5805 17012 5839
rect 16978 5737 17012 5771
rect 16978 5669 17012 5703
rect 16978 5601 17012 5635
rect 16978 5533 17012 5567
rect 16978 5465 17012 5499
rect 16978 5397 17012 5431
rect 16978 5329 17012 5363
rect 16978 5261 17012 5295
rect 16978 5193 17012 5227
rect 17064 6145 17098 6179
rect 17064 6077 17098 6111
rect 17064 6009 17098 6043
rect 17064 5941 17098 5975
rect 17064 5873 17098 5907
rect 17064 5805 17098 5839
rect 17064 5737 17098 5771
rect 17064 5669 17098 5703
rect 17064 5601 17098 5635
rect 17064 5533 17098 5567
rect 17064 5465 17098 5499
rect 17064 5397 17098 5431
rect 17064 5329 17098 5363
rect 17064 5261 17098 5295
rect 17064 5193 17098 5227
rect 17150 6145 17184 6179
rect 17150 6077 17184 6111
rect 17150 6009 17184 6043
rect 17150 5941 17184 5975
rect 17150 5873 17184 5907
rect 17150 5805 17184 5839
rect 17150 5737 17184 5771
rect 17150 5669 17184 5703
rect 17150 5601 17184 5635
rect 17150 5533 17184 5567
rect 17150 5465 17184 5499
rect 17150 5397 17184 5431
rect 17150 5329 17184 5363
rect 17150 5261 17184 5295
rect 17150 5193 17184 5227
<< pdiffc >>
rect 17622 7874 17656 7908
rect 17622 7802 17656 7836
rect 17622 7730 17656 7764
rect 17622 7658 17656 7692
rect 17622 7586 17656 7620
rect 17622 7514 17656 7548
rect 17622 7442 17656 7476
rect 17622 7370 17656 7404
rect 17622 7298 17656 7332
rect 17622 7226 17656 7260
rect 17622 7154 17656 7188
rect 17622 7082 17656 7116
rect 17622 7010 17656 7044
rect 17708 7874 17742 7908
rect 17708 7802 17742 7836
rect 17708 7730 17742 7764
rect 17708 7658 17742 7692
rect 17708 7586 17742 7620
rect 17708 7514 17742 7548
rect 17708 7442 17742 7476
rect 17708 7370 17742 7404
rect 17708 7298 17742 7332
rect 17708 7226 17742 7260
rect 17708 7154 17742 7188
rect 17708 7082 17742 7116
rect 17708 7010 17742 7044
rect 17794 7874 17828 7908
rect 17794 7802 17828 7836
rect 17794 7730 17828 7764
rect 17794 7658 17828 7692
rect 17794 7586 17828 7620
rect 17794 7514 17828 7548
rect 17794 7442 17828 7476
rect 17794 7370 17828 7404
rect 17794 7298 17828 7332
rect 17794 7226 17828 7260
rect 17794 7154 17828 7188
rect 17794 7082 17828 7116
rect 17794 7010 17828 7044
rect 17880 7874 17914 7908
rect 17880 7802 17914 7836
rect 17880 7730 17914 7764
rect 17880 7658 17914 7692
rect 17880 7586 17914 7620
rect 17880 7514 17914 7548
rect 17880 7442 17914 7476
rect 17880 7370 17914 7404
rect 17880 7298 17914 7332
rect 17880 7226 17914 7260
rect 17880 7154 17914 7188
rect 17880 7082 17914 7116
rect 17880 7010 17914 7044
rect 17966 7874 18000 7908
rect 17966 7802 18000 7836
rect 17966 7730 18000 7764
rect 17966 7658 18000 7692
rect 17966 7586 18000 7620
rect 17966 7514 18000 7548
rect 17966 7442 18000 7476
rect 17966 7370 18000 7404
rect 17966 7298 18000 7332
rect 17966 7226 18000 7260
rect 17966 7154 18000 7188
rect 17966 7082 18000 7116
rect 17966 7010 18000 7044
rect 18052 7874 18086 7908
rect 18052 7802 18086 7836
rect 18052 7730 18086 7764
rect 18052 7658 18086 7692
rect 18052 7586 18086 7620
rect 18052 7514 18086 7548
rect 18052 7442 18086 7476
rect 18052 7370 18086 7404
rect 18052 7298 18086 7332
rect 18052 7226 18086 7260
rect 18052 7154 18086 7188
rect 18052 7082 18086 7116
rect 18052 7010 18086 7044
rect 18138 7874 18172 7908
rect 18138 7802 18172 7836
rect 18138 7730 18172 7764
rect 18138 7658 18172 7692
rect 18138 7586 18172 7620
rect 18138 7514 18172 7548
rect 18138 7442 18172 7476
rect 18138 7370 18172 7404
rect 18138 7298 18172 7332
rect 18138 7226 18172 7260
rect 18138 7154 18172 7188
rect 18138 7082 18172 7116
rect 18138 7010 18172 7044
rect 18224 7874 18258 7908
rect 18224 7802 18258 7836
rect 18224 7730 18258 7764
rect 18224 7658 18258 7692
rect 18224 7586 18258 7620
rect 18224 7514 18258 7548
rect 18224 7442 18258 7476
rect 18224 7370 18258 7404
rect 18224 7298 18258 7332
rect 18224 7226 18258 7260
rect 18224 7154 18258 7188
rect 18224 7082 18258 7116
rect 18224 7010 18258 7044
rect 18310 7874 18344 7908
rect 18310 7802 18344 7836
rect 18310 7730 18344 7764
rect 18310 7658 18344 7692
rect 18310 7586 18344 7620
rect 18310 7514 18344 7548
rect 18310 7442 18344 7476
rect 18310 7370 18344 7404
rect 18310 7298 18344 7332
rect 18310 7226 18344 7260
rect 18310 7154 18344 7188
rect 18310 7082 18344 7116
rect 18310 7010 18344 7044
rect 18396 7874 18430 7908
rect 18396 7802 18430 7836
rect 18396 7730 18430 7764
rect 18396 7658 18430 7692
rect 18396 7586 18430 7620
rect 18396 7514 18430 7548
rect 18396 7442 18430 7476
rect 18396 7370 18430 7404
rect 18396 7298 18430 7332
rect 18396 7226 18430 7260
rect 18396 7154 18430 7188
rect 18396 7082 18430 7116
rect 18396 7010 18430 7044
rect 18482 7874 18516 7908
rect 18482 7802 18516 7836
rect 18482 7730 18516 7764
rect 18482 7658 18516 7692
rect 18482 7586 18516 7620
rect 18482 7514 18516 7548
rect 18482 7442 18516 7476
rect 18482 7370 18516 7404
rect 18482 7298 18516 7332
rect 18482 7226 18516 7260
rect 18482 7154 18516 7188
rect 18482 7082 18516 7116
rect 18482 7010 18516 7044
rect 18568 7874 18602 7908
rect 18568 7802 18602 7836
rect 18568 7730 18602 7764
rect 18568 7658 18602 7692
rect 18568 7586 18602 7620
rect 18568 7514 18602 7548
rect 18568 7442 18602 7476
rect 18568 7370 18602 7404
rect 18568 7298 18602 7332
rect 18568 7226 18602 7260
rect 18568 7154 18602 7188
rect 18568 7082 18602 7116
rect 18568 7010 18602 7044
rect 18654 7874 18688 7908
rect 18654 7802 18688 7836
rect 18654 7730 18688 7764
rect 18654 7658 18688 7692
rect 18654 7586 18688 7620
rect 18654 7514 18688 7548
rect 18654 7442 18688 7476
rect 18654 7370 18688 7404
rect 18654 7298 18688 7332
rect 18654 7226 18688 7260
rect 18654 7154 18688 7188
rect 18654 7082 18688 7116
rect 18654 7010 18688 7044
rect 18740 7874 18774 7908
rect 18740 7802 18774 7836
rect 18740 7730 18774 7764
rect 18740 7658 18774 7692
rect 18740 7586 18774 7620
rect 18740 7514 18774 7548
rect 18740 7442 18774 7476
rect 18740 7370 18774 7404
rect 18740 7298 18774 7332
rect 18740 7226 18774 7260
rect 18740 7154 18774 7188
rect 18740 7082 18774 7116
rect 18740 7010 18774 7044
rect 18826 7874 18860 7908
rect 18826 7802 18860 7836
rect 18826 7730 18860 7764
rect 18826 7658 18860 7692
rect 18826 7586 18860 7620
rect 18826 7514 18860 7548
rect 18826 7442 18860 7476
rect 18826 7370 18860 7404
rect 18826 7298 18860 7332
rect 18826 7226 18860 7260
rect 18826 7154 18860 7188
rect 18826 7082 18860 7116
rect 18826 7010 18860 7044
rect 18912 7874 18946 7908
rect 18912 7802 18946 7836
rect 18912 7730 18946 7764
rect 18912 7658 18946 7692
rect 18912 7586 18946 7620
rect 18912 7514 18946 7548
rect 18912 7442 18946 7476
rect 18912 7370 18946 7404
rect 18912 7298 18946 7332
rect 18912 7226 18946 7260
rect 18912 7154 18946 7188
rect 18912 7082 18946 7116
rect 18912 7010 18946 7044
rect 18998 7874 19032 7908
rect 18998 7802 19032 7836
rect 18998 7730 19032 7764
rect 18998 7658 19032 7692
rect 18998 7586 19032 7620
rect 18998 7514 19032 7548
rect 18998 7442 19032 7476
rect 18998 7370 19032 7404
rect 18998 7298 19032 7332
rect 18998 7226 19032 7260
rect 18998 7154 19032 7188
rect 18998 7082 19032 7116
rect 18998 7010 19032 7044
rect 19084 7874 19118 7908
rect 19084 7802 19118 7836
rect 19084 7730 19118 7764
rect 19084 7658 19118 7692
rect 19084 7586 19118 7620
rect 19084 7514 19118 7548
rect 19084 7442 19118 7476
rect 19084 7370 19118 7404
rect 19084 7298 19118 7332
rect 19084 7226 19118 7260
rect 19084 7154 19118 7188
rect 19084 7082 19118 7116
rect 19084 7010 19118 7044
rect 19170 7874 19204 7908
rect 19170 7802 19204 7836
rect 19170 7730 19204 7764
rect 19170 7658 19204 7692
rect 19170 7586 19204 7620
rect 19170 7514 19204 7548
rect 19170 7442 19204 7476
rect 19170 7370 19204 7404
rect 19170 7298 19204 7332
rect 19170 7226 19204 7260
rect 19170 7154 19204 7188
rect 19170 7082 19204 7116
rect 19170 7010 19204 7044
rect 19256 7874 19290 7908
rect 19256 7802 19290 7836
rect 19256 7730 19290 7764
rect 19256 7658 19290 7692
rect 19256 7586 19290 7620
rect 19256 7514 19290 7548
rect 19256 7442 19290 7476
rect 19256 7370 19290 7404
rect 19256 7298 19290 7332
rect 19256 7226 19290 7260
rect 19256 7154 19290 7188
rect 19256 7082 19290 7116
rect 19256 7010 19290 7044
rect 19342 7874 19376 7908
rect 19342 7802 19376 7836
rect 19342 7730 19376 7764
rect 19342 7658 19376 7692
rect 19342 7586 19376 7620
rect 19342 7514 19376 7548
rect 19342 7442 19376 7476
rect 19342 7370 19376 7404
rect 19342 7298 19376 7332
rect 19342 7226 19376 7260
rect 19342 7154 19376 7188
rect 19342 7082 19376 7116
rect 19342 7010 19376 7044
rect 19428 7874 19462 7908
rect 19428 7802 19462 7836
rect 19428 7730 19462 7764
rect 19428 7658 19462 7692
rect 19428 7586 19462 7620
rect 19428 7514 19462 7548
rect 19428 7442 19462 7476
rect 19428 7370 19462 7404
rect 19428 7298 19462 7332
rect 19428 7226 19462 7260
rect 19428 7154 19462 7188
rect 19428 7082 19462 7116
rect 19428 7010 19462 7044
rect 19514 7874 19548 7908
rect 19514 7802 19548 7836
rect 19514 7730 19548 7764
rect 19514 7658 19548 7692
rect 19514 7586 19548 7620
rect 19514 7514 19548 7548
rect 19514 7442 19548 7476
rect 19514 7370 19548 7404
rect 19514 7298 19548 7332
rect 19514 7226 19548 7260
rect 19514 7154 19548 7188
rect 19514 7082 19548 7116
rect 19514 7010 19548 7044
rect 19600 7874 19634 7908
rect 19600 7802 19634 7836
rect 19600 7730 19634 7764
rect 19600 7658 19634 7692
rect 19600 7586 19634 7620
rect 19600 7514 19634 7548
rect 19600 7442 19634 7476
rect 19600 7370 19634 7404
rect 19600 7298 19634 7332
rect 19600 7226 19634 7260
rect 19600 7154 19634 7188
rect 19600 7082 19634 7116
rect 19600 7010 19634 7044
rect 19686 7874 19720 7908
rect 19686 7802 19720 7836
rect 19686 7730 19720 7764
rect 19686 7658 19720 7692
rect 19686 7586 19720 7620
rect 19686 7514 19720 7548
rect 19686 7442 19720 7476
rect 19686 7370 19720 7404
rect 19686 7298 19720 7332
rect 19686 7226 19720 7260
rect 19686 7154 19720 7188
rect 19686 7082 19720 7116
rect 19686 7010 19720 7044
rect 19772 7874 19806 7908
rect 19772 7802 19806 7836
rect 19772 7730 19806 7764
rect 19772 7658 19806 7692
rect 19772 7586 19806 7620
rect 19772 7514 19806 7548
rect 19772 7442 19806 7476
rect 19772 7370 19806 7404
rect 19772 7298 19806 7332
rect 19772 7226 19806 7260
rect 19772 7154 19806 7188
rect 19772 7082 19806 7116
rect 19772 7010 19806 7044
rect 19858 7874 19892 7908
rect 19858 7802 19892 7836
rect 19858 7730 19892 7764
rect 19858 7658 19892 7692
rect 19858 7586 19892 7620
rect 19858 7514 19892 7548
rect 19858 7442 19892 7476
rect 19858 7370 19892 7404
rect 19858 7298 19892 7332
rect 19858 7226 19892 7260
rect 19858 7154 19892 7188
rect 19858 7082 19892 7116
rect 19858 7010 19892 7044
rect 19944 7874 19978 7908
rect 19944 7802 19978 7836
rect 19944 7730 19978 7764
rect 19944 7658 19978 7692
rect 19944 7586 19978 7620
rect 19944 7514 19978 7548
rect 19944 7442 19978 7476
rect 19944 7370 19978 7404
rect 19944 7298 19978 7332
rect 19944 7226 19978 7260
rect 19944 7154 19978 7188
rect 19944 7082 19978 7116
rect 19944 7010 19978 7044
rect 20030 7874 20064 7908
rect 20030 7802 20064 7836
rect 20030 7730 20064 7764
rect 20030 7658 20064 7692
rect 20030 7586 20064 7620
rect 20030 7514 20064 7548
rect 20030 7442 20064 7476
rect 20030 7370 20064 7404
rect 20030 7298 20064 7332
rect 20030 7226 20064 7260
rect 20030 7154 20064 7188
rect 20030 7082 20064 7116
rect 20030 7010 20064 7044
rect 17604 6146 17638 6180
rect 17604 6074 17638 6108
rect 17604 6002 17638 6036
rect 17604 5930 17638 5964
rect 17604 5858 17638 5892
rect 17604 5786 17638 5820
rect 17604 5714 17638 5748
rect 17604 5642 17638 5676
rect 17604 5570 17638 5604
rect 17604 5498 17638 5532
rect 17604 5426 17638 5460
rect 17604 5354 17638 5388
rect 17604 5282 17638 5316
rect 17690 6146 17724 6180
rect 17690 6074 17724 6108
rect 17690 6002 17724 6036
rect 17690 5930 17724 5964
rect 17690 5858 17724 5892
rect 17690 5786 17724 5820
rect 17690 5714 17724 5748
rect 17690 5642 17724 5676
rect 17690 5570 17724 5604
rect 17690 5498 17724 5532
rect 17690 5426 17724 5460
rect 17690 5354 17724 5388
rect 17690 5282 17724 5316
rect 17776 6146 17810 6180
rect 17776 6074 17810 6108
rect 17776 6002 17810 6036
rect 17776 5930 17810 5964
rect 17776 5858 17810 5892
rect 17776 5786 17810 5820
rect 17776 5714 17810 5748
rect 17776 5642 17810 5676
rect 17776 5570 17810 5604
rect 17776 5498 17810 5532
rect 17776 5426 17810 5460
rect 17776 5354 17810 5388
rect 17776 5282 17810 5316
rect 17862 6146 17896 6180
rect 17862 6074 17896 6108
rect 17862 6002 17896 6036
rect 17862 5930 17896 5964
rect 17862 5858 17896 5892
rect 17862 5786 17896 5820
rect 17862 5714 17896 5748
rect 17862 5642 17896 5676
rect 17862 5570 17896 5604
rect 17862 5498 17896 5532
rect 17862 5426 17896 5460
rect 17862 5354 17896 5388
rect 17862 5282 17896 5316
rect 17948 6146 17982 6180
rect 17948 6074 17982 6108
rect 17948 6002 17982 6036
rect 17948 5930 17982 5964
rect 17948 5858 17982 5892
rect 17948 5786 17982 5820
rect 17948 5714 17982 5748
rect 17948 5642 17982 5676
rect 17948 5570 17982 5604
rect 17948 5498 17982 5532
rect 17948 5426 17982 5460
rect 17948 5354 17982 5388
rect 17948 5282 17982 5316
rect 18034 6146 18068 6180
rect 18034 6074 18068 6108
rect 18034 6002 18068 6036
rect 18034 5930 18068 5964
rect 18034 5858 18068 5892
rect 18034 5786 18068 5820
rect 18034 5714 18068 5748
rect 18034 5642 18068 5676
rect 18034 5570 18068 5604
rect 18034 5498 18068 5532
rect 18034 5426 18068 5460
rect 18034 5354 18068 5388
rect 18034 5282 18068 5316
rect 18120 6146 18154 6180
rect 18120 6074 18154 6108
rect 18120 6002 18154 6036
rect 18120 5930 18154 5964
rect 18120 5858 18154 5892
rect 18120 5786 18154 5820
rect 18120 5714 18154 5748
rect 18120 5642 18154 5676
rect 18120 5570 18154 5604
rect 18120 5498 18154 5532
rect 18120 5426 18154 5460
rect 18120 5354 18154 5388
rect 18120 5282 18154 5316
rect 18206 6146 18240 6180
rect 18206 6074 18240 6108
rect 18206 6002 18240 6036
rect 18206 5930 18240 5964
rect 18206 5858 18240 5892
rect 18206 5786 18240 5820
rect 18206 5714 18240 5748
rect 18206 5642 18240 5676
rect 18206 5570 18240 5604
rect 18206 5498 18240 5532
rect 18206 5426 18240 5460
rect 18206 5354 18240 5388
rect 18206 5282 18240 5316
rect 18292 6146 18326 6180
rect 18292 6074 18326 6108
rect 18292 6002 18326 6036
rect 18292 5930 18326 5964
rect 18292 5858 18326 5892
rect 18292 5786 18326 5820
rect 18292 5714 18326 5748
rect 18292 5642 18326 5676
rect 18292 5570 18326 5604
rect 18292 5498 18326 5532
rect 18292 5426 18326 5460
rect 18292 5354 18326 5388
rect 18292 5282 18326 5316
rect 18378 6146 18412 6180
rect 18378 6074 18412 6108
rect 18378 6002 18412 6036
rect 18378 5930 18412 5964
rect 18378 5858 18412 5892
rect 18378 5786 18412 5820
rect 18378 5714 18412 5748
rect 18378 5642 18412 5676
rect 18378 5570 18412 5604
rect 18378 5498 18412 5532
rect 18378 5426 18412 5460
rect 18378 5354 18412 5388
rect 18378 5282 18412 5316
rect 18464 6146 18498 6180
rect 18464 6074 18498 6108
rect 18464 6002 18498 6036
rect 18464 5930 18498 5964
rect 18464 5858 18498 5892
rect 18464 5786 18498 5820
rect 18464 5714 18498 5748
rect 18464 5642 18498 5676
rect 18464 5570 18498 5604
rect 18464 5498 18498 5532
rect 18464 5426 18498 5460
rect 18464 5354 18498 5388
rect 18464 5282 18498 5316
rect 18550 6146 18584 6180
rect 18550 6074 18584 6108
rect 18550 6002 18584 6036
rect 18550 5930 18584 5964
rect 18550 5858 18584 5892
rect 18550 5786 18584 5820
rect 18550 5714 18584 5748
rect 18550 5642 18584 5676
rect 18550 5570 18584 5604
rect 18550 5498 18584 5532
rect 18550 5426 18584 5460
rect 18550 5354 18584 5388
rect 18550 5282 18584 5316
rect 18636 6146 18670 6180
rect 18636 6074 18670 6108
rect 18636 6002 18670 6036
rect 18636 5930 18670 5964
rect 18636 5858 18670 5892
rect 18636 5786 18670 5820
rect 18636 5714 18670 5748
rect 18636 5642 18670 5676
rect 18636 5570 18670 5604
rect 18636 5498 18670 5532
rect 18636 5426 18670 5460
rect 18636 5354 18670 5388
rect 18636 5282 18670 5316
rect 18722 6146 18756 6180
rect 18722 6074 18756 6108
rect 18722 6002 18756 6036
rect 18722 5930 18756 5964
rect 18722 5858 18756 5892
rect 18722 5786 18756 5820
rect 18722 5714 18756 5748
rect 18722 5642 18756 5676
rect 18722 5570 18756 5604
rect 18722 5498 18756 5532
rect 18722 5426 18756 5460
rect 18722 5354 18756 5388
rect 18722 5282 18756 5316
rect 18808 6146 18842 6180
rect 18808 6074 18842 6108
rect 18808 6002 18842 6036
rect 18808 5930 18842 5964
rect 18808 5858 18842 5892
rect 18808 5786 18842 5820
rect 18808 5714 18842 5748
rect 18808 5642 18842 5676
rect 18808 5570 18842 5604
rect 18808 5498 18842 5532
rect 18808 5426 18842 5460
rect 18808 5354 18842 5388
rect 18808 5282 18842 5316
rect 18894 6146 18928 6180
rect 18894 6074 18928 6108
rect 18894 6002 18928 6036
rect 18894 5930 18928 5964
rect 18894 5858 18928 5892
rect 18894 5786 18928 5820
rect 18894 5714 18928 5748
rect 18894 5642 18928 5676
rect 18894 5570 18928 5604
rect 18894 5498 18928 5532
rect 18894 5426 18928 5460
rect 18894 5354 18928 5388
rect 18894 5282 18928 5316
rect 18980 6146 19014 6180
rect 18980 6074 19014 6108
rect 18980 6002 19014 6036
rect 18980 5930 19014 5964
rect 18980 5858 19014 5892
rect 18980 5786 19014 5820
rect 18980 5714 19014 5748
rect 18980 5642 19014 5676
rect 18980 5570 19014 5604
rect 18980 5498 19014 5532
rect 18980 5426 19014 5460
rect 18980 5354 19014 5388
rect 18980 5282 19014 5316
rect 19066 6146 19100 6180
rect 19066 6074 19100 6108
rect 19066 6002 19100 6036
rect 19066 5930 19100 5964
rect 19066 5858 19100 5892
rect 19066 5786 19100 5820
rect 19066 5714 19100 5748
rect 19066 5642 19100 5676
rect 19066 5570 19100 5604
rect 19066 5498 19100 5532
rect 19066 5426 19100 5460
rect 19066 5354 19100 5388
rect 19066 5282 19100 5316
rect 19152 6146 19186 6180
rect 19152 6074 19186 6108
rect 19152 6002 19186 6036
rect 19152 5930 19186 5964
rect 19152 5858 19186 5892
rect 19152 5786 19186 5820
rect 19152 5714 19186 5748
rect 19152 5642 19186 5676
rect 19152 5570 19186 5604
rect 19152 5498 19186 5532
rect 19152 5426 19186 5460
rect 19152 5354 19186 5388
rect 19152 5282 19186 5316
rect 19238 6146 19272 6180
rect 19238 6074 19272 6108
rect 19238 6002 19272 6036
rect 19238 5930 19272 5964
rect 19238 5858 19272 5892
rect 19238 5786 19272 5820
rect 19238 5714 19272 5748
rect 19238 5642 19272 5676
rect 19238 5570 19272 5604
rect 19238 5498 19272 5532
rect 19238 5426 19272 5460
rect 19238 5354 19272 5388
rect 19238 5282 19272 5316
rect 19324 6146 19358 6180
rect 19324 6074 19358 6108
rect 19324 6002 19358 6036
rect 19324 5930 19358 5964
rect 19324 5858 19358 5892
rect 19324 5786 19358 5820
rect 19324 5714 19358 5748
rect 19324 5642 19358 5676
rect 19324 5570 19358 5604
rect 19324 5498 19358 5532
rect 19324 5426 19358 5460
rect 19324 5354 19358 5388
rect 19324 5282 19358 5316
rect 19410 6146 19444 6180
rect 19410 6074 19444 6108
rect 19410 6002 19444 6036
rect 19410 5930 19444 5964
rect 19410 5858 19444 5892
rect 19410 5786 19444 5820
rect 19410 5714 19444 5748
rect 19410 5642 19444 5676
rect 19410 5570 19444 5604
rect 19410 5498 19444 5532
rect 19410 5426 19444 5460
rect 19410 5354 19444 5388
rect 19410 5282 19444 5316
rect 19496 6146 19530 6180
rect 19496 6074 19530 6108
rect 19496 6002 19530 6036
rect 19496 5930 19530 5964
rect 19496 5858 19530 5892
rect 19496 5786 19530 5820
rect 19496 5714 19530 5748
rect 19496 5642 19530 5676
rect 19496 5570 19530 5604
rect 19496 5498 19530 5532
rect 19496 5426 19530 5460
rect 19496 5354 19530 5388
rect 19496 5282 19530 5316
rect 19582 6146 19616 6180
rect 19582 6074 19616 6108
rect 19582 6002 19616 6036
rect 19582 5930 19616 5964
rect 19582 5858 19616 5892
rect 19582 5786 19616 5820
rect 19582 5714 19616 5748
rect 19582 5642 19616 5676
rect 19582 5570 19616 5604
rect 19582 5498 19616 5532
rect 19582 5426 19616 5460
rect 19582 5354 19616 5388
rect 19582 5282 19616 5316
rect 19668 6146 19702 6180
rect 19668 6074 19702 6108
rect 19668 6002 19702 6036
rect 19668 5930 19702 5964
rect 19668 5858 19702 5892
rect 19668 5786 19702 5820
rect 19668 5714 19702 5748
rect 19668 5642 19702 5676
rect 19668 5570 19702 5604
rect 19668 5498 19702 5532
rect 19668 5426 19702 5460
rect 19668 5354 19702 5388
rect 19668 5282 19702 5316
rect 19754 6146 19788 6180
rect 19754 6074 19788 6108
rect 19754 6002 19788 6036
rect 19754 5930 19788 5964
rect 19754 5858 19788 5892
rect 19754 5786 19788 5820
rect 19754 5714 19788 5748
rect 19754 5642 19788 5676
rect 19754 5570 19788 5604
rect 19754 5498 19788 5532
rect 19754 5426 19788 5460
rect 19754 5354 19788 5388
rect 19754 5282 19788 5316
rect 19840 6146 19874 6180
rect 19840 6074 19874 6108
rect 19840 6002 19874 6036
rect 19840 5930 19874 5964
rect 19840 5858 19874 5892
rect 19840 5786 19874 5820
rect 19840 5714 19874 5748
rect 19840 5642 19874 5676
rect 19840 5570 19874 5604
rect 19840 5498 19874 5532
rect 19840 5426 19874 5460
rect 19840 5354 19874 5388
rect 19840 5282 19874 5316
rect 19926 6146 19960 6180
rect 19926 6074 19960 6108
rect 19926 6002 19960 6036
rect 19926 5930 19960 5964
rect 19926 5858 19960 5892
rect 19926 5786 19960 5820
rect 19926 5714 19960 5748
rect 19926 5642 19960 5676
rect 19926 5570 19960 5604
rect 19926 5498 19960 5532
rect 19926 5426 19960 5460
rect 19926 5354 19960 5388
rect 19926 5282 19960 5316
rect 20012 6146 20046 6180
rect 20012 6074 20046 6108
rect 20012 6002 20046 6036
rect 20012 5930 20046 5964
rect 20012 5858 20046 5892
rect 20012 5786 20046 5820
rect 20012 5714 20046 5748
rect 20012 5642 20046 5676
rect 20012 5570 20046 5604
rect 20012 5498 20046 5532
rect 20012 5426 20046 5460
rect 20012 5354 20046 5388
rect 20012 5282 20046 5316
<< psubdiff >>
rect 15970 8110 17340 8130
rect 15970 8076 16070 8110
rect 16104 8076 16140 8110
rect 16174 8076 16210 8110
rect 16244 8076 16280 8110
rect 16314 8076 16350 8110
rect 16384 8076 16420 8110
rect 16454 8076 16490 8110
rect 16524 8076 16560 8110
rect 16594 8076 16630 8110
rect 16664 8076 16700 8110
rect 16734 8076 16770 8110
rect 16804 8076 16840 8110
rect 16874 8076 16910 8110
rect 16944 8076 16980 8110
rect 17014 8076 17050 8110
rect 17084 8076 17120 8110
rect 17154 8076 17190 8110
rect 17224 8076 17340 8110
rect 15970 8050 17340 8076
rect 15970 8020 16040 8050
rect 15970 7986 15990 8020
rect 16024 7986 16040 8020
rect 15970 7950 16040 7986
rect 17260 8020 17340 8050
rect 17260 7986 17280 8020
rect 17314 7986 17340 8020
rect 15970 7916 15990 7950
rect 16024 7916 16040 7950
rect 15970 7880 16040 7916
rect 15970 7846 15990 7880
rect 16024 7846 16040 7880
rect 15970 7810 16040 7846
rect 15970 7776 15990 7810
rect 16024 7776 16040 7810
rect 15970 7740 16040 7776
rect 15970 7706 15990 7740
rect 16024 7706 16040 7740
rect 15970 7670 16040 7706
rect 15970 7636 15990 7670
rect 16024 7636 16040 7670
rect 15970 7600 16040 7636
rect 15970 7566 15990 7600
rect 16024 7566 16040 7600
rect 15970 7530 16040 7566
rect 15970 7496 15990 7530
rect 16024 7496 16040 7530
rect 15970 7460 16040 7496
rect 15970 7426 15990 7460
rect 16024 7426 16040 7460
rect 15970 7390 16040 7426
rect 15970 7356 15990 7390
rect 16024 7356 16040 7390
rect 15970 7320 16040 7356
rect 15970 7286 15990 7320
rect 16024 7286 16040 7320
rect 15970 7250 16040 7286
rect 15970 7216 15990 7250
rect 16024 7216 16040 7250
rect 15970 7180 16040 7216
rect 15970 7146 15990 7180
rect 16024 7146 16040 7180
rect 15970 7110 16040 7146
rect 15970 7076 15990 7110
rect 16024 7076 16040 7110
rect 15970 7040 16040 7076
rect 15970 7006 15990 7040
rect 16024 7006 16040 7040
rect 15970 6970 16040 7006
rect 17260 7950 17340 7986
rect 17260 7916 17280 7950
rect 17314 7916 17340 7950
rect 17260 7880 17340 7916
rect 17260 7846 17280 7880
rect 17314 7846 17340 7880
rect 17260 7810 17340 7846
rect 17260 7776 17280 7810
rect 17314 7776 17340 7810
rect 17260 7740 17340 7776
rect 17260 7706 17280 7740
rect 17314 7706 17340 7740
rect 17260 7670 17340 7706
rect 17260 7636 17280 7670
rect 17314 7636 17340 7670
rect 17260 7600 17340 7636
rect 17260 7566 17280 7600
rect 17314 7566 17340 7600
rect 17260 7530 17340 7566
rect 17260 7496 17280 7530
rect 17314 7496 17340 7530
rect 17260 7460 17340 7496
rect 17260 7426 17280 7460
rect 17314 7426 17340 7460
rect 17260 7390 17340 7426
rect 17260 7356 17280 7390
rect 17314 7356 17340 7390
rect 17260 7320 17340 7356
rect 17260 7286 17280 7320
rect 17314 7286 17340 7320
rect 17260 7250 17340 7286
rect 17260 7216 17280 7250
rect 17314 7216 17340 7250
rect 17260 7180 17340 7216
rect 17260 7146 17280 7180
rect 17314 7146 17340 7180
rect 17260 7110 17340 7146
rect 17260 7076 17280 7110
rect 17314 7076 17340 7110
rect 17260 7040 17340 7076
rect 17260 7006 17280 7040
rect 17314 7006 17340 7040
rect 17260 6970 17340 7006
rect 11662 6812 11720 6858
rect 11662 6778 11674 6812
rect 11708 6778 11720 6812
rect 11662 6744 11720 6778
rect 11662 6710 11674 6744
rect 11708 6710 11720 6744
rect 11662 6676 11720 6710
rect 11662 6642 11674 6676
rect 11708 6642 11720 6676
rect 11662 6608 11720 6642
rect 11662 6574 11674 6608
rect 11708 6574 11720 6608
rect 11662 6540 11720 6574
rect 11662 6506 11674 6540
rect 11708 6506 11720 6540
rect 11662 6472 11720 6506
rect 11662 6438 11674 6472
rect 11708 6438 11720 6472
rect 11662 6404 11720 6438
rect 11662 6370 11674 6404
rect 11708 6370 11720 6404
rect 11662 6336 11720 6370
rect 11662 6302 11674 6336
rect 11708 6302 11720 6336
rect 11662 6268 11720 6302
rect 11662 6234 11674 6268
rect 11708 6234 11720 6268
rect 11662 6200 11720 6234
rect 11662 6166 11674 6200
rect 11708 6166 11720 6200
rect 11662 6132 11720 6166
rect 11662 6098 11674 6132
rect 11708 6098 11720 6132
rect 11662 6064 11720 6098
rect 11662 6030 11674 6064
rect 11708 6030 11720 6064
rect 11662 5996 11720 6030
rect 11662 5962 11674 5996
rect 11708 5962 11720 5996
rect 11662 5928 11720 5962
rect 11662 5894 11674 5928
rect 11708 5894 11720 5928
rect 11662 5848 11720 5894
rect 12228 6812 12286 6858
rect 12228 6778 12240 6812
rect 12274 6778 12286 6812
rect 12228 6744 12286 6778
rect 12228 6710 12240 6744
rect 12274 6710 12286 6744
rect 12228 6676 12286 6710
rect 12228 6642 12240 6676
rect 12274 6642 12286 6676
rect 12228 6608 12286 6642
rect 12228 6574 12240 6608
rect 12274 6574 12286 6608
rect 12228 6540 12286 6574
rect 12228 6506 12240 6540
rect 12274 6506 12286 6540
rect 12228 6472 12286 6506
rect 12228 6438 12240 6472
rect 12274 6438 12286 6472
rect 12228 6404 12286 6438
rect 12228 6370 12240 6404
rect 12274 6370 12286 6404
rect 12228 6336 12286 6370
rect 12228 6302 12240 6336
rect 12274 6302 12286 6336
rect 12228 6268 12286 6302
rect 12228 6234 12240 6268
rect 12274 6234 12286 6268
rect 12228 6200 12286 6234
rect 12228 6166 12240 6200
rect 12274 6166 12286 6200
rect 12228 6132 12286 6166
rect 12228 6098 12240 6132
rect 12274 6098 12286 6132
rect 12228 6064 12286 6098
rect 12228 6030 12240 6064
rect 12274 6030 12286 6064
rect 12228 5996 12286 6030
rect 12228 5962 12240 5996
rect 12274 5962 12286 5996
rect 12228 5928 12286 5962
rect 12228 5894 12240 5928
rect 12274 5894 12286 5928
rect 12228 5848 12286 5894
rect 12794 6812 12852 6858
rect 12794 6778 12806 6812
rect 12840 6778 12852 6812
rect 12794 6744 12852 6778
rect 12794 6710 12806 6744
rect 12840 6710 12852 6744
rect 12794 6676 12852 6710
rect 12794 6642 12806 6676
rect 12840 6642 12852 6676
rect 12794 6608 12852 6642
rect 12794 6574 12806 6608
rect 12840 6574 12852 6608
rect 12794 6540 12852 6574
rect 12794 6506 12806 6540
rect 12840 6506 12852 6540
rect 12794 6472 12852 6506
rect 12794 6438 12806 6472
rect 12840 6438 12852 6472
rect 12794 6404 12852 6438
rect 12794 6370 12806 6404
rect 12840 6370 12852 6404
rect 12794 6336 12852 6370
rect 12794 6302 12806 6336
rect 12840 6302 12852 6336
rect 12794 6268 12852 6302
rect 12794 6234 12806 6268
rect 12840 6234 12852 6268
rect 12794 6200 12852 6234
rect 12794 6166 12806 6200
rect 12840 6166 12852 6200
rect 12794 6132 12852 6166
rect 12794 6098 12806 6132
rect 12840 6098 12852 6132
rect 12794 6064 12852 6098
rect 12794 6030 12806 6064
rect 12840 6030 12852 6064
rect 12794 5996 12852 6030
rect 12794 5962 12806 5996
rect 12840 5962 12852 5996
rect 12794 5928 12852 5962
rect 12794 5894 12806 5928
rect 12840 5894 12852 5928
rect 12794 5848 12852 5894
rect 13360 6812 13418 6858
rect 13360 6778 13372 6812
rect 13406 6778 13418 6812
rect 13360 6744 13418 6778
rect 13360 6710 13372 6744
rect 13406 6710 13418 6744
rect 13360 6676 13418 6710
rect 13360 6642 13372 6676
rect 13406 6642 13418 6676
rect 13360 6608 13418 6642
rect 13360 6574 13372 6608
rect 13406 6574 13418 6608
rect 13360 6540 13418 6574
rect 13360 6506 13372 6540
rect 13406 6506 13418 6540
rect 13360 6472 13418 6506
rect 13360 6438 13372 6472
rect 13406 6438 13418 6472
rect 13360 6404 13418 6438
rect 13360 6370 13372 6404
rect 13406 6370 13418 6404
rect 13360 6336 13418 6370
rect 13360 6302 13372 6336
rect 13406 6302 13418 6336
rect 13360 6268 13418 6302
rect 13360 6234 13372 6268
rect 13406 6234 13418 6268
rect 13360 6200 13418 6234
rect 13360 6166 13372 6200
rect 13406 6166 13418 6200
rect 13360 6132 13418 6166
rect 13360 6098 13372 6132
rect 13406 6098 13418 6132
rect 13360 6064 13418 6098
rect 13360 6030 13372 6064
rect 13406 6030 13418 6064
rect 13360 5996 13418 6030
rect 13360 5962 13372 5996
rect 13406 5962 13418 5996
rect 13360 5928 13418 5962
rect 13360 5894 13372 5928
rect 13406 5894 13418 5928
rect 13360 5848 13418 5894
rect 13926 6812 13984 6858
rect 13926 6778 13938 6812
rect 13972 6778 13984 6812
rect 13926 6744 13984 6778
rect 13926 6710 13938 6744
rect 13972 6710 13984 6744
rect 13926 6676 13984 6710
rect 13926 6642 13938 6676
rect 13972 6642 13984 6676
rect 13926 6608 13984 6642
rect 13926 6574 13938 6608
rect 13972 6574 13984 6608
rect 13926 6540 13984 6574
rect 13926 6506 13938 6540
rect 13972 6506 13984 6540
rect 13926 6472 13984 6506
rect 13926 6438 13938 6472
rect 13972 6438 13984 6472
rect 13926 6404 13984 6438
rect 13926 6370 13938 6404
rect 13972 6370 13984 6404
rect 13926 6336 13984 6370
rect 13926 6302 13938 6336
rect 13972 6302 13984 6336
rect 13926 6268 13984 6302
rect 13926 6234 13938 6268
rect 13972 6234 13984 6268
rect 13926 6200 13984 6234
rect 13926 6166 13938 6200
rect 13972 6166 13984 6200
rect 13926 6132 13984 6166
rect 13926 6098 13938 6132
rect 13972 6098 13984 6132
rect 13926 6064 13984 6098
rect 13926 6030 13938 6064
rect 13972 6030 13984 6064
rect 13926 5996 13984 6030
rect 13926 5962 13938 5996
rect 13972 5962 13984 5996
rect 13926 5928 13984 5962
rect 13926 5894 13938 5928
rect 13972 5894 13984 5928
rect 13926 5848 13984 5894
rect 14492 6812 14550 6858
rect 14492 6778 14504 6812
rect 14538 6778 14550 6812
rect 14492 6744 14550 6778
rect 14492 6710 14504 6744
rect 14538 6710 14550 6744
rect 14492 6676 14550 6710
rect 14492 6642 14504 6676
rect 14538 6642 14550 6676
rect 14492 6608 14550 6642
rect 14492 6574 14504 6608
rect 14538 6574 14550 6608
rect 14492 6540 14550 6574
rect 14492 6506 14504 6540
rect 14538 6506 14550 6540
rect 14492 6472 14550 6506
rect 14492 6438 14504 6472
rect 14538 6438 14550 6472
rect 14492 6404 14550 6438
rect 14492 6370 14504 6404
rect 14538 6370 14550 6404
rect 14492 6336 14550 6370
rect 14492 6302 14504 6336
rect 14538 6302 14550 6336
rect 14492 6268 14550 6302
rect 14492 6234 14504 6268
rect 14538 6234 14550 6268
rect 14492 6200 14550 6234
rect 14492 6166 14504 6200
rect 14538 6166 14550 6200
rect 14492 6132 14550 6166
rect 14492 6098 14504 6132
rect 14538 6098 14550 6132
rect 14492 6064 14550 6098
rect 14492 6030 14504 6064
rect 14538 6030 14550 6064
rect 14492 5996 14550 6030
rect 14492 5962 14504 5996
rect 14538 5962 14550 5996
rect 14492 5928 14550 5962
rect 14492 5894 14504 5928
rect 14538 5894 14550 5928
rect 14492 5848 14550 5894
rect 15058 6812 15116 6858
rect 15058 6778 15070 6812
rect 15104 6778 15116 6812
rect 15058 6744 15116 6778
rect 15058 6710 15070 6744
rect 15104 6710 15116 6744
rect 15058 6676 15116 6710
rect 15058 6642 15070 6676
rect 15104 6642 15116 6676
rect 15058 6608 15116 6642
rect 15058 6574 15070 6608
rect 15104 6574 15116 6608
rect 15058 6540 15116 6574
rect 15058 6506 15070 6540
rect 15104 6506 15116 6540
rect 15058 6472 15116 6506
rect 15058 6438 15070 6472
rect 15104 6438 15116 6472
rect 15058 6404 15116 6438
rect 15058 6370 15070 6404
rect 15104 6370 15116 6404
rect 15058 6336 15116 6370
rect 15058 6302 15070 6336
rect 15104 6302 15116 6336
rect 15058 6268 15116 6302
rect 15058 6234 15070 6268
rect 15104 6234 15116 6268
rect 15058 6200 15116 6234
rect 15058 6166 15070 6200
rect 15104 6166 15116 6200
rect 15058 6132 15116 6166
rect 15058 6098 15070 6132
rect 15104 6098 15116 6132
rect 15058 6064 15116 6098
rect 15058 6030 15070 6064
rect 15104 6030 15116 6064
rect 15058 5996 15116 6030
rect 15058 5962 15070 5996
rect 15104 5962 15116 5996
rect 15058 5928 15116 5962
rect 15058 5894 15070 5928
rect 15104 5894 15116 5928
rect 15058 5848 15116 5894
rect 15624 6812 15682 6858
rect 15624 6778 15636 6812
rect 15670 6778 15682 6812
rect 15624 6744 15682 6778
rect 15624 6710 15636 6744
rect 15670 6710 15682 6744
rect 15624 6676 15682 6710
rect 15624 6642 15636 6676
rect 15670 6642 15682 6676
rect 15624 6608 15682 6642
rect 15624 6574 15636 6608
rect 15670 6574 15682 6608
rect 15624 6540 15682 6574
rect 15624 6506 15636 6540
rect 15670 6506 15682 6540
rect 15624 6472 15682 6506
rect 15624 6438 15636 6472
rect 15670 6438 15682 6472
rect 15624 6404 15682 6438
rect 15624 6370 15636 6404
rect 15670 6370 15682 6404
rect 15624 6336 15682 6370
rect 15624 6302 15636 6336
rect 15670 6302 15682 6336
rect 15624 6268 15682 6302
rect 15624 6234 15636 6268
rect 15670 6234 15682 6268
rect 15624 6200 15682 6234
rect 15624 6166 15636 6200
rect 15670 6166 15682 6200
rect 15624 6132 15682 6166
rect 15624 6098 15636 6132
rect 15670 6098 15682 6132
rect 15624 6064 15682 6098
rect 15624 6030 15636 6064
rect 15670 6030 15682 6064
rect 15624 5996 15682 6030
rect 15624 5962 15636 5996
rect 15670 5962 15682 5996
rect 15624 5928 15682 5962
rect 15624 5894 15636 5928
rect 15670 5894 15682 5928
rect 15624 5848 15682 5894
rect 15970 6154 16040 6190
rect 15970 6120 15990 6154
rect 16024 6120 16040 6154
rect 15970 6084 16040 6120
rect 15970 6050 15990 6084
rect 16024 6050 16040 6084
rect 15970 6014 16040 6050
rect 15970 5980 15990 6014
rect 16024 5980 16040 6014
rect 15970 5944 16040 5980
rect 15970 5910 15990 5944
rect 16024 5910 16040 5944
rect 15970 5874 16040 5910
rect 15970 5840 15990 5874
rect 16024 5840 16040 5874
rect 15970 5804 16040 5840
rect 15970 5770 15990 5804
rect 16024 5770 16040 5804
rect 15970 5734 16040 5770
rect 15970 5700 15990 5734
rect 16024 5700 16040 5734
rect 15970 5664 16040 5700
rect 15970 5630 15990 5664
rect 16024 5630 16040 5664
rect 15970 5594 16040 5630
rect 15970 5560 15990 5594
rect 16024 5560 16040 5594
rect 15970 5524 16040 5560
rect 15970 5490 15990 5524
rect 16024 5490 16040 5524
rect 15970 5454 16040 5490
rect 15970 5420 15990 5454
rect 16024 5420 16040 5454
rect 15970 5384 16040 5420
rect 15970 5350 15990 5384
rect 16024 5350 16040 5384
rect 15970 5314 16040 5350
rect 15970 5280 15990 5314
rect 16024 5280 16040 5314
rect 15970 5244 16040 5280
rect 15970 5210 15990 5244
rect 16024 5210 16040 5244
rect 15970 5174 16040 5210
rect 17260 6154 17340 6190
rect 17260 6120 17280 6154
rect 17314 6120 17340 6154
rect 17260 6084 17340 6120
rect 17260 6050 17280 6084
rect 17314 6050 17340 6084
rect 17260 6014 17340 6050
rect 17260 5980 17280 6014
rect 17314 5980 17340 6014
rect 17260 5944 17340 5980
rect 17260 5910 17280 5944
rect 17314 5910 17340 5944
rect 17260 5874 17340 5910
rect 17260 5840 17280 5874
rect 17314 5840 17340 5874
rect 17260 5804 17340 5840
rect 17260 5770 17280 5804
rect 17314 5770 17340 5804
rect 17260 5734 17340 5770
rect 17260 5700 17280 5734
rect 17314 5700 17340 5734
rect 17260 5664 17340 5700
rect 17260 5630 17280 5664
rect 17314 5630 17340 5664
rect 17260 5594 17340 5630
rect 17260 5560 17280 5594
rect 17314 5560 17340 5594
rect 17260 5524 17340 5560
rect 17260 5490 17280 5524
rect 17314 5490 17340 5524
rect 17260 5454 17340 5490
rect 17260 5420 17280 5454
rect 17314 5420 17340 5454
rect 17260 5384 17340 5420
rect 17260 5350 17280 5384
rect 17314 5350 17340 5384
rect 17260 5314 17340 5350
rect 17260 5280 17280 5314
rect 17314 5280 17340 5314
rect 17260 5244 17340 5280
rect 17260 5210 17280 5244
rect 17314 5210 17340 5244
rect 15970 5140 15990 5174
rect 16024 5140 16040 5174
rect 15970 5110 16040 5140
rect 17260 5174 17340 5210
rect 17260 5140 17280 5174
rect 17314 5140 17340 5174
rect 17260 5110 17340 5140
rect 15970 5084 17340 5110
rect 15970 5050 16070 5084
rect 16104 5050 16140 5084
rect 16174 5050 16210 5084
rect 16244 5050 16280 5084
rect 16314 5050 16350 5084
rect 16384 5050 16420 5084
rect 16454 5050 16490 5084
rect 16524 5050 16560 5084
rect 16594 5050 16630 5084
rect 16664 5050 16700 5084
rect 16734 5050 16770 5084
rect 16804 5050 16840 5084
rect 16874 5050 16910 5084
rect 16944 5050 16980 5084
rect 17014 5050 17050 5084
rect 17084 5050 17120 5084
rect 17154 5050 17190 5084
rect 17224 5050 17340 5084
rect 15970 5030 17340 5050
<< nsubdiff >>
rect 17478 8090 20218 8110
rect 17478 8050 17678 8090
rect 17718 8050 17758 8090
rect 17798 8050 17838 8090
rect 17878 8050 17918 8090
rect 17958 8050 17998 8090
rect 18038 8050 18078 8090
rect 18118 8050 18158 8090
rect 18198 8050 18238 8090
rect 18278 8050 18318 8090
rect 18358 8050 18398 8090
rect 18438 8050 18478 8090
rect 18518 8050 18558 8090
rect 18598 8050 18638 8090
rect 18678 8050 18718 8090
rect 18758 8050 18798 8090
rect 18838 8050 18878 8090
rect 18918 8050 18958 8090
rect 18998 8050 19038 8090
rect 19078 8050 19118 8090
rect 19158 8050 19198 8090
rect 19238 8050 19278 8090
rect 19318 8050 19358 8090
rect 19398 8050 19438 8090
rect 19478 8050 19518 8090
rect 19558 8050 19598 8090
rect 19638 8050 19678 8090
rect 19718 8050 19758 8090
rect 19798 8050 19838 8090
rect 19878 8050 19918 8090
rect 19958 8050 19998 8090
rect 20038 8050 20218 8090
rect 17478 8030 20218 8050
rect 17478 7930 17558 8030
rect 17478 7890 17498 7930
rect 17538 7890 17558 7930
rect 17478 7850 17558 7890
rect 17478 7810 17498 7850
rect 17538 7810 17558 7850
rect 17478 7770 17558 7810
rect 17478 7730 17498 7770
rect 17538 7730 17558 7770
rect 17478 7690 17558 7730
rect 17478 7650 17498 7690
rect 17538 7650 17558 7690
rect 17478 7610 17558 7650
rect 17478 7570 17498 7610
rect 17538 7570 17558 7610
rect 17478 7530 17558 7570
rect 17478 7490 17498 7530
rect 17538 7490 17558 7530
rect 17478 7450 17558 7490
rect 17478 7410 17498 7450
rect 17538 7410 17558 7450
rect 17478 7370 17558 7410
rect 17478 7330 17498 7370
rect 17538 7330 17558 7370
rect 17478 7290 17558 7330
rect 17478 7250 17498 7290
rect 17538 7250 17558 7290
rect 17478 7210 17558 7250
rect 17478 7170 17498 7210
rect 17538 7170 17558 7210
rect 17478 7130 17558 7170
rect 17478 7090 17498 7130
rect 17538 7090 17558 7130
rect 17478 7050 17558 7090
rect 17478 7010 17498 7050
rect 17538 7010 17558 7050
rect 17478 6970 17558 7010
rect 20138 7930 20218 8030
rect 20138 7890 20158 7930
rect 20198 7890 20218 7930
rect 20138 7850 20218 7890
rect 20138 7810 20158 7850
rect 20198 7810 20218 7850
rect 20138 7770 20218 7810
rect 20138 7730 20158 7770
rect 20198 7730 20218 7770
rect 20138 7690 20218 7730
rect 20138 7650 20158 7690
rect 20198 7650 20218 7690
rect 20138 7610 20218 7650
rect 20138 7570 20158 7610
rect 20198 7570 20218 7610
rect 20138 7530 20218 7570
rect 20138 7490 20158 7530
rect 20198 7490 20218 7530
rect 20138 7450 20218 7490
rect 20138 7410 20158 7450
rect 20198 7410 20218 7450
rect 20138 7370 20218 7410
rect 20138 7330 20158 7370
rect 20198 7330 20218 7370
rect 20138 7290 20218 7330
rect 20138 7250 20158 7290
rect 20198 7250 20218 7290
rect 20138 7210 20218 7250
rect 20138 7170 20158 7210
rect 20198 7170 20218 7210
rect 20138 7130 20218 7170
rect 20138 7090 20158 7130
rect 20198 7090 20218 7130
rect 20138 7050 20218 7090
rect 20138 7010 20158 7050
rect 20198 7010 20218 7050
rect 20138 6970 20218 7010
rect 17460 6180 17540 6220
rect 17460 6140 17480 6180
rect 17520 6140 17540 6180
rect 17460 6100 17540 6140
rect 17460 6060 17480 6100
rect 17520 6060 17540 6100
rect 17460 6020 17540 6060
rect 17460 5980 17480 6020
rect 17520 5980 17540 6020
rect 17460 5940 17540 5980
rect 17460 5900 17480 5940
rect 17520 5900 17540 5940
rect 17460 5860 17540 5900
rect 17460 5820 17480 5860
rect 17520 5820 17540 5860
rect 17460 5780 17540 5820
rect 17460 5740 17480 5780
rect 17520 5740 17540 5780
rect 17460 5700 17540 5740
rect 17460 5660 17480 5700
rect 17520 5660 17540 5700
rect 17460 5620 17540 5660
rect 17460 5580 17480 5620
rect 17520 5580 17540 5620
rect 17460 5540 17540 5580
rect 17460 5500 17480 5540
rect 17520 5500 17540 5540
rect 17460 5460 17540 5500
rect 17460 5420 17480 5460
rect 17520 5420 17540 5460
rect 17460 5380 17540 5420
rect 17460 5340 17480 5380
rect 17520 5340 17540 5380
rect 17460 5300 17540 5340
rect 17460 5260 17480 5300
rect 17520 5260 17540 5300
rect 17460 5160 17540 5260
rect 20120 6180 20200 6220
rect 20120 6140 20140 6180
rect 20180 6140 20200 6180
rect 20120 6100 20200 6140
rect 20120 6060 20140 6100
rect 20180 6060 20200 6100
rect 20120 6020 20200 6060
rect 20120 5980 20140 6020
rect 20180 5980 20200 6020
rect 20120 5940 20200 5980
rect 20120 5900 20140 5940
rect 20180 5900 20200 5940
rect 20120 5860 20200 5900
rect 20120 5820 20140 5860
rect 20180 5820 20200 5860
rect 20120 5780 20200 5820
rect 20120 5740 20140 5780
rect 20180 5740 20200 5780
rect 20120 5700 20200 5740
rect 20120 5660 20140 5700
rect 20180 5660 20200 5700
rect 20120 5620 20200 5660
rect 20120 5580 20140 5620
rect 20180 5580 20200 5620
rect 20120 5540 20200 5580
rect 20120 5500 20140 5540
rect 20180 5500 20200 5540
rect 20120 5460 20200 5500
rect 20120 5420 20140 5460
rect 20180 5420 20200 5460
rect 20120 5380 20200 5420
rect 20120 5340 20140 5380
rect 20180 5340 20200 5380
rect 20120 5300 20200 5340
rect 20120 5260 20140 5300
rect 20180 5260 20200 5300
rect 20120 5160 20200 5260
rect 17460 5140 20200 5160
rect 17460 5100 17660 5140
rect 17700 5100 17740 5140
rect 17780 5100 17820 5140
rect 17860 5100 17900 5140
rect 17940 5100 17980 5140
rect 18020 5100 18060 5140
rect 18100 5100 18140 5140
rect 18180 5100 18220 5140
rect 18260 5100 18300 5140
rect 18340 5100 18380 5140
rect 18420 5100 18460 5140
rect 18500 5100 18540 5140
rect 18580 5100 18620 5140
rect 18660 5100 18700 5140
rect 18740 5100 18780 5140
rect 18820 5100 18860 5140
rect 18900 5100 18940 5140
rect 18980 5100 19020 5140
rect 19060 5100 19100 5140
rect 19140 5100 19180 5140
rect 19220 5100 19260 5140
rect 19300 5100 19340 5140
rect 19380 5100 19420 5140
rect 19460 5100 19500 5140
rect 19540 5100 19580 5140
rect 19620 5100 19660 5140
rect 19700 5100 19740 5140
rect 19780 5100 19820 5140
rect 19860 5100 19900 5140
rect 19940 5100 19980 5140
rect 20020 5100 20200 5140
rect 17460 5080 20200 5100
<< psubdiffcont >>
rect 16070 8076 16104 8110
rect 16140 8076 16174 8110
rect 16210 8076 16244 8110
rect 16280 8076 16314 8110
rect 16350 8076 16384 8110
rect 16420 8076 16454 8110
rect 16490 8076 16524 8110
rect 16560 8076 16594 8110
rect 16630 8076 16664 8110
rect 16700 8076 16734 8110
rect 16770 8076 16804 8110
rect 16840 8076 16874 8110
rect 16910 8076 16944 8110
rect 16980 8076 17014 8110
rect 17050 8076 17084 8110
rect 17120 8076 17154 8110
rect 17190 8076 17224 8110
rect 15990 7986 16024 8020
rect 17280 7986 17314 8020
rect 15990 7916 16024 7950
rect 15990 7846 16024 7880
rect 15990 7776 16024 7810
rect 15990 7706 16024 7740
rect 15990 7636 16024 7670
rect 15990 7566 16024 7600
rect 15990 7496 16024 7530
rect 15990 7426 16024 7460
rect 15990 7356 16024 7390
rect 15990 7286 16024 7320
rect 15990 7216 16024 7250
rect 15990 7146 16024 7180
rect 15990 7076 16024 7110
rect 15990 7006 16024 7040
rect 17280 7916 17314 7950
rect 17280 7846 17314 7880
rect 17280 7776 17314 7810
rect 17280 7706 17314 7740
rect 17280 7636 17314 7670
rect 17280 7566 17314 7600
rect 17280 7496 17314 7530
rect 17280 7426 17314 7460
rect 17280 7356 17314 7390
rect 17280 7286 17314 7320
rect 17280 7216 17314 7250
rect 17280 7146 17314 7180
rect 17280 7076 17314 7110
rect 17280 7006 17314 7040
rect 11674 6778 11708 6812
rect 11674 6710 11708 6744
rect 11674 6642 11708 6676
rect 11674 6574 11708 6608
rect 11674 6506 11708 6540
rect 11674 6438 11708 6472
rect 11674 6370 11708 6404
rect 11674 6302 11708 6336
rect 11674 6234 11708 6268
rect 11674 6166 11708 6200
rect 11674 6098 11708 6132
rect 11674 6030 11708 6064
rect 11674 5962 11708 5996
rect 11674 5894 11708 5928
rect 12240 6778 12274 6812
rect 12240 6710 12274 6744
rect 12240 6642 12274 6676
rect 12240 6574 12274 6608
rect 12240 6506 12274 6540
rect 12240 6438 12274 6472
rect 12240 6370 12274 6404
rect 12240 6302 12274 6336
rect 12240 6234 12274 6268
rect 12240 6166 12274 6200
rect 12240 6098 12274 6132
rect 12240 6030 12274 6064
rect 12240 5962 12274 5996
rect 12240 5894 12274 5928
rect 12806 6778 12840 6812
rect 12806 6710 12840 6744
rect 12806 6642 12840 6676
rect 12806 6574 12840 6608
rect 12806 6506 12840 6540
rect 12806 6438 12840 6472
rect 12806 6370 12840 6404
rect 12806 6302 12840 6336
rect 12806 6234 12840 6268
rect 12806 6166 12840 6200
rect 12806 6098 12840 6132
rect 12806 6030 12840 6064
rect 12806 5962 12840 5996
rect 12806 5894 12840 5928
rect 13372 6778 13406 6812
rect 13372 6710 13406 6744
rect 13372 6642 13406 6676
rect 13372 6574 13406 6608
rect 13372 6506 13406 6540
rect 13372 6438 13406 6472
rect 13372 6370 13406 6404
rect 13372 6302 13406 6336
rect 13372 6234 13406 6268
rect 13372 6166 13406 6200
rect 13372 6098 13406 6132
rect 13372 6030 13406 6064
rect 13372 5962 13406 5996
rect 13372 5894 13406 5928
rect 13938 6778 13972 6812
rect 13938 6710 13972 6744
rect 13938 6642 13972 6676
rect 13938 6574 13972 6608
rect 13938 6506 13972 6540
rect 13938 6438 13972 6472
rect 13938 6370 13972 6404
rect 13938 6302 13972 6336
rect 13938 6234 13972 6268
rect 13938 6166 13972 6200
rect 13938 6098 13972 6132
rect 13938 6030 13972 6064
rect 13938 5962 13972 5996
rect 13938 5894 13972 5928
rect 14504 6778 14538 6812
rect 14504 6710 14538 6744
rect 14504 6642 14538 6676
rect 14504 6574 14538 6608
rect 14504 6506 14538 6540
rect 14504 6438 14538 6472
rect 14504 6370 14538 6404
rect 14504 6302 14538 6336
rect 14504 6234 14538 6268
rect 14504 6166 14538 6200
rect 14504 6098 14538 6132
rect 14504 6030 14538 6064
rect 14504 5962 14538 5996
rect 14504 5894 14538 5928
rect 15070 6778 15104 6812
rect 15070 6710 15104 6744
rect 15070 6642 15104 6676
rect 15070 6574 15104 6608
rect 15070 6506 15104 6540
rect 15070 6438 15104 6472
rect 15070 6370 15104 6404
rect 15070 6302 15104 6336
rect 15070 6234 15104 6268
rect 15070 6166 15104 6200
rect 15070 6098 15104 6132
rect 15070 6030 15104 6064
rect 15070 5962 15104 5996
rect 15070 5894 15104 5928
rect 15636 6778 15670 6812
rect 15636 6710 15670 6744
rect 15636 6642 15670 6676
rect 15636 6574 15670 6608
rect 15636 6506 15670 6540
rect 15636 6438 15670 6472
rect 15636 6370 15670 6404
rect 15636 6302 15670 6336
rect 15636 6234 15670 6268
rect 15636 6166 15670 6200
rect 15636 6098 15670 6132
rect 15636 6030 15670 6064
rect 15636 5962 15670 5996
rect 15636 5894 15670 5928
rect 15990 6120 16024 6154
rect 15990 6050 16024 6084
rect 15990 5980 16024 6014
rect 15990 5910 16024 5944
rect 15990 5840 16024 5874
rect 15990 5770 16024 5804
rect 15990 5700 16024 5734
rect 15990 5630 16024 5664
rect 15990 5560 16024 5594
rect 15990 5490 16024 5524
rect 15990 5420 16024 5454
rect 15990 5350 16024 5384
rect 15990 5280 16024 5314
rect 15990 5210 16024 5244
rect 17280 6120 17314 6154
rect 17280 6050 17314 6084
rect 17280 5980 17314 6014
rect 17280 5910 17314 5944
rect 17280 5840 17314 5874
rect 17280 5770 17314 5804
rect 17280 5700 17314 5734
rect 17280 5630 17314 5664
rect 17280 5560 17314 5594
rect 17280 5490 17314 5524
rect 17280 5420 17314 5454
rect 17280 5350 17314 5384
rect 17280 5280 17314 5314
rect 17280 5210 17314 5244
rect 15990 5140 16024 5174
rect 17280 5140 17314 5174
rect 16070 5050 16104 5084
rect 16140 5050 16174 5084
rect 16210 5050 16244 5084
rect 16280 5050 16314 5084
rect 16350 5050 16384 5084
rect 16420 5050 16454 5084
rect 16490 5050 16524 5084
rect 16560 5050 16594 5084
rect 16630 5050 16664 5084
rect 16700 5050 16734 5084
rect 16770 5050 16804 5084
rect 16840 5050 16874 5084
rect 16910 5050 16944 5084
rect 16980 5050 17014 5084
rect 17050 5050 17084 5084
rect 17120 5050 17154 5084
rect 17190 5050 17224 5084
<< nsubdiffcont >>
rect 17678 8050 17718 8090
rect 17758 8050 17798 8090
rect 17838 8050 17878 8090
rect 17918 8050 17958 8090
rect 17998 8050 18038 8090
rect 18078 8050 18118 8090
rect 18158 8050 18198 8090
rect 18238 8050 18278 8090
rect 18318 8050 18358 8090
rect 18398 8050 18438 8090
rect 18478 8050 18518 8090
rect 18558 8050 18598 8090
rect 18638 8050 18678 8090
rect 18718 8050 18758 8090
rect 18798 8050 18838 8090
rect 18878 8050 18918 8090
rect 18958 8050 18998 8090
rect 19038 8050 19078 8090
rect 19118 8050 19158 8090
rect 19198 8050 19238 8090
rect 19278 8050 19318 8090
rect 19358 8050 19398 8090
rect 19438 8050 19478 8090
rect 19518 8050 19558 8090
rect 19598 8050 19638 8090
rect 19678 8050 19718 8090
rect 19758 8050 19798 8090
rect 19838 8050 19878 8090
rect 19918 8050 19958 8090
rect 19998 8050 20038 8090
rect 17498 7890 17538 7930
rect 17498 7810 17538 7850
rect 17498 7730 17538 7770
rect 17498 7650 17538 7690
rect 17498 7570 17538 7610
rect 17498 7490 17538 7530
rect 17498 7410 17538 7450
rect 17498 7330 17538 7370
rect 17498 7250 17538 7290
rect 17498 7170 17538 7210
rect 17498 7090 17538 7130
rect 17498 7010 17538 7050
rect 20158 7890 20198 7930
rect 20158 7810 20198 7850
rect 20158 7730 20198 7770
rect 20158 7650 20198 7690
rect 20158 7570 20198 7610
rect 20158 7490 20198 7530
rect 20158 7410 20198 7450
rect 20158 7330 20198 7370
rect 20158 7250 20198 7290
rect 20158 7170 20198 7210
rect 20158 7090 20198 7130
rect 20158 7010 20198 7050
rect 17480 6140 17520 6180
rect 17480 6060 17520 6100
rect 17480 5980 17520 6020
rect 17480 5900 17520 5940
rect 17480 5820 17520 5860
rect 17480 5740 17520 5780
rect 17480 5660 17520 5700
rect 17480 5580 17520 5620
rect 17480 5500 17520 5540
rect 17480 5420 17520 5460
rect 17480 5340 17520 5380
rect 17480 5260 17520 5300
rect 20140 6140 20180 6180
rect 20140 6060 20180 6100
rect 20140 5980 20180 6020
rect 20140 5900 20180 5940
rect 20140 5820 20180 5860
rect 20140 5740 20180 5780
rect 20140 5660 20180 5700
rect 20140 5580 20180 5620
rect 20140 5500 20180 5540
rect 20140 5420 20180 5460
rect 20140 5340 20180 5380
rect 20140 5260 20180 5300
rect 17660 5100 17700 5140
rect 17740 5100 17780 5140
rect 17820 5100 17860 5140
rect 17900 5100 17940 5140
rect 17980 5100 18020 5140
rect 18060 5100 18100 5140
rect 18140 5100 18180 5140
rect 18220 5100 18260 5140
rect 18300 5100 18340 5140
rect 18380 5100 18420 5140
rect 18460 5100 18500 5140
rect 18540 5100 18580 5140
rect 18620 5100 18660 5140
rect 18700 5100 18740 5140
rect 18780 5100 18820 5140
rect 18860 5100 18900 5140
rect 18940 5100 18980 5140
rect 19020 5100 19060 5140
rect 19100 5100 19140 5140
rect 19180 5100 19220 5140
rect 19260 5100 19300 5140
rect 19340 5100 19380 5140
rect 19420 5100 19460 5140
rect 19500 5100 19540 5140
rect 19580 5100 19620 5140
rect 19660 5100 19700 5140
rect 19740 5100 19780 5140
rect 19820 5100 19860 5140
rect 19900 5100 19940 5140
rect 19980 5100 20020 5140
<< poly >>
rect 16163 8005 16451 8035
rect 16163 7979 16193 8005
rect 16249 7979 16279 8005
rect 16335 7979 16365 8005
rect 16421 7979 16451 8005
rect 16507 8005 16795 8035
rect 16507 7979 16537 8005
rect 16593 7979 16623 8005
rect 16679 7979 16709 8005
rect 16765 7979 16795 8005
rect 16851 8005 17139 8035
rect 16851 7979 16881 8005
rect 16937 7979 16967 8005
rect 17023 7979 17053 8005
rect 17109 7979 17139 8005
rect 17667 7957 17697 7983
rect 17753 7957 17783 7983
rect 17839 7957 17869 7983
rect 17925 7957 17955 7983
rect 18011 7957 18041 7983
rect 18097 7957 18127 7983
rect 18183 7957 18213 7983
rect 18269 7957 18299 7983
rect 18355 7957 18385 7983
rect 18441 7957 18471 7983
rect 18527 7957 18557 7983
rect 18613 7957 18643 7983
rect 18699 7957 18729 7983
rect 18785 7957 18815 7983
rect 18871 7957 18901 7983
rect 18957 7957 18987 7983
rect 19043 7957 19073 7983
rect 19129 7957 19159 7983
rect 19215 7957 19245 7983
rect 19301 7957 19331 7983
rect 19387 7957 19417 7983
rect 19473 7957 19503 7983
rect 19559 7957 19589 7983
rect 19645 7957 19675 7983
rect 19731 7957 19761 7983
rect 19817 7957 19847 7983
rect 19903 7957 19933 7983
rect 19989 7957 20019 7983
rect 11805 6930 12143 6950
rect 11805 6896 11821 6930
rect 11855 6896 11889 6930
rect 11923 6896 11957 6930
rect 11991 6896 12025 6930
rect 12059 6896 12093 6930
rect 12127 6896 12143 6930
rect 11805 6880 12143 6896
rect 12371 6930 12709 6950
rect 12371 6896 12387 6930
rect 12421 6896 12455 6930
rect 12489 6896 12523 6930
rect 12557 6896 12591 6930
rect 12625 6896 12659 6930
rect 12693 6896 12709 6930
rect 12371 6880 12709 6896
rect 12937 6930 13275 6950
rect 12937 6896 12953 6930
rect 12987 6896 13021 6930
rect 13055 6896 13089 6930
rect 13123 6896 13157 6930
rect 13191 6896 13225 6930
rect 13259 6896 13275 6930
rect 12937 6880 13275 6896
rect 13503 6930 13841 6950
rect 13503 6896 13519 6930
rect 13553 6896 13587 6930
rect 13621 6896 13655 6930
rect 13689 6896 13723 6930
rect 13757 6896 13791 6930
rect 13825 6896 13841 6930
rect 13503 6880 13841 6896
rect 14069 6930 14407 6950
rect 14069 6896 14085 6930
rect 14119 6896 14153 6930
rect 14187 6896 14221 6930
rect 14255 6896 14289 6930
rect 14323 6896 14357 6930
rect 14391 6896 14407 6930
rect 14069 6880 14407 6896
rect 14635 6930 14973 6950
rect 14635 6896 14651 6930
rect 14685 6896 14719 6930
rect 14753 6896 14787 6930
rect 14821 6896 14855 6930
rect 14889 6896 14923 6930
rect 14957 6896 14973 6930
rect 14635 6880 14973 6896
rect 15201 6930 15539 6950
rect 16163 6947 16193 6969
rect 16249 6947 16279 6969
rect 16335 6947 16365 6969
rect 16421 6947 16451 6969
rect 16507 6947 16537 6969
rect 16593 6947 16623 6969
rect 16679 6947 16709 6969
rect 16765 6947 16795 6969
rect 16851 6947 16881 6969
rect 16937 6947 16967 6969
rect 17023 6947 17053 6969
rect 17109 6947 17139 6969
rect 15201 6896 15217 6930
rect 15251 6896 15285 6930
rect 15319 6896 15353 6930
rect 15387 6896 15421 6930
rect 15455 6896 15489 6930
rect 15523 6896 15539 6930
rect 15201 6880 15539 6896
rect 16138 6931 17185 6947
rect 16138 6897 16154 6931
rect 16188 6897 16222 6931
rect 16256 6897 16290 6931
rect 16324 6897 16358 6931
rect 16392 6897 16426 6931
rect 16460 6897 16494 6931
rect 16528 6897 16566 6931
rect 16600 6897 16634 6931
rect 16668 6897 16702 6931
rect 16736 6897 16770 6931
rect 16804 6897 16838 6931
rect 16872 6897 16910 6931
rect 16944 6897 16978 6931
rect 17012 6897 17046 6931
rect 17080 6897 17185 6931
rect 11830 6858 11860 6880
rect 11916 6858 11946 6880
rect 12002 6858 12032 6880
rect 12088 6858 12118 6880
rect 12396 6858 12426 6880
rect 12482 6858 12512 6880
rect 12568 6858 12598 6880
rect 12654 6858 12684 6880
rect 12962 6858 12992 6880
rect 13048 6858 13078 6880
rect 13134 6858 13164 6880
rect 13220 6858 13250 6880
rect 13528 6858 13558 6880
rect 13614 6858 13644 6880
rect 13700 6858 13730 6880
rect 13786 6858 13816 6880
rect 14094 6858 14124 6880
rect 14180 6858 14210 6880
rect 14266 6858 14296 6880
rect 14352 6858 14382 6880
rect 14660 6858 14690 6880
rect 14746 6858 14776 6880
rect 14832 6858 14862 6880
rect 14918 6858 14948 6880
rect 15226 6858 15256 6880
rect 15312 6858 15342 6880
rect 15398 6858 15428 6880
rect 15484 6858 15514 6880
rect 16138 6877 17185 6897
rect 17667 6931 17697 6957
rect 17753 6931 17783 6957
rect 17839 6931 17869 6957
rect 17925 6931 17955 6957
rect 17667 6908 17955 6931
rect 17667 6874 17692 6908
rect 17726 6874 17760 6908
rect 17794 6874 17828 6908
rect 17862 6874 17896 6908
rect 17930 6874 17955 6908
rect 17667 6858 17955 6874
rect 18011 6931 18041 6957
rect 18097 6931 18127 6957
rect 18183 6931 18213 6957
rect 18269 6931 18299 6957
rect 18011 6908 18299 6931
rect 18011 6874 18036 6908
rect 18070 6874 18104 6908
rect 18138 6874 18172 6908
rect 18206 6874 18240 6908
rect 18274 6874 18299 6908
rect 18011 6858 18299 6874
rect 18355 6931 18385 6957
rect 18441 6931 18471 6957
rect 18527 6931 18557 6957
rect 18613 6931 18643 6957
rect 18355 6908 18643 6931
rect 18355 6874 18380 6908
rect 18414 6874 18448 6908
rect 18482 6874 18516 6908
rect 18550 6874 18584 6908
rect 18618 6874 18643 6908
rect 18355 6858 18643 6874
rect 18699 6931 18729 6957
rect 18785 6931 18815 6957
rect 18871 6931 18901 6957
rect 18957 6931 18987 6957
rect 18699 6908 18987 6931
rect 18699 6874 18724 6908
rect 18758 6874 18792 6908
rect 18826 6874 18860 6908
rect 18894 6874 18928 6908
rect 18962 6874 18987 6908
rect 18699 6858 18987 6874
rect 19043 6931 19073 6957
rect 19129 6931 19159 6957
rect 19215 6931 19245 6957
rect 19301 6931 19331 6957
rect 19043 6908 19331 6931
rect 19043 6874 19068 6908
rect 19102 6874 19136 6908
rect 19170 6874 19204 6908
rect 19238 6874 19272 6908
rect 19306 6874 19331 6908
rect 19043 6858 19331 6874
rect 19387 6931 19417 6957
rect 19473 6931 19503 6957
rect 19559 6931 19589 6957
rect 19645 6931 19675 6957
rect 19387 6908 19675 6931
rect 19387 6874 19412 6908
rect 19446 6874 19480 6908
rect 19514 6874 19548 6908
rect 19582 6874 19616 6908
rect 19650 6874 19675 6908
rect 19387 6858 19675 6874
rect 19731 6931 19761 6957
rect 19817 6931 19847 6957
rect 19903 6931 19933 6957
rect 19989 6931 20019 6957
rect 19731 6908 20019 6931
rect 19731 6874 19756 6908
rect 19790 6874 19824 6908
rect 19858 6874 19892 6908
rect 19926 6874 19960 6908
rect 19994 6874 20019 6908
rect 19731 6858 20019 6874
rect 17649 6316 17937 6332
rect 16138 6263 17185 6283
rect 16138 6229 16154 6263
rect 16188 6229 16222 6263
rect 16256 6229 16290 6263
rect 16324 6229 16358 6263
rect 16392 6229 16426 6263
rect 16460 6229 16494 6263
rect 16528 6229 16566 6263
rect 16600 6229 16634 6263
rect 16668 6229 16702 6263
rect 16736 6229 16770 6263
rect 16804 6229 16838 6263
rect 16872 6229 16910 6263
rect 16944 6229 16978 6263
rect 17012 6229 17046 6263
rect 17080 6229 17185 6263
rect 17649 6282 17674 6316
rect 17708 6282 17742 6316
rect 17776 6282 17810 6316
rect 17844 6282 17878 6316
rect 17912 6282 17937 6316
rect 17649 6259 17937 6282
rect 17649 6233 17679 6259
rect 17735 6233 17765 6259
rect 17821 6233 17851 6259
rect 17907 6233 17937 6259
rect 17993 6316 18281 6332
rect 17993 6282 18018 6316
rect 18052 6282 18086 6316
rect 18120 6282 18154 6316
rect 18188 6282 18222 6316
rect 18256 6282 18281 6316
rect 17993 6259 18281 6282
rect 17993 6233 18023 6259
rect 18079 6233 18109 6259
rect 18165 6233 18195 6259
rect 18251 6233 18281 6259
rect 18337 6316 18625 6332
rect 18337 6282 18362 6316
rect 18396 6282 18430 6316
rect 18464 6282 18498 6316
rect 18532 6282 18566 6316
rect 18600 6282 18625 6316
rect 18337 6259 18625 6282
rect 18337 6233 18367 6259
rect 18423 6233 18453 6259
rect 18509 6233 18539 6259
rect 18595 6233 18625 6259
rect 18681 6316 18969 6332
rect 18681 6282 18706 6316
rect 18740 6282 18774 6316
rect 18808 6282 18842 6316
rect 18876 6282 18910 6316
rect 18944 6282 18969 6316
rect 18681 6259 18969 6282
rect 18681 6233 18711 6259
rect 18767 6233 18797 6259
rect 18853 6233 18883 6259
rect 18939 6233 18969 6259
rect 19025 6316 19313 6332
rect 19025 6282 19050 6316
rect 19084 6282 19118 6316
rect 19152 6282 19186 6316
rect 19220 6282 19254 6316
rect 19288 6282 19313 6316
rect 19025 6259 19313 6282
rect 19025 6233 19055 6259
rect 19111 6233 19141 6259
rect 19197 6233 19227 6259
rect 19283 6233 19313 6259
rect 19369 6316 19657 6332
rect 19369 6282 19394 6316
rect 19428 6282 19462 6316
rect 19496 6282 19530 6316
rect 19564 6282 19598 6316
rect 19632 6282 19657 6316
rect 19369 6259 19657 6282
rect 19369 6233 19399 6259
rect 19455 6233 19485 6259
rect 19541 6233 19571 6259
rect 19627 6233 19657 6259
rect 19713 6316 20001 6332
rect 19713 6282 19738 6316
rect 19772 6282 19806 6316
rect 19840 6282 19874 6316
rect 19908 6282 19942 6316
rect 19976 6282 20001 6316
rect 19713 6259 20001 6282
rect 19713 6233 19743 6259
rect 19799 6233 19829 6259
rect 19885 6233 19915 6259
rect 19971 6233 20001 6259
rect 16138 6213 17185 6229
rect 16163 6191 16193 6213
rect 16249 6191 16279 6213
rect 16335 6191 16365 6213
rect 16421 6191 16451 6213
rect 16507 6191 16537 6213
rect 16593 6191 16623 6213
rect 16679 6191 16709 6213
rect 16765 6191 16795 6213
rect 16851 6191 16881 6213
rect 16937 6191 16967 6213
rect 17023 6191 17053 6213
rect 17109 6191 17139 6213
rect 11830 5826 11860 5848
rect 11916 5826 11946 5848
rect 12002 5826 12032 5848
rect 12088 5826 12118 5848
rect 12396 5826 12426 5848
rect 12482 5826 12512 5848
rect 12568 5826 12598 5848
rect 12654 5826 12684 5848
rect 12962 5826 12992 5848
rect 13048 5826 13078 5848
rect 13134 5826 13164 5848
rect 13220 5826 13250 5848
rect 13528 5826 13558 5848
rect 13614 5826 13644 5848
rect 13700 5826 13730 5848
rect 13786 5826 13816 5848
rect 14094 5826 14124 5848
rect 14180 5826 14210 5848
rect 14266 5826 14296 5848
rect 14352 5826 14382 5848
rect 14660 5826 14690 5848
rect 14746 5826 14776 5848
rect 14832 5826 14862 5848
rect 14918 5826 14948 5848
rect 15226 5826 15256 5848
rect 15312 5826 15342 5848
rect 15398 5826 15428 5848
rect 15484 5826 15514 5848
rect 11805 5810 12143 5826
rect 11805 5776 11821 5810
rect 11855 5776 11889 5810
rect 11923 5776 11957 5810
rect 11991 5776 12025 5810
rect 12059 5776 12093 5810
rect 12127 5776 12143 5810
rect 11805 5756 12143 5776
rect 12371 5810 12709 5826
rect 12371 5776 12387 5810
rect 12421 5776 12455 5810
rect 12489 5776 12523 5810
rect 12557 5776 12591 5810
rect 12625 5776 12659 5810
rect 12693 5776 12709 5810
rect 12371 5756 12709 5776
rect 12937 5810 13275 5826
rect 12937 5776 12953 5810
rect 12987 5776 13021 5810
rect 13055 5776 13089 5810
rect 13123 5776 13157 5810
rect 13191 5776 13225 5810
rect 13259 5776 13275 5810
rect 12937 5756 13275 5776
rect 13503 5810 13841 5826
rect 13503 5776 13519 5810
rect 13553 5776 13587 5810
rect 13621 5776 13655 5810
rect 13689 5776 13723 5810
rect 13757 5776 13791 5810
rect 13825 5776 13841 5810
rect 13503 5756 13841 5776
rect 14069 5810 14407 5826
rect 14069 5776 14085 5810
rect 14119 5776 14153 5810
rect 14187 5776 14221 5810
rect 14255 5776 14289 5810
rect 14323 5776 14357 5810
rect 14391 5776 14407 5810
rect 14069 5756 14407 5776
rect 14635 5810 14973 5826
rect 14635 5776 14651 5810
rect 14685 5776 14719 5810
rect 14753 5776 14787 5810
rect 14821 5776 14855 5810
rect 14889 5776 14923 5810
rect 14957 5776 14973 5810
rect 14635 5756 14973 5776
rect 15201 5810 15539 5826
rect 15201 5776 15217 5810
rect 15251 5776 15285 5810
rect 15319 5776 15353 5810
rect 15387 5776 15421 5810
rect 15455 5776 15489 5810
rect 15523 5776 15539 5810
rect 15201 5756 15539 5776
rect 16163 5155 16193 5181
rect 16249 5155 16279 5181
rect 16335 5155 16365 5181
rect 16421 5155 16451 5181
rect 16163 5125 16451 5155
rect 16507 5155 16537 5181
rect 16593 5155 16623 5181
rect 16679 5155 16709 5181
rect 16765 5155 16795 5181
rect 16507 5125 16795 5155
rect 16851 5155 16881 5181
rect 16937 5155 16967 5181
rect 17023 5155 17053 5181
rect 17109 5155 17139 5181
rect 16851 5125 17139 5155
rect 17649 5207 17679 5233
rect 17735 5207 17765 5233
rect 17821 5207 17851 5233
rect 17907 5207 17937 5233
rect 17993 5207 18023 5233
rect 18079 5207 18109 5233
rect 18165 5207 18195 5233
rect 18251 5207 18281 5233
rect 18337 5207 18367 5233
rect 18423 5207 18453 5233
rect 18509 5207 18539 5233
rect 18595 5207 18625 5233
rect 18681 5207 18711 5233
rect 18767 5207 18797 5233
rect 18853 5207 18883 5233
rect 18939 5207 18969 5233
rect 19025 5207 19055 5233
rect 19111 5207 19141 5233
rect 19197 5207 19227 5233
rect 19283 5207 19313 5233
rect 19369 5207 19399 5233
rect 19455 5207 19485 5233
rect 19541 5207 19571 5233
rect 19627 5207 19657 5233
rect 19713 5207 19743 5233
rect 19799 5207 19829 5233
rect 19885 5207 19915 5233
rect 19971 5207 20001 5233
<< polycont >>
rect 11821 6896 11855 6930
rect 11889 6896 11923 6930
rect 11957 6896 11991 6930
rect 12025 6896 12059 6930
rect 12093 6896 12127 6930
rect 12387 6896 12421 6930
rect 12455 6896 12489 6930
rect 12523 6896 12557 6930
rect 12591 6896 12625 6930
rect 12659 6896 12693 6930
rect 12953 6896 12987 6930
rect 13021 6896 13055 6930
rect 13089 6896 13123 6930
rect 13157 6896 13191 6930
rect 13225 6896 13259 6930
rect 13519 6896 13553 6930
rect 13587 6896 13621 6930
rect 13655 6896 13689 6930
rect 13723 6896 13757 6930
rect 13791 6896 13825 6930
rect 14085 6896 14119 6930
rect 14153 6896 14187 6930
rect 14221 6896 14255 6930
rect 14289 6896 14323 6930
rect 14357 6896 14391 6930
rect 14651 6896 14685 6930
rect 14719 6896 14753 6930
rect 14787 6896 14821 6930
rect 14855 6896 14889 6930
rect 14923 6896 14957 6930
rect 15217 6896 15251 6930
rect 15285 6896 15319 6930
rect 15353 6896 15387 6930
rect 15421 6896 15455 6930
rect 15489 6896 15523 6930
rect 16154 6897 16188 6931
rect 16222 6897 16256 6931
rect 16290 6897 16324 6931
rect 16358 6897 16392 6931
rect 16426 6897 16460 6931
rect 16494 6897 16528 6931
rect 16566 6897 16600 6931
rect 16634 6897 16668 6931
rect 16702 6897 16736 6931
rect 16770 6897 16804 6931
rect 16838 6897 16872 6931
rect 16910 6897 16944 6931
rect 16978 6897 17012 6931
rect 17046 6897 17080 6931
rect 17692 6874 17726 6908
rect 17760 6874 17794 6908
rect 17828 6874 17862 6908
rect 17896 6874 17930 6908
rect 18036 6874 18070 6908
rect 18104 6874 18138 6908
rect 18172 6874 18206 6908
rect 18240 6874 18274 6908
rect 18380 6874 18414 6908
rect 18448 6874 18482 6908
rect 18516 6874 18550 6908
rect 18584 6874 18618 6908
rect 18724 6874 18758 6908
rect 18792 6874 18826 6908
rect 18860 6874 18894 6908
rect 18928 6874 18962 6908
rect 19068 6874 19102 6908
rect 19136 6874 19170 6908
rect 19204 6874 19238 6908
rect 19272 6874 19306 6908
rect 19412 6874 19446 6908
rect 19480 6874 19514 6908
rect 19548 6874 19582 6908
rect 19616 6874 19650 6908
rect 19756 6874 19790 6908
rect 19824 6874 19858 6908
rect 19892 6874 19926 6908
rect 19960 6874 19994 6908
rect 16154 6229 16188 6263
rect 16222 6229 16256 6263
rect 16290 6229 16324 6263
rect 16358 6229 16392 6263
rect 16426 6229 16460 6263
rect 16494 6229 16528 6263
rect 16566 6229 16600 6263
rect 16634 6229 16668 6263
rect 16702 6229 16736 6263
rect 16770 6229 16804 6263
rect 16838 6229 16872 6263
rect 16910 6229 16944 6263
rect 16978 6229 17012 6263
rect 17046 6229 17080 6263
rect 17674 6282 17708 6316
rect 17742 6282 17776 6316
rect 17810 6282 17844 6316
rect 17878 6282 17912 6316
rect 18018 6282 18052 6316
rect 18086 6282 18120 6316
rect 18154 6282 18188 6316
rect 18222 6282 18256 6316
rect 18362 6282 18396 6316
rect 18430 6282 18464 6316
rect 18498 6282 18532 6316
rect 18566 6282 18600 6316
rect 18706 6282 18740 6316
rect 18774 6282 18808 6316
rect 18842 6282 18876 6316
rect 18910 6282 18944 6316
rect 19050 6282 19084 6316
rect 19118 6282 19152 6316
rect 19186 6282 19220 6316
rect 19254 6282 19288 6316
rect 19394 6282 19428 6316
rect 19462 6282 19496 6316
rect 19530 6282 19564 6316
rect 19598 6282 19632 6316
rect 19738 6282 19772 6316
rect 19806 6282 19840 6316
rect 19874 6282 19908 6316
rect 19942 6282 19976 6316
rect 11821 5776 11855 5810
rect 11889 5776 11923 5810
rect 11957 5776 11991 5810
rect 12025 5776 12059 5810
rect 12093 5776 12127 5810
rect 12387 5776 12421 5810
rect 12455 5776 12489 5810
rect 12523 5776 12557 5810
rect 12591 5776 12625 5810
rect 12659 5776 12693 5810
rect 12953 5776 12987 5810
rect 13021 5776 13055 5810
rect 13089 5776 13123 5810
rect 13157 5776 13191 5810
rect 13225 5776 13259 5810
rect 13519 5776 13553 5810
rect 13587 5776 13621 5810
rect 13655 5776 13689 5810
rect 13723 5776 13757 5810
rect 13791 5776 13825 5810
rect 14085 5776 14119 5810
rect 14153 5776 14187 5810
rect 14221 5776 14255 5810
rect 14289 5776 14323 5810
rect 14357 5776 14391 5810
rect 14651 5776 14685 5810
rect 14719 5776 14753 5810
rect 14787 5776 14821 5810
rect 14855 5776 14889 5810
rect 14923 5776 14957 5810
rect 15217 5776 15251 5810
rect 15285 5776 15319 5810
rect 15353 5776 15387 5810
rect 15421 5776 15455 5810
rect 15489 5776 15523 5810
<< locali >>
rect 16550 9852 18266 9868
rect 16550 9818 16635 9852
rect 16669 9818 16707 9852
rect 16741 9818 16779 9852
rect 16813 9818 16851 9852
rect 16885 9818 16923 9852
rect 16957 9818 16995 9852
rect 17029 9818 17067 9852
rect 17101 9818 17139 9852
rect 17173 9818 17211 9852
rect 17245 9818 17283 9852
rect 17317 9818 17355 9852
rect 17389 9818 17427 9852
rect 17461 9818 17499 9852
rect 17533 9818 17571 9852
rect 17605 9818 17643 9852
rect 17677 9818 17715 9852
rect 17749 9818 17787 9852
rect 17821 9818 17859 9852
rect 17893 9818 17931 9852
rect 17965 9818 18003 9852
rect 18037 9818 18075 9852
rect 18109 9818 18147 9852
rect 18181 9818 18266 9852
rect 16550 9785 18266 9818
rect 16550 9751 16566 9785
rect 16600 9751 18216 9785
rect 18250 9751 18266 9785
rect 16550 9713 18266 9751
rect 16550 9679 16566 9713
rect 16600 9679 18216 9713
rect 18250 9679 18266 9713
rect 16550 9641 18266 9679
rect 16550 9607 16566 9641
rect 16600 9607 18216 9641
rect 18250 9607 18266 9641
rect 16550 9569 18266 9607
rect 16550 9535 16566 9569
rect 16600 9535 18216 9569
rect 18250 9535 18266 9569
rect 16550 9497 18266 9535
rect 16550 9463 16566 9497
rect 16600 9463 18216 9497
rect 18250 9463 18266 9497
rect 16550 9425 18266 9463
rect 16550 9391 16566 9425
rect 16600 9391 18216 9425
rect 18250 9391 18266 9425
rect 16550 9353 18266 9391
rect 16550 9319 16566 9353
rect 16600 9319 18216 9353
rect 18250 9319 18266 9353
rect 16550 9281 18266 9319
rect 16550 9247 16566 9281
rect 16600 9247 18216 9281
rect 18250 9247 18266 9281
rect 16550 9209 18266 9247
rect 16550 9175 16566 9209
rect 16600 9175 18216 9209
rect 18250 9175 18266 9209
rect 16550 9137 18266 9175
rect 16550 9103 16566 9137
rect 16600 9103 18216 9137
rect 18250 9103 18266 9137
rect 16550 9065 18266 9103
rect 16550 9031 16566 9065
rect 16600 9031 18216 9065
rect 18250 9031 18266 9065
rect 16550 8993 18266 9031
rect 16550 8959 16566 8993
rect 16600 8959 18216 8993
rect 18250 8959 18266 8993
rect 16550 8921 18266 8959
rect 16550 8887 16566 8921
rect 16600 8887 18216 8921
rect 18250 8887 18266 8921
rect 16550 8849 18266 8887
rect 16550 8815 16566 8849
rect 16600 8815 18216 8849
rect 18250 8815 18266 8849
rect 16550 8777 18266 8815
rect 16550 8743 16566 8777
rect 16600 8743 18216 8777
rect 18250 8743 18266 8777
rect 16550 8705 18266 8743
rect 16550 8671 16566 8705
rect 16600 8671 18216 8705
rect 18250 8671 18266 8705
rect 16550 8633 18266 8671
rect 16550 8599 16566 8633
rect 16600 8599 18216 8633
rect 18250 8599 18266 8633
rect 16550 8561 18266 8599
rect 16550 8527 16566 8561
rect 16600 8527 18216 8561
rect 18250 8527 18266 8561
rect 16550 8489 18266 8527
rect 16550 8455 16566 8489
rect 16600 8455 18216 8489
rect 18250 8455 18266 8489
rect 16550 8417 18266 8455
rect 16550 8383 16566 8417
rect 16600 8383 18216 8417
rect 18250 8383 18266 8417
rect 16550 8350 18266 8383
rect 16550 8316 16635 8350
rect 16669 8316 16707 8350
rect 16741 8316 16779 8350
rect 16813 8316 16851 8350
rect 16885 8316 16923 8350
rect 16957 8316 16995 8350
rect 17029 8316 17067 8350
rect 17101 8316 17139 8350
rect 17173 8316 17211 8350
rect 17245 8316 17283 8350
rect 17317 8316 17355 8350
rect 17389 8316 17427 8350
rect 17461 8316 17499 8350
rect 17533 8316 17571 8350
rect 17605 8316 17643 8350
rect 17677 8316 17715 8350
rect 17749 8316 17787 8350
rect 17821 8316 17859 8350
rect 17893 8316 17931 8350
rect 17965 8316 18003 8350
rect 18037 8316 18075 8350
rect 18109 8316 18147 8350
rect 18181 8316 18266 8350
rect 16550 8300 18266 8316
rect 18400 9852 20116 9868
rect 18400 9818 18485 9852
rect 18519 9818 18557 9852
rect 18591 9818 18629 9852
rect 18663 9818 18701 9852
rect 18735 9818 18773 9852
rect 18807 9818 18845 9852
rect 18879 9818 18917 9852
rect 18951 9818 18989 9852
rect 19023 9818 19061 9852
rect 19095 9818 19133 9852
rect 19167 9818 19205 9852
rect 19239 9818 19277 9852
rect 19311 9818 19349 9852
rect 19383 9818 19421 9852
rect 19455 9818 19493 9852
rect 19527 9818 19565 9852
rect 19599 9818 19637 9852
rect 19671 9818 19709 9852
rect 19743 9818 19781 9852
rect 19815 9818 19853 9852
rect 19887 9818 19925 9852
rect 19959 9818 19997 9852
rect 20031 9818 20116 9852
rect 18400 9785 20116 9818
rect 18400 9751 18416 9785
rect 18450 9751 20066 9785
rect 20100 9751 20116 9785
rect 18400 9713 20116 9751
rect 18400 9679 18416 9713
rect 18450 9679 20066 9713
rect 20100 9679 20116 9713
rect 18400 9641 20116 9679
rect 18400 9607 18416 9641
rect 18450 9607 20066 9641
rect 20100 9607 20116 9641
rect 18400 9569 20116 9607
rect 18400 9535 18416 9569
rect 18450 9535 20066 9569
rect 20100 9535 20116 9569
rect 18400 9497 20116 9535
rect 18400 9463 18416 9497
rect 18450 9463 20066 9497
rect 20100 9463 20116 9497
rect 18400 9425 20116 9463
rect 18400 9391 18416 9425
rect 18450 9391 20066 9425
rect 20100 9391 20116 9425
rect 18400 9353 20116 9391
rect 18400 9319 18416 9353
rect 18450 9319 20066 9353
rect 20100 9319 20116 9353
rect 18400 9281 20116 9319
rect 18400 9247 18416 9281
rect 18450 9247 20066 9281
rect 20100 9247 20116 9281
rect 18400 9209 20116 9247
rect 18400 9175 18416 9209
rect 18450 9175 20066 9209
rect 20100 9175 20116 9209
rect 18400 9137 20116 9175
rect 18400 9103 18416 9137
rect 18450 9103 20066 9137
rect 20100 9103 20116 9137
rect 18400 9065 20116 9103
rect 18400 9031 18416 9065
rect 18450 9031 20066 9065
rect 20100 9031 20116 9065
rect 18400 8993 20116 9031
rect 18400 8959 18416 8993
rect 18450 8959 20066 8993
rect 20100 8959 20116 8993
rect 18400 8921 20116 8959
rect 18400 8887 18416 8921
rect 18450 8887 20066 8921
rect 20100 8887 20116 8921
rect 18400 8849 20116 8887
rect 18400 8815 18416 8849
rect 18450 8815 20066 8849
rect 20100 8815 20116 8849
rect 18400 8777 20116 8815
rect 18400 8743 18416 8777
rect 18450 8743 20066 8777
rect 20100 8743 20116 8777
rect 18400 8705 20116 8743
rect 18400 8671 18416 8705
rect 18450 8671 20066 8705
rect 20100 8671 20116 8705
rect 18400 8633 20116 8671
rect 18400 8599 18416 8633
rect 18450 8599 20066 8633
rect 20100 8599 20116 8633
rect 18400 8561 20116 8599
rect 18400 8527 18416 8561
rect 18450 8527 20066 8561
rect 20100 8527 20116 8561
rect 18400 8489 20116 8527
rect 18400 8455 18416 8489
rect 18450 8455 20066 8489
rect 20100 8455 20116 8489
rect 18400 8417 20116 8455
rect 18400 8383 18416 8417
rect 18450 8383 20066 8417
rect 20100 8383 20116 8417
rect 18400 8350 20116 8383
rect 18400 8316 18485 8350
rect 18519 8316 18557 8350
rect 18591 8316 18629 8350
rect 18663 8316 18701 8350
rect 18735 8316 18773 8350
rect 18807 8316 18845 8350
rect 18879 8316 18917 8350
rect 18951 8316 18989 8350
rect 19023 8316 19061 8350
rect 19095 8316 19133 8350
rect 19167 8316 19205 8350
rect 19239 8316 19277 8350
rect 19311 8316 19349 8350
rect 19383 8316 19421 8350
rect 19455 8316 19493 8350
rect 19527 8316 19565 8350
rect 19599 8316 19637 8350
rect 19671 8316 19709 8350
rect 19743 8316 19781 8350
rect 19815 8316 19853 8350
rect 19887 8316 19925 8350
rect 19959 8316 19997 8350
rect 20031 8316 20116 8350
rect 18400 8300 20116 8316
rect 15980 8110 17330 8120
rect 15980 8076 16070 8110
rect 16114 8076 16140 8110
rect 16194 8076 16210 8110
rect 16274 8076 16280 8110
rect 16314 8076 16320 8110
rect 16384 8076 16400 8110
rect 16454 8076 16480 8110
rect 16524 8076 16560 8110
rect 16594 8076 16630 8110
rect 16674 8076 16700 8110
rect 16754 8076 16770 8110
rect 16834 8076 16840 8110
rect 16874 8076 16880 8110
rect 16944 8076 16960 8110
rect 17014 8076 17040 8110
rect 17084 8076 17120 8110
rect 17154 8076 17190 8110
rect 17224 8076 17330 8110
rect 15980 8060 17330 8076
rect 15980 8020 16030 8060
rect 15980 7966 15990 8020
rect 16024 7966 16030 8020
rect 17270 8020 17330 8060
rect 17618 8090 20078 8110
rect 17618 8050 17638 8090
rect 20058 8050 20078 8090
rect 17618 8030 20078 8050
rect 15980 7950 16030 7966
rect 15980 7886 15990 7950
rect 16024 7886 16030 7950
rect 15980 7880 16030 7886
rect 15980 7846 15990 7880
rect 16024 7846 16030 7880
rect 15980 7840 16030 7846
rect 15980 7776 15990 7840
rect 16024 7776 16030 7840
rect 15980 7760 16030 7776
rect 15980 7706 15990 7760
rect 16024 7706 16030 7760
rect 15980 7680 16030 7706
rect 15980 7636 15990 7680
rect 16024 7636 16030 7680
rect 15980 7600 16030 7636
rect 15980 7566 15990 7600
rect 16024 7566 16030 7600
rect 15980 7530 16030 7566
rect 15980 7486 15990 7530
rect 16024 7486 16030 7530
rect 15980 7460 16030 7486
rect 15980 7406 15990 7460
rect 16024 7406 16030 7460
rect 15980 7390 16030 7406
rect 15980 7326 15990 7390
rect 16024 7326 16030 7390
rect 15980 7320 16030 7326
rect 15980 7286 15990 7320
rect 16024 7286 16030 7320
rect 15980 7280 16030 7286
rect 15980 7216 15990 7280
rect 16024 7216 16030 7280
rect 15980 7200 16030 7216
rect 15980 7146 15990 7200
rect 16024 7146 16030 7200
rect 15980 7120 16030 7146
rect 15980 7076 15990 7120
rect 16024 7076 16030 7120
rect 15980 7040 16030 7076
rect 15980 7006 15990 7040
rect 16024 7006 16030 7040
rect 15980 6990 16030 7006
rect 16118 7967 16152 7983
rect 16118 7899 16152 7925
rect 16118 7831 16152 7853
rect 16118 7763 16152 7781
rect 16118 7695 16152 7709
rect 16118 7627 16152 7637
rect 16118 7559 16152 7565
rect 16118 7491 16152 7493
rect 16118 7455 16152 7457
rect 16118 7383 16152 7389
rect 16118 7311 16152 7321
rect 16118 7239 16152 7253
rect 16118 7167 16152 7185
rect 16118 7095 16152 7117
rect 16118 7023 16152 7049
rect 16118 6965 16152 6981
rect 16204 7967 16238 7983
rect 16204 7899 16238 7925
rect 16204 7831 16238 7853
rect 16204 7763 16238 7781
rect 16204 7695 16238 7709
rect 16204 7627 16238 7637
rect 16204 7559 16238 7565
rect 16204 7491 16238 7493
rect 16204 7455 16238 7457
rect 16204 7383 16238 7389
rect 16204 7311 16238 7321
rect 16204 7239 16238 7253
rect 16204 7167 16238 7185
rect 16204 7095 16238 7117
rect 16204 7023 16238 7049
rect 16204 6965 16238 6981
rect 16290 7967 16324 7983
rect 16290 7899 16324 7925
rect 16290 7831 16324 7853
rect 16290 7763 16324 7781
rect 16290 7695 16324 7709
rect 16290 7627 16324 7637
rect 16290 7559 16324 7565
rect 16290 7491 16324 7493
rect 16290 7455 16324 7457
rect 16290 7383 16324 7389
rect 16290 7311 16324 7321
rect 16290 7239 16324 7253
rect 16290 7167 16324 7185
rect 16290 7095 16324 7117
rect 16290 7023 16324 7049
rect 16290 6965 16324 6981
rect 16376 7967 16410 7983
rect 16376 7899 16410 7925
rect 16376 7831 16410 7853
rect 16376 7763 16410 7781
rect 16376 7695 16410 7709
rect 16376 7627 16410 7637
rect 16376 7559 16410 7565
rect 16376 7491 16410 7493
rect 16376 7455 16410 7457
rect 16376 7383 16410 7389
rect 16376 7311 16410 7321
rect 16376 7239 16410 7253
rect 16376 7167 16410 7185
rect 16376 7095 16410 7117
rect 16376 7023 16410 7049
rect 16376 6965 16410 6981
rect 16462 7967 16496 7983
rect 16462 7899 16496 7925
rect 16462 7831 16496 7853
rect 16462 7763 16496 7781
rect 16462 7695 16496 7709
rect 16462 7627 16496 7637
rect 16462 7559 16496 7565
rect 16462 7491 16496 7493
rect 16462 7455 16496 7457
rect 16462 7383 16496 7389
rect 16462 7311 16496 7321
rect 16462 7239 16496 7253
rect 16462 7167 16496 7185
rect 16462 7095 16496 7117
rect 16462 7023 16496 7049
rect 16462 6965 16496 6981
rect 16548 7967 16582 7983
rect 16548 7899 16582 7925
rect 16548 7831 16582 7853
rect 16548 7763 16582 7781
rect 16548 7695 16582 7709
rect 16548 7627 16582 7637
rect 16548 7559 16582 7565
rect 16548 7491 16582 7493
rect 16548 7455 16582 7457
rect 16548 7383 16582 7389
rect 16548 7311 16582 7321
rect 16548 7239 16582 7253
rect 16548 7167 16582 7185
rect 16548 7095 16582 7117
rect 16548 7023 16582 7049
rect 16548 6965 16582 6981
rect 16634 7967 16668 7983
rect 16634 7899 16668 7925
rect 16634 7831 16668 7853
rect 16634 7763 16668 7781
rect 16634 7695 16668 7709
rect 16634 7627 16668 7637
rect 16634 7559 16668 7565
rect 16634 7491 16668 7493
rect 16634 7455 16668 7457
rect 16634 7383 16668 7389
rect 16634 7311 16668 7321
rect 16634 7239 16668 7253
rect 16634 7167 16668 7185
rect 16634 7095 16668 7117
rect 16634 7023 16668 7049
rect 16634 6965 16668 6981
rect 16720 7967 16754 7983
rect 16720 7899 16754 7925
rect 16720 7831 16754 7853
rect 16720 7763 16754 7781
rect 16720 7695 16754 7709
rect 16720 7627 16754 7637
rect 16720 7559 16754 7565
rect 16720 7491 16754 7493
rect 16720 7455 16754 7457
rect 16720 7383 16754 7389
rect 16720 7311 16754 7321
rect 16720 7239 16754 7253
rect 16720 7167 16754 7185
rect 16720 7095 16754 7117
rect 16720 7023 16754 7049
rect 16720 6965 16754 6981
rect 16806 7967 16840 7983
rect 16806 7899 16840 7925
rect 16806 7831 16840 7853
rect 16806 7763 16840 7781
rect 16806 7695 16840 7709
rect 16806 7627 16840 7637
rect 16806 7559 16840 7565
rect 16806 7491 16840 7493
rect 16806 7455 16840 7457
rect 16806 7383 16840 7389
rect 16806 7311 16840 7321
rect 16806 7239 16840 7253
rect 16806 7167 16840 7185
rect 16806 7095 16840 7117
rect 16806 7023 16840 7049
rect 16806 6965 16840 6981
rect 16892 7967 16926 7983
rect 16892 7899 16926 7925
rect 16892 7831 16926 7853
rect 16892 7763 16926 7781
rect 16892 7695 16926 7709
rect 16892 7627 16926 7637
rect 16892 7559 16926 7565
rect 16892 7491 16926 7493
rect 16892 7455 16926 7457
rect 16892 7383 16926 7389
rect 16892 7311 16926 7321
rect 16892 7239 16926 7253
rect 16892 7167 16926 7185
rect 16892 7095 16926 7117
rect 16892 7023 16926 7049
rect 16892 6965 16926 6981
rect 16978 7967 17012 7983
rect 16978 7899 17012 7925
rect 16978 7831 17012 7853
rect 16978 7763 17012 7781
rect 16978 7695 17012 7709
rect 16978 7627 17012 7637
rect 16978 7559 17012 7565
rect 16978 7491 17012 7493
rect 16978 7455 17012 7457
rect 16978 7383 17012 7389
rect 16978 7311 17012 7321
rect 16978 7239 17012 7253
rect 16978 7167 17012 7185
rect 16978 7095 17012 7117
rect 16978 7023 17012 7049
rect 16978 6965 17012 6981
rect 17064 7967 17098 7983
rect 17064 7899 17098 7925
rect 17064 7831 17098 7853
rect 17064 7763 17098 7781
rect 17064 7695 17098 7709
rect 17064 7627 17098 7637
rect 17064 7559 17098 7565
rect 17064 7491 17098 7493
rect 17064 7455 17098 7457
rect 17064 7383 17098 7389
rect 17064 7311 17098 7321
rect 17064 7239 17098 7253
rect 17064 7167 17098 7185
rect 17064 7095 17098 7117
rect 17064 7023 17098 7049
rect 17064 6965 17098 6981
rect 17150 7967 17184 7983
rect 17150 7899 17184 7925
rect 17150 7831 17184 7853
rect 17150 7763 17184 7781
rect 17150 7695 17184 7709
rect 17150 7627 17184 7637
rect 17150 7559 17184 7565
rect 17150 7491 17184 7493
rect 17150 7455 17184 7457
rect 17150 7383 17184 7389
rect 17150 7311 17184 7321
rect 17150 7239 17184 7253
rect 17150 7167 17184 7185
rect 17150 7095 17184 7117
rect 17150 7023 17184 7049
rect 17270 7966 17280 8020
rect 17314 7966 17330 8020
rect 17270 7950 17330 7966
rect 17270 7886 17280 7950
rect 17314 7886 17330 7950
rect 17270 7880 17330 7886
rect 17270 7846 17280 7880
rect 17314 7846 17330 7880
rect 17270 7840 17330 7846
rect 17270 7776 17280 7840
rect 17314 7776 17330 7840
rect 17270 7760 17330 7776
rect 17270 7706 17280 7760
rect 17314 7706 17330 7760
rect 17270 7680 17330 7706
rect 17270 7636 17280 7680
rect 17314 7636 17330 7680
rect 17270 7600 17330 7636
rect 17270 7566 17280 7600
rect 17314 7566 17330 7600
rect 17270 7530 17330 7566
rect 17270 7486 17280 7530
rect 17314 7486 17330 7530
rect 17270 7460 17330 7486
rect 17270 7406 17280 7460
rect 17314 7406 17330 7460
rect 17270 7390 17330 7406
rect 17270 7326 17280 7390
rect 17314 7326 17330 7390
rect 17270 7320 17330 7326
rect 17270 7286 17280 7320
rect 17314 7286 17330 7320
rect 17270 7280 17330 7286
rect 17270 7216 17280 7280
rect 17314 7216 17330 7280
rect 17270 7200 17330 7216
rect 17270 7146 17280 7200
rect 17314 7146 17330 7200
rect 17270 7120 17330 7146
rect 17270 7076 17280 7120
rect 17314 7076 17330 7120
rect 17270 7040 17330 7076
rect 17270 7006 17280 7040
rect 17314 7006 17330 7040
rect 17270 6990 17330 7006
rect 17498 7930 17578 7950
rect 17498 7850 17518 7890
rect 17498 7770 17518 7810
rect 17498 7690 17518 7730
rect 17498 7610 17518 7650
rect 17498 7530 17518 7570
rect 17498 7450 17518 7490
rect 17498 7370 17518 7410
rect 17498 7290 17518 7330
rect 17498 7210 17518 7250
rect 17498 7130 17518 7170
rect 17498 7050 17518 7090
rect 17498 6990 17518 7010
rect 17558 6990 17578 7930
rect 17150 6965 17184 6981
rect 17498 6970 17578 6990
rect 17622 7908 17656 7942
rect 17622 7836 17656 7874
rect 17622 7764 17656 7802
rect 17622 7692 17656 7730
rect 17622 7620 17656 7658
rect 17622 7548 17656 7586
rect 17622 7476 17656 7514
rect 17622 7404 17656 7442
rect 17622 7332 17656 7370
rect 17622 7260 17656 7298
rect 17622 7188 17656 7226
rect 17622 7116 17656 7154
rect 17622 7044 17656 7082
rect 17622 6972 17656 7010
rect 17708 7908 17742 7942
rect 17708 7836 17742 7874
rect 17708 7764 17742 7802
rect 17708 7692 17742 7730
rect 17708 7620 17742 7658
rect 17708 7548 17742 7586
rect 17708 7476 17742 7514
rect 17708 7404 17742 7442
rect 17708 7332 17742 7370
rect 17708 7260 17742 7298
rect 17708 7188 17742 7226
rect 17708 7116 17742 7154
rect 17708 7044 17742 7082
rect 17708 6972 17742 7010
rect 17794 7908 17828 7942
rect 17794 7836 17828 7874
rect 17794 7764 17828 7802
rect 17794 7692 17828 7730
rect 17794 7620 17828 7658
rect 17794 7548 17828 7586
rect 17794 7476 17828 7514
rect 17794 7404 17828 7442
rect 17794 7332 17828 7370
rect 17794 7260 17828 7298
rect 17794 7188 17828 7226
rect 17794 7116 17828 7154
rect 17794 7044 17828 7082
rect 17794 6972 17828 7010
rect 17880 7908 17914 7942
rect 17880 7836 17914 7874
rect 17880 7764 17914 7802
rect 17880 7692 17914 7730
rect 17880 7620 17914 7658
rect 17880 7548 17914 7586
rect 17880 7476 17914 7514
rect 17880 7404 17914 7442
rect 17880 7332 17914 7370
rect 17880 7260 17914 7298
rect 17880 7188 17914 7226
rect 17880 7116 17914 7154
rect 17880 7044 17914 7082
rect 17880 6972 17914 7010
rect 17966 7908 18000 7942
rect 17966 7836 18000 7874
rect 17966 7764 18000 7802
rect 17966 7692 18000 7730
rect 17966 7620 18000 7658
rect 17966 7548 18000 7586
rect 17966 7476 18000 7514
rect 17966 7404 18000 7442
rect 17966 7332 18000 7370
rect 17966 7260 18000 7298
rect 17966 7188 18000 7226
rect 17966 7116 18000 7154
rect 17966 7044 18000 7082
rect 17966 6972 18000 7010
rect 18052 7908 18086 7942
rect 18052 7836 18086 7874
rect 18052 7764 18086 7802
rect 18052 7692 18086 7730
rect 18052 7620 18086 7658
rect 18052 7548 18086 7586
rect 18052 7476 18086 7514
rect 18052 7404 18086 7442
rect 18052 7332 18086 7370
rect 18052 7260 18086 7298
rect 18052 7188 18086 7226
rect 18052 7116 18086 7154
rect 18052 7044 18086 7082
rect 18052 6972 18086 7010
rect 18138 7908 18172 7942
rect 18138 7836 18172 7874
rect 18138 7764 18172 7802
rect 18138 7692 18172 7730
rect 18138 7620 18172 7658
rect 18138 7548 18172 7586
rect 18138 7476 18172 7514
rect 18138 7404 18172 7442
rect 18138 7332 18172 7370
rect 18138 7260 18172 7298
rect 18138 7188 18172 7226
rect 18138 7116 18172 7154
rect 18138 7044 18172 7082
rect 18138 6972 18172 7010
rect 18224 7908 18258 7942
rect 18224 7836 18258 7874
rect 18224 7764 18258 7802
rect 18224 7692 18258 7730
rect 18224 7620 18258 7658
rect 18224 7548 18258 7586
rect 18224 7476 18258 7514
rect 18224 7404 18258 7442
rect 18224 7332 18258 7370
rect 18224 7260 18258 7298
rect 18224 7188 18258 7226
rect 18224 7116 18258 7154
rect 18224 7044 18258 7082
rect 18224 6972 18258 7010
rect 18310 7908 18344 7942
rect 18310 7836 18344 7874
rect 18310 7764 18344 7802
rect 18310 7692 18344 7730
rect 18310 7620 18344 7658
rect 18310 7548 18344 7586
rect 18310 7476 18344 7514
rect 18310 7404 18344 7442
rect 18310 7332 18344 7370
rect 18310 7260 18344 7298
rect 18310 7188 18344 7226
rect 18310 7116 18344 7154
rect 18310 7044 18344 7082
rect 18310 6972 18344 7010
rect 18396 7908 18430 7942
rect 18396 7836 18430 7874
rect 18396 7764 18430 7802
rect 18396 7692 18430 7730
rect 18396 7620 18430 7658
rect 18396 7548 18430 7586
rect 18396 7476 18430 7514
rect 18396 7404 18430 7442
rect 18396 7332 18430 7370
rect 18396 7260 18430 7298
rect 18396 7188 18430 7226
rect 18396 7116 18430 7154
rect 18396 7044 18430 7082
rect 18396 6972 18430 7010
rect 18482 7908 18516 7942
rect 18482 7836 18516 7874
rect 18482 7764 18516 7802
rect 18482 7692 18516 7730
rect 18482 7620 18516 7658
rect 18482 7548 18516 7586
rect 18482 7476 18516 7514
rect 18482 7404 18516 7442
rect 18482 7332 18516 7370
rect 18482 7260 18516 7298
rect 18482 7188 18516 7226
rect 18482 7116 18516 7154
rect 18482 7044 18516 7082
rect 18482 6972 18516 7010
rect 18568 7908 18602 7942
rect 18568 7836 18602 7874
rect 18568 7764 18602 7802
rect 18568 7692 18602 7730
rect 18568 7620 18602 7658
rect 18568 7548 18602 7586
rect 18568 7476 18602 7514
rect 18568 7404 18602 7442
rect 18568 7332 18602 7370
rect 18568 7260 18602 7298
rect 18568 7188 18602 7226
rect 18568 7116 18602 7154
rect 18568 7044 18602 7082
rect 18568 6972 18602 7010
rect 18654 7908 18688 7942
rect 18654 7836 18688 7874
rect 18654 7764 18688 7802
rect 18654 7692 18688 7730
rect 18654 7620 18688 7658
rect 18654 7548 18688 7586
rect 18654 7476 18688 7514
rect 18654 7404 18688 7442
rect 18654 7332 18688 7370
rect 18654 7260 18688 7298
rect 18654 7188 18688 7226
rect 18654 7116 18688 7154
rect 18654 7044 18688 7082
rect 18654 6972 18688 7010
rect 18740 7908 18774 7942
rect 18740 7836 18774 7874
rect 18740 7764 18774 7802
rect 18740 7692 18774 7730
rect 18740 7620 18774 7658
rect 18740 7548 18774 7586
rect 18740 7476 18774 7514
rect 18740 7404 18774 7442
rect 18740 7332 18774 7370
rect 18740 7260 18774 7298
rect 18740 7188 18774 7226
rect 18740 7116 18774 7154
rect 18740 7044 18774 7082
rect 18740 6972 18774 7010
rect 18826 7908 18860 7942
rect 18826 7836 18860 7874
rect 18826 7764 18860 7802
rect 18826 7692 18860 7730
rect 18826 7620 18860 7658
rect 18826 7548 18860 7586
rect 18826 7476 18860 7514
rect 18826 7404 18860 7442
rect 18826 7332 18860 7370
rect 18826 7260 18860 7298
rect 18826 7188 18860 7226
rect 18826 7116 18860 7154
rect 18826 7044 18860 7082
rect 18826 6972 18860 7010
rect 18912 7908 18946 7942
rect 18912 7836 18946 7874
rect 18912 7764 18946 7802
rect 18912 7692 18946 7730
rect 18912 7620 18946 7658
rect 18912 7548 18946 7586
rect 18912 7476 18946 7514
rect 18912 7404 18946 7442
rect 18912 7332 18946 7370
rect 18912 7260 18946 7298
rect 18912 7188 18946 7226
rect 18912 7116 18946 7154
rect 18912 7044 18946 7082
rect 18912 6972 18946 7010
rect 18998 7908 19032 7942
rect 18998 7836 19032 7874
rect 18998 7764 19032 7802
rect 18998 7692 19032 7730
rect 18998 7620 19032 7658
rect 18998 7548 19032 7586
rect 18998 7476 19032 7514
rect 18998 7404 19032 7442
rect 18998 7332 19032 7370
rect 18998 7260 19032 7298
rect 18998 7188 19032 7226
rect 18998 7116 19032 7154
rect 18998 7044 19032 7082
rect 18998 6972 19032 7010
rect 19084 7908 19118 7942
rect 19084 7836 19118 7874
rect 19084 7764 19118 7802
rect 19084 7692 19118 7730
rect 19084 7620 19118 7658
rect 19084 7548 19118 7586
rect 19084 7476 19118 7514
rect 19084 7404 19118 7442
rect 19084 7332 19118 7370
rect 19084 7260 19118 7298
rect 19084 7188 19118 7226
rect 19084 7116 19118 7154
rect 19084 7044 19118 7082
rect 19084 6972 19118 7010
rect 19170 7908 19204 7942
rect 19170 7836 19204 7874
rect 19170 7764 19204 7802
rect 19170 7692 19204 7730
rect 19170 7620 19204 7658
rect 19170 7548 19204 7586
rect 19170 7476 19204 7514
rect 19170 7404 19204 7442
rect 19170 7332 19204 7370
rect 19170 7260 19204 7298
rect 19170 7188 19204 7226
rect 19170 7116 19204 7154
rect 19170 7044 19204 7082
rect 19170 6972 19204 7010
rect 19256 7908 19290 7942
rect 19256 7836 19290 7874
rect 19256 7764 19290 7802
rect 19256 7692 19290 7730
rect 19256 7620 19290 7658
rect 19256 7548 19290 7586
rect 19256 7476 19290 7514
rect 19256 7404 19290 7442
rect 19256 7332 19290 7370
rect 19256 7260 19290 7298
rect 19256 7188 19290 7226
rect 19256 7116 19290 7154
rect 19256 7044 19290 7082
rect 19256 6972 19290 7010
rect 19342 7908 19376 7942
rect 19342 7836 19376 7874
rect 19342 7764 19376 7802
rect 19342 7692 19376 7730
rect 19342 7620 19376 7658
rect 19342 7548 19376 7586
rect 19342 7476 19376 7514
rect 19342 7404 19376 7442
rect 19342 7332 19376 7370
rect 19342 7260 19376 7298
rect 19342 7188 19376 7226
rect 19342 7116 19376 7154
rect 19342 7044 19376 7082
rect 19342 6972 19376 7010
rect 19428 7908 19462 7942
rect 19428 7836 19462 7874
rect 19428 7764 19462 7802
rect 19428 7692 19462 7730
rect 19428 7620 19462 7658
rect 19428 7548 19462 7586
rect 19428 7476 19462 7514
rect 19428 7404 19462 7442
rect 19428 7332 19462 7370
rect 19428 7260 19462 7298
rect 19428 7188 19462 7226
rect 19428 7116 19462 7154
rect 19428 7044 19462 7082
rect 19428 6972 19462 7010
rect 19514 7908 19548 7942
rect 19514 7836 19548 7874
rect 19514 7764 19548 7802
rect 19514 7692 19548 7730
rect 19514 7620 19548 7658
rect 19514 7548 19548 7586
rect 19514 7476 19548 7514
rect 19514 7404 19548 7442
rect 19514 7332 19548 7370
rect 19514 7260 19548 7298
rect 19514 7188 19548 7226
rect 19514 7116 19548 7154
rect 19514 7044 19548 7082
rect 19514 6972 19548 7010
rect 19600 7908 19634 7942
rect 19600 7836 19634 7874
rect 19600 7764 19634 7802
rect 19600 7692 19634 7730
rect 19600 7620 19634 7658
rect 19600 7548 19634 7586
rect 19600 7476 19634 7514
rect 19600 7404 19634 7442
rect 19600 7332 19634 7370
rect 19600 7260 19634 7298
rect 19600 7188 19634 7226
rect 19600 7116 19634 7154
rect 19600 7044 19634 7082
rect 19600 6972 19634 7010
rect 19686 7908 19720 7942
rect 19686 7836 19720 7874
rect 19686 7764 19720 7802
rect 19686 7692 19720 7730
rect 19686 7620 19720 7658
rect 19686 7548 19720 7586
rect 19686 7476 19720 7514
rect 19686 7404 19720 7442
rect 19686 7332 19720 7370
rect 19686 7260 19720 7298
rect 19686 7188 19720 7226
rect 19686 7116 19720 7154
rect 19686 7044 19720 7082
rect 19686 6972 19720 7010
rect 19772 7908 19806 7942
rect 19772 7836 19806 7874
rect 19772 7764 19806 7802
rect 19772 7692 19806 7730
rect 19772 7620 19806 7658
rect 19772 7548 19806 7586
rect 19772 7476 19806 7514
rect 19772 7404 19806 7442
rect 19772 7332 19806 7370
rect 19772 7260 19806 7298
rect 19772 7188 19806 7226
rect 19772 7116 19806 7154
rect 19772 7044 19806 7082
rect 19772 6972 19806 7010
rect 19858 7908 19892 7942
rect 19858 7836 19892 7874
rect 19858 7764 19892 7802
rect 19858 7692 19892 7730
rect 19858 7620 19892 7658
rect 19858 7548 19892 7586
rect 19858 7476 19892 7514
rect 19858 7404 19892 7442
rect 19858 7332 19892 7370
rect 19858 7260 19892 7298
rect 19858 7188 19892 7226
rect 19858 7116 19892 7154
rect 19858 7044 19892 7082
rect 19858 6972 19892 7010
rect 19944 7908 19978 7942
rect 19944 7836 19978 7874
rect 19944 7764 19978 7802
rect 19944 7692 19978 7730
rect 19944 7620 19978 7658
rect 19944 7548 19978 7586
rect 19944 7476 19978 7514
rect 19944 7404 19978 7442
rect 19944 7332 19978 7370
rect 19944 7260 19978 7298
rect 19944 7188 19978 7226
rect 19944 7116 19978 7154
rect 19944 7044 19978 7082
rect 19944 6972 19978 7010
rect 20030 7908 20064 7942
rect 20030 7836 20064 7874
rect 20030 7764 20064 7802
rect 20030 7692 20064 7730
rect 20030 7620 20064 7658
rect 20030 7548 20064 7586
rect 20030 7476 20064 7514
rect 20030 7404 20064 7442
rect 20030 7332 20064 7370
rect 20030 7260 20064 7298
rect 20030 7188 20064 7226
rect 20030 7116 20064 7154
rect 20030 7044 20064 7082
rect 20030 6972 20064 7010
rect 20118 7930 20198 7950
rect 20118 6990 20138 7930
rect 20178 7850 20198 7890
rect 20178 7770 20198 7810
rect 20178 7690 20198 7730
rect 20178 7610 20198 7650
rect 20178 7530 20198 7570
rect 20178 7450 20198 7490
rect 20178 7370 20198 7410
rect 20178 7290 20198 7330
rect 20178 7210 20198 7250
rect 20178 7130 20198 7170
rect 20178 7050 20198 7090
rect 20178 6990 20198 7010
rect 20118 6970 20198 6990
rect 11805 6896 11813 6930
rect 11855 6896 11885 6930
rect 11923 6896 11957 6930
rect 11991 6896 12025 6930
rect 12063 6896 12093 6930
rect 12135 6896 12143 6930
rect 12371 6896 12379 6930
rect 12421 6896 12451 6930
rect 12489 6896 12523 6930
rect 12557 6896 12591 6930
rect 12629 6896 12659 6930
rect 12701 6896 12709 6930
rect 12937 6896 12945 6930
rect 12987 6896 13017 6930
rect 13055 6896 13089 6930
rect 13123 6896 13157 6930
rect 13195 6896 13225 6930
rect 13267 6896 13275 6930
rect 13503 6896 13511 6930
rect 13553 6896 13583 6930
rect 13621 6896 13655 6930
rect 13689 6896 13723 6930
rect 13761 6896 13791 6930
rect 13833 6896 13841 6930
rect 14069 6896 14077 6930
rect 14119 6896 14149 6930
rect 14187 6896 14221 6930
rect 14255 6896 14289 6930
rect 14327 6896 14357 6930
rect 14399 6896 14407 6930
rect 14635 6896 14643 6930
rect 14685 6896 14715 6930
rect 14753 6896 14787 6930
rect 14821 6896 14855 6930
rect 14893 6896 14923 6930
rect 14965 6896 14973 6930
rect 15201 6896 15209 6930
rect 15251 6896 15281 6930
rect 15319 6896 15353 6930
rect 15387 6896 15421 6930
rect 15459 6896 15489 6930
rect 15531 6896 15539 6930
rect 16138 6897 16154 6931
rect 16188 6897 16218 6931
rect 16256 6897 16290 6931
rect 16324 6897 16358 6931
rect 16396 6897 16426 6931
rect 16460 6897 16494 6931
rect 16528 6897 16562 6931
rect 16600 6897 16634 6931
rect 16668 6897 16702 6931
rect 16740 6897 16770 6931
rect 16804 6897 16838 6931
rect 16872 6897 16906 6931
rect 16944 6897 16978 6931
rect 17012 6897 17046 6931
rect 17084 6897 17184 6931
rect 17676 6908 17946 6926
rect 17676 6874 17686 6908
rect 17726 6874 17758 6908
rect 17794 6874 17828 6908
rect 17864 6874 17896 6908
rect 17936 6874 17946 6908
rect 11785 6846 11819 6862
rect 11674 6766 11708 6778
rect 11674 6694 11708 6710
rect 11674 6622 11708 6642
rect 11674 6550 11708 6574
rect 11674 6478 11708 6506
rect 11674 6406 11708 6438
rect 11674 6336 11708 6370
rect 11674 6268 11708 6300
rect 11674 6200 11708 6228
rect 11674 6132 11708 6156
rect 11674 6064 11708 6084
rect 11674 5996 11708 6012
rect 11674 5928 11708 5940
rect 11785 6778 11819 6804
rect 11785 6710 11819 6732
rect 11785 6642 11819 6660
rect 11785 6574 11819 6588
rect 11785 6506 11819 6516
rect 11785 6438 11819 6444
rect 11785 6370 11819 6372
rect 11785 6334 11819 6336
rect 11785 6262 11819 6268
rect 11785 6190 11819 6200
rect 11785 6118 11819 6132
rect 11785 6046 11819 6064
rect 11785 5974 11819 5996
rect 11785 5902 11819 5928
rect 11785 5844 11819 5860
rect 11871 6846 11905 6862
rect 11871 6778 11905 6804
rect 11871 6710 11905 6732
rect 11871 6642 11905 6660
rect 11871 6574 11905 6588
rect 11871 6506 11905 6516
rect 11871 6438 11905 6444
rect 11871 6370 11905 6372
rect 11871 6334 11905 6336
rect 11871 6262 11905 6268
rect 11871 6190 11905 6200
rect 11871 6118 11905 6132
rect 11871 6046 11905 6064
rect 11871 5974 11905 5996
rect 11871 5902 11905 5928
rect 11871 5844 11905 5860
rect 11957 6846 11991 6862
rect 11957 6778 11991 6804
rect 11957 6710 11991 6732
rect 11957 6642 11991 6660
rect 11957 6574 11991 6588
rect 11957 6506 11991 6516
rect 11957 6438 11991 6444
rect 11957 6370 11991 6372
rect 11957 6334 11991 6336
rect 11957 6262 11991 6268
rect 11957 6190 11991 6200
rect 11957 6118 11991 6132
rect 11957 6046 11991 6064
rect 11957 5974 11991 5996
rect 11957 5902 11991 5928
rect 11957 5844 11991 5860
rect 12043 6846 12077 6862
rect 12043 6778 12077 6804
rect 12043 6710 12077 6732
rect 12043 6642 12077 6660
rect 12043 6574 12077 6588
rect 12043 6506 12077 6516
rect 12043 6438 12077 6444
rect 12043 6370 12077 6372
rect 12043 6334 12077 6336
rect 12043 6262 12077 6268
rect 12043 6190 12077 6200
rect 12043 6118 12077 6132
rect 12043 6046 12077 6064
rect 12043 5974 12077 5996
rect 12043 5902 12077 5928
rect 12043 5844 12077 5860
rect 12129 6846 12163 6862
rect 12351 6846 12385 6862
rect 12129 6778 12163 6804
rect 12129 6710 12163 6732
rect 12129 6642 12163 6660
rect 12129 6574 12163 6588
rect 12129 6506 12163 6516
rect 12129 6438 12163 6444
rect 12129 6370 12163 6372
rect 12129 6334 12163 6336
rect 12129 6262 12163 6268
rect 12129 6190 12163 6200
rect 12129 6118 12163 6132
rect 12129 6046 12163 6064
rect 12129 5974 12163 5996
rect 12129 5902 12163 5928
rect 12240 6766 12274 6778
rect 12240 6694 12274 6710
rect 12240 6622 12274 6642
rect 12240 6550 12274 6574
rect 12240 6478 12274 6506
rect 12240 6406 12274 6438
rect 12240 6336 12274 6370
rect 12240 6268 12274 6300
rect 12240 6200 12274 6228
rect 12240 6132 12274 6156
rect 12240 6064 12274 6084
rect 12240 5996 12274 6012
rect 12240 5928 12274 5940
rect 12351 6778 12385 6804
rect 12351 6710 12385 6732
rect 12351 6642 12385 6660
rect 12351 6574 12385 6588
rect 12351 6506 12385 6516
rect 12351 6438 12385 6444
rect 12351 6370 12385 6372
rect 12351 6334 12385 6336
rect 12351 6262 12385 6268
rect 12351 6190 12385 6200
rect 12351 6118 12385 6132
rect 12351 6046 12385 6064
rect 12351 5974 12385 5996
rect 12351 5902 12385 5928
rect 12129 5844 12163 5860
rect 12351 5844 12385 5860
rect 12437 6846 12471 6862
rect 12437 6778 12471 6804
rect 12437 6710 12471 6732
rect 12437 6642 12471 6660
rect 12437 6574 12471 6588
rect 12437 6506 12471 6516
rect 12437 6438 12471 6444
rect 12437 6370 12471 6372
rect 12437 6334 12471 6336
rect 12437 6262 12471 6268
rect 12437 6190 12471 6200
rect 12437 6118 12471 6132
rect 12437 6046 12471 6064
rect 12437 5974 12471 5996
rect 12437 5902 12471 5928
rect 12437 5844 12471 5860
rect 12523 6846 12557 6862
rect 12523 6778 12557 6804
rect 12523 6710 12557 6732
rect 12523 6642 12557 6660
rect 12523 6574 12557 6588
rect 12523 6506 12557 6516
rect 12523 6438 12557 6444
rect 12523 6370 12557 6372
rect 12523 6334 12557 6336
rect 12523 6262 12557 6268
rect 12523 6190 12557 6200
rect 12523 6118 12557 6132
rect 12523 6046 12557 6064
rect 12523 5974 12557 5996
rect 12523 5902 12557 5928
rect 12523 5844 12557 5860
rect 12609 6846 12643 6862
rect 12609 6778 12643 6804
rect 12609 6710 12643 6732
rect 12609 6642 12643 6660
rect 12609 6574 12643 6588
rect 12609 6506 12643 6516
rect 12609 6438 12643 6444
rect 12609 6370 12643 6372
rect 12609 6334 12643 6336
rect 12609 6262 12643 6268
rect 12609 6190 12643 6200
rect 12609 6118 12643 6132
rect 12609 6046 12643 6064
rect 12609 5974 12643 5996
rect 12609 5902 12643 5928
rect 12609 5844 12643 5860
rect 12695 6846 12729 6862
rect 12917 6846 12951 6862
rect 12695 6778 12729 6804
rect 12695 6710 12729 6732
rect 12695 6642 12729 6660
rect 12695 6574 12729 6588
rect 12695 6506 12729 6516
rect 12695 6438 12729 6444
rect 12695 6370 12729 6372
rect 12695 6334 12729 6336
rect 12695 6262 12729 6268
rect 12695 6190 12729 6200
rect 12695 6118 12729 6132
rect 12695 6046 12729 6064
rect 12695 5974 12729 5996
rect 12695 5902 12729 5928
rect 12806 6766 12840 6778
rect 12806 6694 12840 6710
rect 12806 6622 12840 6642
rect 12806 6550 12840 6574
rect 12806 6478 12840 6506
rect 12806 6406 12840 6438
rect 12806 6336 12840 6370
rect 12806 6268 12840 6300
rect 12806 6200 12840 6228
rect 12806 6132 12840 6156
rect 12806 6064 12840 6084
rect 12806 5996 12840 6012
rect 12806 5928 12840 5940
rect 12917 6778 12951 6804
rect 12917 6710 12951 6732
rect 12917 6642 12951 6660
rect 12917 6574 12951 6588
rect 12917 6506 12951 6516
rect 12917 6438 12951 6444
rect 12917 6370 12951 6372
rect 12917 6334 12951 6336
rect 12917 6262 12951 6268
rect 12917 6190 12951 6200
rect 12917 6118 12951 6132
rect 12917 6046 12951 6064
rect 12917 5974 12951 5996
rect 12917 5902 12951 5928
rect 12695 5844 12729 5860
rect 12917 5844 12951 5860
rect 13003 6846 13037 6862
rect 13003 6778 13037 6804
rect 13003 6710 13037 6732
rect 13003 6642 13037 6660
rect 13003 6574 13037 6588
rect 13003 6506 13037 6516
rect 13003 6438 13037 6444
rect 13003 6370 13037 6372
rect 13003 6334 13037 6336
rect 13003 6262 13037 6268
rect 13003 6190 13037 6200
rect 13003 6118 13037 6132
rect 13003 6046 13037 6064
rect 13003 5974 13037 5996
rect 13003 5902 13037 5928
rect 13003 5844 13037 5860
rect 13089 6846 13123 6862
rect 13089 6778 13123 6804
rect 13089 6710 13123 6732
rect 13089 6642 13123 6660
rect 13089 6574 13123 6588
rect 13089 6506 13123 6516
rect 13089 6438 13123 6444
rect 13089 6370 13123 6372
rect 13089 6334 13123 6336
rect 13089 6262 13123 6268
rect 13089 6190 13123 6200
rect 13089 6118 13123 6132
rect 13089 6046 13123 6064
rect 13089 5974 13123 5996
rect 13089 5902 13123 5928
rect 13089 5844 13123 5860
rect 13175 6846 13209 6862
rect 13175 6778 13209 6804
rect 13175 6710 13209 6732
rect 13175 6642 13209 6660
rect 13175 6574 13209 6588
rect 13175 6506 13209 6516
rect 13175 6438 13209 6444
rect 13175 6370 13209 6372
rect 13175 6334 13209 6336
rect 13175 6262 13209 6268
rect 13175 6190 13209 6200
rect 13175 6118 13209 6132
rect 13175 6046 13209 6064
rect 13175 5974 13209 5996
rect 13175 5902 13209 5928
rect 13175 5844 13209 5860
rect 13261 6846 13295 6862
rect 13483 6846 13517 6862
rect 13261 6778 13295 6804
rect 13261 6710 13295 6732
rect 13261 6642 13295 6660
rect 13261 6574 13295 6588
rect 13261 6506 13295 6516
rect 13261 6438 13295 6444
rect 13261 6370 13295 6372
rect 13261 6334 13295 6336
rect 13261 6262 13295 6268
rect 13261 6190 13295 6200
rect 13261 6118 13295 6132
rect 13261 6046 13295 6064
rect 13261 5974 13295 5996
rect 13261 5902 13295 5928
rect 13372 6766 13406 6778
rect 13372 6694 13406 6710
rect 13372 6622 13406 6642
rect 13372 6550 13406 6574
rect 13372 6478 13406 6506
rect 13372 6406 13406 6438
rect 13372 6336 13406 6370
rect 13372 6268 13406 6300
rect 13372 6200 13406 6228
rect 13372 6132 13406 6156
rect 13372 6064 13406 6084
rect 13372 5996 13406 6012
rect 13372 5928 13406 5940
rect 13483 6778 13517 6804
rect 13483 6710 13517 6732
rect 13483 6642 13517 6660
rect 13483 6574 13517 6588
rect 13483 6506 13517 6516
rect 13483 6438 13517 6444
rect 13483 6370 13517 6372
rect 13483 6334 13517 6336
rect 13483 6262 13517 6268
rect 13483 6190 13517 6200
rect 13483 6118 13517 6132
rect 13483 6046 13517 6064
rect 13483 5974 13517 5996
rect 13483 5902 13517 5928
rect 13261 5844 13295 5860
rect 13483 5844 13517 5860
rect 13569 6846 13603 6862
rect 13569 6778 13603 6804
rect 13569 6710 13603 6732
rect 13569 6642 13603 6660
rect 13569 6574 13603 6588
rect 13569 6506 13603 6516
rect 13569 6438 13603 6444
rect 13569 6370 13603 6372
rect 13569 6334 13603 6336
rect 13569 6262 13603 6268
rect 13569 6190 13603 6200
rect 13569 6118 13603 6132
rect 13569 6046 13603 6064
rect 13569 5974 13603 5996
rect 13569 5902 13603 5928
rect 13569 5844 13603 5860
rect 13655 6846 13689 6862
rect 13655 6778 13689 6804
rect 13655 6710 13689 6732
rect 13655 6642 13689 6660
rect 13655 6574 13689 6588
rect 13655 6506 13689 6516
rect 13655 6438 13689 6444
rect 13655 6370 13689 6372
rect 13655 6334 13689 6336
rect 13655 6262 13689 6268
rect 13655 6190 13689 6200
rect 13655 6118 13689 6132
rect 13655 6046 13689 6064
rect 13655 5974 13689 5996
rect 13655 5902 13689 5928
rect 13655 5844 13689 5860
rect 13741 6846 13775 6862
rect 13741 6778 13775 6804
rect 13741 6710 13775 6732
rect 13741 6642 13775 6660
rect 13741 6574 13775 6588
rect 13741 6506 13775 6516
rect 13741 6438 13775 6444
rect 13741 6370 13775 6372
rect 13741 6334 13775 6336
rect 13741 6262 13775 6268
rect 13741 6190 13775 6200
rect 13741 6118 13775 6132
rect 13741 6046 13775 6064
rect 13741 5974 13775 5996
rect 13741 5902 13775 5928
rect 13741 5844 13775 5860
rect 13827 6846 13861 6862
rect 14049 6846 14083 6862
rect 13827 6778 13861 6804
rect 13827 6710 13861 6732
rect 13827 6642 13861 6660
rect 13827 6574 13861 6588
rect 13827 6506 13861 6516
rect 13827 6438 13861 6444
rect 13827 6370 13861 6372
rect 13827 6334 13861 6336
rect 13827 6262 13861 6268
rect 13827 6190 13861 6200
rect 13827 6118 13861 6132
rect 13827 6046 13861 6064
rect 13827 5974 13861 5996
rect 13827 5902 13861 5928
rect 13938 6766 13972 6778
rect 13938 6694 13972 6710
rect 13938 6622 13972 6642
rect 13938 6550 13972 6574
rect 13938 6478 13972 6506
rect 13938 6406 13972 6438
rect 13938 6336 13972 6370
rect 13938 6268 13972 6300
rect 13938 6200 13972 6228
rect 13938 6132 13972 6156
rect 13938 6064 13972 6084
rect 13938 5996 13972 6012
rect 13938 5928 13972 5940
rect 14049 6778 14083 6804
rect 14049 6710 14083 6732
rect 14049 6642 14083 6660
rect 14049 6574 14083 6588
rect 14049 6506 14083 6516
rect 14049 6438 14083 6444
rect 14049 6370 14083 6372
rect 14049 6334 14083 6336
rect 14049 6262 14083 6268
rect 14049 6190 14083 6200
rect 14049 6118 14083 6132
rect 14049 6046 14083 6064
rect 14049 5974 14083 5996
rect 14049 5902 14083 5928
rect 13827 5844 13861 5860
rect 14049 5844 14083 5860
rect 14135 6846 14169 6862
rect 14135 6778 14169 6804
rect 14135 6710 14169 6732
rect 14135 6642 14169 6660
rect 14135 6574 14169 6588
rect 14135 6506 14169 6516
rect 14135 6438 14169 6444
rect 14135 6370 14169 6372
rect 14135 6334 14169 6336
rect 14135 6262 14169 6268
rect 14135 6190 14169 6200
rect 14135 6118 14169 6132
rect 14135 6046 14169 6064
rect 14135 5974 14169 5996
rect 14135 5902 14169 5928
rect 14135 5844 14169 5860
rect 14221 6846 14255 6862
rect 14221 6778 14255 6804
rect 14221 6710 14255 6732
rect 14221 6642 14255 6660
rect 14221 6574 14255 6588
rect 14221 6506 14255 6516
rect 14221 6438 14255 6444
rect 14221 6370 14255 6372
rect 14221 6334 14255 6336
rect 14221 6262 14255 6268
rect 14221 6190 14255 6200
rect 14221 6118 14255 6132
rect 14221 6046 14255 6064
rect 14221 5974 14255 5996
rect 14221 5902 14255 5928
rect 14221 5844 14255 5860
rect 14307 6846 14341 6862
rect 14307 6778 14341 6804
rect 14307 6710 14341 6732
rect 14307 6642 14341 6660
rect 14307 6574 14341 6588
rect 14307 6506 14341 6516
rect 14307 6438 14341 6444
rect 14307 6370 14341 6372
rect 14307 6334 14341 6336
rect 14307 6262 14341 6268
rect 14307 6190 14341 6200
rect 14307 6118 14341 6132
rect 14307 6046 14341 6064
rect 14307 5974 14341 5996
rect 14307 5902 14341 5928
rect 14307 5844 14341 5860
rect 14393 6846 14427 6862
rect 14615 6846 14649 6862
rect 14393 6778 14427 6804
rect 14393 6710 14427 6732
rect 14393 6642 14427 6660
rect 14393 6574 14427 6588
rect 14393 6506 14427 6516
rect 14393 6438 14427 6444
rect 14393 6370 14427 6372
rect 14393 6334 14427 6336
rect 14393 6262 14427 6268
rect 14393 6190 14427 6200
rect 14393 6118 14427 6132
rect 14393 6046 14427 6064
rect 14393 5974 14427 5996
rect 14393 5902 14427 5928
rect 14504 6766 14538 6778
rect 14504 6694 14538 6710
rect 14504 6622 14538 6642
rect 14504 6550 14538 6574
rect 14504 6478 14538 6506
rect 14504 6406 14538 6438
rect 14504 6336 14538 6370
rect 14504 6268 14538 6300
rect 14504 6200 14538 6228
rect 14504 6132 14538 6156
rect 14504 6064 14538 6084
rect 14504 5996 14538 6012
rect 14504 5928 14538 5940
rect 14615 6778 14649 6804
rect 14615 6710 14649 6732
rect 14615 6642 14649 6660
rect 14615 6574 14649 6588
rect 14615 6506 14649 6516
rect 14615 6438 14649 6444
rect 14615 6370 14649 6372
rect 14615 6334 14649 6336
rect 14615 6262 14649 6268
rect 14615 6190 14649 6200
rect 14615 6118 14649 6132
rect 14615 6046 14649 6064
rect 14615 5974 14649 5996
rect 14615 5902 14649 5928
rect 14393 5844 14427 5860
rect 14615 5844 14649 5860
rect 14701 6846 14735 6862
rect 14701 6778 14735 6804
rect 14701 6710 14735 6732
rect 14701 6642 14735 6660
rect 14701 6574 14735 6588
rect 14701 6506 14735 6516
rect 14701 6438 14735 6444
rect 14701 6370 14735 6372
rect 14701 6334 14735 6336
rect 14701 6262 14735 6268
rect 14701 6190 14735 6200
rect 14701 6118 14735 6132
rect 14701 6046 14735 6064
rect 14701 5974 14735 5996
rect 14701 5902 14735 5928
rect 14701 5844 14735 5860
rect 14787 6846 14821 6862
rect 14787 6778 14821 6804
rect 14787 6710 14821 6732
rect 14787 6642 14821 6660
rect 14787 6574 14821 6588
rect 14787 6506 14821 6516
rect 14787 6438 14821 6444
rect 14787 6370 14821 6372
rect 14787 6334 14821 6336
rect 14787 6262 14821 6268
rect 14787 6190 14821 6200
rect 14787 6118 14821 6132
rect 14787 6046 14821 6064
rect 14787 5974 14821 5996
rect 14787 5902 14821 5928
rect 14787 5844 14821 5860
rect 14873 6846 14907 6862
rect 14873 6778 14907 6804
rect 14873 6710 14907 6732
rect 14873 6642 14907 6660
rect 14873 6574 14907 6588
rect 14873 6506 14907 6516
rect 14873 6438 14907 6444
rect 14873 6370 14907 6372
rect 14873 6334 14907 6336
rect 14873 6262 14907 6268
rect 14873 6190 14907 6200
rect 14873 6118 14907 6132
rect 14873 6046 14907 6064
rect 14873 5974 14907 5996
rect 14873 5902 14907 5928
rect 14873 5844 14907 5860
rect 14959 6846 14993 6862
rect 15181 6846 15215 6862
rect 14959 6778 14993 6804
rect 14959 6710 14993 6732
rect 14959 6642 14993 6660
rect 14959 6574 14993 6588
rect 14959 6506 14993 6516
rect 14959 6438 14993 6444
rect 14959 6370 14993 6372
rect 14959 6334 14993 6336
rect 14959 6262 14993 6268
rect 14959 6190 14993 6200
rect 14959 6118 14993 6132
rect 14959 6046 14993 6064
rect 14959 5974 14993 5996
rect 14959 5902 14993 5928
rect 15070 6766 15104 6778
rect 15070 6694 15104 6710
rect 15070 6622 15104 6642
rect 15070 6550 15104 6574
rect 15070 6478 15104 6506
rect 15070 6406 15104 6438
rect 15070 6336 15104 6370
rect 15070 6268 15104 6300
rect 15070 6200 15104 6228
rect 15070 6132 15104 6156
rect 15070 6064 15104 6084
rect 15070 5996 15104 6012
rect 15070 5928 15104 5940
rect 15181 6778 15215 6804
rect 15181 6710 15215 6732
rect 15181 6642 15215 6660
rect 15181 6574 15215 6588
rect 15181 6506 15215 6516
rect 15181 6438 15215 6444
rect 15181 6370 15215 6372
rect 15181 6334 15215 6336
rect 15181 6262 15215 6268
rect 15181 6190 15215 6200
rect 15181 6118 15215 6132
rect 15181 6046 15215 6064
rect 15181 5974 15215 5996
rect 15181 5902 15215 5928
rect 14959 5844 14993 5860
rect 15181 5844 15215 5860
rect 15267 6846 15301 6862
rect 15267 6778 15301 6804
rect 15267 6710 15301 6732
rect 15267 6642 15301 6660
rect 15267 6574 15301 6588
rect 15267 6506 15301 6516
rect 15267 6438 15301 6444
rect 15267 6370 15301 6372
rect 15267 6334 15301 6336
rect 15267 6262 15301 6268
rect 15267 6190 15301 6200
rect 15267 6118 15301 6132
rect 15267 6046 15301 6064
rect 15267 5974 15301 5996
rect 15267 5902 15301 5928
rect 15267 5844 15301 5860
rect 15353 6846 15387 6862
rect 15353 6778 15387 6804
rect 15353 6710 15387 6732
rect 15353 6642 15387 6660
rect 15353 6574 15387 6588
rect 15353 6506 15387 6516
rect 15353 6438 15387 6444
rect 15353 6370 15387 6372
rect 15353 6334 15387 6336
rect 15353 6262 15387 6268
rect 15353 6190 15387 6200
rect 15353 6118 15387 6132
rect 15353 6046 15387 6064
rect 15353 5974 15387 5996
rect 15353 5902 15387 5928
rect 15353 5844 15387 5860
rect 15439 6846 15473 6862
rect 15439 6778 15473 6804
rect 15439 6710 15473 6732
rect 15439 6642 15473 6660
rect 15439 6574 15473 6588
rect 15439 6506 15473 6516
rect 15439 6438 15473 6444
rect 15439 6370 15473 6372
rect 15439 6334 15473 6336
rect 15439 6262 15473 6268
rect 15439 6190 15473 6200
rect 15439 6118 15473 6132
rect 15439 6046 15473 6064
rect 15439 5974 15473 5996
rect 15439 5902 15473 5928
rect 15439 5844 15473 5860
rect 15525 6846 15559 6862
rect 17676 6858 17946 6874
rect 18020 6908 18290 6926
rect 18020 6874 18030 6908
rect 18070 6874 18102 6908
rect 18138 6874 18172 6908
rect 18208 6874 18240 6908
rect 18280 6874 18290 6908
rect 18020 6858 18290 6874
rect 18364 6908 18634 6926
rect 18364 6874 18374 6908
rect 18414 6874 18446 6908
rect 18482 6874 18516 6908
rect 18552 6874 18584 6908
rect 18624 6874 18634 6908
rect 18364 6858 18634 6874
rect 18708 6908 18978 6926
rect 18708 6874 18718 6908
rect 18758 6874 18790 6908
rect 18826 6874 18860 6908
rect 18896 6874 18928 6908
rect 18968 6874 18978 6908
rect 18708 6858 18978 6874
rect 19052 6908 19322 6926
rect 19052 6874 19062 6908
rect 19102 6874 19134 6908
rect 19170 6874 19204 6908
rect 19240 6874 19272 6908
rect 19312 6874 19322 6908
rect 19052 6858 19322 6874
rect 19396 6908 19666 6926
rect 19396 6874 19406 6908
rect 19446 6874 19478 6908
rect 19514 6874 19548 6908
rect 19584 6874 19616 6908
rect 19656 6874 19666 6908
rect 19396 6858 19666 6874
rect 19740 6908 20010 6926
rect 19740 6874 19750 6908
rect 19790 6874 19822 6908
rect 19858 6874 19892 6908
rect 19928 6874 19960 6908
rect 20000 6874 20010 6908
rect 19740 6858 20010 6874
rect 15525 6778 15559 6804
rect 15525 6710 15559 6732
rect 15525 6642 15559 6660
rect 15525 6574 15559 6588
rect 15525 6506 15559 6516
rect 15525 6438 15559 6444
rect 15525 6370 15559 6372
rect 15525 6334 15559 6336
rect 15525 6262 15559 6268
rect 15525 6190 15559 6200
rect 15525 6118 15559 6132
rect 15525 6046 15559 6064
rect 15525 5974 15559 5996
rect 15525 5902 15559 5928
rect 15636 6766 15670 6778
rect 15636 6694 15670 6710
rect 15636 6622 15670 6642
rect 15636 6550 15670 6574
rect 15636 6478 15670 6506
rect 15636 6406 15670 6438
rect 15636 6336 15670 6370
rect 15636 6268 15670 6300
rect 17658 6316 17928 6332
rect 17658 6282 17668 6316
rect 17708 6282 17740 6316
rect 17776 6282 17810 6316
rect 17846 6282 17878 6316
rect 17918 6282 17928 6316
rect 17658 6264 17928 6282
rect 18002 6316 18272 6332
rect 18002 6282 18012 6316
rect 18052 6282 18084 6316
rect 18120 6282 18154 6316
rect 18190 6282 18222 6316
rect 18262 6282 18272 6316
rect 18002 6264 18272 6282
rect 18346 6316 18616 6332
rect 18346 6282 18356 6316
rect 18396 6282 18428 6316
rect 18464 6282 18498 6316
rect 18534 6282 18566 6316
rect 18606 6282 18616 6316
rect 18346 6264 18616 6282
rect 18690 6316 18960 6332
rect 18690 6282 18700 6316
rect 18740 6282 18772 6316
rect 18808 6282 18842 6316
rect 18878 6282 18910 6316
rect 18950 6282 18960 6316
rect 18690 6264 18960 6282
rect 19034 6316 19304 6332
rect 19034 6282 19044 6316
rect 19084 6282 19116 6316
rect 19152 6282 19186 6316
rect 19222 6282 19254 6316
rect 19294 6282 19304 6316
rect 19034 6264 19304 6282
rect 19378 6316 19648 6332
rect 19378 6282 19388 6316
rect 19428 6282 19460 6316
rect 19496 6282 19530 6316
rect 19566 6282 19598 6316
rect 19638 6282 19648 6316
rect 19378 6264 19648 6282
rect 19722 6316 19992 6332
rect 19722 6282 19732 6316
rect 19772 6282 19804 6316
rect 19840 6282 19874 6316
rect 19910 6282 19942 6316
rect 19982 6282 19992 6316
rect 19722 6264 19992 6282
rect 16138 6229 16154 6263
rect 16188 6229 16218 6263
rect 16256 6229 16290 6263
rect 16324 6229 16358 6263
rect 16396 6229 16426 6263
rect 16460 6229 16494 6263
rect 16528 6229 16562 6263
rect 16600 6229 16634 6263
rect 16668 6229 16702 6263
rect 16740 6229 16770 6263
rect 16804 6229 16838 6263
rect 16872 6229 16906 6263
rect 16944 6229 16978 6263
rect 17012 6229 17046 6263
rect 17084 6229 17184 6263
rect 15636 6200 15670 6228
rect 17480 6200 17560 6220
rect 16118 6179 16152 6195
rect 15636 6132 15670 6156
rect 15636 6064 15670 6084
rect 15636 5996 15670 6012
rect 15636 5928 15670 5940
rect 15980 6154 16030 6170
rect 15980 6120 15990 6154
rect 16024 6120 16030 6154
rect 15980 6084 16030 6120
rect 15980 6040 15990 6084
rect 16024 6040 16030 6084
rect 15980 6014 16030 6040
rect 15980 5960 15990 6014
rect 16024 5960 16030 6014
rect 15980 5944 16030 5960
rect 15980 5880 15990 5944
rect 16024 5880 16030 5944
rect 15980 5874 16030 5880
rect 15525 5844 15559 5860
rect 15980 5840 15990 5874
rect 16024 5840 16030 5874
rect 15980 5834 16030 5840
rect 11805 5776 11813 5810
rect 11855 5776 11885 5810
rect 11923 5776 11957 5810
rect 11991 5776 12025 5810
rect 12063 5776 12093 5810
rect 12135 5776 12143 5810
rect 12371 5776 12379 5810
rect 12421 5776 12451 5810
rect 12489 5776 12523 5810
rect 12557 5776 12591 5810
rect 12629 5776 12659 5810
rect 12701 5776 12709 5810
rect 12937 5776 12945 5810
rect 12987 5776 13017 5810
rect 13055 5776 13089 5810
rect 13123 5776 13157 5810
rect 13195 5776 13225 5810
rect 13267 5776 13275 5810
rect 13503 5776 13511 5810
rect 13553 5776 13583 5810
rect 13621 5776 13655 5810
rect 13689 5776 13723 5810
rect 13761 5776 13791 5810
rect 13833 5776 13841 5810
rect 14069 5776 14077 5810
rect 14119 5776 14149 5810
rect 14187 5776 14221 5810
rect 14255 5776 14289 5810
rect 14327 5776 14357 5810
rect 14399 5776 14407 5810
rect 14635 5776 14643 5810
rect 14685 5776 14715 5810
rect 14753 5776 14787 5810
rect 14821 5776 14855 5810
rect 14893 5776 14923 5810
rect 14965 5776 14973 5810
rect 15201 5776 15209 5810
rect 15251 5776 15281 5810
rect 15319 5776 15353 5810
rect 15387 5776 15421 5810
rect 15459 5776 15489 5810
rect 15531 5776 15539 5810
rect 15980 5770 15990 5834
rect 16024 5770 16030 5834
rect 15980 5754 16030 5770
rect 15980 5700 15990 5754
rect 16024 5700 16030 5754
rect 15980 5674 16030 5700
rect 15980 5630 15990 5674
rect 16024 5630 16030 5674
rect 15980 5594 16030 5630
rect 15980 5560 15990 5594
rect 16024 5560 16030 5594
rect 15980 5524 16030 5560
rect 15980 5480 15990 5524
rect 16024 5480 16030 5524
rect 15980 5454 16030 5480
rect 15980 5400 15990 5454
rect 16024 5400 16030 5454
rect 15980 5384 16030 5400
rect 15980 5320 15990 5384
rect 16024 5320 16030 5384
rect 15980 5314 16030 5320
rect 15980 5280 15990 5314
rect 16024 5280 16030 5314
rect 15980 5274 16030 5280
rect 15980 5210 15990 5274
rect 16024 5210 16030 5274
rect 15980 5194 16030 5210
rect 15980 5140 15990 5194
rect 16024 5140 16030 5194
rect 16118 6111 16152 6137
rect 16118 6043 16152 6065
rect 16118 5975 16152 5993
rect 16118 5907 16152 5921
rect 16118 5839 16152 5849
rect 16118 5771 16152 5777
rect 16118 5703 16152 5705
rect 16118 5667 16152 5669
rect 16118 5595 16152 5601
rect 16118 5523 16152 5533
rect 16118 5451 16152 5465
rect 16118 5379 16152 5397
rect 16118 5307 16152 5329
rect 16118 5235 16152 5261
rect 16118 5177 16152 5193
rect 16204 6179 16238 6195
rect 16204 6111 16238 6137
rect 16204 6043 16238 6065
rect 16204 5975 16238 5993
rect 16204 5907 16238 5921
rect 16204 5839 16238 5849
rect 16204 5771 16238 5777
rect 16204 5703 16238 5705
rect 16204 5667 16238 5669
rect 16204 5595 16238 5601
rect 16204 5523 16238 5533
rect 16204 5451 16238 5465
rect 16204 5379 16238 5397
rect 16204 5307 16238 5329
rect 16204 5235 16238 5261
rect 16204 5177 16238 5193
rect 16290 6179 16324 6195
rect 16290 6111 16324 6137
rect 16290 6043 16324 6065
rect 16290 5975 16324 5993
rect 16290 5907 16324 5921
rect 16290 5839 16324 5849
rect 16290 5771 16324 5777
rect 16290 5703 16324 5705
rect 16290 5667 16324 5669
rect 16290 5595 16324 5601
rect 16290 5523 16324 5533
rect 16290 5451 16324 5465
rect 16290 5379 16324 5397
rect 16290 5307 16324 5329
rect 16290 5235 16324 5261
rect 16290 5177 16324 5193
rect 16376 6179 16410 6195
rect 16376 6111 16410 6137
rect 16376 6043 16410 6065
rect 16376 5975 16410 5993
rect 16376 5907 16410 5921
rect 16376 5839 16410 5849
rect 16376 5771 16410 5777
rect 16376 5703 16410 5705
rect 16376 5667 16410 5669
rect 16376 5595 16410 5601
rect 16376 5523 16410 5533
rect 16376 5451 16410 5465
rect 16376 5379 16410 5397
rect 16376 5307 16410 5329
rect 16376 5235 16410 5261
rect 16376 5177 16410 5193
rect 16462 6179 16496 6195
rect 16462 6111 16496 6137
rect 16462 6043 16496 6065
rect 16462 5975 16496 5993
rect 16462 5907 16496 5921
rect 16462 5839 16496 5849
rect 16462 5771 16496 5777
rect 16462 5703 16496 5705
rect 16462 5667 16496 5669
rect 16462 5595 16496 5601
rect 16462 5523 16496 5533
rect 16462 5451 16496 5465
rect 16462 5379 16496 5397
rect 16462 5307 16496 5329
rect 16462 5235 16496 5261
rect 16462 5177 16496 5193
rect 16548 6179 16582 6195
rect 16548 6111 16582 6137
rect 16548 6043 16582 6065
rect 16548 5975 16582 5993
rect 16548 5907 16582 5921
rect 16548 5839 16582 5849
rect 16548 5771 16582 5777
rect 16548 5703 16582 5705
rect 16548 5667 16582 5669
rect 16548 5595 16582 5601
rect 16548 5523 16582 5533
rect 16548 5451 16582 5465
rect 16548 5379 16582 5397
rect 16548 5307 16582 5329
rect 16548 5235 16582 5261
rect 16548 5177 16582 5193
rect 16634 6179 16668 6195
rect 16634 6111 16668 6137
rect 16634 6043 16668 6065
rect 16634 5975 16668 5993
rect 16634 5907 16668 5921
rect 16634 5839 16668 5849
rect 16634 5771 16668 5777
rect 16634 5703 16668 5705
rect 16634 5667 16668 5669
rect 16634 5595 16668 5601
rect 16634 5523 16668 5533
rect 16634 5451 16668 5465
rect 16634 5379 16668 5397
rect 16634 5307 16668 5329
rect 16634 5235 16668 5261
rect 16634 5177 16668 5193
rect 16720 6179 16754 6195
rect 16720 6111 16754 6137
rect 16720 6043 16754 6065
rect 16720 5975 16754 5993
rect 16720 5907 16754 5921
rect 16720 5839 16754 5849
rect 16720 5771 16754 5777
rect 16720 5703 16754 5705
rect 16720 5667 16754 5669
rect 16720 5595 16754 5601
rect 16720 5523 16754 5533
rect 16720 5451 16754 5465
rect 16720 5379 16754 5397
rect 16720 5307 16754 5329
rect 16720 5235 16754 5261
rect 16720 5177 16754 5193
rect 16806 6179 16840 6195
rect 16806 6111 16840 6137
rect 16806 6043 16840 6065
rect 16806 5975 16840 5993
rect 16806 5907 16840 5921
rect 16806 5839 16840 5849
rect 16806 5771 16840 5777
rect 16806 5703 16840 5705
rect 16806 5667 16840 5669
rect 16806 5595 16840 5601
rect 16806 5523 16840 5533
rect 16806 5451 16840 5465
rect 16806 5379 16840 5397
rect 16806 5307 16840 5329
rect 16806 5235 16840 5261
rect 16806 5177 16840 5193
rect 16892 6179 16926 6195
rect 16892 6111 16926 6137
rect 16892 6043 16926 6065
rect 16892 5975 16926 5993
rect 16892 5907 16926 5921
rect 16892 5839 16926 5849
rect 16892 5771 16926 5777
rect 16892 5703 16926 5705
rect 16892 5667 16926 5669
rect 16892 5595 16926 5601
rect 16892 5523 16926 5533
rect 16892 5451 16926 5465
rect 16892 5379 16926 5397
rect 16892 5307 16926 5329
rect 16892 5235 16926 5261
rect 16892 5177 16926 5193
rect 16978 6179 17012 6195
rect 16978 6111 17012 6137
rect 16978 6043 17012 6065
rect 16978 5975 17012 5993
rect 16978 5907 17012 5921
rect 16978 5839 17012 5849
rect 16978 5771 17012 5777
rect 16978 5703 17012 5705
rect 16978 5667 17012 5669
rect 16978 5595 17012 5601
rect 16978 5523 17012 5533
rect 16978 5451 17012 5465
rect 16978 5379 17012 5397
rect 16978 5307 17012 5329
rect 16978 5235 17012 5261
rect 16978 5177 17012 5193
rect 17064 6179 17098 6195
rect 17064 6111 17098 6137
rect 17064 6043 17098 6065
rect 17064 5975 17098 5993
rect 17064 5907 17098 5921
rect 17064 5839 17098 5849
rect 17064 5771 17098 5777
rect 17064 5703 17098 5705
rect 17064 5667 17098 5669
rect 17064 5595 17098 5601
rect 17064 5523 17098 5533
rect 17064 5451 17098 5465
rect 17064 5379 17098 5397
rect 17064 5307 17098 5329
rect 17064 5235 17098 5261
rect 17064 5177 17098 5193
rect 17150 6179 17184 6195
rect 17480 6180 17500 6200
rect 17150 6111 17184 6137
rect 17150 6043 17184 6065
rect 17150 5975 17184 5993
rect 17150 5907 17184 5921
rect 17150 5839 17184 5849
rect 17150 5771 17184 5777
rect 17150 5703 17184 5705
rect 17150 5667 17184 5669
rect 17150 5595 17184 5601
rect 17150 5523 17184 5533
rect 17150 5451 17184 5465
rect 17150 5379 17184 5397
rect 17150 5307 17184 5329
rect 17150 5235 17184 5261
rect 17150 5177 17184 5193
rect 17270 6154 17330 6170
rect 17270 6120 17280 6154
rect 17314 6120 17330 6154
rect 17270 6084 17330 6120
rect 17270 6040 17280 6084
rect 17314 6040 17330 6084
rect 17270 6014 17330 6040
rect 17270 5960 17280 6014
rect 17314 5960 17330 6014
rect 17270 5944 17330 5960
rect 17270 5880 17280 5944
rect 17314 5880 17330 5944
rect 17270 5874 17330 5880
rect 17270 5840 17280 5874
rect 17314 5840 17330 5874
rect 17270 5834 17330 5840
rect 17270 5770 17280 5834
rect 17314 5770 17330 5834
rect 17270 5754 17330 5770
rect 17270 5700 17280 5754
rect 17314 5700 17330 5754
rect 17270 5674 17330 5700
rect 17270 5630 17280 5674
rect 17314 5630 17330 5674
rect 17270 5594 17330 5630
rect 17270 5560 17280 5594
rect 17314 5560 17330 5594
rect 17270 5524 17330 5560
rect 17270 5480 17280 5524
rect 17314 5480 17330 5524
rect 17270 5454 17330 5480
rect 17270 5400 17280 5454
rect 17314 5400 17330 5454
rect 17270 5384 17330 5400
rect 17270 5320 17280 5384
rect 17314 5320 17330 5384
rect 17270 5314 17330 5320
rect 17270 5280 17280 5314
rect 17314 5280 17330 5314
rect 17270 5274 17330 5280
rect 17270 5210 17280 5274
rect 17314 5210 17330 5274
rect 17480 6100 17500 6140
rect 17480 6020 17500 6060
rect 17480 5940 17500 5980
rect 17480 5860 17500 5900
rect 17480 5780 17500 5820
rect 17480 5700 17500 5740
rect 17480 5620 17500 5660
rect 17480 5540 17500 5580
rect 17480 5460 17500 5500
rect 17480 5380 17500 5420
rect 17480 5300 17500 5340
rect 17540 5260 17560 6200
rect 17480 5240 17560 5260
rect 17604 6180 17638 6218
rect 17604 6108 17638 6146
rect 17604 6036 17638 6074
rect 17604 5964 17638 6002
rect 17604 5892 17638 5930
rect 17604 5820 17638 5858
rect 17604 5748 17638 5786
rect 17604 5676 17638 5714
rect 17604 5604 17638 5642
rect 17604 5532 17638 5570
rect 17604 5460 17638 5498
rect 17604 5388 17638 5426
rect 17604 5316 17638 5354
rect 17604 5248 17638 5282
rect 17690 6180 17724 6218
rect 17690 6108 17724 6146
rect 17690 6036 17724 6074
rect 17690 5964 17724 6002
rect 17690 5892 17724 5930
rect 17690 5820 17724 5858
rect 17690 5748 17724 5786
rect 17690 5676 17724 5714
rect 17690 5604 17724 5642
rect 17690 5532 17724 5570
rect 17690 5460 17724 5498
rect 17690 5388 17724 5426
rect 17690 5316 17724 5354
rect 17690 5248 17724 5282
rect 17776 6180 17810 6218
rect 17776 6108 17810 6146
rect 17776 6036 17810 6074
rect 17776 5964 17810 6002
rect 17776 5892 17810 5930
rect 17776 5820 17810 5858
rect 17776 5748 17810 5786
rect 17776 5676 17810 5714
rect 17776 5604 17810 5642
rect 17776 5532 17810 5570
rect 17776 5460 17810 5498
rect 17776 5388 17810 5426
rect 17776 5316 17810 5354
rect 17776 5248 17810 5282
rect 17862 6180 17896 6218
rect 17862 6108 17896 6146
rect 17862 6036 17896 6074
rect 17862 5964 17896 6002
rect 17862 5892 17896 5930
rect 17862 5820 17896 5858
rect 17862 5748 17896 5786
rect 17862 5676 17896 5714
rect 17862 5604 17896 5642
rect 17862 5532 17896 5570
rect 17862 5460 17896 5498
rect 17862 5388 17896 5426
rect 17862 5316 17896 5354
rect 17862 5248 17896 5282
rect 17948 6180 17982 6218
rect 17948 6108 17982 6146
rect 17948 6036 17982 6074
rect 17948 5964 17982 6002
rect 17948 5892 17982 5930
rect 17948 5820 17982 5858
rect 17948 5748 17982 5786
rect 17948 5676 17982 5714
rect 17948 5604 17982 5642
rect 17948 5532 17982 5570
rect 17948 5460 17982 5498
rect 17948 5388 17982 5426
rect 17948 5316 17982 5354
rect 17948 5248 17982 5282
rect 18034 6180 18068 6218
rect 18034 6108 18068 6146
rect 18034 6036 18068 6074
rect 18034 5964 18068 6002
rect 18034 5892 18068 5930
rect 18034 5820 18068 5858
rect 18034 5748 18068 5786
rect 18034 5676 18068 5714
rect 18034 5604 18068 5642
rect 18034 5532 18068 5570
rect 18034 5460 18068 5498
rect 18034 5388 18068 5426
rect 18034 5316 18068 5354
rect 18034 5248 18068 5282
rect 18120 6180 18154 6218
rect 18120 6108 18154 6146
rect 18120 6036 18154 6074
rect 18120 5964 18154 6002
rect 18120 5892 18154 5930
rect 18120 5820 18154 5858
rect 18120 5748 18154 5786
rect 18120 5676 18154 5714
rect 18120 5604 18154 5642
rect 18120 5532 18154 5570
rect 18120 5460 18154 5498
rect 18120 5388 18154 5426
rect 18120 5316 18154 5354
rect 18120 5248 18154 5282
rect 18206 6180 18240 6218
rect 18206 6108 18240 6146
rect 18206 6036 18240 6074
rect 18206 5964 18240 6002
rect 18206 5892 18240 5930
rect 18206 5820 18240 5858
rect 18206 5748 18240 5786
rect 18206 5676 18240 5714
rect 18206 5604 18240 5642
rect 18206 5532 18240 5570
rect 18206 5460 18240 5498
rect 18206 5388 18240 5426
rect 18206 5316 18240 5354
rect 18206 5248 18240 5282
rect 18292 6180 18326 6218
rect 18292 6108 18326 6146
rect 18292 6036 18326 6074
rect 18292 5964 18326 6002
rect 18292 5892 18326 5930
rect 18292 5820 18326 5858
rect 18292 5748 18326 5786
rect 18292 5676 18326 5714
rect 18292 5604 18326 5642
rect 18292 5532 18326 5570
rect 18292 5460 18326 5498
rect 18292 5388 18326 5426
rect 18292 5316 18326 5354
rect 18292 5248 18326 5282
rect 18378 6180 18412 6218
rect 18378 6108 18412 6146
rect 18378 6036 18412 6074
rect 18378 5964 18412 6002
rect 18378 5892 18412 5930
rect 18378 5820 18412 5858
rect 18378 5748 18412 5786
rect 18378 5676 18412 5714
rect 18378 5604 18412 5642
rect 18378 5532 18412 5570
rect 18378 5460 18412 5498
rect 18378 5388 18412 5426
rect 18378 5316 18412 5354
rect 18378 5248 18412 5282
rect 18464 6180 18498 6218
rect 18464 6108 18498 6146
rect 18464 6036 18498 6074
rect 18464 5964 18498 6002
rect 18464 5892 18498 5930
rect 18464 5820 18498 5858
rect 18464 5748 18498 5786
rect 18464 5676 18498 5714
rect 18464 5604 18498 5642
rect 18464 5532 18498 5570
rect 18464 5460 18498 5498
rect 18464 5388 18498 5426
rect 18464 5316 18498 5354
rect 18464 5248 18498 5282
rect 18550 6180 18584 6218
rect 18550 6108 18584 6146
rect 18550 6036 18584 6074
rect 18550 5964 18584 6002
rect 18550 5892 18584 5930
rect 18550 5820 18584 5858
rect 18550 5748 18584 5786
rect 18550 5676 18584 5714
rect 18550 5604 18584 5642
rect 18550 5532 18584 5570
rect 18550 5460 18584 5498
rect 18550 5388 18584 5426
rect 18550 5316 18584 5354
rect 18550 5248 18584 5282
rect 18636 6180 18670 6218
rect 18636 6108 18670 6146
rect 18636 6036 18670 6074
rect 18636 5964 18670 6002
rect 18636 5892 18670 5930
rect 18636 5820 18670 5858
rect 18636 5748 18670 5786
rect 18636 5676 18670 5714
rect 18636 5604 18670 5642
rect 18636 5532 18670 5570
rect 18636 5460 18670 5498
rect 18636 5388 18670 5426
rect 18636 5316 18670 5354
rect 18636 5248 18670 5282
rect 18722 6180 18756 6218
rect 18722 6108 18756 6146
rect 18722 6036 18756 6074
rect 18722 5964 18756 6002
rect 18722 5892 18756 5930
rect 18722 5820 18756 5858
rect 18722 5748 18756 5786
rect 18722 5676 18756 5714
rect 18722 5604 18756 5642
rect 18722 5532 18756 5570
rect 18722 5460 18756 5498
rect 18722 5388 18756 5426
rect 18722 5316 18756 5354
rect 18722 5248 18756 5282
rect 18808 6180 18842 6218
rect 18808 6108 18842 6146
rect 18808 6036 18842 6074
rect 18808 5964 18842 6002
rect 18808 5892 18842 5930
rect 18808 5820 18842 5858
rect 18808 5748 18842 5786
rect 18808 5676 18842 5714
rect 18808 5604 18842 5642
rect 18808 5532 18842 5570
rect 18808 5460 18842 5498
rect 18808 5388 18842 5426
rect 18808 5316 18842 5354
rect 18808 5248 18842 5282
rect 18894 6180 18928 6218
rect 18894 6108 18928 6146
rect 18894 6036 18928 6074
rect 18894 5964 18928 6002
rect 18894 5892 18928 5930
rect 18894 5820 18928 5858
rect 18894 5748 18928 5786
rect 18894 5676 18928 5714
rect 18894 5604 18928 5642
rect 18894 5532 18928 5570
rect 18894 5460 18928 5498
rect 18894 5388 18928 5426
rect 18894 5316 18928 5354
rect 18894 5248 18928 5282
rect 18980 6180 19014 6218
rect 18980 6108 19014 6146
rect 18980 6036 19014 6074
rect 18980 5964 19014 6002
rect 18980 5892 19014 5930
rect 18980 5820 19014 5858
rect 18980 5748 19014 5786
rect 18980 5676 19014 5714
rect 18980 5604 19014 5642
rect 18980 5532 19014 5570
rect 18980 5460 19014 5498
rect 18980 5388 19014 5426
rect 18980 5316 19014 5354
rect 18980 5248 19014 5282
rect 19066 6180 19100 6218
rect 19066 6108 19100 6146
rect 19066 6036 19100 6074
rect 19066 5964 19100 6002
rect 19066 5892 19100 5930
rect 19066 5820 19100 5858
rect 19066 5748 19100 5786
rect 19066 5676 19100 5714
rect 19066 5604 19100 5642
rect 19066 5532 19100 5570
rect 19066 5460 19100 5498
rect 19066 5388 19100 5426
rect 19066 5316 19100 5354
rect 19066 5248 19100 5282
rect 19152 6180 19186 6218
rect 19152 6108 19186 6146
rect 19152 6036 19186 6074
rect 19152 5964 19186 6002
rect 19152 5892 19186 5930
rect 19152 5820 19186 5858
rect 19152 5748 19186 5786
rect 19152 5676 19186 5714
rect 19152 5604 19186 5642
rect 19152 5532 19186 5570
rect 19152 5460 19186 5498
rect 19152 5388 19186 5426
rect 19152 5316 19186 5354
rect 19152 5248 19186 5282
rect 19238 6180 19272 6218
rect 19238 6108 19272 6146
rect 19238 6036 19272 6074
rect 19238 5964 19272 6002
rect 19238 5892 19272 5930
rect 19238 5820 19272 5858
rect 19238 5748 19272 5786
rect 19238 5676 19272 5714
rect 19238 5604 19272 5642
rect 19238 5532 19272 5570
rect 19238 5460 19272 5498
rect 19238 5388 19272 5426
rect 19238 5316 19272 5354
rect 19238 5248 19272 5282
rect 19324 6180 19358 6218
rect 19324 6108 19358 6146
rect 19324 6036 19358 6074
rect 19324 5964 19358 6002
rect 19324 5892 19358 5930
rect 19324 5820 19358 5858
rect 19324 5748 19358 5786
rect 19324 5676 19358 5714
rect 19324 5604 19358 5642
rect 19324 5532 19358 5570
rect 19324 5460 19358 5498
rect 19324 5388 19358 5426
rect 19324 5316 19358 5354
rect 19324 5248 19358 5282
rect 19410 6180 19444 6218
rect 19410 6108 19444 6146
rect 19410 6036 19444 6074
rect 19410 5964 19444 6002
rect 19410 5892 19444 5930
rect 19410 5820 19444 5858
rect 19410 5748 19444 5786
rect 19410 5676 19444 5714
rect 19410 5604 19444 5642
rect 19410 5532 19444 5570
rect 19410 5460 19444 5498
rect 19410 5388 19444 5426
rect 19410 5316 19444 5354
rect 19410 5248 19444 5282
rect 19496 6180 19530 6218
rect 19496 6108 19530 6146
rect 19496 6036 19530 6074
rect 19496 5964 19530 6002
rect 19496 5892 19530 5930
rect 19496 5820 19530 5858
rect 19496 5748 19530 5786
rect 19496 5676 19530 5714
rect 19496 5604 19530 5642
rect 19496 5532 19530 5570
rect 19496 5460 19530 5498
rect 19496 5388 19530 5426
rect 19496 5316 19530 5354
rect 19496 5248 19530 5282
rect 19582 6180 19616 6218
rect 19582 6108 19616 6146
rect 19582 6036 19616 6074
rect 19582 5964 19616 6002
rect 19582 5892 19616 5930
rect 19582 5820 19616 5858
rect 19582 5748 19616 5786
rect 19582 5676 19616 5714
rect 19582 5604 19616 5642
rect 19582 5532 19616 5570
rect 19582 5460 19616 5498
rect 19582 5388 19616 5426
rect 19582 5316 19616 5354
rect 19582 5248 19616 5282
rect 19668 6180 19702 6218
rect 19668 6108 19702 6146
rect 19668 6036 19702 6074
rect 19668 5964 19702 6002
rect 19668 5892 19702 5930
rect 19668 5820 19702 5858
rect 19668 5748 19702 5786
rect 19668 5676 19702 5714
rect 19668 5604 19702 5642
rect 19668 5532 19702 5570
rect 19668 5460 19702 5498
rect 19668 5388 19702 5426
rect 19668 5316 19702 5354
rect 19668 5248 19702 5282
rect 19754 6180 19788 6218
rect 19754 6108 19788 6146
rect 19754 6036 19788 6074
rect 19754 5964 19788 6002
rect 19754 5892 19788 5930
rect 19754 5820 19788 5858
rect 19754 5748 19788 5786
rect 19754 5676 19788 5714
rect 19754 5604 19788 5642
rect 19754 5532 19788 5570
rect 19754 5460 19788 5498
rect 19754 5388 19788 5426
rect 19754 5316 19788 5354
rect 19754 5248 19788 5282
rect 19840 6180 19874 6218
rect 19840 6108 19874 6146
rect 19840 6036 19874 6074
rect 19840 5964 19874 6002
rect 19840 5892 19874 5930
rect 19840 5820 19874 5858
rect 19840 5748 19874 5786
rect 19840 5676 19874 5714
rect 19840 5604 19874 5642
rect 19840 5532 19874 5570
rect 19840 5460 19874 5498
rect 19840 5388 19874 5426
rect 19840 5316 19874 5354
rect 19840 5248 19874 5282
rect 19926 6180 19960 6218
rect 19926 6108 19960 6146
rect 19926 6036 19960 6074
rect 19926 5964 19960 6002
rect 19926 5892 19960 5930
rect 19926 5820 19960 5858
rect 19926 5748 19960 5786
rect 19926 5676 19960 5714
rect 19926 5604 19960 5642
rect 19926 5532 19960 5570
rect 19926 5460 19960 5498
rect 19926 5388 19960 5426
rect 19926 5316 19960 5354
rect 19926 5248 19960 5282
rect 20012 6180 20046 6218
rect 20012 6108 20046 6146
rect 20012 6036 20046 6074
rect 20012 5964 20046 6002
rect 20012 5892 20046 5930
rect 20012 5820 20046 5858
rect 20012 5748 20046 5786
rect 20012 5676 20046 5714
rect 20012 5604 20046 5642
rect 20012 5532 20046 5570
rect 20012 5460 20046 5498
rect 20012 5388 20046 5426
rect 20012 5316 20046 5354
rect 20012 5248 20046 5282
rect 20100 6200 20180 6220
rect 20100 5260 20120 6200
rect 20160 6180 20180 6200
rect 20160 6100 20180 6140
rect 20160 6020 20180 6060
rect 20160 5940 20180 5980
rect 20160 5860 20180 5900
rect 20160 5780 20180 5820
rect 20160 5700 20180 5740
rect 20160 5620 20180 5660
rect 20160 5540 20180 5580
rect 20160 5460 20180 5500
rect 20160 5380 20180 5420
rect 20160 5300 20180 5340
rect 20100 5240 20180 5260
rect 17270 5194 17330 5210
rect 15980 5100 16030 5140
rect 17270 5140 17280 5194
rect 17314 5140 17330 5194
rect 17270 5100 17330 5140
rect 15980 5084 17330 5100
rect 15980 5050 16070 5084
rect 16114 5050 16140 5084
rect 16194 5050 16210 5084
rect 16274 5050 16280 5084
rect 16314 5050 16320 5084
rect 16384 5050 16400 5084
rect 16454 5050 16480 5084
rect 16524 5050 16560 5084
rect 16594 5050 16630 5084
rect 16674 5050 16700 5084
rect 16754 5050 16770 5084
rect 16834 5050 16840 5084
rect 16874 5050 16880 5084
rect 16944 5050 16960 5084
rect 17014 5050 17040 5084
rect 17084 5050 17120 5084
rect 17154 5050 17190 5084
rect 17224 5050 17330 5084
rect 17600 5140 20060 5160
rect 17600 5100 17620 5140
rect 20040 5100 20060 5140
rect 17600 5080 20060 5100
rect 15980 5040 17330 5050
rect 16550 4802 18266 4818
rect 16550 4768 16635 4802
rect 16669 4768 16707 4802
rect 16741 4768 16779 4802
rect 16813 4768 16851 4802
rect 16885 4768 16923 4802
rect 16957 4768 16995 4802
rect 17029 4768 17067 4802
rect 17101 4768 17139 4802
rect 17173 4768 17211 4802
rect 17245 4768 17283 4802
rect 17317 4768 17355 4802
rect 17389 4768 17427 4802
rect 17461 4768 17499 4802
rect 17533 4768 17571 4802
rect 17605 4768 17643 4802
rect 17677 4768 17715 4802
rect 17749 4768 17787 4802
rect 17821 4768 17859 4802
rect 17893 4768 17931 4802
rect 17965 4768 18003 4802
rect 18037 4768 18075 4802
rect 18109 4768 18147 4802
rect 18181 4768 18266 4802
rect 16550 4735 18266 4768
rect 16550 4701 16566 4735
rect 16600 4701 18216 4735
rect 18250 4701 18266 4735
rect 16550 4663 18266 4701
rect 16550 4629 16566 4663
rect 16600 4629 18216 4663
rect 18250 4629 18266 4663
rect 16550 4591 18266 4629
rect 16550 4557 16566 4591
rect 16600 4557 18216 4591
rect 18250 4557 18266 4591
rect 16550 4519 18266 4557
rect 16550 4485 16566 4519
rect 16600 4485 18216 4519
rect 18250 4485 18266 4519
rect 16550 4447 18266 4485
rect 16550 4413 16566 4447
rect 16600 4413 18216 4447
rect 18250 4413 18266 4447
rect 16550 4375 18266 4413
rect 16550 4341 16566 4375
rect 16600 4341 18216 4375
rect 18250 4341 18266 4375
rect 16550 4303 18266 4341
rect 16550 4269 16566 4303
rect 16600 4269 18216 4303
rect 18250 4269 18266 4303
rect 16550 4231 18266 4269
rect 16550 4197 16566 4231
rect 16600 4197 18216 4231
rect 18250 4197 18266 4231
rect 16550 4159 18266 4197
rect 16550 4125 16566 4159
rect 16600 4125 18216 4159
rect 18250 4125 18266 4159
rect 16550 4087 18266 4125
rect 16550 4053 16566 4087
rect 16600 4053 18216 4087
rect 18250 4053 18266 4087
rect 16550 4015 18266 4053
rect 16550 3981 16566 4015
rect 16600 3981 18216 4015
rect 18250 3981 18266 4015
rect 16550 3943 18266 3981
rect 16550 3909 16566 3943
rect 16600 3909 18216 3943
rect 18250 3909 18266 3943
rect 16550 3871 18266 3909
rect 16550 3837 16566 3871
rect 16600 3837 18216 3871
rect 18250 3837 18266 3871
rect 16550 3799 18266 3837
rect 16550 3765 16566 3799
rect 16600 3765 18216 3799
rect 18250 3765 18266 3799
rect 16550 3727 18266 3765
rect 16550 3693 16566 3727
rect 16600 3693 18216 3727
rect 18250 3693 18266 3727
rect 16550 3655 18266 3693
rect 16550 3621 16566 3655
rect 16600 3621 18216 3655
rect 18250 3621 18266 3655
rect 16550 3583 18266 3621
rect 16550 3549 16566 3583
rect 16600 3549 18216 3583
rect 18250 3549 18266 3583
rect 16550 3511 18266 3549
rect 16550 3477 16566 3511
rect 16600 3477 18216 3511
rect 18250 3477 18266 3511
rect 16550 3439 18266 3477
rect 16550 3405 16566 3439
rect 16600 3405 18216 3439
rect 18250 3405 18266 3439
rect 16550 3367 18266 3405
rect 16550 3333 16566 3367
rect 16600 3333 18216 3367
rect 18250 3333 18266 3367
rect 16550 3300 18266 3333
rect 16550 3266 16635 3300
rect 16669 3266 16707 3300
rect 16741 3266 16779 3300
rect 16813 3266 16851 3300
rect 16885 3266 16923 3300
rect 16957 3266 16995 3300
rect 17029 3266 17067 3300
rect 17101 3266 17139 3300
rect 17173 3266 17211 3300
rect 17245 3266 17283 3300
rect 17317 3266 17355 3300
rect 17389 3266 17427 3300
rect 17461 3266 17499 3300
rect 17533 3266 17571 3300
rect 17605 3266 17643 3300
rect 17677 3266 17715 3300
rect 17749 3266 17787 3300
rect 17821 3266 17859 3300
rect 17893 3266 17931 3300
rect 17965 3266 18003 3300
rect 18037 3266 18075 3300
rect 18109 3266 18147 3300
rect 18181 3266 18266 3300
rect 16550 3250 18266 3266
rect 18400 4802 20116 4818
rect 18400 4768 18485 4802
rect 18519 4768 18557 4802
rect 18591 4768 18629 4802
rect 18663 4768 18701 4802
rect 18735 4768 18773 4802
rect 18807 4768 18845 4802
rect 18879 4768 18917 4802
rect 18951 4768 18989 4802
rect 19023 4768 19061 4802
rect 19095 4768 19133 4802
rect 19167 4768 19205 4802
rect 19239 4768 19277 4802
rect 19311 4768 19349 4802
rect 19383 4768 19421 4802
rect 19455 4768 19493 4802
rect 19527 4768 19565 4802
rect 19599 4768 19637 4802
rect 19671 4768 19709 4802
rect 19743 4768 19781 4802
rect 19815 4768 19853 4802
rect 19887 4768 19925 4802
rect 19959 4768 19997 4802
rect 20031 4768 20116 4802
rect 18400 4735 20116 4768
rect 18400 4701 18416 4735
rect 18450 4701 20066 4735
rect 20100 4701 20116 4735
rect 18400 4663 20116 4701
rect 18400 4629 18416 4663
rect 18450 4629 20066 4663
rect 20100 4629 20116 4663
rect 18400 4591 20116 4629
rect 18400 4557 18416 4591
rect 18450 4557 20066 4591
rect 20100 4557 20116 4591
rect 18400 4519 20116 4557
rect 18400 4485 18416 4519
rect 18450 4485 20066 4519
rect 20100 4485 20116 4519
rect 18400 4447 20116 4485
rect 18400 4413 18416 4447
rect 18450 4413 20066 4447
rect 20100 4413 20116 4447
rect 18400 4375 20116 4413
rect 18400 4341 18416 4375
rect 18450 4341 20066 4375
rect 20100 4341 20116 4375
rect 18400 4303 20116 4341
rect 18400 4269 18416 4303
rect 18450 4269 20066 4303
rect 20100 4269 20116 4303
rect 18400 4231 20116 4269
rect 18400 4197 18416 4231
rect 18450 4197 20066 4231
rect 20100 4197 20116 4231
rect 18400 4159 20116 4197
rect 18400 4125 18416 4159
rect 18450 4125 20066 4159
rect 20100 4125 20116 4159
rect 18400 4087 20116 4125
rect 18400 4053 18416 4087
rect 18450 4053 20066 4087
rect 20100 4053 20116 4087
rect 18400 4015 20116 4053
rect 18400 3981 18416 4015
rect 18450 3981 20066 4015
rect 20100 3981 20116 4015
rect 18400 3943 20116 3981
rect 18400 3909 18416 3943
rect 18450 3909 20066 3943
rect 20100 3909 20116 3943
rect 18400 3871 20116 3909
rect 18400 3837 18416 3871
rect 18450 3837 20066 3871
rect 20100 3837 20116 3871
rect 18400 3799 20116 3837
rect 18400 3765 18416 3799
rect 18450 3765 20066 3799
rect 20100 3765 20116 3799
rect 18400 3727 20116 3765
rect 18400 3693 18416 3727
rect 18450 3693 20066 3727
rect 20100 3693 20116 3727
rect 18400 3655 20116 3693
rect 18400 3621 18416 3655
rect 18450 3621 20066 3655
rect 20100 3621 20116 3655
rect 18400 3583 20116 3621
rect 18400 3549 18416 3583
rect 18450 3549 20066 3583
rect 20100 3549 20116 3583
rect 18400 3511 20116 3549
rect 18400 3477 18416 3511
rect 18450 3477 20066 3511
rect 20100 3477 20116 3511
rect 18400 3439 20116 3477
rect 18400 3405 18416 3439
rect 18450 3405 20066 3439
rect 20100 3405 20116 3439
rect 18400 3367 20116 3405
rect 18400 3333 18416 3367
rect 18450 3333 20066 3367
rect 20100 3333 20116 3367
rect 18400 3300 20116 3333
rect 18400 3266 18485 3300
rect 18519 3266 18557 3300
rect 18591 3266 18629 3300
rect 18663 3266 18701 3300
rect 18735 3266 18773 3300
rect 18807 3266 18845 3300
rect 18879 3266 18917 3300
rect 18951 3266 18989 3300
rect 19023 3266 19061 3300
rect 19095 3266 19133 3300
rect 19167 3266 19205 3300
rect 19239 3266 19277 3300
rect 19311 3266 19349 3300
rect 19383 3266 19421 3300
rect 19455 3266 19493 3300
rect 19527 3266 19565 3300
rect 19599 3266 19637 3300
rect 19671 3266 19709 3300
rect 19743 3266 19781 3300
rect 19815 3266 19853 3300
rect 19887 3266 19925 3300
rect 19959 3266 19997 3300
rect 20031 3266 20116 3300
rect 18400 3250 20116 3266
<< viali >>
rect 16635 9818 16669 9852
rect 16707 9818 16741 9852
rect 16779 9818 16813 9852
rect 16851 9818 16885 9852
rect 16923 9818 16957 9852
rect 16995 9818 17029 9852
rect 17067 9818 17101 9852
rect 17139 9818 17173 9852
rect 17211 9818 17245 9852
rect 17283 9818 17317 9852
rect 17355 9818 17389 9852
rect 17427 9818 17461 9852
rect 17499 9818 17533 9852
rect 17571 9818 17605 9852
rect 17643 9818 17677 9852
rect 17715 9818 17749 9852
rect 17787 9818 17821 9852
rect 17859 9818 17893 9852
rect 17931 9818 17965 9852
rect 18003 9818 18037 9852
rect 18075 9818 18109 9852
rect 18147 9818 18181 9852
rect 16566 9751 16600 9785
rect 18216 9751 18250 9785
rect 16566 9679 16600 9713
rect 18216 9679 18250 9713
rect 16566 9607 16600 9641
rect 18216 9607 18250 9641
rect 16566 9535 16600 9569
rect 18216 9535 18250 9569
rect 16566 9463 16600 9497
rect 18216 9463 18250 9497
rect 16566 9391 16600 9425
rect 18216 9391 18250 9425
rect 16566 9319 16600 9353
rect 18216 9319 18250 9353
rect 16566 9247 16600 9281
rect 18216 9247 18250 9281
rect 16566 9175 16600 9209
rect 18216 9175 18250 9209
rect 16566 9103 16600 9137
rect 18216 9103 18250 9137
rect 16566 9031 16600 9065
rect 18216 9031 18250 9065
rect 16566 8959 16600 8993
rect 18216 8959 18250 8993
rect 16566 8887 16600 8921
rect 18216 8887 18250 8921
rect 16566 8815 16600 8849
rect 18216 8815 18250 8849
rect 16566 8743 16600 8777
rect 18216 8743 18250 8777
rect 16566 8671 16600 8705
rect 18216 8671 18250 8705
rect 16566 8599 16600 8633
rect 18216 8599 18250 8633
rect 16566 8527 16600 8561
rect 18216 8527 18250 8561
rect 16566 8455 16600 8489
rect 18216 8455 18250 8489
rect 16566 8383 16600 8417
rect 18216 8383 18250 8417
rect 16635 8316 16669 8350
rect 16707 8316 16741 8350
rect 16779 8316 16813 8350
rect 16851 8316 16885 8350
rect 16923 8316 16957 8350
rect 16995 8316 17029 8350
rect 17067 8316 17101 8350
rect 17139 8316 17173 8350
rect 17211 8316 17245 8350
rect 17283 8316 17317 8350
rect 17355 8316 17389 8350
rect 17427 8316 17461 8350
rect 17499 8316 17533 8350
rect 17571 8316 17605 8350
rect 17643 8316 17677 8350
rect 17715 8316 17749 8350
rect 17787 8316 17821 8350
rect 17859 8316 17893 8350
rect 17931 8316 17965 8350
rect 18003 8316 18037 8350
rect 18075 8316 18109 8350
rect 18147 8316 18181 8350
rect 18485 9818 18519 9852
rect 18557 9818 18591 9852
rect 18629 9818 18663 9852
rect 18701 9818 18735 9852
rect 18773 9818 18807 9852
rect 18845 9818 18879 9852
rect 18917 9818 18951 9852
rect 18989 9818 19023 9852
rect 19061 9818 19095 9852
rect 19133 9818 19167 9852
rect 19205 9818 19239 9852
rect 19277 9818 19311 9852
rect 19349 9818 19383 9852
rect 19421 9818 19455 9852
rect 19493 9818 19527 9852
rect 19565 9818 19599 9852
rect 19637 9818 19671 9852
rect 19709 9818 19743 9852
rect 19781 9818 19815 9852
rect 19853 9818 19887 9852
rect 19925 9818 19959 9852
rect 19997 9818 20031 9852
rect 18416 9751 18450 9785
rect 20066 9751 20100 9785
rect 18416 9679 18450 9713
rect 20066 9679 20100 9713
rect 18416 9607 18450 9641
rect 20066 9607 20100 9641
rect 18416 9535 18450 9569
rect 20066 9535 20100 9569
rect 18416 9463 18450 9497
rect 20066 9463 20100 9497
rect 18416 9391 18450 9425
rect 20066 9391 20100 9425
rect 18416 9319 18450 9353
rect 20066 9319 20100 9353
rect 18416 9247 18450 9281
rect 20066 9247 20100 9281
rect 18416 9175 18450 9209
rect 20066 9175 20100 9209
rect 18416 9103 18450 9137
rect 20066 9103 20100 9137
rect 18416 9031 18450 9065
rect 20066 9031 20100 9065
rect 18416 8959 18450 8993
rect 20066 8959 20100 8993
rect 18416 8887 18450 8921
rect 20066 8887 20100 8921
rect 18416 8815 18450 8849
rect 20066 8815 20100 8849
rect 18416 8743 18450 8777
rect 20066 8743 20100 8777
rect 18416 8671 18450 8705
rect 20066 8671 20100 8705
rect 18416 8599 18450 8633
rect 20066 8599 20100 8633
rect 18416 8527 18450 8561
rect 20066 8527 20100 8561
rect 18416 8455 18450 8489
rect 20066 8455 20100 8489
rect 18416 8383 18450 8417
rect 20066 8383 20100 8417
rect 18485 8316 18519 8350
rect 18557 8316 18591 8350
rect 18629 8316 18663 8350
rect 18701 8316 18735 8350
rect 18773 8316 18807 8350
rect 18845 8316 18879 8350
rect 18917 8316 18951 8350
rect 18989 8316 19023 8350
rect 19061 8316 19095 8350
rect 19133 8316 19167 8350
rect 19205 8316 19239 8350
rect 19277 8316 19311 8350
rect 19349 8316 19383 8350
rect 19421 8316 19455 8350
rect 19493 8316 19527 8350
rect 19565 8316 19599 8350
rect 19637 8316 19671 8350
rect 19709 8316 19743 8350
rect 19781 8316 19815 8350
rect 19853 8316 19887 8350
rect 19925 8316 19959 8350
rect 19997 8316 20031 8350
rect 16080 8076 16104 8110
rect 16104 8076 16114 8110
rect 16160 8076 16174 8110
rect 16174 8076 16194 8110
rect 16240 8076 16244 8110
rect 16244 8076 16274 8110
rect 16320 8076 16350 8110
rect 16350 8076 16354 8110
rect 16400 8076 16420 8110
rect 16420 8076 16434 8110
rect 16480 8076 16490 8110
rect 16490 8076 16514 8110
rect 16560 8076 16594 8110
rect 16640 8076 16664 8110
rect 16664 8076 16674 8110
rect 16720 8076 16734 8110
rect 16734 8076 16754 8110
rect 16800 8076 16804 8110
rect 16804 8076 16834 8110
rect 16880 8076 16910 8110
rect 16910 8076 16914 8110
rect 16960 8076 16980 8110
rect 16980 8076 16994 8110
rect 17040 8076 17050 8110
rect 17050 8076 17074 8110
rect 17120 8076 17154 8110
rect 15990 7986 16024 8000
rect 15990 7966 16024 7986
rect 17638 8050 17678 8090
rect 17678 8050 17718 8090
rect 17718 8050 17758 8090
rect 17758 8050 17798 8090
rect 17798 8050 17838 8090
rect 17838 8050 17878 8090
rect 17878 8050 17918 8090
rect 17918 8050 17958 8090
rect 17958 8050 17998 8090
rect 17998 8050 18038 8090
rect 18038 8050 18078 8090
rect 18078 8050 18118 8090
rect 18118 8050 18158 8090
rect 18158 8050 18198 8090
rect 18198 8050 18238 8090
rect 18238 8050 18278 8090
rect 18278 8050 18318 8090
rect 18318 8050 18358 8090
rect 18358 8050 18398 8090
rect 18398 8050 18438 8090
rect 18438 8050 18478 8090
rect 18478 8050 18518 8090
rect 18518 8050 18558 8090
rect 18558 8050 18598 8090
rect 18598 8050 18638 8090
rect 18638 8050 18678 8090
rect 18678 8050 18718 8090
rect 18718 8050 18758 8090
rect 18758 8050 18798 8090
rect 18798 8050 18838 8090
rect 18838 8050 18878 8090
rect 18878 8050 18918 8090
rect 18918 8050 18958 8090
rect 18958 8050 18998 8090
rect 18998 8050 19038 8090
rect 19038 8050 19078 8090
rect 19078 8050 19118 8090
rect 19118 8050 19158 8090
rect 19158 8050 19198 8090
rect 19198 8050 19238 8090
rect 19238 8050 19278 8090
rect 19278 8050 19318 8090
rect 19318 8050 19358 8090
rect 19358 8050 19398 8090
rect 19398 8050 19438 8090
rect 19438 8050 19478 8090
rect 19478 8050 19518 8090
rect 19518 8050 19558 8090
rect 19558 8050 19598 8090
rect 19598 8050 19638 8090
rect 19638 8050 19678 8090
rect 19678 8050 19718 8090
rect 19718 8050 19758 8090
rect 19758 8050 19798 8090
rect 19798 8050 19838 8090
rect 19838 8050 19878 8090
rect 19878 8050 19918 8090
rect 19918 8050 19958 8090
rect 19958 8050 19998 8090
rect 19998 8050 20038 8090
rect 20038 8050 20058 8090
rect 15990 7916 16024 7920
rect 15990 7886 16024 7916
rect 15990 7810 16024 7840
rect 15990 7806 16024 7810
rect 15990 7740 16024 7760
rect 15990 7726 16024 7740
rect 15990 7670 16024 7680
rect 15990 7646 16024 7670
rect 15990 7566 16024 7600
rect 15990 7496 16024 7520
rect 15990 7486 16024 7496
rect 15990 7426 16024 7440
rect 15990 7406 16024 7426
rect 15990 7356 16024 7360
rect 15990 7326 16024 7356
rect 15990 7250 16024 7280
rect 15990 7246 16024 7250
rect 15990 7180 16024 7200
rect 15990 7166 16024 7180
rect 15990 7110 16024 7120
rect 15990 7086 16024 7110
rect 15990 7006 16024 7040
rect 16118 7933 16152 7959
rect 16118 7925 16152 7933
rect 16118 7865 16152 7887
rect 16118 7853 16152 7865
rect 16118 7797 16152 7815
rect 16118 7781 16152 7797
rect 16118 7729 16152 7743
rect 16118 7709 16152 7729
rect 16118 7661 16152 7671
rect 16118 7637 16152 7661
rect 16118 7593 16152 7599
rect 16118 7565 16152 7593
rect 16118 7525 16152 7527
rect 16118 7493 16152 7525
rect 16118 7423 16152 7455
rect 16118 7421 16152 7423
rect 16118 7355 16152 7383
rect 16118 7349 16152 7355
rect 16118 7287 16152 7311
rect 16118 7277 16152 7287
rect 16118 7219 16152 7239
rect 16118 7205 16152 7219
rect 16118 7151 16152 7167
rect 16118 7133 16152 7151
rect 16118 7083 16152 7095
rect 16118 7061 16152 7083
rect 16118 7015 16152 7023
rect 16118 6989 16152 7015
rect 16204 7933 16238 7959
rect 16204 7925 16238 7933
rect 16204 7865 16238 7887
rect 16204 7853 16238 7865
rect 16204 7797 16238 7815
rect 16204 7781 16238 7797
rect 16204 7729 16238 7743
rect 16204 7709 16238 7729
rect 16204 7661 16238 7671
rect 16204 7637 16238 7661
rect 16204 7593 16238 7599
rect 16204 7565 16238 7593
rect 16204 7525 16238 7527
rect 16204 7493 16238 7525
rect 16204 7423 16238 7455
rect 16204 7421 16238 7423
rect 16204 7355 16238 7383
rect 16204 7349 16238 7355
rect 16204 7287 16238 7311
rect 16204 7277 16238 7287
rect 16204 7219 16238 7239
rect 16204 7205 16238 7219
rect 16204 7151 16238 7167
rect 16204 7133 16238 7151
rect 16204 7083 16238 7095
rect 16204 7061 16238 7083
rect 16204 7015 16238 7023
rect 16204 6989 16238 7015
rect 16290 7933 16324 7959
rect 16290 7925 16324 7933
rect 16290 7865 16324 7887
rect 16290 7853 16324 7865
rect 16290 7797 16324 7815
rect 16290 7781 16324 7797
rect 16290 7729 16324 7743
rect 16290 7709 16324 7729
rect 16290 7661 16324 7671
rect 16290 7637 16324 7661
rect 16290 7593 16324 7599
rect 16290 7565 16324 7593
rect 16290 7525 16324 7527
rect 16290 7493 16324 7525
rect 16290 7423 16324 7455
rect 16290 7421 16324 7423
rect 16290 7355 16324 7383
rect 16290 7349 16324 7355
rect 16290 7287 16324 7311
rect 16290 7277 16324 7287
rect 16290 7219 16324 7239
rect 16290 7205 16324 7219
rect 16290 7151 16324 7167
rect 16290 7133 16324 7151
rect 16290 7083 16324 7095
rect 16290 7061 16324 7083
rect 16290 7015 16324 7023
rect 16290 6989 16324 7015
rect 16376 7933 16410 7959
rect 16376 7925 16410 7933
rect 16376 7865 16410 7887
rect 16376 7853 16410 7865
rect 16376 7797 16410 7815
rect 16376 7781 16410 7797
rect 16376 7729 16410 7743
rect 16376 7709 16410 7729
rect 16376 7661 16410 7671
rect 16376 7637 16410 7661
rect 16376 7593 16410 7599
rect 16376 7565 16410 7593
rect 16376 7525 16410 7527
rect 16376 7493 16410 7525
rect 16376 7423 16410 7455
rect 16376 7421 16410 7423
rect 16376 7355 16410 7383
rect 16376 7349 16410 7355
rect 16376 7287 16410 7311
rect 16376 7277 16410 7287
rect 16376 7219 16410 7239
rect 16376 7205 16410 7219
rect 16376 7151 16410 7167
rect 16376 7133 16410 7151
rect 16376 7083 16410 7095
rect 16376 7061 16410 7083
rect 16376 7015 16410 7023
rect 16376 6989 16410 7015
rect 16462 7933 16496 7959
rect 16462 7925 16496 7933
rect 16462 7865 16496 7887
rect 16462 7853 16496 7865
rect 16462 7797 16496 7815
rect 16462 7781 16496 7797
rect 16462 7729 16496 7743
rect 16462 7709 16496 7729
rect 16462 7661 16496 7671
rect 16462 7637 16496 7661
rect 16462 7593 16496 7599
rect 16462 7565 16496 7593
rect 16462 7525 16496 7527
rect 16462 7493 16496 7525
rect 16462 7423 16496 7455
rect 16462 7421 16496 7423
rect 16462 7355 16496 7383
rect 16462 7349 16496 7355
rect 16462 7287 16496 7311
rect 16462 7277 16496 7287
rect 16462 7219 16496 7239
rect 16462 7205 16496 7219
rect 16462 7151 16496 7167
rect 16462 7133 16496 7151
rect 16462 7083 16496 7095
rect 16462 7061 16496 7083
rect 16462 7015 16496 7023
rect 16462 6989 16496 7015
rect 16548 7933 16582 7959
rect 16548 7925 16582 7933
rect 16548 7865 16582 7887
rect 16548 7853 16582 7865
rect 16548 7797 16582 7815
rect 16548 7781 16582 7797
rect 16548 7729 16582 7743
rect 16548 7709 16582 7729
rect 16548 7661 16582 7671
rect 16548 7637 16582 7661
rect 16548 7593 16582 7599
rect 16548 7565 16582 7593
rect 16548 7525 16582 7527
rect 16548 7493 16582 7525
rect 16548 7423 16582 7455
rect 16548 7421 16582 7423
rect 16548 7355 16582 7383
rect 16548 7349 16582 7355
rect 16548 7287 16582 7311
rect 16548 7277 16582 7287
rect 16548 7219 16582 7239
rect 16548 7205 16582 7219
rect 16548 7151 16582 7167
rect 16548 7133 16582 7151
rect 16548 7083 16582 7095
rect 16548 7061 16582 7083
rect 16548 7015 16582 7023
rect 16548 6989 16582 7015
rect 16634 7933 16668 7959
rect 16634 7925 16668 7933
rect 16634 7865 16668 7887
rect 16634 7853 16668 7865
rect 16634 7797 16668 7815
rect 16634 7781 16668 7797
rect 16634 7729 16668 7743
rect 16634 7709 16668 7729
rect 16634 7661 16668 7671
rect 16634 7637 16668 7661
rect 16634 7593 16668 7599
rect 16634 7565 16668 7593
rect 16634 7525 16668 7527
rect 16634 7493 16668 7525
rect 16634 7423 16668 7455
rect 16634 7421 16668 7423
rect 16634 7355 16668 7383
rect 16634 7349 16668 7355
rect 16634 7287 16668 7311
rect 16634 7277 16668 7287
rect 16634 7219 16668 7239
rect 16634 7205 16668 7219
rect 16634 7151 16668 7167
rect 16634 7133 16668 7151
rect 16634 7083 16668 7095
rect 16634 7061 16668 7083
rect 16634 7015 16668 7023
rect 16634 6989 16668 7015
rect 16720 7933 16754 7959
rect 16720 7925 16754 7933
rect 16720 7865 16754 7887
rect 16720 7853 16754 7865
rect 16720 7797 16754 7815
rect 16720 7781 16754 7797
rect 16720 7729 16754 7743
rect 16720 7709 16754 7729
rect 16720 7661 16754 7671
rect 16720 7637 16754 7661
rect 16720 7593 16754 7599
rect 16720 7565 16754 7593
rect 16720 7525 16754 7527
rect 16720 7493 16754 7525
rect 16720 7423 16754 7455
rect 16720 7421 16754 7423
rect 16720 7355 16754 7383
rect 16720 7349 16754 7355
rect 16720 7287 16754 7311
rect 16720 7277 16754 7287
rect 16720 7219 16754 7239
rect 16720 7205 16754 7219
rect 16720 7151 16754 7167
rect 16720 7133 16754 7151
rect 16720 7083 16754 7095
rect 16720 7061 16754 7083
rect 16720 7015 16754 7023
rect 16720 6989 16754 7015
rect 16806 7933 16840 7959
rect 16806 7925 16840 7933
rect 16806 7865 16840 7887
rect 16806 7853 16840 7865
rect 16806 7797 16840 7815
rect 16806 7781 16840 7797
rect 16806 7729 16840 7743
rect 16806 7709 16840 7729
rect 16806 7661 16840 7671
rect 16806 7637 16840 7661
rect 16806 7593 16840 7599
rect 16806 7565 16840 7593
rect 16806 7525 16840 7527
rect 16806 7493 16840 7525
rect 16806 7423 16840 7455
rect 16806 7421 16840 7423
rect 16806 7355 16840 7383
rect 16806 7349 16840 7355
rect 16806 7287 16840 7311
rect 16806 7277 16840 7287
rect 16806 7219 16840 7239
rect 16806 7205 16840 7219
rect 16806 7151 16840 7167
rect 16806 7133 16840 7151
rect 16806 7083 16840 7095
rect 16806 7061 16840 7083
rect 16806 7015 16840 7023
rect 16806 6989 16840 7015
rect 16892 7933 16926 7959
rect 16892 7925 16926 7933
rect 16892 7865 16926 7887
rect 16892 7853 16926 7865
rect 16892 7797 16926 7815
rect 16892 7781 16926 7797
rect 16892 7729 16926 7743
rect 16892 7709 16926 7729
rect 16892 7661 16926 7671
rect 16892 7637 16926 7661
rect 16892 7593 16926 7599
rect 16892 7565 16926 7593
rect 16892 7525 16926 7527
rect 16892 7493 16926 7525
rect 16892 7423 16926 7455
rect 16892 7421 16926 7423
rect 16892 7355 16926 7383
rect 16892 7349 16926 7355
rect 16892 7287 16926 7311
rect 16892 7277 16926 7287
rect 16892 7219 16926 7239
rect 16892 7205 16926 7219
rect 16892 7151 16926 7167
rect 16892 7133 16926 7151
rect 16892 7083 16926 7095
rect 16892 7061 16926 7083
rect 16892 7015 16926 7023
rect 16892 6989 16926 7015
rect 16978 7933 17012 7959
rect 16978 7925 17012 7933
rect 16978 7865 17012 7887
rect 16978 7853 17012 7865
rect 16978 7797 17012 7815
rect 16978 7781 17012 7797
rect 16978 7729 17012 7743
rect 16978 7709 17012 7729
rect 16978 7661 17012 7671
rect 16978 7637 17012 7661
rect 16978 7593 17012 7599
rect 16978 7565 17012 7593
rect 16978 7525 17012 7527
rect 16978 7493 17012 7525
rect 16978 7423 17012 7455
rect 16978 7421 17012 7423
rect 16978 7355 17012 7383
rect 16978 7349 17012 7355
rect 16978 7287 17012 7311
rect 16978 7277 17012 7287
rect 16978 7219 17012 7239
rect 16978 7205 17012 7219
rect 16978 7151 17012 7167
rect 16978 7133 17012 7151
rect 16978 7083 17012 7095
rect 16978 7061 17012 7083
rect 16978 7015 17012 7023
rect 16978 6989 17012 7015
rect 17064 7933 17098 7959
rect 17064 7925 17098 7933
rect 17064 7865 17098 7887
rect 17064 7853 17098 7865
rect 17064 7797 17098 7815
rect 17064 7781 17098 7797
rect 17064 7729 17098 7743
rect 17064 7709 17098 7729
rect 17064 7661 17098 7671
rect 17064 7637 17098 7661
rect 17064 7593 17098 7599
rect 17064 7565 17098 7593
rect 17064 7525 17098 7527
rect 17064 7493 17098 7525
rect 17064 7423 17098 7455
rect 17064 7421 17098 7423
rect 17064 7355 17098 7383
rect 17064 7349 17098 7355
rect 17064 7287 17098 7311
rect 17064 7277 17098 7287
rect 17064 7219 17098 7239
rect 17064 7205 17098 7219
rect 17064 7151 17098 7167
rect 17064 7133 17098 7151
rect 17064 7083 17098 7095
rect 17064 7061 17098 7083
rect 17064 7015 17098 7023
rect 17064 6989 17098 7015
rect 17150 7933 17184 7959
rect 17150 7925 17184 7933
rect 17150 7865 17184 7887
rect 17150 7853 17184 7865
rect 17150 7797 17184 7815
rect 17150 7781 17184 7797
rect 17150 7729 17184 7743
rect 17150 7709 17184 7729
rect 17150 7661 17184 7671
rect 17150 7637 17184 7661
rect 17150 7593 17184 7599
rect 17150 7565 17184 7593
rect 17150 7525 17184 7527
rect 17150 7493 17184 7525
rect 17150 7423 17184 7455
rect 17150 7421 17184 7423
rect 17150 7355 17184 7383
rect 17150 7349 17184 7355
rect 17150 7287 17184 7311
rect 17150 7277 17184 7287
rect 17150 7219 17184 7239
rect 17150 7205 17184 7219
rect 17150 7151 17184 7167
rect 17150 7133 17184 7151
rect 17150 7083 17184 7095
rect 17150 7061 17184 7083
rect 17150 7015 17184 7023
rect 17150 6989 17184 7015
rect 17280 7986 17314 8000
rect 17280 7966 17314 7986
rect 17280 7916 17314 7920
rect 17280 7886 17314 7916
rect 17280 7810 17314 7840
rect 17280 7806 17314 7810
rect 17280 7740 17314 7760
rect 17280 7726 17314 7740
rect 17280 7670 17314 7680
rect 17280 7646 17314 7670
rect 17280 7566 17314 7600
rect 17280 7496 17314 7520
rect 17280 7486 17314 7496
rect 17280 7426 17314 7440
rect 17280 7406 17314 7426
rect 17280 7356 17314 7360
rect 17280 7326 17314 7356
rect 17280 7250 17314 7280
rect 17280 7246 17314 7250
rect 17280 7180 17314 7200
rect 17280 7166 17314 7180
rect 17280 7110 17314 7120
rect 17280 7086 17314 7110
rect 17280 7006 17314 7040
rect 17518 7890 17538 7930
rect 17538 7890 17558 7930
rect 17518 7850 17558 7890
rect 17518 7810 17538 7850
rect 17538 7810 17558 7850
rect 17518 7770 17558 7810
rect 17518 7730 17538 7770
rect 17538 7730 17558 7770
rect 17518 7690 17558 7730
rect 17518 7650 17538 7690
rect 17538 7650 17558 7690
rect 17518 7610 17558 7650
rect 17518 7570 17538 7610
rect 17538 7570 17558 7610
rect 17518 7530 17558 7570
rect 17518 7490 17538 7530
rect 17538 7490 17558 7530
rect 17518 7450 17558 7490
rect 17518 7410 17538 7450
rect 17538 7410 17558 7450
rect 17518 7370 17558 7410
rect 17518 7330 17538 7370
rect 17538 7330 17558 7370
rect 17518 7290 17558 7330
rect 17518 7250 17538 7290
rect 17538 7250 17558 7290
rect 17518 7210 17558 7250
rect 17518 7170 17538 7210
rect 17538 7170 17558 7210
rect 17518 7130 17558 7170
rect 17518 7090 17538 7130
rect 17538 7090 17558 7130
rect 17518 7050 17558 7090
rect 17518 7010 17538 7050
rect 17538 7010 17558 7050
rect 17518 6990 17558 7010
rect 17622 7874 17656 7908
rect 17622 7802 17656 7836
rect 17622 7730 17656 7764
rect 17622 7658 17656 7692
rect 17622 7586 17656 7620
rect 17622 7514 17656 7548
rect 17622 7442 17656 7476
rect 17622 7370 17656 7404
rect 17622 7298 17656 7332
rect 17622 7226 17656 7260
rect 17622 7154 17656 7188
rect 17622 7082 17656 7116
rect 17622 7010 17656 7044
rect 17708 7874 17742 7908
rect 17708 7802 17742 7836
rect 17708 7730 17742 7764
rect 17708 7658 17742 7692
rect 17708 7586 17742 7620
rect 17708 7514 17742 7548
rect 17708 7442 17742 7476
rect 17708 7370 17742 7404
rect 17708 7298 17742 7332
rect 17708 7226 17742 7260
rect 17708 7154 17742 7188
rect 17708 7082 17742 7116
rect 17708 7010 17742 7044
rect 17794 7874 17828 7908
rect 17794 7802 17828 7836
rect 17794 7730 17828 7764
rect 17794 7658 17828 7692
rect 17794 7586 17828 7620
rect 17794 7514 17828 7548
rect 17794 7442 17828 7476
rect 17794 7370 17828 7404
rect 17794 7298 17828 7332
rect 17794 7226 17828 7260
rect 17794 7154 17828 7188
rect 17794 7082 17828 7116
rect 17794 7010 17828 7044
rect 17880 7874 17914 7908
rect 17880 7802 17914 7836
rect 17880 7730 17914 7764
rect 17880 7658 17914 7692
rect 17880 7586 17914 7620
rect 17880 7514 17914 7548
rect 17880 7442 17914 7476
rect 17880 7370 17914 7404
rect 17880 7298 17914 7332
rect 17880 7226 17914 7260
rect 17880 7154 17914 7188
rect 17880 7082 17914 7116
rect 17880 7010 17914 7044
rect 17966 7874 18000 7908
rect 17966 7802 18000 7836
rect 17966 7730 18000 7764
rect 17966 7658 18000 7692
rect 17966 7586 18000 7620
rect 17966 7514 18000 7548
rect 17966 7442 18000 7476
rect 17966 7370 18000 7404
rect 17966 7298 18000 7332
rect 17966 7226 18000 7260
rect 17966 7154 18000 7188
rect 17966 7082 18000 7116
rect 17966 7010 18000 7044
rect 18052 7874 18086 7908
rect 18052 7802 18086 7836
rect 18052 7730 18086 7764
rect 18052 7658 18086 7692
rect 18052 7586 18086 7620
rect 18052 7514 18086 7548
rect 18052 7442 18086 7476
rect 18052 7370 18086 7404
rect 18052 7298 18086 7332
rect 18052 7226 18086 7260
rect 18052 7154 18086 7188
rect 18052 7082 18086 7116
rect 18052 7010 18086 7044
rect 18138 7874 18172 7908
rect 18138 7802 18172 7836
rect 18138 7730 18172 7764
rect 18138 7658 18172 7692
rect 18138 7586 18172 7620
rect 18138 7514 18172 7548
rect 18138 7442 18172 7476
rect 18138 7370 18172 7404
rect 18138 7298 18172 7332
rect 18138 7226 18172 7260
rect 18138 7154 18172 7188
rect 18138 7082 18172 7116
rect 18138 7010 18172 7044
rect 18224 7874 18258 7908
rect 18224 7802 18258 7836
rect 18224 7730 18258 7764
rect 18224 7658 18258 7692
rect 18224 7586 18258 7620
rect 18224 7514 18258 7548
rect 18224 7442 18258 7476
rect 18224 7370 18258 7404
rect 18224 7298 18258 7332
rect 18224 7226 18258 7260
rect 18224 7154 18258 7188
rect 18224 7082 18258 7116
rect 18224 7010 18258 7044
rect 18310 7874 18344 7908
rect 18310 7802 18344 7836
rect 18310 7730 18344 7764
rect 18310 7658 18344 7692
rect 18310 7586 18344 7620
rect 18310 7514 18344 7548
rect 18310 7442 18344 7476
rect 18310 7370 18344 7404
rect 18310 7298 18344 7332
rect 18310 7226 18344 7260
rect 18310 7154 18344 7188
rect 18310 7082 18344 7116
rect 18310 7010 18344 7044
rect 18396 7874 18430 7908
rect 18396 7802 18430 7836
rect 18396 7730 18430 7764
rect 18396 7658 18430 7692
rect 18396 7586 18430 7620
rect 18396 7514 18430 7548
rect 18396 7442 18430 7476
rect 18396 7370 18430 7404
rect 18396 7298 18430 7332
rect 18396 7226 18430 7260
rect 18396 7154 18430 7188
rect 18396 7082 18430 7116
rect 18396 7010 18430 7044
rect 18482 7874 18516 7908
rect 18482 7802 18516 7836
rect 18482 7730 18516 7764
rect 18482 7658 18516 7692
rect 18482 7586 18516 7620
rect 18482 7514 18516 7548
rect 18482 7442 18516 7476
rect 18482 7370 18516 7404
rect 18482 7298 18516 7332
rect 18482 7226 18516 7260
rect 18482 7154 18516 7188
rect 18482 7082 18516 7116
rect 18482 7010 18516 7044
rect 18568 7874 18602 7908
rect 18568 7802 18602 7836
rect 18568 7730 18602 7764
rect 18568 7658 18602 7692
rect 18568 7586 18602 7620
rect 18568 7514 18602 7548
rect 18568 7442 18602 7476
rect 18568 7370 18602 7404
rect 18568 7298 18602 7332
rect 18568 7226 18602 7260
rect 18568 7154 18602 7188
rect 18568 7082 18602 7116
rect 18568 7010 18602 7044
rect 18654 7874 18688 7908
rect 18654 7802 18688 7836
rect 18654 7730 18688 7764
rect 18654 7658 18688 7692
rect 18654 7586 18688 7620
rect 18654 7514 18688 7548
rect 18654 7442 18688 7476
rect 18654 7370 18688 7404
rect 18654 7298 18688 7332
rect 18654 7226 18688 7260
rect 18654 7154 18688 7188
rect 18654 7082 18688 7116
rect 18654 7010 18688 7044
rect 18740 7874 18774 7908
rect 18740 7802 18774 7836
rect 18740 7730 18774 7764
rect 18740 7658 18774 7692
rect 18740 7586 18774 7620
rect 18740 7514 18774 7548
rect 18740 7442 18774 7476
rect 18740 7370 18774 7404
rect 18740 7298 18774 7332
rect 18740 7226 18774 7260
rect 18740 7154 18774 7188
rect 18740 7082 18774 7116
rect 18740 7010 18774 7044
rect 18826 7874 18860 7908
rect 18826 7802 18860 7836
rect 18826 7730 18860 7764
rect 18826 7658 18860 7692
rect 18826 7586 18860 7620
rect 18826 7514 18860 7548
rect 18826 7442 18860 7476
rect 18826 7370 18860 7404
rect 18826 7298 18860 7332
rect 18826 7226 18860 7260
rect 18826 7154 18860 7188
rect 18826 7082 18860 7116
rect 18826 7010 18860 7044
rect 18912 7874 18946 7908
rect 18912 7802 18946 7836
rect 18912 7730 18946 7764
rect 18912 7658 18946 7692
rect 18912 7586 18946 7620
rect 18912 7514 18946 7548
rect 18912 7442 18946 7476
rect 18912 7370 18946 7404
rect 18912 7298 18946 7332
rect 18912 7226 18946 7260
rect 18912 7154 18946 7188
rect 18912 7082 18946 7116
rect 18912 7010 18946 7044
rect 18998 7874 19032 7908
rect 18998 7802 19032 7836
rect 18998 7730 19032 7764
rect 18998 7658 19032 7692
rect 18998 7586 19032 7620
rect 18998 7514 19032 7548
rect 18998 7442 19032 7476
rect 18998 7370 19032 7404
rect 18998 7298 19032 7332
rect 18998 7226 19032 7260
rect 18998 7154 19032 7188
rect 18998 7082 19032 7116
rect 18998 7010 19032 7044
rect 19084 7874 19118 7908
rect 19084 7802 19118 7836
rect 19084 7730 19118 7764
rect 19084 7658 19118 7692
rect 19084 7586 19118 7620
rect 19084 7514 19118 7548
rect 19084 7442 19118 7476
rect 19084 7370 19118 7404
rect 19084 7298 19118 7332
rect 19084 7226 19118 7260
rect 19084 7154 19118 7188
rect 19084 7082 19118 7116
rect 19084 7010 19118 7044
rect 19170 7874 19204 7908
rect 19170 7802 19204 7836
rect 19170 7730 19204 7764
rect 19170 7658 19204 7692
rect 19170 7586 19204 7620
rect 19170 7514 19204 7548
rect 19170 7442 19204 7476
rect 19170 7370 19204 7404
rect 19170 7298 19204 7332
rect 19170 7226 19204 7260
rect 19170 7154 19204 7188
rect 19170 7082 19204 7116
rect 19170 7010 19204 7044
rect 19256 7874 19290 7908
rect 19256 7802 19290 7836
rect 19256 7730 19290 7764
rect 19256 7658 19290 7692
rect 19256 7586 19290 7620
rect 19256 7514 19290 7548
rect 19256 7442 19290 7476
rect 19256 7370 19290 7404
rect 19256 7298 19290 7332
rect 19256 7226 19290 7260
rect 19256 7154 19290 7188
rect 19256 7082 19290 7116
rect 19256 7010 19290 7044
rect 19342 7874 19376 7908
rect 19342 7802 19376 7836
rect 19342 7730 19376 7764
rect 19342 7658 19376 7692
rect 19342 7586 19376 7620
rect 19342 7514 19376 7548
rect 19342 7442 19376 7476
rect 19342 7370 19376 7404
rect 19342 7298 19376 7332
rect 19342 7226 19376 7260
rect 19342 7154 19376 7188
rect 19342 7082 19376 7116
rect 19342 7010 19376 7044
rect 19428 7874 19462 7908
rect 19428 7802 19462 7836
rect 19428 7730 19462 7764
rect 19428 7658 19462 7692
rect 19428 7586 19462 7620
rect 19428 7514 19462 7548
rect 19428 7442 19462 7476
rect 19428 7370 19462 7404
rect 19428 7298 19462 7332
rect 19428 7226 19462 7260
rect 19428 7154 19462 7188
rect 19428 7082 19462 7116
rect 19428 7010 19462 7044
rect 19514 7874 19548 7908
rect 19514 7802 19548 7836
rect 19514 7730 19548 7764
rect 19514 7658 19548 7692
rect 19514 7586 19548 7620
rect 19514 7514 19548 7548
rect 19514 7442 19548 7476
rect 19514 7370 19548 7404
rect 19514 7298 19548 7332
rect 19514 7226 19548 7260
rect 19514 7154 19548 7188
rect 19514 7082 19548 7116
rect 19514 7010 19548 7044
rect 19600 7874 19634 7908
rect 19600 7802 19634 7836
rect 19600 7730 19634 7764
rect 19600 7658 19634 7692
rect 19600 7586 19634 7620
rect 19600 7514 19634 7548
rect 19600 7442 19634 7476
rect 19600 7370 19634 7404
rect 19600 7298 19634 7332
rect 19600 7226 19634 7260
rect 19600 7154 19634 7188
rect 19600 7082 19634 7116
rect 19600 7010 19634 7044
rect 19686 7874 19720 7908
rect 19686 7802 19720 7836
rect 19686 7730 19720 7764
rect 19686 7658 19720 7692
rect 19686 7586 19720 7620
rect 19686 7514 19720 7548
rect 19686 7442 19720 7476
rect 19686 7370 19720 7404
rect 19686 7298 19720 7332
rect 19686 7226 19720 7260
rect 19686 7154 19720 7188
rect 19686 7082 19720 7116
rect 19686 7010 19720 7044
rect 19772 7874 19806 7908
rect 19772 7802 19806 7836
rect 19772 7730 19806 7764
rect 19772 7658 19806 7692
rect 19772 7586 19806 7620
rect 19772 7514 19806 7548
rect 19772 7442 19806 7476
rect 19772 7370 19806 7404
rect 19772 7298 19806 7332
rect 19772 7226 19806 7260
rect 19772 7154 19806 7188
rect 19772 7082 19806 7116
rect 19772 7010 19806 7044
rect 19858 7874 19892 7908
rect 19858 7802 19892 7836
rect 19858 7730 19892 7764
rect 19858 7658 19892 7692
rect 19858 7586 19892 7620
rect 19858 7514 19892 7548
rect 19858 7442 19892 7476
rect 19858 7370 19892 7404
rect 19858 7298 19892 7332
rect 19858 7226 19892 7260
rect 19858 7154 19892 7188
rect 19858 7082 19892 7116
rect 19858 7010 19892 7044
rect 19944 7874 19978 7908
rect 19944 7802 19978 7836
rect 19944 7730 19978 7764
rect 19944 7658 19978 7692
rect 19944 7586 19978 7620
rect 19944 7514 19978 7548
rect 19944 7442 19978 7476
rect 19944 7370 19978 7404
rect 19944 7298 19978 7332
rect 19944 7226 19978 7260
rect 19944 7154 19978 7188
rect 19944 7082 19978 7116
rect 19944 7010 19978 7044
rect 20030 7874 20064 7908
rect 20030 7802 20064 7836
rect 20030 7730 20064 7764
rect 20030 7658 20064 7692
rect 20030 7586 20064 7620
rect 20030 7514 20064 7548
rect 20030 7442 20064 7476
rect 20030 7370 20064 7404
rect 20030 7298 20064 7332
rect 20030 7226 20064 7260
rect 20030 7154 20064 7188
rect 20030 7082 20064 7116
rect 20030 7010 20064 7044
rect 20138 7890 20158 7930
rect 20158 7890 20178 7930
rect 20138 7850 20178 7890
rect 20138 7810 20158 7850
rect 20158 7810 20178 7850
rect 20138 7770 20178 7810
rect 20138 7730 20158 7770
rect 20158 7730 20178 7770
rect 20138 7690 20178 7730
rect 20138 7650 20158 7690
rect 20158 7650 20178 7690
rect 20138 7610 20178 7650
rect 20138 7570 20158 7610
rect 20158 7570 20178 7610
rect 20138 7530 20178 7570
rect 20138 7490 20158 7530
rect 20158 7490 20178 7530
rect 20138 7450 20178 7490
rect 20138 7410 20158 7450
rect 20158 7410 20178 7450
rect 20138 7370 20178 7410
rect 20138 7330 20158 7370
rect 20158 7330 20178 7370
rect 20138 7290 20178 7330
rect 20138 7250 20158 7290
rect 20158 7250 20178 7290
rect 20138 7210 20178 7250
rect 20138 7170 20158 7210
rect 20158 7170 20178 7210
rect 20138 7130 20178 7170
rect 20138 7090 20158 7130
rect 20158 7090 20178 7130
rect 20138 7050 20178 7090
rect 20138 7010 20158 7050
rect 20158 7010 20178 7050
rect 20138 6990 20178 7010
rect 11813 6896 11821 6930
rect 11821 6896 11847 6930
rect 11885 6896 11889 6930
rect 11889 6896 11919 6930
rect 11957 6896 11991 6930
rect 12029 6896 12059 6930
rect 12059 6896 12063 6930
rect 12101 6896 12127 6930
rect 12127 6896 12135 6930
rect 12379 6896 12387 6930
rect 12387 6896 12413 6930
rect 12451 6896 12455 6930
rect 12455 6896 12485 6930
rect 12523 6896 12557 6930
rect 12595 6896 12625 6930
rect 12625 6896 12629 6930
rect 12667 6896 12693 6930
rect 12693 6896 12701 6930
rect 12945 6896 12953 6930
rect 12953 6896 12979 6930
rect 13017 6896 13021 6930
rect 13021 6896 13051 6930
rect 13089 6896 13123 6930
rect 13161 6896 13191 6930
rect 13191 6896 13195 6930
rect 13233 6896 13259 6930
rect 13259 6896 13267 6930
rect 13511 6896 13519 6930
rect 13519 6896 13545 6930
rect 13583 6896 13587 6930
rect 13587 6896 13617 6930
rect 13655 6896 13689 6930
rect 13727 6896 13757 6930
rect 13757 6896 13761 6930
rect 13799 6896 13825 6930
rect 13825 6896 13833 6930
rect 14077 6896 14085 6930
rect 14085 6896 14111 6930
rect 14149 6896 14153 6930
rect 14153 6896 14183 6930
rect 14221 6896 14255 6930
rect 14293 6896 14323 6930
rect 14323 6896 14327 6930
rect 14365 6896 14391 6930
rect 14391 6896 14399 6930
rect 14643 6896 14651 6930
rect 14651 6896 14677 6930
rect 14715 6896 14719 6930
rect 14719 6896 14749 6930
rect 14787 6896 14821 6930
rect 14859 6896 14889 6930
rect 14889 6896 14893 6930
rect 14931 6896 14957 6930
rect 14957 6896 14965 6930
rect 15209 6896 15217 6930
rect 15217 6896 15243 6930
rect 15281 6896 15285 6930
rect 15285 6896 15315 6930
rect 15353 6896 15387 6930
rect 15425 6896 15455 6930
rect 15455 6896 15459 6930
rect 15497 6896 15523 6930
rect 15523 6896 15531 6930
rect 16218 6897 16222 6931
rect 16222 6897 16252 6931
rect 16290 6897 16324 6931
rect 16362 6897 16392 6931
rect 16392 6897 16396 6931
rect 16562 6897 16566 6931
rect 16566 6897 16596 6931
rect 16634 6897 16668 6931
rect 16706 6897 16736 6931
rect 16736 6897 16740 6931
rect 16906 6897 16910 6931
rect 16910 6897 16940 6931
rect 16978 6897 17012 6931
rect 17050 6897 17080 6931
rect 17080 6897 17084 6931
rect 17686 6874 17692 6908
rect 17692 6874 17720 6908
rect 17758 6874 17760 6908
rect 17760 6874 17792 6908
rect 17830 6874 17862 6908
rect 17862 6874 17864 6908
rect 17902 6874 17930 6908
rect 17930 6874 17936 6908
rect 11674 6812 11708 6838
rect 11674 6804 11708 6812
rect 11674 6744 11708 6766
rect 11674 6732 11708 6744
rect 11674 6676 11708 6694
rect 11674 6660 11708 6676
rect 11674 6608 11708 6622
rect 11674 6588 11708 6608
rect 11674 6540 11708 6550
rect 11674 6516 11708 6540
rect 11674 6472 11708 6478
rect 11674 6444 11708 6472
rect 11674 6404 11708 6406
rect 11674 6372 11708 6404
rect 11674 6302 11708 6334
rect 11674 6300 11708 6302
rect 11674 6234 11708 6262
rect 11674 6228 11708 6234
rect 11674 6166 11708 6190
rect 11674 6156 11708 6166
rect 11674 6098 11708 6118
rect 11674 6084 11708 6098
rect 11674 6030 11708 6046
rect 11674 6012 11708 6030
rect 11674 5962 11708 5974
rect 11674 5940 11708 5962
rect 11674 5894 11708 5902
rect 11674 5868 11708 5894
rect 11785 6812 11819 6838
rect 11785 6804 11819 6812
rect 11785 6744 11819 6766
rect 11785 6732 11819 6744
rect 11785 6676 11819 6694
rect 11785 6660 11819 6676
rect 11785 6608 11819 6622
rect 11785 6588 11819 6608
rect 11785 6540 11819 6550
rect 11785 6516 11819 6540
rect 11785 6472 11819 6478
rect 11785 6444 11819 6472
rect 11785 6404 11819 6406
rect 11785 6372 11819 6404
rect 11785 6302 11819 6334
rect 11785 6300 11819 6302
rect 11785 6234 11819 6262
rect 11785 6228 11819 6234
rect 11785 6166 11819 6190
rect 11785 6156 11819 6166
rect 11785 6098 11819 6118
rect 11785 6084 11819 6098
rect 11785 6030 11819 6046
rect 11785 6012 11819 6030
rect 11785 5962 11819 5974
rect 11785 5940 11819 5962
rect 11785 5894 11819 5902
rect 11785 5868 11819 5894
rect 11871 6812 11905 6838
rect 11871 6804 11905 6812
rect 11871 6744 11905 6766
rect 11871 6732 11905 6744
rect 11871 6676 11905 6694
rect 11871 6660 11905 6676
rect 11871 6608 11905 6622
rect 11871 6588 11905 6608
rect 11871 6540 11905 6550
rect 11871 6516 11905 6540
rect 11871 6472 11905 6478
rect 11871 6444 11905 6472
rect 11871 6404 11905 6406
rect 11871 6372 11905 6404
rect 11871 6302 11905 6334
rect 11871 6300 11905 6302
rect 11871 6234 11905 6262
rect 11871 6228 11905 6234
rect 11871 6166 11905 6190
rect 11871 6156 11905 6166
rect 11871 6098 11905 6118
rect 11871 6084 11905 6098
rect 11871 6030 11905 6046
rect 11871 6012 11905 6030
rect 11871 5962 11905 5974
rect 11871 5940 11905 5962
rect 11871 5894 11905 5902
rect 11871 5868 11905 5894
rect 11957 6812 11991 6838
rect 11957 6804 11991 6812
rect 11957 6744 11991 6766
rect 11957 6732 11991 6744
rect 11957 6676 11991 6694
rect 11957 6660 11991 6676
rect 11957 6608 11991 6622
rect 11957 6588 11991 6608
rect 11957 6540 11991 6550
rect 11957 6516 11991 6540
rect 11957 6472 11991 6478
rect 11957 6444 11991 6472
rect 11957 6404 11991 6406
rect 11957 6372 11991 6404
rect 11957 6302 11991 6334
rect 11957 6300 11991 6302
rect 11957 6234 11991 6262
rect 11957 6228 11991 6234
rect 11957 6166 11991 6190
rect 11957 6156 11991 6166
rect 11957 6098 11991 6118
rect 11957 6084 11991 6098
rect 11957 6030 11991 6046
rect 11957 6012 11991 6030
rect 11957 5962 11991 5974
rect 11957 5940 11991 5962
rect 11957 5894 11991 5902
rect 11957 5868 11991 5894
rect 12043 6812 12077 6838
rect 12043 6804 12077 6812
rect 12043 6744 12077 6766
rect 12043 6732 12077 6744
rect 12043 6676 12077 6694
rect 12043 6660 12077 6676
rect 12043 6608 12077 6622
rect 12043 6588 12077 6608
rect 12043 6540 12077 6550
rect 12043 6516 12077 6540
rect 12043 6472 12077 6478
rect 12043 6444 12077 6472
rect 12043 6404 12077 6406
rect 12043 6372 12077 6404
rect 12043 6302 12077 6334
rect 12043 6300 12077 6302
rect 12043 6234 12077 6262
rect 12043 6228 12077 6234
rect 12043 6166 12077 6190
rect 12043 6156 12077 6166
rect 12043 6098 12077 6118
rect 12043 6084 12077 6098
rect 12043 6030 12077 6046
rect 12043 6012 12077 6030
rect 12043 5962 12077 5974
rect 12043 5940 12077 5962
rect 12043 5894 12077 5902
rect 12043 5868 12077 5894
rect 12129 6812 12163 6838
rect 12129 6804 12163 6812
rect 12129 6744 12163 6766
rect 12129 6732 12163 6744
rect 12129 6676 12163 6694
rect 12129 6660 12163 6676
rect 12129 6608 12163 6622
rect 12129 6588 12163 6608
rect 12129 6540 12163 6550
rect 12129 6516 12163 6540
rect 12129 6472 12163 6478
rect 12129 6444 12163 6472
rect 12129 6404 12163 6406
rect 12129 6372 12163 6404
rect 12129 6302 12163 6334
rect 12129 6300 12163 6302
rect 12129 6234 12163 6262
rect 12129 6228 12163 6234
rect 12129 6166 12163 6190
rect 12129 6156 12163 6166
rect 12129 6098 12163 6118
rect 12129 6084 12163 6098
rect 12129 6030 12163 6046
rect 12129 6012 12163 6030
rect 12129 5962 12163 5974
rect 12129 5940 12163 5962
rect 12129 5894 12163 5902
rect 12129 5868 12163 5894
rect 12240 6812 12274 6838
rect 12240 6804 12274 6812
rect 12240 6744 12274 6766
rect 12240 6732 12274 6744
rect 12240 6676 12274 6694
rect 12240 6660 12274 6676
rect 12240 6608 12274 6622
rect 12240 6588 12274 6608
rect 12240 6540 12274 6550
rect 12240 6516 12274 6540
rect 12240 6472 12274 6478
rect 12240 6444 12274 6472
rect 12240 6404 12274 6406
rect 12240 6372 12274 6404
rect 12240 6302 12274 6334
rect 12240 6300 12274 6302
rect 12240 6234 12274 6262
rect 12240 6228 12274 6234
rect 12240 6166 12274 6190
rect 12240 6156 12274 6166
rect 12240 6098 12274 6118
rect 12240 6084 12274 6098
rect 12240 6030 12274 6046
rect 12240 6012 12274 6030
rect 12240 5962 12274 5974
rect 12240 5940 12274 5962
rect 12240 5894 12274 5902
rect 12240 5868 12274 5894
rect 12351 6812 12385 6838
rect 12351 6804 12385 6812
rect 12351 6744 12385 6766
rect 12351 6732 12385 6744
rect 12351 6676 12385 6694
rect 12351 6660 12385 6676
rect 12351 6608 12385 6622
rect 12351 6588 12385 6608
rect 12351 6540 12385 6550
rect 12351 6516 12385 6540
rect 12351 6472 12385 6478
rect 12351 6444 12385 6472
rect 12351 6404 12385 6406
rect 12351 6372 12385 6404
rect 12351 6302 12385 6334
rect 12351 6300 12385 6302
rect 12351 6234 12385 6262
rect 12351 6228 12385 6234
rect 12351 6166 12385 6190
rect 12351 6156 12385 6166
rect 12351 6098 12385 6118
rect 12351 6084 12385 6098
rect 12351 6030 12385 6046
rect 12351 6012 12385 6030
rect 12351 5962 12385 5974
rect 12351 5940 12385 5962
rect 12351 5894 12385 5902
rect 12351 5868 12385 5894
rect 12437 6812 12471 6838
rect 12437 6804 12471 6812
rect 12437 6744 12471 6766
rect 12437 6732 12471 6744
rect 12437 6676 12471 6694
rect 12437 6660 12471 6676
rect 12437 6608 12471 6622
rect 12437 6588 12471 6608
rect 12437 6540 12471 6550
rect 12437 6516 12471 6540
rect 12437 6472 12471 6478
rect 12437 6444 12471 6472
rect 12437 6404 12471 6406
rect 12437 6372 12471 6404
rect 12437 6302 12471 6334
rect 12437 6300 12471 6302
rect 12437 6234 12471 6262
rect 12437 6228 12471 6234
rect 12437 6166 12471 6190
rect 12437 6156 12471 6166
rect 12437 6098 12471 6118
rect 12437 6084 12471 6098
rect 12437 6030 12471 6046
rect 12437 6012 12471 6030
rect 12437 5962 12471 5974
rect 12437 5940 12471 5962
rect 12437 5894 12471 5902
rect 12437 5868 12471 5894
rect 12523 6812 12557 6838
rect 12523 6804 12557 6812
rect 12523 6744 12557 6766
rect 12523 6732 12557 6744
rect 12523 6676 12557 6694
rect 12523 6660 12557 6676
rect 12523 6608 12557 6622
rect 12523 6588 12557 6608
rect 12523 6540 12557 6550
rect 12523 6516 12557 6540
rect 12523 6472 12557 6478
rect 12523 6444 12557 6472
rect 12523 6404 12557 6406
rect 12523 6372 12557 6404
rect 12523 6302 12557 6334
rect 12523 6300 12557 6302
rect 12523 6234 12557 6262
rect 12523 6228 12557 6234
rect 12523 6166 12557 6190
rect 12523 6156 12557 6166
rect 12523 6098 12557 6118
rect 12523 6084 12557 6098
rect 12523 6030 12557 6046
rect 12523 6012 12557 6030
rect 12523 5962 12557 5974
rect 12523 5940 12557 5962
rect 12523 5894 12557 5902
rect 12523 5868 12557 5894
rect 12609 6812 12643 6838
rect 12609 6804 12643 6812
rect 12609 6744 12643 6766
rect 12609 6732 12643 6744
rect 12609 6676 12643 6694
rect 12609 6660 12643 6676
rect 12609 6608 12643 6622
rect 12609 6588 12643 6608
rect 12609 6540 12643 6550
rect 12609 6516 12643 6540
rect 12609 6472 12643 6478
rect 12609 6444 12643 6472
rect 12609 6404 12643 6406
rect 12609 6372 12643 6404
rect 12609 6302 12643 6334
rect 12609 6300 12643 6302
rect 12609 6234 12643 6262
rect 12609 6228 12643 6234
rect 12609 6166 12643 6190
rect 12609 6156 12643 6166
rect 12609 6098 12643 6118
rect 12609 6084 12643 6098
rect 12609 6030 12643 6046
rect 12609 6012 12643 6030
rect 12609 5962 12643 5974
rect 12609 5940 12643 5962
rect 12609 5894 12643 5902
rect 12609 5868 12643 5894
rect 12695 6812 12729 6838
rect 12695 6804 12729 6812
rect 12695 6744 12729 6766
rect 12695 6732 12729 6744
rect 12695 6676 12729 6694
rect 12695 6660 12729 6676
rect 12695 6608 12729 6622
rect 12695 6588 12729 6608
rect 12695 6540 12729 6550
rect 12695 6516 12729 6540
rect 12695 6472 12729 6478
rect 12695 6444 12729 6472
rect 12695 6404 12729 6406
rect 12695 6372 12729 6404
rect 12695 6302 12729 6334
rect 12695 6300 12729 6302
rect 12695 6234 12729 6262
rect 12695 6228 12729 6234
rect 12695 6166 12729 6190
rect 12695 6156 12729 6166
rect 12695 6098 12729 6118
rect 12695 6084 12729 6098
rect 12695 6030 12729 6046
rect 12695 6012 12729 6030
rect 12695 5962 12729 5974
rect 12695 5940 12729 5962
rect 12695 5894 12729 5902
rect 12695 5868 12729 5894
rect 12806 6812 12840 6838
rect 12806 6804 12840 6812
rect 12806 6744 12840 6766
rect 12806 6732 12840 6744
rect 12806 6676 12840 6694
rect 12806 6660 12840 6676
rect 12806 6608 12840 6622
rect 12806 6588 12840 6608
rect 12806 6540 12840 6550
rect 12806 6516 12840 6540
rect 12806 6472 12840 6478
rect 12806 6444 12840 6472
rect 12806 6404 12840 6406
rect 12806 6372 12840 6404
rect 12806 6302 12840 6334
rect 12806 6300 12840 6302
rect 12806 6234 12840 6262
rect 12806 6228 12840 6234
rect 12806 6166 12840 6190
rect 12806 6156 12840 6166
rect 12806 6098 12840 6118
rect 12806 6084 12840 6098
rect 12806 6030 12840 6046
rect 12806 6012 12840 6030
rect 12806 5962 12840 5974
rect 12806 5940 12840 5962
rect 12806 5894 12840 5902
rect 12806 5868 12840 5894
rect 12917 6812 12951 6838
rect 12917 6804 12951 6812
rect 12917 6744 12951 6766
rect 12917 6732 12951 6744
rect 12917 6676 12951 6694
rect 12917 6660 12951 6676
rect 12917 6608 12951 6622
rect 12917 6588 12951 6608
rect 12917 6540 12951 6550
rect 12917 6516 12951 6540
rect 12917 6472 12951 6478
rect 12917 6444 12951 6472
rect 12917 6404 12951 6406
rect 12917 6372 12951 6404
rect 12917 6302 12951 6334
rect 12917 6300 12951 6302
rect 12917 6234 12951 6262
rect 12917 6228 12951 6234
rect 12917 6166 12951 6190
rect 12917 6156 12951 6166
rect 12917 6098 12951 6118
rect 12917 6084 12951 6098
rect 12917 6030 12951 6046
rect 12917 6012 12951 6030
rect 12917 5962 12951 5974
rect 12917 5940 12951 5962
rect 12917 5894 12951 5902
rect 12917 5868 12951 5894
rect 13003 6812 13037 6838
rect 13003 6804 13037 6812
rect 13003 6744 13037 6766
rect 13003 6732 13037 6744
rect 13003 6676 13037 6694
rect 13003 6660 13037 6676
rect 13003 6608 13037 6622
rect 13003 6588 13037 6608
rect 13003 6540 13037 6550
rect 13003 6516 13037 6540
rect 13003 6472 13037 6478
rect 13003 6444 13037 6472
rect 13003 6404 13037 6406
rect 13003 6372 13037 6404
rect 13003 6302 13037 6334
rect 13003 6300 13037 6302
rect 13003 6234 13037 6262
rect 13003 6228 13037 6234
rect 13003 6166 13037 6190
rect 13003 6156 13037 6166
rect 13003 6098 13037 6118
rect 13003 6084 13037 6098
rect 13003 6030 13037 6046
rect 13003 6012 13037 6030
rect 13003 5962 13037 5974
rect 13003 5940 13037 5962
rect 13003 5894 13037 5902
rect 13003 5868 13037 5894
rect 13089 6812 13123 6838
rect 13089 6804 13123 6812
rect 13089 6744 13123 6766
rect 13089 6732 13123 6744
rect 13089 6676 13123 6694
rect 13089 6660 13123 6676
rect 13089 6608 13123 6622
rect 13089 6588 13123 6608
rect 13089 6540 13123 6550
rect 13089 6516 13123 6540
rect 13089 6472 13123 6478
rect 13089 6444 13123 6472
rect 13089 6404 13123 6406
rect 13089 6372 13123 6404
rect 13089 6302 13123 6334
rect 13089 6300 13123 6302
rect 13089 6234 13123 6262
rect 13089 6228 13123 6234
rect 13089 6166 13123 6190
rect 13089 6156 13123 6166
rect 13089 6098 13123 6118
rect 13089 6084 13123 6098
rect 13089 6030 13123 6046
rect 13089 6012 13123 6030
rect 13089 5962 13123 5974
rect 13089 5940 13123 5962
rect 13089 5894 13123 5902
rect 13089 5868 13123 5894
rect 13175 6812 13209 6838
rect 13175 6804 13209 6812
rect 13175 6744 13209 6766
rect 13175 6732 13209 6744
rect 13175 6676 13209 6694
rect 13175 6660 13209 6676
rect 13175 6608 13209 6622
rect 13175 6588 13209 6608
rect 13175 6540 13209 6550
rect 13175 6516 13209 6540
rect 13175 6472 13209 6478
rect 13175 6444 13209 6472
rect 13175 6404 13209 6406
rect 13175 6372 13209 6404
rect 13175 6302 13209 6334
rect 13175 6300 13209 6302
rect 13175 6234 13209 6262
rect 13175 6228 13209 6234
rect 13175 6166 13209 6190
rect 13175 6156 13209 6166
rect 13175 6098 13209 6118
rect 13175 6084 13209 6098
rect 13175 6030 13209 6046
rect 13175 6012 13209 6030
rect 13175 5962 13209 5974
rect 13175 5940 13209 5962
rect 13175 5894 13209 5902
rect 13175 5868 13209 5894
rect 13261 6812 13295 6838
rect 13261 6804 13295 6812
rect 13261 6744 13295 6766
rect 13261 6732 13295 6744
rect 13261 6676 13295 6694
rect 13261 6660 13295 6676
rect 13261 6608 13295 6622
rect 13261 6588 13295 6608
rect 13261 6540 13295 6550
rect 13261 6516 13295 6540
rect 13261 6472 13295 6478
rect 13261 6444 13295 6472
rect 13261 6404 13295 6406
rect 13261 6372 13295 6404
rect 13261 6302 13295 6334
rect 13261 6300 13295 6302
rect 13261 6234 13295 6262
rect 13261 6228 13295 6234
rect 13261 6166 13295 6190
rect 13261 6156 13295 6166
rect 13261 6098 13295 6118
rect 13261 6084 13295 6098
rect 13261 6030 13295 6046
rect 13261 6012 13295 6030
rect 13261 5962 13295 5974
rect 13261 5940 13295 5962
rect 13261 5894 13295 5902
rect 13261 5868 13295 5894
rect 13372 6812 13406 6838
rect 13372 6804 13406 6812
rect 13372 6744 13406 6766
rect 13372 6732 13406 6744
rect 13372 6676 13406 6694
rect 13372 6660 13406 6676
rect 13372 6608 13406 6622
rect 13372 6588 13406 6608
rect 13372 6540 13406 6550
rect 13372 6516 13406 6540
rect 13372 6472 13406 6478
rect 13372 6444 13406 6472
rect 13372 6404 13406 6406
rect 13372 6372 13406 6404
rect 13372 6302 13406 6334
rect 13372 6300 13406 6302
rect 13372 6234 13406 6262
rect 13372 6228 13406 6234
rect 13372 6166 13406 6190
rect 13372 6156 13406 6166
rect 13372 6098 13406 6118
rect 13372 6084 13406 6098
rect 13372 6030 13406 6046
rect 13372 6012 13406 6030
rect 13372 5962 13406 5974
rect 13372 5940 13406 5962
rect 13372 5894 13406 5902
rect 13372 5868 13406 5894
rect 13483 6812 13517 6838
rect 13483 6804 13517 6812
rect 13483 6744 13517 6766
rect 13483 6732 13517 6744
rect 13483 6676 13517 6694
rect 13483 6660 13517 6676
rect 13483 6608 13517 6622
rect 13483 6588 13517 6608
rect 13483 6540 13517 6550
rect 13483 6516 13517 6540
rect 13483 6472 13517 6478
rect 13483 6444 13517 6472
rect 13483 6404 13517 6406
rect 13483 6372 13517 6404
rect 13483 6302 13517 6334
rect 13483 6300 13517 6302
rect 13483 6234 13517 6262
rect 13483 6228 13517 6234
rect 13483 6166 13517 6190
rect 13483 6156 13517 6166
rect 13483 6098 13517 6118
rect 13483 6084 13517 6098
rect 13483 6030 13517 6046
rect 13483 6012 13517 6030
rect 13483 5962 13517 5974
rect 13483 5940 13517 5962
rect 13483 5894 13517 5902
rect 13483 5868 13517 5894
rect 13569 6812 13603 6838
rect 13569 6804 13603 6812
rect 13569 6744 13603 6766
rect 13569 6732 13603 6744
rect 13569 6676 13603 6694
rect 13569 6660 13603 6676
rect 13569 6608 13603 6622
rect 13569 6588 13603 6608
rect 13569 6540 13603 6550
rect 13569 6516 13603 6540
rect 13569 6472 13603 6478
rect 13569 6444 13603 6472
rect 13569 6404 13603 6406
rect 13569 6372 13603 6404
rect 13569 6302 13603 6334
rect 13569 6300 13603 6302
rect 13569 6234 13603 6262
rect 13569 6228 13603 6234
rect 13569 6166 13603 6190
rect 13569 6156 13603 6166
rect 13569 6098 13603 6118
rect 13569 6084 13603 6098
rect 13569 6030 13603 6046
rect 13569 6012 13603 6030
rect 13569 5962 13603 5974
rect 13569 5940 13603 5962
rect 13569 5894 13603 5902
rect 13569 5868 13603 5894
rect 13655 6812 13689 6838
rect 13655 6804 13689 6812
rect 13655 6744 13689 6766
rect 13655 6732 13689 6744
rect 13655 6676 13689 6694
rect 13655 6660 13689 6676
rect 13655 6608 13689 6622
rect 13655 6588 13689 6608
rect 13655 6540 13689 6550
rect 13655 6516 13689 6540
rect 13655 6472 13689 6478
rect 13655 6444 13689 6472
rect 13655 6404 13689 6406
rect 13655 6372 13689 6404
rect 13655 6302 13689 6334
rect 13655 6300 13689 6302
rect 13655 6234 13689 6262
rect 13655 6228 13689 6234
rect 13655 6166 13689 6190
rect 13655 6156 13689 6166
rect 13655 6098 13689 6118
rect 13655 6084 13689 6098
rect 13655 6030 13689 6046
rect 13655 6012 13689 6030
rect 13655 5962 13689 5974
rect 13655 5940 13689 5962
rect 13655 5894 13689 5902
rect 13655 5868 13689 5894
rect 13741 6812 13775 6838
rect 13741 6804 13775 6812
rect 13741 6744 13775 6766
rect 13741 6732 13775 6744
rect 13741 6676 13775 6694
rect 13741 6660 13775 6676
rect 13741 6608 13775 6622
rect 13741 6588 13775 6608
rect 13741 6540 13775 6550
rect 13741 6516 13775 6540
rect 13741 6472 13775 6478
rect 13741 6444 13775 6472
rect 13741 6404 13775 6406
rect 13741 6372 13775 6404
rect 13741 6302 13775 6334
rect 13741 6300 13775 6302
rect 13741 6234 13775 6262
rect 13741 6228 13775 6234
rect 13741 6166 13775 6190
rect 13741 6156 13775 6166
rect 13741 6098 13775 6118
rect 13741 6084 13775 6098
rect 13741 6030 13775 6046
rect 13741 6012 13775 6030
rect 13741 5962 13775 5974
rect 13741 5940 13775 5962
rect 13741 5894 13775 5902
rect 13741 5868 13775 5894
rect 13827 6812 13861 6838
rect 13827 6804 13861 6812
rect 13827 6744 13861 6766
rect 13827 6732 13861 6744
rect 13827 6676 13861 6694
rect 13827 6660 13861 6676
rect 13827 6608 13861 6622
rect 13827 6588 13861 6608
rect 13827 6540 13861 6550
rect 13827 6516 13861 6540
rect 13827 6472 13861 6478
rect 13827 6444 13861 6472
rect 13827 6404 13861 6406
rect 13827 6372 13861 6404
rect 13827 6302 13861 6334
rect 13827 6300 13861 6302
rect 13827 6234 13861 6262
rect 13827 6228 13861 6234
rect 13827 6166 13861 6190
rect 13827 6156 13861 6166
rect 13827 6098 13861 6118
rect 13827 6084 13861 6098
rect 13827 6030 13861 6046
rect 13827 6012 13861 6030
rect 13827 5962 13861 5974
rect 13827 5940 13861 5962
rect 13827 5894 13861 5902
rect 13827 5868 13861 5894
rect 13938 6812 13972 6838
rect 13938 6804 13972 6812
rect 13938 6744 13972 6766
rect 13938 6732 13972 6744
rect 13938 6676 13972 6694
rect 13938 6660 13972 6676
rect 13938 6608 13972 6622
rect 13938 6588 13972 6608
rect 13938 6540 13972 6550
rect 13938 6516 13972 6540
rect 13938 6472 13972 6478
rect 13938 6444 13972 6472
rect 13938 6404 13972 6406
rect 13938 6372 13972 6404
rect 13938 6302 13972 6334
rect 13938 6300 13972 6302
rect 13938 6234 13972 6262
rect 13938 6228 13972 6234
rect 13938 6166 13972 6190
rect 13938 6156 13972 6166
rect 13938 6098 13972 6118
rect 13938 6084 13972 6098
rect 13938 6030 13972 6046
rect 13938 6012 13972 6030
rect 13938 5962 13972 5974
rect 13938 5940 13972 5962
rect 13938 5894 13972 5902
rect 13938 5868 13972 5894
rect 14049 6812 14083 6838
rect 14049 6804 14083 6812
rect 14049 6744 14083 6766
rect 14049 6732 14083 6744
rect 14049 6676 14083 6694
rect 14049 6660 14083 6676
rect 14049 6608 14083 6622
rect 14049 6588 14083 6608
rect 14049 6540 14083 6550
rect 14049 6516 14083 6540
rect 14049 6472 14083 6478
rect 14049 6444 14083 6472
rect 14049 6404 14083 6406
rect 14049 6372 14083 6404
rect 14049 6302 14083 6334
rect 14049 6300 14083 6302
rect 14049 6234 14083 6262
rect 14049 6228 14083 6234
rect 14049 6166 14083 6190
rect 14049 6156 14083 6166
rect 14049 6098 14083 6118
rect 14049 6084 14083 6098
rect 14049 6030 14083 6046
rect 14049 6012 14083 6030
rect 14049 5962 14083 5974
rect 14049 5940 14083 5962
rect 14049 5894 14083 5902
rect 14049 5868 14083 5894
rect 14135 6812 14169 6838
rect 14135 6804 14169 6812
rect 14135 6744 14169 6766
rect 14135 6732 14169 6744
rect 14135 6676 14169 6694
rect 14135 6660 14169 6676
rect 14135 6608 14169 6622
rect 14135 6588 14169 6608
rect 14135 6540 14169 6550
rect 14135 6516 14169 6540
rect 14135 6472 14169 6478
rect 14135 6444 14169 6472
rect 14135 6404 14169 6406
rect 14135 6372 14169 6404
rect 14135 6302 14169 6334
rect 14135 6300 14169 6302
rect 14135 6234 14169 6262
rect 14135 6228 14169 6234
rect 14135 6166 14169 6190
rect 14135 6156 14169 6166
rect 14135 6098 14169 6118
rect 14135 6084 14169 6098
rect 14135 6030 14169 6046
rect 14135 6012 14169 6030
rect 14135 5962 14169 5974
rect 14135 5940 14169 5962
rect 14135 5894 14169 5902
rect 14135 5868 14169 5894
rect 14221 6812 14255 6838
rect 14221 6804 14255 6812
rect 14221 6744 14255 6766
rect 14221 6732 14255 6744
rect 14221 6676 14255 6694
rect 14221 6660 14255 6676
rect 14221 6608 14255 6622
rect 14221 6588 14255 6608
rect 14221 6540 14255 6550
rect 14221 6516 14255 6540
rect 14221 6472 14255 6478
rect 14221 6444 14255 6472
rect 14221 6404 14255 6406
rect 14221 6372 14255 6404
rect 14221 6302 14255 6334
rect 14221 6300 14255 6302
rect 14221 6234 14255 6262
rect 14221 6228 14255 6234
rect 14221 6166 14255 6190
rect 14221 6156 14255 6166
rect 14221 6098 14255 6118
rect 14221 6084 14255 6098
rect 14221 6030 14255 6046
rect 14221 6012 14255 6030
rect 14221 5962 14255 5974
rect 14221 5940 14255 5962
rect 14221 5894 14255 5902
rect 14221 5868 14255 5894
rect 14307 6812 14341 6838
rect 14307 6804 14341 6812
rect 14307 6744 14341 6766
rect 14307 6732 14341 6744
rect 14307 6676 14341 6694
rect 14307 6660 14341 6676
rect 14307 6608 14341 6622
rect 14307 6588 14341 6608
rect 14307 6540 14341 6550
rect 14307 6516 14341 6540
rect 14307 6472 14341 6478
rect 14307 6444 14341 6472
rect 14307 6404 14341 6406
rect 14307 6372 14341 6404
rect 14307 6302 14341 6334
rect 14307 6300 14341 6302
rect 14307 6234 14341 6262
rect 14307 6228 14341 6234
rect 14307 6166 14341 6190
rect 14307 6156 14341 6166
rect 14307 6098 14341 6118
rect 14307 6084 14341 6098
rect 14307 6030 14341 6046
rect 14307 6012 14341 6030
rect 14307 5962 14341 5974
rect 14307 5940 14341 5962
rect 14307 5894 14341 5902
rect 14307 5868 14341 5894
rect 14393 6812 14427 6838
rect 14393 6804 14427 6812
rect 14393 6744 14427 6766
rect 14393 6732 14427 6744
rect 14393 6676 14427 6694
rect 14393 6660 14427 6676
rect 14393 6608 14427 6622
rect 14393 6588 14427 6608
rect 14393 6540 14427 6550
rect 14393 6516 14427 6540
rect 14393 6472 14427 6478
rect 14393 6444 14427 6472
rect 14393 6404 14427 6406
rect 14393 6372 14427 6404
rect 14393 6302 14427 6334
rect 14393 6300 14427 6302
rect 14393 6234 14427 6262
rect 14393 6228 14427 6234
rect 14393 6166 14427 6190
rect 14393 6156 14427 6166
rect 14393 6098 14427 6118
rect 14393 6084 14427 6098
rect 14393 6030 14427 6046
rect 14393 6012 14427 6030
rect 14393 5962 14427 5974
rect 14393 5940 14427 5962
rect 14393 5894 14427 5902
rect 14393 5868 14427 5894
rect 14504 6812 14538 6838
rect 14504 6804 14538 6812
rect 14504 6744 14538 6766
rect 14504 6732 14538 6744
rect 14504 6676 14538 6694
rect 14504 6660 14538 6676
rect 14504 6608 14538 6622
rect 14504 6588 14538 6608
rect 14504 6540 14538 6550
rect 14504 6516 14538 6540
rect 14504 6472 14538 6478
rect 14504 6444 14538 6472
rect 14504 6404 14538 6406
rect 14504 6372 14538 6404
rect 14504 6302 14538 6334
rect 14504 6300 14538 6302
rect 14504 6234 14538 6262
rect 14504 6228 14538 6234
rect 14504 6166 14538 6190
rect 14504 6156 14538 6166
rect 14504 6098 14538 6118
rect 14504 6084 14538 6098
rect 14504 6030 14538 6046
rect 14504 6012 14538 6030
rect 14504 5962 14538 5974
rect 14504 5940 14538 5962
rect 14504 5894 14538 5902
rect 14504 5868 14538 5894
rect 14615 6812 14649 6838
rect 14615 6804 14649 6812
rect 14615 6744 14649 6766
rect 14615 6732 14649 6744
rect 14615 6676 14649 6694
rect 14615 6660 14649 6676
rect 14615 6608 14649 6622
rect 14615 6588 14649 6608
rect 14615 6540 14649 6550
rect 14615 6516 14649 6540
rect 14615 6472 14649 6478
rect 14615 6444 14649 6472
rect 14615 6404 14649 6406
rect 14615 6372 14649 6404
rect 14615 6302 14649 6334
rect 14615 6300 14649 6302
rect 14615 6234 14649 6262
rect 14615 6228 14649 6234
rect 14615 6166 14649 6190
rect 14615 6156 14649 6166
rect 14615 6098 14649 6118
rect 14615 6084 14649 6098
rect 14615 6030 14649 6046
rect 14615 6012 14649 6030
rect 14615 5962 14649 5974
rect 14615 5940 14649 5962
rect 14615 5894 14649 5902
rect 14615 5868 14649 5894
rect 14701 6812 14735 6838
rect 14701 6804 14735 6812
rect 14701 6744 14735 6766
rect 14701 6732 14735 6744
rect 14701 6676 14735 6694
rect 14701 6660 14735 6676
rect 14701 6608 14735 6622
rect 14701 6588 14735 6608
rect 14701 6540 14735 6550
rect 14701 6516 14735 6540
rect 14701 6472 14735 6478
rect 14701 6444 14735 6472
rect 14701 6404 14735 6406
rect 14701 6372 14735 6404
rect 14701 6302 14735 6334
rect 14701 6300 14735 6302
rect 14701 6234 14735 6262
rect 14701 6228 14735 6234
rect 14701 6166 14735 6190
rect 14701 6156 14735 6166
rect 14701 6098 14735 6118
rect 14701 6084 14735 6098
rect 14701 6030 14735 6046
rect 14701 6012 14735 6030
rect 14701 5962 14735 5974
rect 14701 5940 14735 5962
rect 14701 5894 14735 5902
rect 14701 5868 14735 5894
rect 14787 6812 14821 6838
rect 14787 6804 14821 6812
rect 14787 6744 14821 6766
rect 14787 6732 14821 6744
rect 14787 6676 14821 6694
rect 14787 6660 14821 6676
rect 14787 6608 14821 6622
rect 14787 6588 14821 6608
rect 14787 6540 14821 6550
rect 14787 6516 14821 6540
rect 14787 6472 14821 6478
rect 14787 6444 14821 6472
rect 14787 6404 14821 6406
rect 14787 6372 14821 6404
rect 14787 6302 14821 6334
rect 14787 6300 14821 6302
rect 14787 6234 14821 6262
rect 14787 6228 14821 6234
rect 14787 6166 14821 6190
rect 14787 6156 14821 6166
rect 14787 6098 14821 6118
rect 14787 6084 14821 6098
rect 14787 6030 14821 6046
rect 14787 6012 14821 6030
rect 14787 5962 14821 5974
rect 14787 5940 14821 5962
rect 14787 5894 14821 5902
rect 14787 5868 14821 5894
rect 14873 6812 14907 6838
rect 14873 6804 14907 6812
rect 14873 6744 14907 6766
rect 14873 6732 14907 6744
rect 14873 6676 14907 6694
rect 14873 6660 14907 6676
rect 14873 6608 14907 6622
rect 14873 6588 14907 6608
rect 14873 6540 14907 6550
rect 14873 6516 14907 6540
rect 14873 6472 14907 6478
rect 14873 6444 14907 6472
rect 14873 6404 14907 6406
rect 14873 6372 14907 6404
rect 14873 6302 14907 6334
rect 14873 6300 14907 6302
rect 14873 6234 14907 6262
rect 14873 6228 14907 6234
rect 14873 6166 14907 6190
rect 14873 6156 14907 6166
rect 14873 6098 14907 6118
rect 14873 6084 14907 6098
rect 14873 6030 14907 6046
rect 14873 6012 14907 6030
rect 14873 5962 14907 5974
rect 14873 5940 14907 5962
rect 14873 5894 14907 5902
rect 14873 5868 14907 5894
rect 14959 6812 14993 6838
rect 14959 6804 14993 6812
rect 14959 6744 14993 6766
rect 14959 6732 14993 6744
rect 14959 6676 14993 6694
rect 14959 6660 14993 6676
rect 14959 6608 14993 6622
rect 14959 6588 14993 6608
rect 14959 6540 14993 6550
rect 14959 6516 14993 6540
rect 14959 6472 14993 6478
rect 14959 6444 14993 6472
rect 14959 6404 14993 6406
rect 14959 6372 14993 6404
rect 14959 6302 14993 6334
rect 14959 6300 14993 6302
rect 14959 6234 14993 6262
rect 14959 6228 14993 6234
rect 14959 6166 14993 6190
rect 14959 6156 14993 6166
rect 14959 6098 14993 6118
rect 14959 6084 14993 6098
rect 14959 6030 14993 6046
rect 14959 6012 14993 6030
rect 14959 5962 14993 5974
rect 14959 5940 14993 5962
rect 14959 5894 14993 5902
rect 14959 5868 14993 5894
rect 15070 6812 15104 6838
rect 15070 6804 15104 6812
rect 15070 6744 15104 6766
rect 15070 6732 15104 6744
rect 15070 6676 15104 6694
rect 15070 6660 15104 6676
rect 15070 6608 15104 6622
rect 15070 6588 15104 6608
rect 15070 6540 15104 6550
rect 15070 6516 15104 6540
rect 15070 6472 15104 6478
rect 15070 6444 15104 6472
rect 15070 6404 15104 6406
rect 15070 6372 15104 6404
rect 15070 6302 15104 6334
rect 15070 6300 15104 6302
rect 15070 6234 15104 6262
rect 15070 6228 15104 6234
rect 15070 6166 15104 6190
rect 15070 6156 15104 6166
rect 15070 6098 15104 6118
rect 15070 6084 15104 6098
rect 15070 6030 15104 6046
rect 15070 6012 15104 6030
rect 15070 5962 15104 5974
rect 15070 5940 15104 5962
rect 15070 5894 15104 5902
rect 15070 5868 15104 5894
rect 15181 6812 15215 6838
rect 15181 6804 15215 6812
rect 15181 6744 15215 6766
rect 15181 6732 15215 6744
rect 15181 6676 15215 6694
rect 15181 6660 15215 6676
rect 15181 6608 15215 6622
rect 15181 6588 15215 6608
rect 15181 6540 15215 6550
rect 15181 6516 15215 6540
rect 15181 6472 15215 6478
rect 15181 6444 15215 6472
rect 15181 6404 15215 6406
rect 15181 6372 15215 6404
rect 15181 6302 15215 6334
rect 15181 6300 15215 6302
rect 15181 6234 15215 6262
rect 15181 6228 15215 6234
rect 15181 6166 15215 6190
rect 15181 6156 15215 6166
rect 15181 6098 15215 6118
rect 15181 6084 15215 6098
rect 15181 6030 15215 6046
rect 15181 6012 15215 6030
rect 15181 5962 15215 5974
rect 15181 5940 15215 5962
rect 15181 5894 15215 5902
rect 15181 5868 15215 5894
rect 15267 6812 15301 6838
rect 15267 6804 15301 6812
rect 15267 6744 15301 6766
rect 15267 6732 15301 6744
rect 15267 6676 15301 6694
rect 15267 6660 15301 6676
rect 15267 6608 15301 6622
rect 15267 6588 15301 6608
rect 15267 6540 15301 6550
rect 15267 6516 15301 6540
rect 15267 6472 15301 6478
rect 15267 6444 15301 6472
rect 15267 6404 15301 6406
rect 15267 6372 15301 6404
rect 15267 6302 15301 6334
rect 15267 6300 15301 6302
rect 15267 6234 15301 6262
rect 15267 6228 15301 6234
rect 15267 6166 15301 6190
rect 15267 6156 15301 6166
rect 15267 6098 15301 6118
rect 15267 6084 15301 6098
rect 15267 6030 15301 6046
rect 15267 6012 15301 6030
rect 15267 5962 15301 5974
rect 15267 5940 15301 5962
rect 15267 5894 15301 5902
rect 15267 5868 15301 5894
rect 15353 6812 15387 6838
rect 15353 6804 15387 6812
rect 15353 6744 15387 6766
rect 15353 6732 15387 6744
rect 15353 6676 15387 6694
rect 15353 6660 15387 6676
rect 15353 6608 15387 6622
rect 15353 6588 15387 6608
rect 15353 6540 15387 6550
rect 15353 6516 15387 6540
rect 15353 6472 15387 6478
rect 15353 6444 15387 6472
rect 15353 6404 15387 6406
rect 15353 6372 15387 6404
rect 15353 6302 15387 6334
rect 15353 6300 15387 6302
rect 15353 6234 15387 6262
rect 15353 6228 15387 6234
rect 15353 6166 15387 6190
rect 15353 6156 15387 6166
rect 15353 6098 15387 6118
rect 15353 6084 15387 6098
rect 15353 6030 15387 6046
rect 15353 6012 15387 6030
rect 15353 5962 15387 5974
rect 15353 5940 15387 5962
rect 15353 5894 15387 5902
rect 15353 5868 15387 5894
rect 15439 6812 15473 6838
rect 15439 6804 15473 6812
rect 15439 6744 15473 6766
rect 15439 6732 15473 6744
rect 15439 6676 15473 6694
rect 15439 6660 15473 6676
rect 15439 6608 15473 6622
rect 15439 6588 15473 6608
rect 15439 6540 15473 6550
rect 15439 6516 15473 6540
rect 15439 6472 15473 6478
rect 15439 6444 15473 6472
rect 15439 6404 15473 6406
rect 15439 6372 15473 6404
rect 15439 6302 15473 6334
rect 15439 6300 15473 6302
rect 15439 6234 15473 6262
rect 15439 6228 15473 6234
rect 15439 6166 15473 6190
rect 15439 6156 15473 6166
rect 15439 6098 15473 6118
rect 15439 6084 15473 6098
rect 15439 6030 15473 6046
rect 15439 6012 15473 6030
rect 15439 5962 15473 5974
rect 15439 5940 15473 5962
rect 15439 5894 15473 5902
rect 15439 5868 15473 5894
rect 18030 6874 18036 6908
rect 18036 6874 18064 6908
rect 18102 6874 18104 6908
rect 18104 6874 18136 6908
rect 18174 6874 18206 6908
rect 18206 6874 18208 6908
rect 18246 6874 18274 6908
rect 18274 6874 18280 6908
rect 18374 6874 18380 6908
rect 18380 6874 18408 6908
rect 18446 6874 18448 6908
rect 18448 6874 18480 6908
rect 18518 6874 18550 6908
rect 18550 6874 18552 6908
rect 18590 6874 18618 6908
rect 18618 6874 18624 6908
rect 18718 6874 18724 6908
rect 18724 6874 18752 6908
rect 18790 6874 18792 6908
rect 18792 6874 18824 6908
rect 18862 6874 18894 6908
rect 18894 6874 18896 6908
rect 18934 6874 18962 6908
rect 18962 6874 18968 6908
rect 19062 6874 19068 6908
rect 19068 6874 19096 6908
rect 19134 6874 19136 6908
rect 19136 6874 19168 6908
rect 19206 6874 19238 6908
rect 19238 6874 19240 6908
rect 19278 6874 19306 6908
rect 19306 6874 19312 6908
rect 19406 6874 19412 6908
rect 19412 6874 19440 6908
rect 19478 6874 19480 6908
rect 19480 6874 19512 6908
rect 19550 6874 19582 6908
rect 19582 6874 19584 6908
rect 19622 6874 19650 6908
rect 19650 6874 19656 6908
rect 19750 6874 19756 6908
rect 19756 6874 19784 6908
rect 19822 6874 19824 6908
rect 19824 6874 19856 6908
rect 19894 6874 19926 6908
rect 19926 6874 19928 6908
rect 19966 6874 19994 6908
rect 19994 6874 20000 6908
rect 15525 6812 15559 6838
rect 15525 6804 15559 6812
rect 15525 6744 15559 6766
rect 15525 6732 15559 6744
rect 15525 6676 15559 6694
rect 15525 6660 15559 6676
rect 15525 6608 15559 6622
rect 15525 6588 15559 6608
rect 15525 6540 15559 6550
rect 15525 6516 15559 6540
rect 15525 6472 15559 6478
rect 15525 6444 15559 6472
rect 15525 6404 15559 6406
rect 15525 6372 15559 6404
rect 15525 6302 15559 6334
rect 15525 6300 15559 6302
rect 15525 6234 15559 6262
rect 15525 6228 15559 6234
rect 15525 6166 15559 6190
rect 15525 6156 15559 6166
rect 15525 6098 15559 6118
rect 15525 6084 15559 6098
rect 15525 6030 15559 6046
rect 15525 6012 15559 6030
rect 15525 5962 15559 5974
rect 15525 5940 15559 5962
rect 15525 5894 15559 5902
rect 15525 5868 15559 5894
rect 15636 6812 15670 6838
rect 15636 6804 15670 6812
rect 15636 6744 15670 6766
rect 15636 6732 15670 6744
rect 15636 6676 15670 6694
rect 15636 6660 15670 6676
rect 15636 6608 15670 6622
rect 15636 6588 15670 6608
rect 15636 6540 15670 6550
rect 15636 6516 15670 6540
rect 15636 6472 15670 6478
rect 15636 6444 15670 6472
rect 15636 6404 15670 6406
rect 15636 6372 15670 6404
rect 15636 6302 15670 6334
rect 15636 6300 15670 6302
rect 17668 6282 17674 6316
rect 17674 6282 17702 6316
rect 17740 6282 17742 6316
rect 17742 6282 17774 6316
rect 17812 6282 17844 6316
rect 17844 6282 17846 6316
rect 17884 6282 17912 6316
rect 17912 6282 17918 6316
rect 18012 6282 18018 6316
rect 18018 6282 18046 6316
rect 18084 6282 18086 6316
rect 18086 6282 18118 6316
rect 18156 6282 18188 6316
rect 18188 6282 18190 6316
rect 18228 6282 18256 6316
rect 18256 6282 18262 6316
rect 18356 6282 18362 6316
rect 18362 6282 18390 6316
rect 18428 6282 18430 6316
rect 18430 6282 18462 6316
rect 18500 6282 18532 6316
rect 18532 6282 18534 6316
rect 18572 6282 18600 6316
rect 18600 6282 18606 6316
rect 18700 6282 18706 6316
rect 18706 6282 18734 6316
rect 18772 6282 18774 6316
rect 18774 6282 18806 6316
rect 18844 6282 18876 6316
rect 18876 6282 18878 6316
rect 18916 6282 18944 6316
rect 18944 6282 18950 6316
rect 19044 6282 19050 6316
rect 19050 6282 19078 6316
rect 19116 6282 19118 6316
rect 19118 6282 19150 6316
rect 19188 6282 19220 6316
rect 19220 6282 19222 6316
rect 19260 6282 19288 6316
rect 19288 6282 19294 6316
rect 19388 6282 19394 6316
rect 19394 6282 19422 6316
rect 19460 6282 19462 6316
rect 19462 6282 19494 6316
rect 19532 6282 19564 6316
rect 19564 6282 19566 6316
rect 19604 6282 19632 6316
rect 19632 6282 19638 6316
rect 19732 6282 19738 6316
rect 19738 6282 19766 6316
rect 19804 6282 19806 6316
rect 19806 6282 19838 6316
rect 19876 6282 19908 6316
rect 19908 6282 19910 6316
rect 19948 6282 19976 6316
rect 19976 6282 19982 6316
rect 15636 6234 15670 6262
rect 15636 6228 15670 6234
rect 16218 6229 16222 6263
rect 16222 6229 16252 6263
rect 16290 6229 16324 6263
rect 16362 6229 16392 6263
rect 16392 6229 16396 6263
rect 16562 6229 16566 6263
rect 16566 6229 16596 6263
rect 16634 6229 16668 6263
rect 16706 6229 16736 6263
rect 16736 6229 16740 6263
rect 16906 6229 16910 6263
rect 16910 6229 16940 6263
rect 16978 6229 17012 6263
rect 17050 6229 17080 6263
rect 17080 6229 17084 6263
rect 15636 6166 15670 6190
rect 15636 6156 15670 6166
rect 15636 6098 15670 6118
rect 15636 6084 15670 6098
rect 15636 6030 15670 6046
rect 15636 6012 15670 6030
rect 15636 5962 15670 5974
rect 15636 5940 15670 5962
rect 15636 5894 15670 5902
rect 15636 5868 15670 5894
rect 15990 6120 16024 6154
rect 15990 6050 16024 6074
rect 15990 6040 16024 6050
rect 15990 5980 16024 5994
rect 15990 5960 16024 5980
rect 15990 5910 16024 5914
rect 15990 5880 16024 5910
rect 11813 5776 11821 5810
rect 11821 5776 11847 5810
rect 11885 5776 11889 5810
rect 11889 5776 11919 5810
rect 11957 5776 11991 5810
rect 12029 5776 12059 5810
rect 12059 5776 12063 5810
rect 12101 5776 12127 5810
rect 12127 5776 12135 5810
rect 12379 5776 12387 5810
rect 12387 5776 12413 5810
rect 12451 5776 12455 5810
rect 12455 5776 12485 5810
rect 12523 5776 12557 5810
rect 12595 5776 12625 5810
rect 12625 5776 12629 5810
rect 12667 5776 12693 5810
rect 12693 5776 12701 5810
rect 12945 5776 12953 5810
rect 12953 5776 12979 5810
rect 13017 5776 13021 5810
rect 13021 5776 13051 5810
rect 13089 5776 13123 5810
rect 13161 5776 13191 5810
rect 13191 5776 13195 5810
rect 13233 5776 13259 5810
rect 13259 5776 13267 5810
rect 13511 5776 13519 5810
rect 13519 5776 13545 5810
rect 13583 5776 13587 5810
rect 13587 5776 13617 5810
rect 13655 5776 13689 5810
rect 13727 5776 13757 5810
rect 13757 5776 13761 5810
rect 13799 5776 13825 5810
rect 13825 5776 13833 5810
rect 14077 5776 14085 5810
rect 14085 5776 14111 5810
rect 14149 5776 14153 5810
rect 14153 5776 14183 5810
rect 14221 5776 14255 5810
rect 14293 5776 14323 5810
rect 14323 5776 14327 5810
rect 14365 5776 14391 5810
rect 14391 5776 14399 5810
rect 14643 5776 14651 5810
rect 14651 5776 14677 5810
rect 14715 5776 14719 5810
rect 14719 5776 14749 5810
rect 14787 5776 14821 5810
rect 14859 5776 14889 5810
rect 14889 5776 14893 5810
rect 14931 5776 14957 5810
rect 14957 5776 14965 5810
rect 15209 5776 15217 5810
rect 15217 5776 15243 5810
rect 15281 5776 15285 5810
rect 15285 5776 15315 5810
rect 15353 5776 15387 5810
rect 15425 5776 15455 5810
rect 15455 5776 15459 5810
rect 15497 5776 15523 5810
rect 15523 5776 15531 5810
rect 15990 5804 16024 5834
rect 15990 5800 16024 5804
rect 15990 5734 16024 5754
rect 15990 5720 16024 5734
rect 15990 5664 16024 5674
rect 15990 5640 16024 5664
rect 15990 5560 16024 5594
rect 15990 5490 16024 5514
rect 15990 5480 16024 5490
rect 15990 5420 16024 5434
rect 15990 5400 16024 5420
rect 15990 5350 16024 5354
rect 15990 5320 16024 5350
rect 15990 5244 16024 5274
rect 15990 5240 16024 5244
rect 15990 5174 16024 5194
rect 15990 5160 16024 5174
rect 16118 6145 16152 6171
rect 16118 6137 16152 6145
rect 16118 6077 16152 6099
rect 16118 6065 16152 6077
rect 16118 6009 16152 6027
rect 16118 5993 16152 6009
rect 16118 5941 16152 5955
rect 16118 5921 16152 5941
rect 16118 5873 16152 5883
rect 16118 5849 16152 5873
rect 16118 5805 16152 5811
rect 16118 5777 16152 5805
rect 16118 5737 16152 5739
rect 16118 5705 16152 5737
rect 16118 5635 16152 5667
rect 16118 5633 16152 5635
rect 16118 5567 16152 5595
rect 16118 5561 16152 5567
rect 16118 5499 16152 5523
rect 16118 5489 16152 5499
rect 16118 5431 16152 5451
rect 16118 5417 16152 5431
rect 16118 5363 16152 5379
rect 16118 5345 16152 5363
rect 16118 5295 16152 5307
rect 16118 5273 16152 5295
rect 16118 5227 16152 5235
rect 16118 5201 16152 5227
rect 16204 6145 16238 6171
rect 16204 6137 16238 6145
rect 16204 6077 16238 6099
rect 16204 6065 16238 6077
rect 16204 6009 16238 6027
rect 16204 5993 16238 6009
rect 16204 5941 16238 5955
rect 16204 5921 16238 5941
rect 16204 5873 16238 5883
rect 16204 5849 16238 5873
rect 16204 5805 16238 5811
rect 16204 5777 16238 5805
rect 16204 5737 16238 5739
rect 16204 5705 16238 5737
rect 16204 5635 16238 5667
rect 16204 5633 16238 5635
rect 16204 5567 16238 5595
rect 16204 5561 16238 5567
rect 16204 5499 16238 5523
rect 16204 5489 16238 5499
rect 16204 5431 16238 5451
rect 16204 5417 16238 5431
rect 16204 5363 16238 5379
rect 16204 5345 16238 5363
rect 16204 5295 16238 5307
rect 16204 5273 16238 5295
rect 16204 5227 16238 5235
rect 16204 5201 16238 5227
rect 16290 6145 16324 6171
rect 16290 6137 16324 6145
rect 16290 6077 16324 6099
rect 16290 6065 16324 6077
rect 16290 6009 16324 6027
rect 16290 5993 16324 6009
rect 16290 5941 16324 5955
rect 16290 5921 16324 5941
rect 16290 5873 16324 5883
rect 16290 5849 16324 5873
rect 16290 5805 16324 5811
rect 16290 5777 16324 5805
rect 16290 5737 16324 5739
rect 16290 5705 16324 5737
rect 16290 5635 16324 5667
rect 16290 5633 16324 5635
rect 16290 5567 16324 5595
rect 16290 5561 16324 5567
rect 16290 5499 16324 5523
rect 16290 5489 16324 5499
rect 16290 5431 16324 5451
rect 16290 5417 16324 5431
rect 16290 5363 16324 5379
rect 16290 5345 16324 5363
rect 16290 5295 16324 5307
rect 16290 5273 16324 5295
rect 16290 5227 16324 5235
rect 16290 5201 16324 5227
rect 16376 6145 16410 6171
rect 16376 6137 16410 6145
rect 16376 6077 16410 6099
rect 16376 6065 16410 6077
rect 16376 6009 16410 6027
rect 16376 5993 16410 6009
rect 16376 5941 16410 5955
rect 16376 5921 16410 5941
rect 16376 5873 16410 5883
rect 16376 5849 16410 5873
rect 16376 5805 16410 5811
rect 16376 5777 16410 5805
rect 16376 5737 16410 5739
rect 16376 5705 16410 5737
rect 16376 5635 16410 5667
rect 16376 5633 16410 5635
rect 16376 5567 16410 5595
rect 16376 5561 16410 5567
rect 16376 5499 16410 5523
rect 16376 5489 16410 5499
rect 16376 5431 16410 5451
rect 16376 5417 16410 5431
rect 16376 5363 16410 5379
rect 16376 5345 16410 5363
rect 16376 5295 16410 5307
rect 16376 5273 16410 5295
rect 16376 5227 16410 5235
rect 16376 5201 16410 5227
rect 16462 6145 16496 6171
rect 16462 6137 16496 6145
rect 16462 6077 16496 6099
rect 16462 6065 16496 6077
rect 16462 6009 16496 6027
rect 16462 5993 16496 6009
rect 16462 5941 16496 5955
rect 16462 5921 16496 5941
rect 16462 5873 16496 5883
rect 16462 5849 16496 5873
rect 16462 5805 16496 5811
rect 16462 5777 16496 5805
rect 16462 5737 16496 5739
rect 16462 5705 16496 5737
rect 16462 5635 16496 5667
rect 16462 5633 16496 5635
rect 16462 5567 16496 5595
rect 16462 5561 16496 5567
rect 16462 5499 16496 5523
rect 16462 5489 16496 5499
rect 16462 5431 16496 5451
rect 16462 5417 16496 5431
rect 16462 5363 16496 5379
rect 16462 5345 16496 5363
rect 16462 5295 16496 5307
rect 16462 5273 16496 5295
rect 16462 5227 16496 5235
rect 16462 5201 16496 5227
rect 16548 6145 16582 6171
rect 16548 6137 16582 6145
rect 16548 6077 16582 6099
rect 16548 6065 16582 6077
rect 16548 6009 16582 6027
rect 16548 5993 16582 6009
rect 16548 5941 16582 5955
rect 16548 5921 16582 5941
rect 16548 5873 16582 5883
rect 16548 5849 16582 5873
rect 16548 5805 16582 5811
rect 16548 5777 16582 5805
rect 16548 5737 16582 5739
rect 16548 5705 16582 5737
rect 16548 5635 16582 5667
rect 16548 5633 16582 5635
rect 16548 5567 16582 5595
rect 16548 5561 16582 5567
rect 16548 5499 16582 5523
rect 16548 5489 16582 5499
rect 16548 5431 16582 5451
rect 16548 5417 16582 5431
rect 16548 5363 16582 5379
rect 16548 5345 16582 5363
rect 16548 5295 16582 5307
rect 16548 5273 16582 5295
rect 16548 5227 16582 5235
rect 16548 5201 16582 5227
rect 16634 6145 16668 6171
rect 16634 6137 16668 6145
rect 16634 6077 16668 6099
rect 16634 6065 16668 6077
rect 16634 6009 16668 6027
rect 16634 5993 16668 6009
rect 16634 5941 16668 5955
rect 16634 5921 16668 5941
rect 16634 5873 16668 5883
rect 16634 5849 16668 5873
rect 16634 5805 16668 5811
rect 16634 5777 16668 5805
rect 16634 5737 16668 5739
rect 16634 5705 16668 5737
rect 16634 5635 16668 5667
rect 16634 5633 16668 5635
rect 16634 5567 16668 5595
rect 16634 5561 16668 5567
rect 16634 5499 16668 5523
rect 16634 5489 16668 5499
rect 16634 5431 16668 5451
rect 16634 5417 16668 5431
rect 16634 5363 16668 5379
rect 16634 5345 16668 5363
rect 16634 5295 16668 5307
rect 16634 5273 16668 5295
rect 16634 5227 16668 5235
rect 16634 5201 16668 5227
rect 16720 6145 16754 6171
rect 16720 6137 16754 6145
rect 16720 6077 16754 6099
rect 16720 6065 16754 6077
rect 16720 6009 16754 6027
rect 16720 5993 16754 6009
rect 16720 5941 16754 5955
rect 16720 5921 16754 5941
rect 16720 5873 16754 5883
rect 16720 5849 16754 5873
rect 16720 5805 16754 5811
rect 16720 5777 16754 5805
rect 16720 5737 16754 5739
rect 16720 5705 16754 5737
rect 16720 5635 16754 5667
rect 16720 5633 16754 5635
rect 16720 5567 16754 5595
rect 16720 5561 16754 5567
rect 16720 5499 16754 5523
rect 16720 5489 16754 5499
rect 16720 5431 16754 5451
rect 16720 5417 16754 5431
rect 16720 5363 16754 5379
rect 16720 5345 16754 5363
rect 16720 5295 16754 5307
rect 16720 5273 16754 5295
rect 16720 5227 16754 5235
rect 16720 5201 16754 5227
rect 16806 6145 16840 6171
rect 16806 6137 16840 6145
rect 16806 6077 16840 6099
rect 16806 6065 16840 6077
rect 16806 6009 16840 6027
rect 16806 5993 16840 6009
rect 16806 5941 16840 5955
rect 16806 5921 16840 5941
rect 16806 5873 16840 5883
rect 16806 5849 16840 5873
rect 16806 5805 16840 5811
rect 16806 5777 16840 5805
rect 16806 5737 16840 5739
rect 16806 5705 16840 5737
rect 16806 5635 16840 5667
rect 16806 5633 16840 5635
rect 16806 5567 16840 5595
rect 16806 5561 16840 5567
rect 16806 5499 16840 5523
rect 16806 5489 16840 5499
rect 16806 5431 16840 5451
rect 16806 5417 16840 5431
rect 16806 5363 16840 5379
rect 16806 5345 16840 5363
rect 16806 5295 16840 5307
rect 16806 5273 16840 5295
rect 16806 5227 16840 5235
rect 16806 5201 16840 5227
rect 16892 6145 16926 6171
rect 16892 6137 16926 6145
rect 16892 6077 16926 6099
rect 16892 6065 16926 6077
rect 16892 6009 16926 6027
rect 16892 5993 16926 6009
rect 16892 5941 16926 5955
rect 16892 5921 16926 5941
rect 16892 5873 16926 5883
rect 16892 5849 16926 5873
rect 16892 5805 16926 5811
rect 16892 5777 16926 5805
rect 16892 5737 16926 5739
rect 16892 5705 16926 5737
rect 16892 5635 16926 5667
rect 16892 5633 16926 5635
rect 16892 5567 16926 5595
rect 16892 5561 16926 5567
rect 16892 5499 16926 5523
rect 16892 5489 16926 5499
rect 16892 5431 16926 5451
rect 16892 5417 16926 5431
rect 16892 5363 16926 5379
rect 16892 5345 16926 5363
rect 16892 5295 16926 5307
rect 16892 5273 16926 5295
rect 16892 5227 16926 5235
rect 16892 5201 16926 5227
rect 16978 6145 17012 6171
rect 16978 6137 17012 6145
rect 16978 6077 17012 6099
rect 16978 6065 17012 6077
rect 16978 6009 17012 6027
rect 16978 5993 17012 6009
rect 16978 5941 17012 5955
rect 16978 5921 17012 5941
rect 16978 5873 17012 5883
rect 16978 5849 17012 5873
rect 16978 5805 17012 5811
rect 16978 5777 17012 5805
rect 16978 5737 17012 5739
rect 16978 5705 17012 5737
rect 16978 5635 17012 5667
rect 16978 5633 17012 5635
rect 16978 5567 17012 5595
rect 16978 5561 17012 5567
rect 16978 5499 17012 5523
rect 16978 5489 17012 5499
rect 16978 5431 17012 5451
rect 16978 5417 17012 5431
rect 16978 5363 17012 5379
rect 16978 5345 17012 5363
rect 16978 5295 17012 5307
rect 16978 5273 17012 5295
rect 16978 5227 17012 5235
rect 16978 5201 17012 5227
rect 17064 6145 17098 6171
rect 17064 6137 17098 6145
rect 17064 6077 17098 6099
rect 17064 6065 17098 6077
rect 17064 6009 17098 6027
rect 17064 5993 17098 6009
rect 17064 5941 17098 5955
rect 17064 5921 17098 5941
rect 17064 5873 17098 5883
rect 17064 5849 17098 5873
rect 17064 5805 17098 5811
rect 17064 5777 17098 5805
rect 17064 5737 17098 5739
rect 17064 5705 17098 5737
rect 17064 5635 17098 5667
rect 17064 5633 17098 5635
rect 17064 5567 17098 5595
rect 17064 5561 17098 5567
rect 17064 5499 17098 5523
rect 17064 5489 17098 5499
rect 17064 5431 17098 5451
rect 17064 5417 17098 5431
rect 17064 5363 17098 5379
rect 17064 5345 17098 5363
rect 17064 5295 17098 5307
rect 17064 5273 17098 5295
rect 17064 5227 17098 5235
rect 17064 5201 17098 5227
rect 17150 6145 17184 6171
rect 17500 6180 17540 6200
rect 17150 6137 17184 6145
rect 17150 6077 17184 6099
rect 17150 6065 17184 6077
rect 17150 6009 17184 6027
rect 17150 5993 17184 6009
rect 17150 5941 17184 5955
rect 17150 5921 17184 5941
rect 17150 5873 17184 5883
rect 17150 5849 17184 5873
rect 17150 5805 17184 5811
rect 17150 5777 17184 5805
rect 17150 5737 17184 5739
rect 17150 5705 17184 5737
rect 17150 5635 17184 5667
rect 17150 5633 17184 5635
rect 17150 5567 17184 5595
rect 17150 5561 17184 5567
rect 17150 5499 17184 5523
rect 17150 5489 17184 5499
rect 17150 5431 17184 5451
rect 17150 5417 17184 5431
rect 17150 5363 17184 5379
rect 17150 5345 17184 5363
rect 17150 5295 17184 5307
rect 17150 5273 17184 5295
rect 17150 5227 17184 5235
rect 17150 5201 17184 5227
rect 17280 6120 17314 6154
rect 17280 6050 17314 6074
rect 17280 6040 17314 6050
rect 17280 5980 17314 5994
rect 17280 5960 17314 5980
rect 17280 5910 17314 5914
rect 17280 5880 17314 5910
rect 17280 5804 17314 5834
rect 17280 5800 17314 5804
rect 17280 5734 17314 5754
rect 17280 5720 17314 5734
rect 17280 5664 17314 5674
rect 17280 5640 17314 5664
rect 17280 5560 17314 5594
rect 17280 5490 17314 5514
rect 17280 5480 17314 5490
rect 17280 5420 17314 5434
rect 17280 5400 17314 5420
rect 17280 5350 17314 5354
rect 17280 5320 17314 5350
rect 17280 5244 17314 5274
rect 17280 5240 17314 5244
rect 17500 6140 17520 6180
rect 17520 6140 17540 6180
rect 17500 6100 17540 6140
rect 17500 6060 17520 6100
rect 17520 6060 17540 6100
rect 17500 6020 17540 6060
rect 17500 5980 17520 6020
rect 17520 5980 17540 6020
rect 17500 5940 17540 5980
rect 17500 5900 17520 5940
rect 17520 5900 17540 5940
rect 17500 5860 17540 5900
rect 17500 5820 17520 5860
rect 17520 5820 17540 5860
rect 17500 5780 17540 5820
rect 17500 5740 17520 5780
rect 17520 5740 17540 5780
rect 17500 5700 17540 5740
rect 17500 5660 17520 5700
rect 17520 5660 17540 5700
rect 17500 5620 17540 5660
rect 17500 5580 17520 5620
rect 17520 5580 17540 5620
rect 17500 5540 17540 5580
rect 17500 5500 17520 5540
rect 17520 5500 17540 5540
rect 17500 5460 17540 5500
rect 17500 5420 17520 5460
rect 17520 5420 17540 5460
rect 17500 5380 17540 5420
rect 17500 5340 17520 5380
rect 17520 5340 17540 5380
rect 17500 5300 17540 5340
rect 17500 5260 17520 5300
rect 17520 5260 17540 5300
rect 17604 6146 17638 6180
rect 17604 6074 17638 6108
rect 17604 6002 17638 6036
rect 17604 5930 17638 5964
rect 17604 5858 17638 5892
rect 17604 5786 17638 5820
rect 17604 5714 17638 5748
rect 17604 5642 17638 5676
rect 17604 5570 17638 5604
rect 17604 5498 17638 5532
rect 17604 5426 17638 5460
rect 17604 5354 17638 5388
rect 17604 5282 17638 5316
rect 17690 6146 17724 6180
rect 17690 6074 17724 6108
rect 17690 6002 17724 6036
rect 17690 5930 17724 5964
rect 17690 5858 17724 5892
rect 17690 5786 17724 5820
rect 17690 5714 17724 5748
rect 17690 5642 17724 5676
rect 17690 5570 17724 5604
rect 17690 5498 17724 5532
rect 17690 5426 17724 5460
rect 17690 5354 17724 5388
rect 17690 5282 17724 5316
rect 17776 6146 17810 6180
rect 17776 6074 17810 6108
rect 17776 6002 17810 6036
rect 17776 5930 17810 5964
rect 17776 5858 17810 5892
rect 17776 5786 17810 5820
rect 17776 5714 17810 5748
rect 17776 5642 17810 5676
rect 17776 5570 17810 5604
rect 17776 5498 17810 5532
rect 17776 5426 17810 5460
rect 17776 5354 17810 5388
rect 17776 5282 17810 5316
rect 17862 6146 17896 6180
rect 17862 6074 17896 6108
rect 17862 6002 17896 6036
rect 17862 5930 17896 5964
rect 17862 5858 17896 5892
rect 17862 5786 17896 5820
rect 17862 5714 17896 5748
rect 17862 5642 17896 5676
rect 17862 5570 17896 5604
rect 17862 5498 17896 5532
rect 17862 5426 17896 5460
rect 17862 5354 17896 5388
rect 17862 5282 17896 5316
rect 17948 6146 17982 6180
rect 17948 6074 17982 6108
rect 17948 6002 17982 6036
rect 17948 5930 17982 5964
rect 17948 5858 17982 5892
rect 17948 5786 17982 5820
rect 17948 5714 17982 5748
rect 17948 5642 17982 5676
rect 17948 5570 17982 5604
rect 17948 5498 17982 5532
rect 17948 5426 17982 5460
rect 17948 5354 17982 5388
rect 17948 5282 17982 5316
rect 18034 6146 18068 6180
rect 18034 6074 18068 6108
rect 18034 6002 18068 6036
rect 18034 5930 18068 5964
rect 18034 5858 18068 5892
rect 18034 5786 18068 5820
rect 18034 5714 18068 5748
rect 18034 5642 18068 5676
rect 18034 5570 18068 5604
rect 18034 5498 18068 5532
rect 18034 5426 18068 5460
rect 18034 5354 18068 5388
rect 18034 5282 18068 5316
rect 18120 6146 18154 6180
rect 18120 6074 18154 6108
rect 18120 6002 18154 6036
rect 18120 5930 18154 5964
rect 18120 5858 18154 5892
rect 18120 5786 18154 5820
rect 18120 5714 18154 5748
rect 18120 5642 18154 5676
rect 18120 5570 18154 5604
rect 18120 5498 18154 5532
rect 18120 5426 18154 5460
rect 18120 5354 18154 5388
rect 18120 5282 18154 5316
rect 18206 6146 18240 6180
rect 18206 6074 18240 6108
rect 18206 6002 18240 6036
rect 18206 5930 18240 5964
rect 18206 5858 18240 5892
rect 18206 5786 18240 5820
rect 18206 5714 18240 5748
rect 18206 5642 18240 5676
rect 18206 5570 18240 5604
rect 18206 5498 18240 5532
rect 18206 5426 18240 5460
rect 18206 5354 18240 5388
rect 18206 5282 18240 5316
rect 18292 6146 18326 6180
rect 18292 6074 18326 6108
rect 18292 6002 18326 6036
rect 18292 5930 18326 5964
rect 18292 5858 18326 5892
rect 18292 5786 18326 5820
rect 18292 5714 18326 5748
rect 18292 5642 18326 5676
rect 18292 5570 18326 5604
rect 18292 5498 18326 5532
rect 18292 5426 18326 5460
rect 18292 5354 18326 5388
rect 18292 5282 18326 5316
rect 18378 6146 18412 6180
rect 18378 6074 18412 6108
rect 18378 6002 18412 6036
rect 18378 5930 18412 5964
rect 18378 5858 18412 5892
rect 18378 5786 18412 5820
rect 18378 5714 18412 5748
rect 18378 5642 18412 5676
rect 18378 5570 18412 5604
rect 18378 5498 18412 5532
rect 18378 5426 18412 5460
rect 18378 5354 18412 5388
rect 18378 5282 18412 5316
rect 18464 6146 18498 6180
rect 18464 6074 18498 6108
rect 18464 6002 18498 6036
rect 18464 5930 18498 5964
rect 18464 5858 18498 5892
rect 18464 5786 18498 5820
rect 18464 5714 18498 5748
rect 18464 5642 18498 5676
rect 18464 5570 18498 5604
rect 18464 5498 18498 5532
rect 18464 5426 18498 5460
rect 18464 5354 18498 5388
rect 18464 5282 18498 5316
rect 18550 6146 18584 6180
rect 18550 6074 18584 6108
rect 18550 6002 18584 6036
rect 18550 5930 18584 5964
rect 18550 5858 18584 5892
rect 18550 5786 18584 5820
rect 18550 5714 18584 5748
rect 18550 5642 18584 5676
rect 18550 5570 18584 5604
rect 18550 5498 18584 5532
rect 18550 5426 18584 5460
rect 18550 5354 18584 5388
rect 18550 5282 18584 5316
rect 18636 6146 18670 6180
rect 18636 6074 18670 6108
rect 18636 6002 18670 6036
rect 18636 5930 18670 5964
rect 18636 5858 18670 5892
rect 18636 5786 18670 5820
rect 18636 5714 18670 5748
rect 18636 5642 18670 5676
rect 18636 5570 18670 5604
rect 18636 5498 18670 5532
rect 18636 5426 18670 5460
rect 18636 5354 18670 5388
rect 18636 5282 18670 5316
rect 18722 6146 18756 6180
rect 18722 6074 18756 6108
rect 18722 6002 18756 6036
rect 18722 5930 18756 5964
rect 18722 5858 18756 5892
rect 18722 5786 18756 5820
rect 18722 5714 18756 5748
rect 18722 5642 18756 5676
rect 18722 5570 18756 5604
rect 18722 5498 18756 5532
rect 18722 5426 18756 5460
rect 18722 5354 18756 5388
rect 18722 5282 18756 5316
rect 18808 6146 18842 6180
rect 18808 6074 18842 6108
rect 18808 6002 18842 6036
rect 18808 5930 18842 5964
rect 18808 5858 18842 5892
rect 18808 5786 18842 5820
rect 18808 5714 18842 5748
rect 18808 5642 18842 5676
rect 18808 5570 18842 5604
rect 18808 5498 18842 5532
rect 18808 5426 18842 5460
rect 18808 5354 18842 5388
rect 18808 5282 18842 5316
rect 18894 6146 18928 6180
rect 18894 6074 18928 6108
rect 18894 6002 18928 6036
rect 18894 5930 18928 5964
rect 18894 5858 18928 5892
rect 18894 5786 18928 5820
rect 18894 5714 18928 5748
rect 18894 5642 18928 5676
rect 18894 5570 18928 5604
rect 18894 5498 18928 5532
rect 18894 5426 18928 5460
rect 18894 5354 18928 5388
rect 18894 5282 18928 5316
rect 18980 6146 19014 6180
rect 18980 6074 19014 6108
rect 18980 6002 19014 6036
rect 18980 5930 19014 5964
rect 18980 5858 19014 5892
rect 18980 5786 19014 5820
rect 18980 5714 19014 5748
rect 18980 5642 19014 5676
rect 18980 5570 19014 5604
rect 18980 5498 19014 5532
rect 18980 5426 19014 5460
rect 18980 5354 19014 5388
rect 18980 5282 19014 5316
rect 19066 6146 19100 6180
rect 19066 6074 19100 6108
rect 19066 6002 19100 6036
rect 19066 5930 19100 5964
rect 19066 5858 19100 5892
rect 19066 5786 19100 5820
rect 19066 5714 19100 5748
rect 19066 5642 19100 5676
rect 19066 5570 19100 5604
rect 19066 5498 19100 5532
rect 19066 5426 19100 5460
rect 19066 5354 19100 5388
rect 19066 5282 19100 5316
rect 19152 6146 19186 6180
rect 19152 6074 19186 6108
rect 19152 6002 19186 6036
rect 19152 5930 19186 5964
rect 19152 5858 19186 5892
rect 19152 5786 19186 5820
rect 19152 5714 19186 5748
rect 19152 5642 19186 5676
rect 19152 5570 19186 5604
rect 19152 5498 19186 5532
rect 19152 5426 19186 5460
rect 19152 5354 19186 5388
rect 19152 5282 19186 5316
rect 19238 6146 19272 6180
rect 19238 6074 19272 6108
rect 19238 6002 19272 6036
rect 19238 5930 19272 5964
rect 19238 5858 19272 5892
rect 19238 5786 19272 5820
rect 19238 5714 19272 5748
rect 19238 5642 19272 5676
rect 19238 5570 19272 5604
rect 19238 5498 19272 5532
rect 19238 5426 19272 5460
rect 19238 5354 19272 5388
rect 19238 5282 19272 5316
rect 19324 6146 19358 6180
rect 19324 6074 19358 6108
rect 19324 6002 19358 6036
rect 19324 5930 19358 5964
rect 19324 5858 19358 5892
rect 19324 5786 19358 5820
rect 19324 5714 19358 5748
rect 19324 5642 19358 5676
rect 19324 5570 19358 5604
rect 19324 5498 19358 5532
rect 19324 5426 19358 5460
rect 19324 5354 19358 5388
rect 19324 5282 19358 5316
rect 19410 6146 19444 6180
rect 19410 6074 19444 6108
rect 19410 6002 19444 6036
rect 19410 5930 19444 5964
rect 19410 5858 19444 5892
rect 19410 5786 19444 5820
rect 19410 5714 19444 5748
rect 19410 5642 19444 5676
rect 19410 5570 19444 5604
rect 19410 5498 19444 5532
rect 19410 5426 19444 5460
rect 19410 5354 19444 5388
rect 19410 5282 19444 5316
rect 19496 6146 19530 6180
rect 19496 6074 19530 6108
rect 19496 6002 19530 6036
rect 19496 5930 19530 5964
rect 19496 5858 19530 5892
rect 19496 5786 19530 5820
rect 19496 5714 19530 5748
rect 19496 5642 19530 5676
rect 19496 5570 19530 5604
rect 19496 5498 19530 5532
rect 19496 5426 19530 5460
rect 19496 5354 19530 5388
rect 19496 5282 19530 5316
rect 19582 6146 19616 6180
rect 19582 6074 19616 6108
rect 19582 6002 19616 6036
rect 19582 5930 19616 5964
rect 19582 5858 19616 5892
rect 19582 5786 19616 5820
rect 19582 5714 19616 5748
rect 19582 5642 19616 5676
rect 19582 5570 19616 5604
rect 19582 5498 19616 5532
rect 19582 5426 19616 5460
rect 19582 5354 19616 5388
rect 19582 5282 19616 5316
rect 19668 6146 19702 6180
rect 19668 6074 19702 6108
rect 19668 6002 19702 6036
rect 19668 5930 19702 5964
rect 19668 5858 19702 5892
rect 19668 5786 19702 5820
rect 19668 5714 19702 5748
rect 19668 5642 19702 5676
rect 19668 5570 19702 5604
rect 19668 5498 19702 5532
rect 19668 5426 19702 5460
rect 19668 5354 19702 5388
rect 19668 5282 19702 5316
rect 19754 6146 19788 6180
rect 19754 6074 19788 6108
rect 19754 6002 19788 6036
rect 19754 5930 19788 5964
rect 19754 5858 19788 5892
rect 19754 5786 19788 5820
rect 19754 5714 19788 5748
rect 19754 5642 19788 5676
rect 19754 5570 19788 5604
rect 19754 5498 19788 5532
rect 19754 5426 19788 5460
rect 19754 5354 19788 5388
rect 19754 5282 19788 5316
rect 19840 6146 19874 6180
rect 19840 6074 19874 6108
rect 19840 6002 19874 6036
rect 19840 5930 19874 5964
rect 19840 5858 19874 5892
rect 19840 5786 19874 5820
rect 19840 5714 19874 5748
rect 19840 5642 19874 5676
rect 19840 5570 19874 5604
rect 19840 5498 19874 5532
rect 19840 5426 19874 5460
rect 19840 5354 19874 5388
rect 19840 5282 19874 5316
rect 19926 6146 19960 6180
rect 19926 6074 19960 6108
rect 19926 6002 19960 6036
rect 19926 5930 19960 5964
rect 19926 5858 19960 5892
rect 19926 5786 19960 5820
rect 19926 5714 19960 5748
rect 19926 5642 19960 5676
rect 19926 5570 19960 5604
rect 19926 5498 19960 5532
rect 19926 5426 19960 5460
rect 19926 5354 19960 5388
rect 19926 5282 19960 5316
rect 20012 6146 20046 6180
rect 20012 6074 20046 6108
rect 20012 6002 20046 6036
rect 20012 5930 20046 5964
rect 20012 5858 20046 5892
rect 20012 5786 20046 5820
rect 20012 5714 20046 5748
rect 20012 5642 20046 5676
rect 20012 5570 20046 5604
rect 20012 5498 20046 5532
rect 20012 5426 20046 5460
rect 20012 5354 20046 5388
rect 20012 5282 20046 5316
rect 20120 6180 20160 6200
rect 20120 6140 20140 6180
rect 20140 6140 20160 6180
rect 20120 6100 20160 6140
rect 20120 6060 20140 6100
rect 20140 6060 20160 6100
rect 20120 6020 20160 6060
rect 20120 5980 20140 6020
rect 20140 5980 20160 6020
rect 20120 5940 20160 5980
rect 20120 5900 20140 5940
rect 20140 5900 20160 5940
rect 20120 5860 20160 5900
rect 20120 5820 20140 5860
rect 20140 5820 20160 5860
rect 20120 5780 20160 5820
rect 20120 5740 20140 5780
rect 20140 5740 20160 5780
rect 20120 5700 20160 5740
rect 20120 5660 20140 5700
rect 20140 5660 20160 5700
rect 20120 5620 20160 5660
rect 20120 5580 20140 5620
rect 20140 5580 20160 5620
rect 20120 5540 20160 5580
rect 20120 5500 20140 5540
rect 20140 5500 20160 5540
rect 20120 5460 20160 5500
rect 20120 5420 20140 5460
rect 20140 5420 20160 5460
rect 20120 5380 20160 5420
rect 20120 5340 20140 5380
rect 20140 5340 20160 5380
rect 20120 5300 20160 5340
rect 20120 5260 20140 5300
rect 20140 5260 20160 5300
rect 17280 5174 17314 5194
rect 17280 5160 17314 5174
rect 16080 5050 16104 5084
rect 16104 5050 16114 5084
rect 16160 5050 16174 5084
rect 16174 5050 16194 5084
rect 16240 5050 16244 5084
rect 16244 5050 16274 5084
rect 16320 5050 16350 5084
rect 16350 5050 16354 5084
rect 16400 5050 16420 5084
rect 16420 5050 16434 5084
rect 16480 5050 16490 5084
rect 16490 5050 16514 5084
rect 16560 5050 16594 5084
rect 16640 5050 16664 5084
rect 16664 5050 16674 5084
rect 16720 5050 16734 5084
rect 16734 5050 16754 5084
rect 16800 5050 16804 5084
rect 16804 5050 16834 5084
rect 16880 5050 16910 5084
rect 16910 5050 16914 5084
rect 16960 5050 16980 5084
rect 16980 5050 16994 5084
rect 17040 5050 17050 5084
rect 17050 5050 17074 5084
rect 17120 5050 17154 5084
rect 17620 5100 17660 5140
rect 17660 5100 17700 5140
rect 17700 5100 17740 5140
rect 17740 5100 17780 5140
rect 17780 5100 17820 5140
rect 17820 5100 17860 5140
rect 17860 5100 17900 5140
rect 17900 5100 17940 5140
rect 17940 5100 17980 5140
rect 17980 5100 18020 5140
rect 18020 5100 18060 5140
rect 18060 5100 18100 5140
rect 18100 5100 18140 5140
rect 18140 5100 18180 5140
rect 18180 5100 18220 5140
rect 18220 5100 18260 5140
rect 18260 5100 18300 5140
rect 18300 5100 18340 5140
rect 18340 5100 18380 5140
rect 18380 5100 18420 5140
rect 18420 5100 18460 5140
rect 18460 5100 18500 5140
rect 18500 5100 18540 5140
rect 18540 5100 18580 5140
rect 18580 5100 18620 5140
rect 18620 5100 18660 5140
rect 18660 5100 18700 5140
rect 18700 5100 18740 5140
rect 18740 5100 18780 5140
rect 18780 5100 18820 5140
rect 18820 5100 18860 5140
rect 18860 5100 18900 5140
rect 18900 5100 18940 5140
rect 18940 5100 18980 5140
rect 18980 5100 19020 5140
rect 19020 5100 19060 5140
rect 19060 5100 19100 5140
rect 19100 5100 19140 5140
rect 19140 5100 19180 5140
rect 19180 5100 19220 5140
rect 19220 5100 19260 5140
rect 19260 5100 19300 5140
rect 19300 5100 19340 5140
rect 19340 5100 19380 5140
rect 19380 5100 19420 5140
rect 19420 5100 19460 5140
rect 19460 5100 19500 5140
rect 19500 5100 19540 5140
rect 19540 5100 19580 5140
rect 19580 5100 19620 5140
rect 19620 5100 19660 5140
rect 19660 5100 19700 5140
rect 19700 5100 19740 5140
rect 19740 5100 19780 5140
rect 19780 5100 19820 5140
rect 19820 5100 19860 5140
rect 19860 5100 19900 5140
rect 19900 5100 19940 5140
rect 19940 5100 19980 5140
rect 19980 5100 20020 5140
rect 20020 5100 20040 5140
rect 16635 4768 16669 4802
rect 16707 4768 16741 4802
rect 16779 4768 16813 4802
rect 16851 4768 16885 4802
rect 16923 4768 16957 4802
rect 16995 4768 17029 4802
rect 17067 4768 17101 4802
rect 17139 4768 17173 4802
rect 17211 4768 17245 4802
rect 17283 4768 17317 4802
rect 17355 4768 17389 4802
rect 17427 4768 17461 4802
rect 17499 4768 17533 4802
rect 17571 4768 17605 4802
rect 17643 4768 17677 4802
rect 17715 4768 17749 4802
rect 17787 4768 17821 4802
rect 17859 4768 17893 4802
rect 17931 4768 17965 4802
rect 18003 4768 18037 4802
rect 18075 4768 18109 4802
rect 18147 4768 18181 4802
rect 16566 4701 16600 4735
rect 18216 4701 18250 4735
rect 16566 4629 16600 4663
rect 18216 4629 18250 4663
rect 16566 4557 16600 4591
rect 18216 4557 18250 4591
rect 16566 4485 16600 4519
rect 18216 4485 18250 4519
rect 16566 4413 16600 4447
rect 18216 4413 18250 4447
rect 16566 4341 16600 4375
rect 18216 4341 18250 4375
rect 16566 4269 16600 4303
rect 18216 4269 18250 4303
rect 16566 4197 16600 4231
rect 18216 4197 18250 4231
rect 16566 4125 16600 4159
rect 18216 4125 18250 4159
rect 16566 4053 16600 4087
rect 18216 4053 18250 4087
rect 16566 3981 16600 4015
rect 18216 3981 18250 4015
rect 16566 3909 16600 3943
rect 18216 3909 18250 3943
rect 16566 3837 16600 3871
rect 18216 3837 18250 3871
rect 16566 3765 16600 3799
rect 18216 3765 18250 3799
rect 16566 3693 16600 3727
rect 18216 3693 18250 3727
rect 16566 3621 16600 3655
rect 18216 3621 18250 3655
rect 16566 3549 16600 3583
rect 18216 3549 18250 3583
rect 16566 3477 16600 3511
rect 18216 3477 18250 3511
rect 16566 3405 16600 3439
rect 18216 3405 18250 3439
rect 16566 3333 16600 3367
rect 18216 3333 18250 3367
rect 16635 3266 16669 3300
rect 16707 3266 16741 3300
rect 16779 3266 16813 3300
rect 16851 3266 16885 3300
rect 16923 3266 16957 3300
rect 16995 3266 17029 3300
rect 17067 3266 17101 3300
rect 17139 3266 17173 3300
rect 17211 3266 17245 3300
rect 17283 3266 17317 3300
rect 17355 3266 17389 3300
rect 17427 3266 17461 3300
rect 17499 3266 17533 3300
rect 17571 3266 17605 3300
rect 17643 3266 17677 3300
rect 17715 3266 17749 3300
rect 17787 3266 17821 3300
rect 17859 3266 17893 3300
rect 17931 3266 17965 3300
rect 18003 3266 18037 3300
rect 18075 3266 18109 3300
rect 18147 3266 18181 3300
rect 18485 4768 18519 4802
rect 18557 4768 18591 4802
rect 18629 4768 18663 4802
rect 18701 4768 18735 4802
rect 18773 4768 18807 4802
rect 18845 4768 18879 4802
rect 18917 4768 18951 4802
rect 18989 4768 19023 4802
rect 19061 4768 19095 4802
rect 19133 4768 19167 4802
rect 19205 4768 19239 4802
rect 19277 4768 19311 4802
rect 19349 4768 19383 4802
rect 19421 4768 19455 4802
rect 19493 4768 19527 4802
rect 19565 4768 19599 4802
rect 19637 4768 19671 4802
rect 19709 4768 19743 4802
rect 19781 4768 19815 4802
rect 19853 4768 19887 4802
rect 19925 4768 19959 4802
rect 19997 4768 20031 4802
rect 18416 4701 18450 4735
rect 20066 4701 20100 4735
rect 18416 4629 18450 4663
rect 20066 4629 20100 4663
rect 18416 4557 18450 4591
rect 20066 4557 20100 4591
rect 18416 4485 18450 4519
rect 20066 4485 20100 4519
rect 18416 4413 18450 4447
rect 20066 4413 20100 4447
rect 18416 4341 18450 4375
rect 20066 4341 20100 4375
rect 18416 4269 18450 4303
rect 20066 4269 20100 4303
rect 18416 4197 18450 4231
rect 20066 4197 20100 4231
rect 18416 4125 18450 4159
rect 20066 4125 20100 4159
rect 18416 4053 18450 4087
rect 20066 4053 20100 4087
rect 18416 3981 18450 4015
rect 20066 3981 20100 4015
rect 18416 3909 18450 3943
rect 20066 3909 20100 3943
rect 18416 3837 18450 3871
rect 20066 3837 20100 3871
rect 18416 3765 18450 3799
rect 20066 3765 20100 3799
rect 18416 3693 18450 3727
rect 20066 3693 20100 3727
rect 18416 3621 18450 3655
rect 20066 3621 20100 3655
rect 18416 3549 18450 3583
rect 20066 3549 20100 3583
rect 18416 3477 18450 3511
rect 20066 3477 20100 3511
rect 18416 3405 18450 3439
rect 20066 3405 20100 3439
rect 18416 3333 18450 3367
rect 20066 3333 20100 3367
rect 18485 3266 18519 3300
rect 18557 3266 18591 3300
rect 18629 3266 18663 3300
rect 18701 3266 18735 3300
rect 18773 3266 18807 3300
rect 18845 3266 18879 3300
rect 18917 3266 18951 3300
rect 18989 3266 19023 3300
rect 19061 3266 19095 3300
rect 19133 3266 19167 3300
rect 19205 3266 19239 3300
rect 19277 3266 19311 3300
rect 19349 3266 19383 3300
rect 19421 3266 19455 3300
rect 19493 3266 19527 3300
rect 19565 3266 19599 3300
rect 19637 3266 19671 3300
rect 19709 3266 19743 3300
rect 19781 3266 19815 3300
rect 19853 3266 19887 3300
rect 19925 3266 19959 3300
rect 19997 3266 20031 3300
<< metal1 >>
rect 16550 9861 18266 9868
rect 16550 9852 16638 9861
rect 16550 9818 16635 9852
rect 16550 9815 16638 9818
rect 16550 9763 16557 9815
rect 16609 9809 16638 9815
rect 16690 9809 16702 9861
rect 16754 9809 16766 9861
rect 16818 9809 16830 9861
rect 16882 9852 16894 9861
rect 16946 9852 16958 9861
rect 17010 9852 17022 9861
rect 17074 9852 17086 9861
rect 17138 9852 17150 9861
rect 17202 9852 17214 9861
rect 16885 9818 16894 9852
rect 16957 9818 16958 9852
rect 17138 9818 17139 9852
rect 17202 9818 17211 9852
rect 16882 9809 16894 9818
rect 16946 9809 16958 9818
rect 17010 9809 17022 9818
rect 17074 9809 17086 9818
rect 17138 9809 17150 9818
rect 17202 9809 17214 9818
rect 17266 9809 17278 9861
rect 17330 9852 17492 9861
rect 17330 9818 17355 9852
rect 17389 9818 17427 9852
rect 17461 9818 17492 9852
rect 17330 9809 17492 9818
rect 17544 9809 17556 9861
rect 17608 9809 17620 9861
rect 17672 9852 17684 9861
rect 17736 9852 17748 9861
rect 17800 9852 17812 9861
rect 17864 9852 17876 9861
rect 17928 9852 17940 9861
rect 17992 9852 18004 9861
rect 17677 9818 17684 9852
rect 17928 9818 17931 9852
rect 17992 9818 18003 9852
rect 17672 9809 17684 9818
rect 17736 9809 17748 9818
rect 17800 9809 17812 9818
rect 17864 9809 17876 9818
rect 17928 9809 17940 9818
rect 17992 9809 18004 9818
rect 18056 9809 18068 9861
rect 18120 9809 18132 9861
rect 18184 9860 18266 9861
rect 18400 9861 20116 9868
rect 18400 9860 18488 9861
rect 18184 9852 18488 9860
rect 18184 9818 18485 9852
rect 18184 9815 18488 9818
rect 18184 9809 18207 9815
rect 16609 9802 18207 9809
rect 16609 9763 16616 9802
rect 16550 9751 16566 9763
rect 16600 9751 16616 9763
rect 16550 9699 16557 9751
rect 16609 9699 16616 9751
rect 16550 9687 16566 9699
rect 16600 9687 16616 9699
rect 16550 9635 16557 9687
rect 16609 9635 16616 9687
rect 16550 9623 16566 9635
rect 16600 9623 16616 9635
rect 16550 9571 16557 9623
rect 16609 9571 16616 9623
rect 16550 9569 16616 9571
rect 16550 9559 16566 9569
rect 16600 9559 16616 9569
rect 16550 9507 16557 9559
rect 16609 9507 16616 9559
rect 16550 9497 16616 9507
rect 16550 9495 16566 9497
rect 16600 9495 16616 9497
rect 16550 9443 16557 9495
rect 16609 9443 16616 9495
rect 16550 9431 16616 9443
rect 16550 9379 16557 9431
rect 16609 9379 16616 9431
rect 16550 9367 16616 9379
rect 16550 9315 16557 9367
rect 16609 9315 16616 9367
rect 16550 9303 16616 9315
rect 16550 9251 16557 9303
rect 16609 9251 16616 9303
rect 16550 9247 16566 9251
rect 16600 9247 16616 9251
rect 16550 9239 16616 9247
rect 16550 9187 16557 9239
rect 16609 9187 16616 9239
rect 16550 9175 16566 9187
rect 16600 9175 16616 9187
rect 16550 9137 16616 9175
rect 16550 9103 16566 9137
rect 16600 9103 16616 9137
rect 16550 9065 16616 9103
rect 16550 9031 16566 9065
rect 16600 9031 16616 9065
rect 16550 8993 16616 9031
rect 16550 8981 16566 8993
rect 16600 8981 16616 8993
rect 16550 8929 16557 8981
rect 16609 8929 16616 8981
rect 16550 8921 16616 8929
rect 16550 8917 16566 8921
rect 16600 8917 16616 8921
rect 16550 8865 16557 8917
rect 16609 8865 16616 8917
rect 16550 8853 16616 8865
rect 16550 8801 16557 8853
rect 16609 8801 16616 8853
rect 16550 8789 16616 8801
rect 16550 8737 16557 8789
rect 16609 8737 16616 8789
rect 16550 8725 16616 8737
rect 16550 8673 16557 8725
rect 16609 8673 16616 8725
rect 16550 8671 16566 8673
rect 16600 8671 16616 8673
rect 16550 8661 16616 8671
rect 16550 8609 16557 8661
rect 16609 8609 16616 8661
rect 16550 8599 16566 8609
rect 16600 8599 16616 8609
rect 16550 8597 16616 8599
rect 16550 8545 16557 8597
rect 16609 8545 16616 8597
rect 16550 8533 16566 8545
rect 16600 8533 16616 8545
rect 16550 8481 16557 8533
rect 16609 8481 16616 8533
rect 16550 8469 16566 8481
rect 16600 8469 16616 8481
rect 16550 8417 16557 8469
rect 16609 8417 16616 8469
rect 16550 8405 16566 8417
rect 16600 8405 16616 8417
rect 16550 8359 16557 8405
rect 16480 8353 16557 8359
rect 16609 8366 16616 8405
rect 16649 9116 16677 9774
rect 16705 9144 16733 9802
rect 16761 9116 16789 9774
rect 16817 9144 16845 9802
rect 16873 9116 16901 9774
rect 16929 9144 16957 9802
rect 16985 9116 17013 9774
rect 17041 9144 17069 9802
rect 17097 9116 17125 9774
rect 17153 9144 17181 9802
rect 17209 9116 17237 9774
rect 17265 9144 17293 9802
rect 17321 9116 17349 9774
rect 17381 9768 17435 9774
rect 17381 9716 17382 9768
rect 17434 9716 17435 9768
rect 17381 9704 17435 9716
rect 17381 9652 17382 9704
rect 17434 9652 17435 9704
rect 17381 9640 17435 9652
rect 17381 9588 17382 9640
rect 17434 9588 17435 9640
rect 17381 9576 17435 9588
rect 17381 9524 17382 9576
rect 17434 9524 17435 9576
rect 17381 9512 17435 9524
rect 17381 9460 17382 9512
rect 17434 9460 17435 9512
rect 17381 9448 17435 9460
rect 17381 9396 17382 9448
rect 17434 9396 17435 9448
rect 17381 9384 17435 9396
rect 17381 9332 17382 9384
rect 17434 9332 17435 9384
rect 17381 9320 17435 9332
rect 17381 9268 17382 9320
rect 17434 9268 17435 9320
rect 17381 9256 17435 9268
rect 17381 9204 17382 9256
rect 17434 9204 17435 9256
rect 17381 9192 17435 9204
rect 17381 9140 17382 9192
rect 17434 9140 17435 9192
rect 17381 9116 17435 9140
rect 17467 9116 17495 9774
rect 17523 9144 17551 9802
rect 17579 9116 17607 9774
rect 17635 9144 17663 9802
rect 17691 9116 17719 9774
rect 17747 9144 17775 9802
rect 17803 9116 17831 9774
rect 17859 9144 17887 9802
rect 17915 9116 17943 9774
rect 17971 9144 17999 9802
rect 18027 9116 18055 9774
rect 18083 9144 18111 9802
rect 18139 9116 18167 9774
rect 16649 9110 18167 9116
rect 16649 9058 16655 9110
rect 16707 9058 16719 9110
rect 16771 9058 16783 9110
rect 16835 9058 16847 9110
rect 16899 9058 16911 9110
rect 16963 9058 16975 9110
rect 17027 9058 17039 9110
rect 17091 9058 17103 9110
rect 17155 9058 17167 9110
rect 17219 9058 17231 9110
rect 17283 9058 17295 9110
rect 17347 9058 17469 9110
rect 17521 9058 17533 9110
rect 17585 9058 17597 9110
rect 17649 9058 17661 9110
rect 17713 9058 17725 9110
rect 17777 9058 17789 9110
rect 17841 9058 17853 9110
rect 17905 9058 17917 9110
rect 17969 9058 17981 9110
rect 18033 9058 18045 9110
rect 18097 9058 18109 9110
rect 18161 9058 18167 9110
rect 16649 9052 18167 9058
rect 16649 8394 16677 9052
rect 16705 8366 16733 9024
rect 16761 8394 16789 9052
rect 16817 8366 16845 9024
rect 16873 8394 16901 9052
rect 16929 8366 16957 9024
rect 16985 8394 17013 9052
rect 17041 8366 17069 9024
rect 17097 8394 17125 9052
rect 17153 8366 17181 9024
rect 17209 8394 17237 9052
rect 17265 8366 17293 9024
rect 17321 8394 17349 9052
rect 17381 9028 17435 9052
rect 17381 8976 17382 9028
rect 17434 8976 17435 9028
rect 17381 8964 17435 8976
rect 17381 8912 17382 8964
rect 17434 8912 17435 8964
rect 17381 8900 17435 8912
rect 17381 8848 17382 8900
rect 17434 8848 17435 8900
rect 17381 8836 17435 8848
rect 17381 8784 17382 8836
rect 17434 8784 17435 8836
rect 17381 8772 17435 8784
rect 17381 8720 17382 8772
rect 17434 8720 17435 8772
rect 17381 8708 17435 8720
rect 17381 8656 17382 8708
rect 17434 8656 17435 8708
rect 17381 8644 17435 8656
rect 17381 8592 17382 8644
rect 17434 8592 17435 8644
rect 17381 8580 17435 8592
rect 17381 8528 17382 8580
rect 17434 8528 17435 8580
rect 17381 8516 17435 8528
rect 17381 8464 17382 8516
rect 17434 8464 17435 8516
rect 17381 8452 17435 8464
rect 17381 8400 17382 8452
rect 17434 8400 17435 8452
rect 17381 8394 17435 8400
rect 17467 8394 17495 9052
rect 17523 8366 17551 9024
rect 17579 8394 17607 9052
rect 17635 8366 17663 9024
rect 17691 8394 17719 9052
rect 17747 8366 17775 9024
rect 17803 8394 17831 9052
rect 17859 8366 17887 9024
rect 17915 8394 17943 9052
rect 17971 8366 17999 9024
rect 18027 8394 18055 9052
rect 18083 8366 18111 9024
rect 18139 8394 18167 9052
rect 18200 9763 18207 9802
rect 18259 9763 18407 9815
rect 18459 9809 18488 9815
rect 18540 9809 18552 9861
rect 18604 9809 18616 9861
rect 18668 9809 18680 9861
rect 18732 9852 18744 9861
rect 18796 9852 18808 9861
rect 18860 9852 18872 9861
rect 18924 9852 18936 9861
rect 18988 9852 19000 9861
rect 19052 9852 19064 9861
rect 18735 9818 18744 9852
rect 18807 9818 18808 9852
rect 18988 9818 18989 9852
rect 19052 9818 19061 9852
rect 18732 9809 18744 9818
rect 18796 9809 18808 9818
rect 18860 9809 18872 9818
rect 18924 9809 18936 9818
rect 18988 9809 19000 9818
rect 19052 9809 19064 9818
rect 19116 9809 19128 9861
rect 19180 9852 19342 9861
rect 19180 9818 19205 9852
rect 19239 9818 19277 9852
rect 19311 9818 19342 9852
rect 19180 9809 19342 9818
rect 19394 9809 19406 9861
rect 19458 9809 19470 9861
rect 19522 9852 19534 9861
rect 19586 9852 19598 9861
rect 19650 9852 19662 9861
rect 19714 9852 19726 9861
rect 19778 9852 19790 9861
rect 19842 9852 19854 9861
rect 19527 9818 19534 9852
rect 19778 9818 19781 9852
rect 19842 9818 19853 9852
rect 19522 9809 19534 9818
rect 19586 9809 19598 9818
rect 19650 9809 19662 9818
rect 19714 9809 19726 9818
rect 19778 9809 19790 9818
rect 19842 9809 19854 9818
rect 19906 9809 19918 9861
rect 19970 9809 19982 9861
rect 20034 9815 20116 9861
rect 20034 9809 20057 9815
rect 18459 9802 20057 9809
rect 18459 9763 18466 9802
rect 18200 9751 18216 9763
rect 18250 9751 18416 9763
rect 18450 9751 18466 9763
rect 18200 9699 18207 9751
rect 18259 9699 18407 9751
rect 18459 9699 18466 9751
rect 18200 9687 18216 9699
rect 18250 9687 18416 9699
rect 18450 9687 18466 9699
rect 18200 9635 18207 9687
rect 18259 9635 18407 9687
rect 18459 9635 18466 9687
rect 18200 9623 18216 9635
rect 18250 9623 18416 9635
rect 18450 9623 18466 9635
rect 18200 9571 18207 9623
rect 18259 9571 18407 9623
rect 18459 9571 18466 9623
rect 18200 9569 18466 9571
rect 18200 9559 18216 9569
rect 18250 9559 18416 9569
rect 18450 9559 18466 9569
rect 18200 9507 18207 9559
rect 18259 9507 18407 9559
rect 18459 9507 18466 9559
rect 18200 9497 18466 9507
rect 18200 9495 18216 9497
rect 18250 9495 18416 9497
rect 18450 9495 18466 9497
rect 18200 9443 18207 9495
rect 18259 9443 18407 9495
rect 18459 9443 18466 9495
rect 18200 9431 18466 9443
rect 18200 9379 18207 9431
rect 18259 9379 18407 9431
rect 18459 9379 18466 9431
rect 18200 9367 18466 9379
rect 18200 9315 18207 9367
rect 18259 9315 18407 9367
rect 18459 9315 18466 9367
rect 18200 9303 18466 9315
rect 18200 9251 18207 9303
rect 18259 9251 18407 9303
rect 18459 9251 18466 9303
rect 18200 9247 18216 9251
rect 18250 9247 18416 9251
rect 18450 9247 18466 9251
rect 18200 9239 18466 9247
rect 18200 9187 18207 9239
rect 18259 9187 18407 9239
rect 18459 9187 18466 9239
rect 18200 9175 18216 9187
rect 18250 9175 18416 9187
rect 18450 9175 18466 9187
rect 18200 9137 18466 9175
rect 18200 9103 18216 9137
rect 18250 9103 18416 9137
rect 18450 9103 18466 9137
rect 18200 9065 18466 9103
rect 18200 9031 18216 9065
rect 18250 9031 18416 9065
rect 18450 9031 18466 9065
rect 18200 8993 18466 9031
rect 18200 8981 18216 8993
rect 18250 8981 18416 8993
rect 18450 8981 18466 8993
rect 18200 8929 18207 8981
rect 18259 8929 18407 8981
rect 18459 8929 18466 8981
rect 18200 8921 18466 8929
rect 18200 8917 18216 8921
rect 18250 8917 18416 8921
rect 18450 8917 18466 8921
rect 18200 8865 18207 8917
rect 18259 8865 18407 8917
rect 18459 8865 18466 8917
rect 18200 8853 18466 8865
rect 18200 8801 18207 8853
rect 18259 8801 18407 8853
rect 18459 8801 18466 8853
rect 18200 8789 18466 8801
rect 18200 8737 18207 8789
rect 18259 8737 18407 8789
rect 18459 8737 18466 8789
rect 18200 8725 18466 8737
rect 18200 8673 18207 8725
rect 18259 8673 18407 8725
rect 18459 8673 18466 8725
rect 18200 8671 18216 8673
rect 18250 8671 18416 8673
rect 18450 8671 18466 8673
rect 18200 8661 18466 8671
rect 18200 8609 18207 8661
rect 18259 8609 18407 8661
rect 18459 8609 18466 8661
rect 18200 8599 18216 8609
rect 18250 8599 18416 8609
rect 18450 8599 18466 8609
rect 18200 8597 18466 8599
rect 18200 8545 18207 8597
rect 18259 8545 18407 8597
rect 18459 8545 18466 8597
rect 18200 8533 18216 8545
rect 18250 8533 18416 8545
rect 18450 8533 18466 8545
rect 18200 8481 18207 8533
rect 18259 8481 18407 8533
rect 18459 8481 18466 8533
rect 18200 8469 18216 8481
rect 18250 8469 18416 8481
rect 18450 8469 18466 8481
rect 18200 8417 18207 8469
rect 18259 8417 18407 8469
rect 18459 8417 18466 8469
rect 18200 8405 18216 8417
rect 18250 8405 18416 8417
rect 18450 8405 18466 8417
rect 18200 8366 18207 8405
rect 16609 8359 18207 8366
rect 16609 8353 16638 8359
rect 16480 8350 16638 8353
rect 16480 8316 16635 8350
rect 16480 8307 16638 8316
rect 16690 8307 16702 8359
rect 16754 8307 16766 8359
rect 16818 8307 16830 8359
rect 16882 8350 16894 8359
rect 16946 8350 16958 8359
rect 17010 8350 17022 8359
rect 17074 8350 17086 8359
rect 17138 8350 17150 8359
rect 17202 8350 17214 8359
rect 16885 8316 16894 8350
rect 16957 8316 16958 8350
rect 17138 8316 17139 8350
rect 17202 8316 17211 8350
rect 16882 8307 16894 8316
rect 16946 8307 16958 8316
rect 17010 8307 17022 8316
rect 17074 8307 17086 8316
rect 17138 8307 17150 8316
rect 17202 8307 17214 8316
rect 17266 8307 17278 8359
rect 17330 8350 17492 8359
rect 17330 8316 17355 8350
rect 17389 8316 17427 8350
rect 17461 8316 17492 8350
rect 17330 8307 17492 8316
rect 17544 8307 17556 8359
rect 17608 8307 17620 8359
rect 17672 8350 17684 8359
rect 17736 8350 17748 8359
rect 17800 8350 17812 8359
rect 17864 8350 17876 8359
rect 17928 8350 17940 8359
rect 17992 8350 18004 8359
rect 17677 8316 17684 8350
rect 17928 8316 17931 8350
rect 17992 8316 18003 8350
rect 17672 8307 17684 8316
rect 17736 8307 17748 8316
rect 17800 8307 17812 8316
rect 17864 8307 17876 8316
rect 17928 8307 17940 8316
rect 17992 8307 18004 8316
rect 18056 8307 18068 8359
rect 18120 8307 18132 8359
rect 18184 8353 18207 8359
rect 18259 8353 18407 8405
rect 18459 8366 18466 8405
rect 18499 9116 18527 9774
rect 18555 9144 18583 9802
rect 18611 9116 18639 9774
rect 18667 9144 18695 9802
rect 18723 9116 18751 9774
rect 18779 9144 18807 9802
rect 18835 9116 18863 9774
rect 18891 9144 18919 9802
rect 18947 9116 18975 9774
rect 19003 9144 19031 9802
rect 19059 9116 19087 9774
rect 19115 9144 19143 9802
rect 19171 9116 19199 9774
rect 19231 9768 19285 9774
rect 19231 9716 19232 9768
rect 19284 9716 19285 9768
rect 19231 9704 19285 9716
rect 19231 9652 19232 9704
rect 19284 9652 19285 9704
rect 19231 9640 19285 9652
rect 19231 9588 19232 9640
rect 19284 9588 19285 9640
rect 19231 9576 19285 9588
rect 19231 9524 19232 9576
rect 19284 9524 19285 9576
rect 19231 9512 19285 9524
rect 19231 9460 19232 9512
rect 19284 9460 19285 9512
rect 19231 9448 19285 9460
rect 19231 9396 19232 9448
rect 19284 9396 19285 9448
rect 19231 9384 19285 9396
rect 19231 9332 19232 9384
rect 19284 9332 19285 9384
rect 19231 9320 19285 9332
rect 19231 9268 19232 9320
rect 19284 9268 19285 9320
rect 19231 9256 19285 9268
rect 19231 9204 19232 9256
rect 19284 9204 19285 9256
rect 19231 9192 19285 9204
rect 19231 9140 19232 9192
rect 19284 9140 19285 9192
rect 19231 9116 19285 9140
rect 19317 9116 19345 9774
rect 19373 9144 19401 9802
rect 19429 9116 19457 9774
rect 19485 9144 19513 9802
rect 19541 9116 19569 9774
rect 19597 9144 19625 9802
rect 19653 9116 19681 9774
rect 19709 9144 19737 9802
rect 19765 9116 19793 9774
rect 19821 9144 19849 9802
rect 19877 9116 19905 9774
rect 19933 9144 19961 9802
rect 19989 9116 20017 9774
rect 18499 9110 20017 9116
rect 18499 9058 18505 9110
rect 18557 9058 18569 9110
rect 18621 9058 18633 9110
rect 18685 9058 18697 9110
rect 18749 9058 18761 9110
rect 18813 9058 18825 9110
rect 18877 9058 18889 9110
rect 18941 9058 18953 9110
rect 19005 9058 19017 9110
rect 19069 9058 19081 9110
rect 19133 9058 19145 9110
rect 19197 9058 19319 9110
rect 19371 9058 19383 9110
rect 19435 9058 19447 9110
rect 19499 9058 19511 9110
rect 19563 9058 19575 9110
rect 19627 9058 19639 9110
rect 19691 9058 19703 9110
rect 19755 9058 19767 9110
rect 19819 9058 19831 9110
rect 19883 9058 19895 9110
rect 19947 9058 19959 9110
rect 20011 9058 20017 9110
rect 18499 9052 20017 9058
rect 18499 8394 18527 9052
rect 18555 8366 18583 9024
rect 18611 8394 18639 9052
rect 18667 8366 18695 9024
rect 18723 8394 18751 9052
rect 18779 8366 18807 9024
rect 18835 8394 18863 9052
rect 18891 8366 18919 9024
rect 18947 8394 18975 9052
rect 19003 8366 19031 9024
rect 19059 8394 19087 9052
rect 19115 8366 19143 9024
rect 19171 8394 19199 9052
rect 19231 9028 19285 9052
rect 19231 8976 19232 9028
rect 19284 8976 19285 9028
rect 19231 8964 19285 8976
rect 19231 8912 19232 8964
rect 19284 8912 19285 8964
rect 19231 8900 19285 8912
rect 19231 8848 19232 8900
rect 19284 8848 19285 8900
rect 19231 8836 19285 8848
rect 19231 8784 19232 8836
rect 19284 8784 19285 8836
rect 19231 8772 19285 8784
rect 19231 8720 19232 8772
rect 19284 8720 19285 8772
rect 19231 8708 19285 8720
rect 19231 8656 19232 8708
rect 19284 8656 19285 8708
rect 19231 8644 19285 8656
rect 19231 8592 19232 8644
rect 19284 8592 19285 8644
rect 19231 8580 19285 8592
rect 19231 8528 19232 8580
rect 19284 8528 19285 8580
rect 19231 8516 19285 8528
rect 19231 8464 19232 8516
rect 19284 8464 19285 8516
rect 19231 8452 19285 8464
rect 19231 8400 19232 8452
rect 19284 8400 19285 8452
rect 19231 8394 19285 8400
rect 19317 8394 19345 9052
rect 19373 8366 19401 9024
rect 19429 8394 19457 9052
rect 19485 8366 19513 9024
rect 19541 8394 19569 9052
rect 19597 8366 19625 9024
rect 19653 8394 19681 9052
rect 19709 8366 19737 9024
rect 19765 8394 19793 9052
rect 19821 8366 19849 9024
rect 19877 8394 19905 9052
rect 19933 8366 19961 9024
rect 19989 8394 20017 9052
rect 20050 9763 20057 9802
rect 20109 9763 20116 9815
rect 20050 9751 20066 9763
rect 20100 9751 20116 9763
rect 20050 9699 20057 9751
rect 20109 9699 20116 9751
rect 20050 9687 20066 9699
rect 20100 9687 20116 9699
rect 20050 9635 20057 9687
rect 20109 9635 20116 9687
rect 20050 9623 20066 9635
rect 20100 9623 20116 9635
rect 20050 9571 20057 9623
rect 20109 9571 20116 9623
rect 20050 9569 20116 9571
rect 20050 9559 20066 9569
rect 20100 9559 20116 9569
rect 20050 9507 20057 9559
rect 20109 9507 20116 9559
rect 20050 9497 20116 9507
rect 20050 9495 20066 9497
rect 20100 9495 20116 9497
rect 20050 9443 20057 9495
rect 20109 9443 20116 9495
rect 20050 9431 20116 9443
rect 20050 9379 20057 9431
rect 20109 9379 20116 9431
rect 20050 9367 20116 9379
rect 20050 9315 20057 9367
rect 20109 9315 20116 9367
rect 20050 9303 20116 9315
rect 20050 9251 20057 9303
rect 20109 9251 20116 9303
rect 20050 9247 20066 9251
rect 20100 9247 20116 9251
rect 20050 9239 20116 9247
rect 20050 9187 20057 9239
rect 20109 9187 20116 9239
rect 20050 9175 20066 9187
rect 20100 9175 20116 9187
rect 20050 9137 20116 9175
rect 20050 9103 20066 9137
rect 20100 9103 20116 9137
rect 20050 9065 20116 9103
rect 20050 9031 20066 9065
rect 20100 9031 20116 9065
rect 20050 8993 20116 9031
rect 20050 8981 20066 8993
rect 20100 8981 20116 8993
rect 20050 8929 20057 8981
rect 20109 8929 20116 8981
rect 20050 8921 20116 8929
rect 20050 8917 20066 8921
rect 20100 8917 20116 8921
rect 20050 8865 20057 8917
rect 20109 8865 20116 8917
rect 20050 8853 20116 8865
rect 20050 8801 20057 8853
rect 20109 8801 20116 8853
rect 20050 8789 20116 8801
rect 20050 8737 20057 8789
rect 20109 8737 20116 8789
rect 20050 8725 20116 8737
rect 20050 8673 20057 8725
rect 20109 8673 20116 8725
rect 20050 8671 20066 8673
rect 20100 8671 20116 8673
rect 20050 8661 20116 8671
rect 20050 8609 20057 8661
rect 20109 8609 20116 8661
rect 20050 8599 20066 8609
rect 20100 8599 20116 8609
rect 20050 8597 20116 8599
rect 20050 8545 20057 8597
rect 20109 8545 20116 8597
rect 20050 8533 20066 8545
rect 20100 8533 20116 8545
rect 20050 8481 20057 8533
rect 20109 8481 20116 8533
rect 20050 8469 20066 8481
rect 20100 8469 20116 8481
rect 20050 8417 20057 8469
rect 20109 8417 20116 8469
rect 20050 8405 20066 8417
rect 20100 8405 20116 8417
rect 20050 8366 20057 8405
rect 18459 8359 20057 8366
rect 18459 8353 18488 8359
rect 18184 8350 18488 8353
rect 18184 8316 18485 8350
rect 18184 8307 18488 8316
rect 18540 8307 18552 8359
rect 18604 8307 18616 8359
rect 18668 8307 18680 8359
rect 18732 8350 18744 8359
rect 18796 8350 18808 8359
rect 18860 8350 18872 8359
rect 18924 8350 18936 8359
rect 18988 8350 19000 8359
rect 19052 8350 19064 8359
rect 18735 8316 18744 8350
rect 18807 8316 18808 8350
rect 18988 8316 18989 8350
rect 19052 8316 19061 8350
rect 18732 8307 18744 8316
rect 18796 8307 18808 8316
rect 18860 8307 18872 8316
rect 18924 8307 18936 8316
rect 18988 8307 19000 8316
rect 19052 8307 19064 8316
rect 19116 8307 19128 8359
rect 19180 8350 19342 8359
rect 19180 8316 19205 8350
rect 19239 8316 19277 8350
rect 19311 8316 19342 8350
rect 19180 8307 19342 8316
rect 19394 8307 19406 8359
rect 19458 8307 19470 8359
rect 19522 8350 19534 8359
rect 19586 8350 19598 8359
rect 19650 8350 19662 8359
rect 19714 8350 19726 8359
rect 19778 8350 19790 8359
rect 19842 8350 19854 8359
rect 19527 8316 19534 8350
rect 19778 8316 19781 8350
rect 19842 8316 19853 8350
rect 19522 8307 19534 8316
rect 19586 8307 19598 8316
rect 19650 8307 19662 8316
rect 19714 8307 19726 8316
rect 19778 8307 19790 8316
rect 19842 8307 19854 8316
rect 19906 8307 19918 8359
rect 19970 8307 19982 8359
rect 20034 8353 20057 8359
rect 20109 8353 20116 8405
rect 20034 8307 20116 8353
rect 16480 8300 20116 8307
rect 16480 8220 17300 8300
rect 15980 8130 16100 8150
rect 16480 8130 16510 8220
rect 15970 8120 16510 8130
rect 17260 8130 17300 8220
rect 17380 8180 20160 8220
rect 17260 8120 17330 8130
rect 15950 8110 17330 8120
rect 15950 7000 15960 8110
rect 16060 8076 16080 8110
rect 16114 8076 16160 8110
rect 16194 8076 16240 8110
rect 16274 8076 16320 8110
rect 16354 8076 16400 8110
rect 16434 8076 16480 8110
rect 16514 8076 16560 8110
rect 16594 8076 16640 8110
rect 16674 8076 16720 8110
rect 16754 8076 16800 8110
rect 16834 8076 16880 8110
rect 16914 8076 16960 8110
rect 16994 8076 17040 8110
rect 17074 8076 17120 8110
rect 17154 8076 17330 8110
rect 16060 8061 17330 8076
rect 16060 7959 16161 8061
rect 16060 7925 16118 7959
rect 16152 7925 16161 7959
rect 16060 7887 16161 7925
rect 16060 7853 16118 7887
rect 16152 7853 16161 7887
rect 16060 7815 16161 7853
rect 16060 7781 16118 7815
rect 16152 7781 16161 7815
rect 16060 7743 16161 7781
rect 16060 7709 16118 7743
rect 16152 7709 16161 7743
rect 16060 7671 16161 7709
rect 16060 7637 16118 7671
rect 16152 7637 16161 7671
rect 16060 7599 16161 7637
rect 16060 7565 16118 7599
rect 16152 7565 16161 7599
rect 16060 7527 16161 7565
rect 16060 7493 16118 7527
rect 16152 7493 16161 7527
rect 16060 7455 16161 7493
rect 16060 7421 16118 7455
rect 16152 7421 16161 7455
rect 16060 7383 16161 7421
rect 16060 7349 16118 7383
rect 16152 7349 16161 7383
rect 16060 7311 16161 7349
rect 16060 7277 16118 7311
rect 16152 7277 16161 7311
rect 16060 7239 16161 7277
rect 16060 7205 16118 7239
rect 16152 7205 16161 7239
rect 16060 7167 16161 7205
rect 16060 7133 16118 7167
rect 16152 7133 16161 7167
rect 16060 7095 16161 7133
rect 16060 7061 16118 7095
rect 16152 7061 16161 7095
rect 16060 7023 16161 7061
rect 16060 7000 16118 7023
rect 15950 6990 16118 7000
rect 15970 6989 16118 6990
rect 16152 6989 16161 7023
rect 15970 6980 16161 6989
rect 15970 6970 16040 6980
rect 16109 6977 16161 6980
rect 16195 7959 16247 7971
rect 16195 7925 16204 7959
rect 16238 7925 16247 7959
rect 16195 7901 16247 7925
rect 16195 7821 16247 7849
rect 16195 7743 16247 7769
rect 16195 7741 16204 7743
rect 16238 7741 16247 7743
rect 16195 7671 16247 7689
rect 16195 7661 16204 7671
rect 16238 7661 16247 7671
rect 16195 7599 16247 7609
rect 16195 7581 16204 7599
rect 16238 7581 16247 7599
rect 16195 7527 16247 7529
rect 16195 7501 16204 7527
rect 16238 7501 16247 7527
rect 16195 7421 16204 7449
rect 16238 7421 16247 7449
rect 16195 7349 16204 7369
rect 16238 7349 16247 7369
rect 16195 7341 16247 7349
rect 16195 7277 16204 7289
rect 16238 7277 16247 7289
rect 16195 7261 16247 7277
rect 16195 7205 16204 7209
rect 16238 7205 16247 7209
rect 16195 7181 16247 7205
rect 16195 7101 16247 7129
rect 16195 7023 16247 7049
rect 16195 6989 16204 7023
rect 16238 6989 16247 7023
rect 16195 6977 16247 6989
rect 16281 7959 16333 8061
rect 16281 7925 16290 7959
rect 16324 7925 16333 7959
rect 16281 7887 16333 7925
rect 16281 7853 16290 7887
rect 16324 7853 16333 7887
rect 16281 7815 16333 7853
rect 16281 7781 16290 7815
rect 16324 7781 16333 7815
rect 16281 7743 16333 7781
rect 16281 7709 16290 7743
rect 16324 7709 16333 7743
rect 16281 7671 16333 7709
rect 16281 7637 16290 7671
rect 16324 7637 16333 7671
rect 16281 7599 16333 7637
rect 16281 7565 16290 7599
rect 16324 7565 16333 7599
rect 16281 7527 16333 7565
rect 16281 7493 16290 7527
rect 16324 7493 16333 7527
rect 16281 7455 16333 7493
rect 16281 7421 16290 7455
rect 16324 7421 16333 7455
rect 16281 7383 16333 7421
rect 16281 7349 16290 7383
rect 16324 7349 16333 7383
rect 16281 7311 16333 7349
rect 16281 7277 16290 7311
rect 16324 7277 16333 7311
rect 16281 7239 16333 7277
rect 16281 7205 16290 7239
rect 16324 7205 16333 7239
rect 16281 7167 16333 7205
rect 16281 7133 16290 7167
rect 16324 7133 16333 7167
rect 16281 7095 16333 7133
rect 16281 7061 16290 7095
rect 16324 7061 16333 7095
rect 16281 7023 16333 7061
rect 16281 6989 16290 7023
rect 16324 6989 16333 7023
rect 16281 6977 16333 6989
rect 16367 7959 16419 7971
rect 16367 7925 16376 7959
rect 16410 7925 16419 7959
rect 16367 7901 16419 7925
rect 16367 7821 16419 7849
rect 16367 7743 16419 7769
rect 16367 7741 16376 7743
rect 16410 7741 16419 7743
rect 16367 7671 16419 7689
rect 16367 7661 16376 7671
rect 16410 7661 16419 7671
rect 16367 7599 16419 7609
rect 16367 7581 16376 7599
rect 16410 7581 16419 7599
rect 16367 7527 16419 7529
rect 16367 7501 16376 7527
rect 16410 7501 16419 7527
rect 16367 7421 16376 7449
rect 16410 7421 16419 7449
rect 16367 7349 16376 7369
rect 16410 7349 16419 7369
rect 16367 7341 16419 7349
rect 16367 7277 16376 7289
rect 16410 7277 16419 7289
rect 16367 7261 16419 7277
rect 16367 7205 16376 7209
rect 16410 7205 16419 7209
rect 16367 7181 16419 7205
rect 16367 7101 16419 7129
rect 16367 7023 16419 7049
rect 16367 6989 16376 7023
rect 16410 6989 16419 7023
rect 16367 6977 16419 6989
rect 16453 7959 16505 8061
rect 16453 7925 16462 7959
rect 16496 7925 16505 7959
rect 16453 7887 16505 7925
rect 16453 7853 16462 7887
rect 16496 7853 16505 7887
rect 16453 7815 16505 7853
rect 16453 7781 16462 7815
rect 16496 7781 16505 7815
rect 16453 7743 16505 7781
rect 16453 7709 16462 7743
rect 16496 7709 16505 7743
rect 16453 7671 16505 7709
rect 16453 7637 16462 7671
rect 16496 7637 16505 7671
rect 16453 7599 16505 7637
rect 16453 7565 16462 7599
rect 16496 7565 16505 7599
rect 16453 7527 16505 7565
rect 16453 7493 16462 7527
rect 16496 7493 16505 7527
rect 16453 7455 16505 7493
rect 16453 7421 16462 7455
rect 16496 7421 16505 7455
rect 16453 7383 16505 7421
rect 16453 7349 16462 7383
rect 16496 7349 16505 7383
rect 16453 7311 16505 7349
rect 16453 7277 16462 7311
rect 16496 7277 16505 7311
rect 16453 7239 16505 7277
rect 16453 7205 16462 7239
rect 16496 7205 16505 7239
rect 16453 7167 16505 7205
rect 16453 7133 16462 7167
rect 16496 7133 16505 7167
rect 16453 7095 16505 7133
rect 16453 7061 16462 7095
rect 16496 7061 16505 7095
rect 16453 7023 16505 7061
rect 16453 6989 16462 7023
rect 16496 6989 16505 7023
rect 16453 6977 16505 6989
rect 16539 7959 16591 7971
rect 16539 7925 16548 7959
rect 16582 7925 16591 7959
rect 16539 7901 16591 7925
rect 16539 7821 16591 7849
rect 16539 7743 16591 7769
rect 16539 7741 16548 7743
rect 16582 7741 16591 7743
rect 16539 7671 16591 7689
rect 16539 7661 16548 7671
rect 16582 7661 16591 7671
rect 16539 7599 16591 7609
rect 16539 7581 16548 7599
rect 16582 7581 16591 7599
rect 16539 7527 16591 7529
rect 16539 7501 16548 7527
rect 16582 7501 16591 7527
rect 16539 7421 16548 7449
rect 16582 7421 16591 7449
rect 16539 7349 16548 7369
rect 16582 7349 16591 7369
rect 16539 7341 16591 7349
rect 16539 7277 16548 7289
rect 16582 7277 16591 7289
rect 16539 7261 16591 7277
rect 16539 7205 16548 7209
rect 16582 7205 16591 7209
rect 16539 7181 16591 7205
rect 16539 7101 16591 7129
rect 16539 7023 16591 7049
rect 16539 6989 16548 7023
rect 16582 6989 16591 7023
rect 16539 6977 16591 6989
rect 16625 7959 16677 8061
rect 16625 7925 16634 7959
rect 16668 7925 16677 7959
rect 16625 7887 16677 7925
rect 16625 7853 16634 7887
rect 16668 7853 16677 7887
rect 16625 7815 16677 7853
rect 16625 7781 16634 7815
rect 16668 7781 16677 7815
rect 16625 7743 16677 7781
rect 16625 7709 16634 7743
rect 16668 7709 16677 7743
rect 16625 7671 16677 7709
rect 16625 7637 16634 7671
rect 16668 7637 16677 7671
rect 16625 7599 16677 7637
rect 16625 7565 16634 7599
rect 16668 7565 16677 7599
rect 16625 7527 16677 7565
rect 16625 7493 16634 7527
rect 16668 7493 16677 7527
rect 16625 7455 16677 7493
rect 16625 7421 16634 7455
rect 16668 7421 16677 7455
rect 16625 7383 16677 7421
rect 16625 7349 16634 7383
rect 16668 7349 16677 7383
rect 16625 7311 16677 7349
rect 16625 7277 16634 7311
rect 16668 7277 16677 7311
rect 16625 7239 16677 7277
rect 16625 7205 16634 7239
rect 16668 7205 16677 7239
rect 16625 7167 16677 7205
rect 16625 7133 16634 7167
rect 16668 7133 16677 7167
rect 16625 7095 16677 7133
rect 16625 7061 16634 7095
rect 16668 7061 16677 7095
rect 16625 7023 16677 7061
rect 16625 6989 16634 7023
rect 16668 6989 16677 7023
rect 16625 6977 16677 6989
rect 16711 7959 16763 7971
rect 16711 7925 16720 7959
rect 16754 7925 16763 7959
rect 16711 7901 16763 7925
rect 16711 7821 16763 7849
rect 16711 7743 16763 7769
rect 16711 7741 16720 7743
rect 16754 7741 16763 7743
rect 16711 7671 16763 7689
rect 16711 7661 16720 7671
rect 16754 7661 16763 7671
rect 16711 7599 16763 7609
rect 16711 7581 16720 7599
rect 16754 7581 16763 7599
rect 16711 7527 16763 7529
rect 16711 7501 16720 7527
rect 16754 7501 16763 7527
rect 16711 7421 16720 7449
rect 16754 7421 16763 7449
rect 16711 7349 16720 7369
rect 16754 7349 16763 7369
rect 16711 7341 16763 7349
rect 16711 7277 16720 7289
rect 16754 7277 16763 7289
rect 16711 7261 16763 7277
rect 16711 7205 16720 7209
rect 16754 7205 16763 7209
rect 16711 7181 16763 7205
rect 16711 7101 16763 7129
rect 16711 7023 16763 7049
rect 16711 6989 16720 7023
rect 16754 6989 16763 7023
rect 16711 6977 16763 6989
rect 16797 7959 16849 8061
rect 16797 7925 16806 7959
rect 16840 7925 16849 7959
rect 16797 7887 16849 7925
rect 16797 7853 16806 7887
rect 16840 7853 16849 7887
rect 16797 7815 16849 7853
rect 16797 7781 16806 7815
rect 16840 7781 16849 7815
rect 16797 7743 16849 7781
rect 16797 7709 16806 7743
rect 16840 7709 16849 7743
rect 16797 7671 16849 7709
rect 16797 7637 16806 7671
rect 16840 7637 16849 7671
rect 16797 7599 16849 7637
rect 16797 7565 16806 7599
rect 16840 7565 16849 7599
rect 16797 7527 16849 7565
rect 16797 7493 16806 7527
rect 16840 7493 16849 7527
rect 16797 7455 16849 7493
rect 16797 7421 16806 7455
rect 16840 7421 16849 7455
rect 16797 7383 16849 7421
rect 16797 7349 16806 7383
rect 16840 7349 16849 7383
rect 16797 7311 16849 7349
rect 16797 7277 16806 7311
rect 16840 7277 16849 7311
rect 16797 7239 16849 7277
rect 16797 7205 16806 7239
rect 16840 7205 16849 7239
rect 16797 7167 16849 7205
rect 16797 7133 16806 7167
rect 16840 7133 16849 7167
rect 16797 7095 16849 7133
rect 16797 7061 16806 7095
rect 16840 7061 16849 7095
rect 16797 7023 16849 7061
rect 16797 6989 16806 7023
rect 16840 6989 16849 7023
rect 16797 6977 16849 6989
rect 16883 7959 16935 7971
rect 16883 7925 16892 7959
rect 16926 7925 16935 7959
rect 16883 7901 16935 7925
rect 16883 7821 16935 7849
rect 16883 7743 16935 7769
rect 16883 7741 16892 7743
rect 16926 7741 16935 7743
rect 16883 7671 16935 7689
rect 16883 7661 16892 7671
rect 16926 7661 16935 7671
rect 16883 7599 16935 7609
rect 16883 7581 16892 7599
rect 16926 7581 16935 7599
rect 16883 7527 16935 7529
rect 16883 7501 16892 7527
rect 16926 7501 16935 7527
rect 16883 7421 16892 7449
rect 16926 7421 16935 7449
rect 16883 7349 16892 7369
rect 16926 7349 16935 7369
rect 16883 7341 16935 7349
rect 16883 7277 16892 7289
rect 16926 7277 16935 7289
rect 16883 7261 16935 7277
rect 16883 7205 16892 7209
rect 16926 7205 16935 7209
rect 16883 7181 16935 7205
rect 16883 7101 16935 7129
rect 16883 7023 16935 7049
rect 16883 6989 16892 7023
rect 16926 6989 16935 7023
rect 16883 6977 16935 6989
rect 16969 7959 17021 8061
rect 17141 8000 17330 8061
rect 17380 8080 17420 8180
rect 20140 8080 20160 8180
rect 17380 8050 17638 8080
rect 20058 8050 20160 8080
rect 17380 8040 20160 8050
rect 16969 7925 16978 7959
rect 17012 7925 17021 7959
rect 16969 7887 17021 7925
rect 16969 7853 16978 7887
rect 17012 7853 17021 7887
rect 16969 7815 17021 7853
rect 16969 7781 16978 7815
rect 17012 7781 17021 7815
rect 16969 7743 17021 7781
rect 16969 7709 16978 7743
rect 17012 7709 17021 7743
rect 16969 7671 17021 7709
rect 16969 7637 16978 7671
rect 17012 7637 17021 7671
rect 16969 7599 17021 7637
rect 16969 7565 16978 7599
rect 17012 7565 17021 7599
rect 16969 7527 17021 7565
rect 16969 7493 16978 7527
rect 17012 7493 17021 7527
rect 16969 7455 17021 7493
rect 16969 7421 16978 7455
rect 17012 7421 17021 7455
rect 16969 7383 17021 7421
rect 16969 7349 16978 7383
rect 17012 7349 17021 7383
rect 16969 7311 17021 7349
rect 16969 7277 16978 7311
rect 17012 7277 17021 7311
rect 16969 7239 17021 7277
rect 16969 7205 16978 7239
rect 17012 7205 17021 7239
rect 16969 7167 17021 7205
rect 16969 7133 16978 7167
rect 17012 7133 17021 7167
rect 16969 7095 17021 7133
rect 16969 7061 16978 7095
rect 17012 7061 17021 7095
rect 16969 7023 17021 7061
rect 16969 6989 16978 7023
rect 17012 6989 17021 7023
rect 16969 6977 17021 6989
rect 17055 7959 17107 7971
rect 17055 7925 17064 7959
rect 17098 7925 17107 7959
rect 17055 7901 17107 7925
rect 17055 7821 17107 7849
rect 17055 7743 17107 7769
rect 17055 7741 17064 7743
rect 17098 7741 17107 7743
rect 17055 7671 17107 7689
rect 17055 7661 17064 7671
rect 17098 7661 17107 7671
rect 17055 7599 17107 7609
rect 17055 7581 17064 7599
rect 17098 7581 17107 7599
rect 17055 7527 17107 7529
rect 17055 7501 17064 7527
rect 17098 7501 17107 7527
rect 17055 7421 17064 7449
rect 17098 7421 17107 7449
rect 17055 7349 17064 7369
rect 17098 7349 17107 7369
rect 17055 7341 17107 7349
rect 17055 7277 17064 7289
rect 17098 7277 17107 7289
rect 17055 7261 17107 7277
rect 17055 7205 17064 7209
rect 17098 7205 17107 7209
rect 17055 7181 17107 7205
rect 17055 7101 17107 7129
rect 17055 7023 17107 7049
rect 17055 6989 17064 7023
rect 17098 6989 17107 7023
rect 17055 6977 17107 6989
rect 17141 7966 17280 8000
rect 17314 7966 17330 8000
rect 17141 7959 17330 7966
rect 17141 7925 17150 7959
rect 17184 7925 17330 7959
rect 17616 8038 20070 8040
rect 17616 7950 17662 8038
rect 17141 7920 17330 7925
rect 17141 7887 17280 7920
rect 17141 7853 17150 7887
rect 17184 7886 17280 7887
rect 17314 7886 17330 7920
rect 17184 7853 17330 7886
rect 17141 7840 17330 7853
rect 17141 7815 17280 7840
rect 17141 7781 17150 7815
rect 17184 7806 17280 7815
rect 17314 7806 17330 7840
rect 17184 7781 17330 7806
rect 17141 7760 17330 7781
rect 17141 7743 17280 7760
rect 17141 7709 17150 7743
rect 17184 7726 17280 7743
rect 17314 7726 17330 7760
rect 17184 7709 17330 7726
rect 17141 7680 17330 7709
rect 17141 7671 17280 7680
rect 17141 7637 17150 7671
rect 17184 7646 17280 7671
rect 17314 7646 17330 7680
rect 17184 7637 17330 7646
rect 17141 7600 17330 7637
rect 17141 7599 17280 7600
rect 17141 7565 17150 7599
rect 17184 7566 17280 7599
rect 17314 7566 17330 7600
rect 17184 7565 17330 7566
rect 17141 7527 17330 7565
rect 17141 7493 17150 7527
rect 17184 7520 17330 7527
rect 17184 7493 17280 7520
rect 17141 7486 17280 7493
rect 17314 7486 17330 7520
rect 17141 7455 17330 7486
rect 17141 7421 17150 7455
rect 17184 7440 17330 7455
rect 17184 7421 17280 7440
rect 17141 7406 17280 7421
rect 17314 7406 17330 7440
rect 17141 7383 17330 7406
rect 17141 7349 17150 7383
rect 17184 7360 17330 7383
rect 17184 7349 17280 7360
rect 17141 7326 17280 7349
rect 17314 7326 17330 7360
rect 17141 7311 17330 7326
rect 17141 7277 17150 7311
rect 17184 7280 17330 7311
rect 17184 7277 17280 7280
rect 17141 7246 17280 7277
rect 17314 7246 17330 7280
rect 17141 7239 17330 7246
rect 17141 7205 17150 7239
rect 17184 7205 17330 7239
rect 17141 7200 17330 7205
rect 17141 7167 17280 7200
rect 17141 7133 17150 7167
rect 17184 7166 17280 7167
rect 17314 7166 17330 7200
rect 17184 7133 17330 7166
rect 17141 7120 17330 7133
rect 17141 7095 17280 7120
rect 17141 7061 17150 7095
rect 17184 7086 17280 7095
rect 17314 7086 17330 7120
rect 17184 7061 17330 7086
rect 17141 7040 17330 7061
rect 17141 7023 17280 7040
rect 17141 6989 17150 7023
rect 17184 7006 17280 7023
rect 17314 7006 17330 7040
rect 17184 6989 17330 7006
rect 17141 6980 17330 6989
rect 17141 6977 17193 6980
rect 17260 6970 17330 6980
rect 17498 7930 17662 7950
rect 17498 6990 17518 7930
rect 17558 7908 17662 7930
rect 17558 7874 17622 7908
rect 17656 7874 17662 7908
rect 17558 7836 17662 7874
rect 17558 7802 17622 7836
rect 17656 7802 17662 7836
rect 17558 7764 17662 7802
rect 17558 7730 17622 7764
rect 17656 7730 17662 7764
rect 17558 7692 17662 7730
rect 17558 7658 17622 7692
rect 17656 7658 17662 7692
rect 17558 7620 17662 7658
rect 17558 7586 17622 7620
rect 17656 7586 17662 7620
rect 17558 7548 17662 7586
rect 17558 7514 17622 7548
rect 17656 7514 17662 7548
rect 17558 7476 17662 7514
rect 17558 7442 17622 7476
rect 17656 7442 17662 7476
rect 17558 7404 17662 7442
rect 17558 7370 17622 7404
rect 17656 7370 17662 7404
rect 17558 7332 17662 7370
rect 17558 7298 17622 7332
rect 17656 7298 17662 7332
rect 17558 7260 17662 7298
rect 17558 7226 17622 7260
rect 17656 7226 17662 7260
rect 17558 7188 17662 7226
rect 17558 7154 17622 7188
rect 17656 7154 17662 7188
rect 17558 7116 17662 7154
rect 17558 7082 17622 7116
rect 17656 7082 17662 7116
rect 17558 7044 17662 7082
rect 17558 7010 17622 7044
rect 17656 7010 17662 7044
rect 17558 6990 17662 7010
rect 17498 6972 17662 6990
rect 17699 7908 17751 7942
rect 17699 7874 17708 7908
rect 17742 7874 17751 7908
rect 17699 7836 17751 7874
rect 17699 7802 17708 7836
rect 17742 7802 17751 7836
rect 17699 7764 17751 7802
rect 17699 7730 17708 7764
rect 17742 7730 17751 7764
rect 17699 7692 17751 7730
rect 17699 7658 17708 7692
rect 17742 7658 17751 7692
rect 17699 7620 17751 7658
rect 17699 7586 17708 7620
rect 17742 7586 17751 7620
rect 17699 7548 17751 7586
rect 17699 7514 17708 7548
rect 17742 7514 17751 7548
rect 17699 7476 17751 7514
rect 17699 7442 17708 7476
rect 17742 7442 17751 7476
rect 17699 7404 17751 7442
rect 17699 7370 17708 7404
rect 17742 7370 17751 7404
rect 17699 7332 17751 7370
rect 17699 7298 17708 7332
rect 17742 7298 17751 7332
rect 17699 7260 17751 7298
rect 17699 7226 17708 7260
rect 17742 7226 17751 7260
rect 17699 7188 17751 7226
rect 17699 7154 17708 7188
rect 17742 7154 17751 7188
rect 17699 7116 17751 7154
rect 17699 7099 17708 7116
rect 17742 7099 17751 7116
rect 17699 7044 17751 7047
rect 17699 7035 17708 7044
rect 17742 7035 17751 7044
rect 17699 6972 17751 6983
rect 17788 7908 17834 8038
rect 17788 7874 17794 7908
rect 17828 7874 17834 7908
rect 17788 7836 17834 7874
rect 17788 7802 17794 7836
rect 17828 7802 17834 7836
rect 17788 7764 17834 7802
rect 17788 7730 17794 7764
rect 17828 7730 17834 7764
rect 17788 7692 17834 7730
rect 17788 7658 17794 7692
rect 17828 7658 17834 7692
rect 17788 7620 17834 7658
rect 17788 7586 17794 7620
rect 17828 7586 17834 7620
rect 17788 7548 17834 7586
rect 17788 7514 17794 7548
rect 17828 7514 17834 7548
rect 17788 7476 17834 7514
rect 17788 7442 17794 7476
rect 17828 7442 17834 7476
rect 17788 7404 17834 7442
rect 17788 7370 17794 7404
rect 17828 7370 17834 7404
rect 17788 7332 17834 7370
rect 17788 7298 17794 7332
rect 17828 7298 17834 7332
rect 17788 7260 17834 7298
rect 17788 7226 17794 7260
rect 17828 7226 17834 7260
rect 17788 7188 17834 7226
rect 17788 7154 17794 7188
rect 17828 7154 17834 7188
rect 17788 7116 17834 7154
rect 17788 7082 17794 7116
rect 17828 7082 17834 7116
rect 17788 7044 17834 7082
rect 17788 7010 17794 7044
rect 17828 7010 17834 7044
rect 17788 6972 17834 7010
rect 17871 7908 17923 7942
rect 17871 7874 17880 7908
rect 17914 7874 17923 7908
rect 17871 7836 17923 7874
rect 17871 7802 17880 7836
rect 17914 7802 17923 7836
rect 17871 7764 17923 7802
rect 17871 7730 17880 7764
rect 17914 7730 17923 7764
rect 17871 7692 17923 7730
rect 17871 7658 17880 7692
rect 17914 7658 17923 7692
rect 17871 7620 17923 7658
rect 17871 7586 17880 7620
rect 17914 7586 17923 7620
rect 17871 7548 17923 7586
rect 17871 7514 17880 7548
rect 17914 7514 17923 7548
rect 17871 7476 17923 7514
rect 17871 7442 17880 7476
rect 17914 7442 17923 7476
rect 17871 7404 17923 7442
rect 17871 7370 17880 7404
rect 17914 7370 17923 7404
rect 17871 7332 17923 7370
rect 17871 7298 17880 7332
rect 17914 7298 17923 7332
rect 17871 7260 17923 7298
rect 17871 7226 17880 7260
rect 17914 7226 17923 7260
rect 17871 7188 17923 7226
rect 17871 7154 17880 7188
rect 17914 7154 17923 7188
rect 17871 7116 17923 7154
rect 17871 7099 17880 7116
rect 17914 7099 17923 7116
rect 17871 7044 17923 7047
rect 17871 7035 17880 7044
rect 17914 7035 17923 7044
rect 17871 6972 17923 6983
rect 17960 7908 18006 8038
rect 17960 7874 17966 7908
rect 18000 7874 18006 7908
rect 17960 7836 18006 7874
rect 17960 7802 17966 7836
rect 18000 7802 18006 7836
rect 17960 7764 18006 7802
rect 17960 7730 17966 7764
rect 18000 7730 18006 7764
rect 17960 7692 18006 7730
rect 17960 7658 17966 7692
rect 18000 7658 18006 7692
rect 17960 7620 18006 7658
rect 17960 7586 17966 7620
rect 18000 7586 18006 7620
rect 17960 7548 18006 7586
rect 17960 7514 17966 7548
rect 18000 7514 18006 7548
rect 17960 7476 18006 7514
rect 17960 7442 17966 7476
rect 18000 7442 18006 7476
rect 17960 7404 18006 7442
rect 17960 7370 17966 7404
rect 18000 7370 18006 7404
rect 17960 7332 18006 7370
rect 17960 7298 17966 7332
rect 18000 7298 18006 7332
rect 17960 7260 18006 7298
rect 17960 7226 17966 7260
rect 18000 7226 18006 7260
rect 17960 7188 18006 7226
rect 17960 7154 17966 7188
rect 18000 7154 18006 7188
rect 17960 7116 18006 7154
rect 17960 7082 17966 7116
rect 18000 7082 18006 7116
rect 17960 7044 18006 7082
rect 17960 7010 17966 7044
rect 18000 7010 18006 7044
rect 17960 6972 18006 7010
rect 18043 7908 18095 7942
rect 18043 7874 18052 7908
rect 18086 7874 18095 7908
rect 18043 7836 18095 7874
rect 18043 7802 18052 7836
rect 18086 7802 18095 7836
rect 18043 7764 18095 7802
rect 18043 7730 18052 7764
rect 18086 7730 18095 7764
rect 18043 7692 18095 7730
rect 18043 7658 18052 7692
rect 18086 7658 18095 7692
rect 18043 7620 18095 7658
rect 18043 7586 18052 7620
rect 18086 7586 18095 7620
rect 18043 7548 18095 7586
rect 18043 7514 18052 7548
rect 18086 7514 18095 7548
rect 18043 7476 18095 7514
rect 18043 7442 18052 7476
rect 18086 7442 18095 7476
rect 18043 7404 18095 7442
rect 18043 7370 18052 7404
rect 18086 7370 18095 7404
rect 18043 7332 18095 7370
rect 18043 7298 18052 7332
rect 18086 7298 18095 7332
rect 18043 7260 18095 7298
rect 18043 7226 18052 7260
rect 18086 7226 18095 7260
rect 18043 7188 18095 7226
rect 18043 7154 18052 7188
rect 18086 7154 18095 7188
rect 18043 7116 18095 7154
rect 18043 7099 18052 7116
rect 18086 7099 18095 7116
rect 18043 7044 18095 7047
rect 18043 7035 18052 7044
rect 18086 7035 18095 7044
rect 18043 6972 18095 6983
rect 18132 7908 18178 8038
rect 18132 7874 18138 7908
rect 18172 7874 18178 7908
rect 18132 7836 18178 7874
rect 18132 7802 18138 7836
rect 18172 7802 18178 7836
rect 18132 7764 18178 7802
rect 18132 7730 18138 7764
rect 18172 7730 18178 7764
rect 18132 7692 18178 7730
rect 18132 7658 18138 7692
rect 18172 7658 18178 7692
rect 18132 7620 18178 7658
rect 18132 7586 18138 7620
rect 18172 7586 18178 7620
rect 18132 7548 18178 7586
rect 18132 7514 18138 7548
rect 18172 7514 18178 7548
rect 18132 7476 18178 7514
rect 18132 7442 18138 7476
rect 18172 7442 18178 7476
rect 18132 7404 18178 7442
rect 18132 7370 18138 7404
rect 18172 7370 18178 7404
rect 18132 7332 18178 7370
rect 18132 7298 18138 7332
rect 18172 7298 18178 7332
rect 18132 7260 18178 7298
rect 18132 7226 18138 7260
rect 18172 7226 18178 7260
rect 18132 7188 18178 7226
rect 18132 7154 18138 7188
rect 18172 7154 18178 7188
rect 18132 7116 18178 7154
rect 18132 7082 18138 7116
rect 18172 7082 18178 7116
rect 18132 7044 18178 7082
rect 18132 7010 18138 7044
rect 18172 7010 18178 7044
rect 18132 6972 18178 7010
rect 18215 7908 18267 7942
rect 18215 7874 18224 7908
rect 18258 7874 18267 7908
rect 18215 7836 18267 7874
rect 18215 7802 18224 7836
rect 18258 7802 18267 7836
rect 18215 7764 18267 7802
rect 18215 7730 18224 7764
rect 18258 7730 18267 7764
rect 18215 7692 18267 7730
rect 18215 7658 18224 7692
rect 18258 7658 18267 7692
rect 18215 7620 18267 7658
rect 18215 7586 18224 7620
rect 18258 7586 18267 7620
rect 18215 7548 18267 7586
rect 18215 7514 18224 7548
rect 18258 7514 18267 7548
rect 18215 7476 18267 7514
rect 18215 7442 18224 7476
rect 18258 7442 18267 7476
rect 18215 7404 18267 7442
rect 18215 7370 18224 7404
rect 18258 7370 18267 7404
rect 18215 7332 18267 7370
rect 18215 7298 18224 7332
rect 18258 7298 18267 7332
rect 18215 7260 18267 7298
rect 18215 7226 18224 7260
rect 18258 7226 18267 7260
rect 18215 7188 18267 7226
rect 18215 7154 18224 7188
rect 18258 7154 18267 7188
rect 18215 7116 18267 7154
rect 18215 7099 18224 7116
rect 18258 7099 18267 7116
rect 18215 7044 18267 7047
rect 18215 7035 18224 7044
rect 18258 7035 18267 7044
rect 18215 6972 18267 6983
rect 18304 7908 18350 8038
rect 18304 7874 18310 7908
rect 18344 7874 18350 7908
rect 18304 7836 18350 7874
rect 18304 7802 18310 7836
rect 18344 7802 18350 7836
rect 18304 7764 18350 7802
rect 18304 7730 18310 7764
rect 18344 7730 18350 7764
rect 18304 7692 18350 7730
rect 18304 7658 18310 7692
rect 18344 7658 18350 7692
rect 18304 7620 18350 7658
rect 18304 7586 18310 7620
rect 18344 7586 18350 7620
rect 18304 7548 18350 7586
rect 18304 7514 18310 7548
rect 18344 7514 18350 7548
rect 18304 7476 18350 7514
rect 18304 7442 18310 7476
rect 18344 7442 18350 7476
rect 18304 7404 18350 7442
rect 18304 7370 18310 7404
rect 18344 7370 18350 7404
rect 18304 7332 18350 7370
rect 18304 7298 18310 7332
rect 18344 7298 18350 7332
rect 18304 7260 18350 7298
rect 18304 7226 18310 7260
rect 18344 7226 18350 7260
rect 18304 7188 18350 7226
rect 18304 7154 18310 7188
rect 18344 7154 18350 7188
rect 18304 7116 18350 7154
rect 18304 7082 18310 7116
rect 18344 7082 18350 7116
rect 18304 7044 18350 7082
rect 18304 7010 18310 7044
rect 18344 7010 18350 7044
rect 18304 6972 18350 7010
rect 18387 7908 18439 7942
rect 18387 7874 18396 7908
rect 18430 7874 18439 7908
rect 18387 7836 18439 7874
rect 18387 7802 18396 7836
rect 18430 7802 18439 7836
rect 18387 7764 18439 7802
rect 18387 7730 18396 7764
rect 18430 7730 18439 7764
rect 18387 7692 18439 7730
rect 18387 7658 18396 7692
rect 18430 7658 18439 7692
rect 18387 7620 18439 7658
rect 18387 7586 18396 7620
rect 18430 7586 18439 7620
rect 18387 7548 18439 7586
rect 18387 7514 18396 7548
rect 18430 7514 18439 7548
rect 18387 7476 18439 7514
rect 18387 7442 18396 7476
rect 18430 7442 18439 7476
rect 18387 7404 18439 7442
rect 18387 7370 18396 7404
rect 18430 7370 18439 7404
rect 18387 7332 18439 7370
rect 18387 7298 18396 7332
rect 18430 7298 18439 7332
rect 18387 7260 18439 7298
rect 18387 7226 18396 7260
rect 18430 7226 18439 7260
rect 18387 7188 18439 7226
rect 18387 7154 18396 7188
rect 18430 7154 18439 7188
rect 18387 7116 18439 7154
rect 18387 7099 18396 7116
rect 18430 7099 18439 7116
rect 18387 7044 18439 7047
rect 18387 7035 18396 7044
rect 18430 7035 18439 7044
rect 18387 6972 18439 6983
rect 18476 7908 18522 8038
rect 18476 7874 18482 7908
rect 18516 7874 18522 7908
rect 18476 7836 18522 7874
rect 18476 7802 18482 7836
rect 18516 7802 18522 7836
rect 18476 7764 18522 7802
rect 18476 7730 18482 7764
rect 18516 7730 18522 7764
rect 18476 7692 18522 7730
rect 18476 7658 18482 7692
rect 18516 7658 18522 7692
rect 18476 7620 18522 7658
rect 18476 7586 18482 7620
rect 18516 7586 18522 7620
rect 18476 7548 18522 7586
rect 18476 7514 18482 7548
rect 18516 7514 18522 7548
rect 18476 7476 18522 7514
rect 18476 7442 18482 7476
rect 18516 7442 18522 7476
rect 18476 7404 18522 7442
rect 18476 7370 18482 7404
rect 18516 7370 18522 7404
rect 18476 7332 18522 7370
rect 18476 7298 18482 7332
rect 18516 7298 18522 7332
rect 18476 7260 18522 7298
rect 18476 7226 18482 7260
rect 18516 7226 18522 7260
rect 18476 7188 18522 7226
rect 18476 7154 18482 7188
rect 18516 7154 18522 7188
rect 18476 7116 18522 7154
rect 18476 7082 18482 7116
rect 18516 7082 18522 7116
rect 18476 7044 18522 7082
rect 18476 7010 18482 7044
rect 18516 7010 18522 7044
rect 18476 6972 18522 7010
rect 18559 7908 18611 7942
rect 18559 7874 18568 7908
rect 18602 7874 18611 7908
rect 18559 7836 18611 7874
rect 18559 7802 18568 7836
rect 18602 7802 18611 7836
rect 18559 7764 18611 7802
rect 18559 7730 18568 7764
rect 18602 7730 18611 7764
rect 18559 7692 18611 7730
rect 18559 7658 18568 7692
rect 18602 7658 18611 7692
rect 18559 7620 18611 7658
rect 18559 7586 18568 7620
rect 18602 7586 18611 7620
rect 18559 7548 18611 7586
rect 18559 7514 18568 7548
rect 18602 7514 18611 7548
rect 18559 7476 18611 7514
rect 18559 7442 18568 7476
rect 18602 7442 18611 7476
rect 18559 7404 18611 7442
rect 18559 7370 18568 7404
rect 18602 7370 18611 7404
rect 18559 7332 18611 7370
rect 18559 7298 18568 7332
rect 18602 7298 18611 7332
rect 18559 7260 18611 7298
rect 18559 7226 18568 7260
rect 18602 7226 18611 7260
rect 18559 7188 18611 7226
rect 18559 7154 18568 7188
rect 18602 7154 18611 7188
rect 18559 7116 18611 7154
rect 18559 7099 18568 7116
rect 18602 7099 18611 7116
rect 18559 7044 18611 7047
rect 18559 7035 18568 7044
rect 18602 7035 18611 7044
rect 18559 6972 18611 6983
rect 18648 7908 18694 8038
rect 18648 7874 18654 7908
rect 18688 7874 18694 7908
rect 18648 7836 18694 7874
rect 18648 7802 18654 7836
rect 18688 7802 18694 7836
rect 18648 7764 18694 7802
rect 18648 7730 18654 7764
rect 18688 7730 18694 7764
rect 18648 7692 18694 7730
rect 18648 7658 18654 7692
rect 18688 7658 18694 7692
rect 18648 7620 18694 7658
rect 18648 7586 18654 7620
rect 18688 7586 18694 7620
rect 18648 7548 18694 7586
rect 18648 7514 18654 7548
rect 18688 7514 18694 7548
rect 18648 7476 18694 7514
rect 18648 7442 18654 7476
rect 18688 7442 18694 7476
rect 18648 7404 18694 7442
rect 18648 7370 18654 7404
rect 18688 7370 18694 7404
rect 18648 7332 18694 7370
rect 18648 7298 18654 7332
rect 18688 7298 18694 7332
rect 18648 7260 18694 7298
rect 18648 7226 18654 7260
rect 18688 7226 18694 7260
rect 18648 7188 18694 7226
rect 18648 7154 18654 7188
rect 18688 7154 18694 7188
rect 18648 7116 18694 7154
rect 18648 7082 18654 7116
rect 18688 7082 18694 7116
rect 18648 7044 18694 7082
rect 18648 7010 18654 7044
rect 18688 7010 18694 7044
rect 18648 6972 18694 7010
rect 18731 7908 18783 7942
rect 18731 7874 18740 7908
rect 18774 7874 18783 7908
rect 18731 7836 18783 7874
rect 18731 7802 18740 7836
rect 18774 7802 18783 7836
rect 18731 7764 18783 7802
rect 18731 7730 18740 7764
rect 18774 7730 18783 7764
rect 18731 7692 18783 7730
rect 18731 7658 18740 7692
rect 18774 7658 18783 7692
rect 18731 7620 18783 7658
rect 18731 7586 18740 7620
rect 18774 7586 18783 7620
rect 18731 7548 18783 7586
rect 18731 7514 18740 7548
rect 18774 7514 18783 7548
rect 18731 7476 18783 7514
rect 18731 7442 18740 7476
rect 18774 7442 18783 7476
rect 18731 7404 18783 7442
rect 18731 7370 18740 7404
rect 18774 7370 18783 7404
rect 18731 7332 18783 7370
rect 18731 7298 18740 7332
rect 18774 7298 18783 7332
rect 18731 7260 18783 7298
rect 18731 7226 18740 7260
rect 18774 7226 18783 7260
rect 18731 7188 18783 7226
rect 18731 7154 18740 7188
rect 18774 7154 18783 7188
rect 18731 7116 18783 7154
rect 18731 7099 18740 7116
rect 18774 7099 18783 7116
rect 18731 7044 18783 7047
rect 18731 7035 18740 7044
rect 18774 7035 18783 7044
rect 18731 6972 18783 6983
rect 18820 7908 18866 8038
rect 18820 7874 18826 7908
rect 18860 7874 18866 7908
rect 18820 7836 18866 7874
rect 18820 7802 18826 7836
rect 18860 7802 18866 7836
rect 18820 7764 18866 7802
rect 18820 7730 18826 7764
rect 18860 7730 18866 7764
rect 18820 7692 18866 7730
rect 18820 7658 18826 7692
rect 18860 7658 18866 7692
rect 18820 7620 18866 7658
rect 18820 7586 18826 7620
rect 18860 7586 18866 7620
rect 18820 7548 18866 7586
rect 18820 7514 18826 7548
rect 18860 7514 18866 7548
rect 18820 7476 18866 7514
rect 18820 7442 18826 7476
rect 18860 7442 18866 7476
rect 18820 7404 18866 7442
rect 18820 7370 18826 7404
rect 18860 7370 18866 7404
rect 18820 7332 18866 7370
rect 18820 7298 18826 7332
rect 18860 7298 18866 7332
rect 18820 7260 18866 7298
rect 18820 7226 18826 7260
rect 18860 7226 18866 7260
rect 18820 7188 18866 7226
rect 18820 7154 18826 7188
rect 18860 7154 18866 7188
rect 18820 7116 18866 7154
rect 18820 7082 18826 7116
rect 18860 7082 18866 7116
rect 18820 7044 18866 7082
rect 18820 7010 18826 7044
rect 18860 7010 18866 7044
rect 18820 6972 18866 7010
rect 18903 7908 18955 7942
rect 18903 7874 18912 7908
rect 18946 7874 18955 7908
rect 18903 7836 18955 7874
rect 18903 7802 18912 7836
rect 18946 7802 18955 7836
rect 18903 7764 18955 7802
rect 18903 7730 18912 7764
rect 18946 7730 18955 7764
rect 18903 7692 18955 7730
rect 18903 7658 18912 7692
rect 18946 7658 18955 7692
rect 18903 7620 18955 7658
rect 18903 7586 18912 7620
rect 18946 7586 18955 7620
rect 18903 7548 18955 7586
rect 18903 7514 18912 7548
rect 18946 7514 18955 7548
rect 18903 7476 18955 7514
rect 18903 7442 18912 7476
rect 18946 7442 18955 7476
rect 18903 7404 18955 7442
rect 18903 7370 18912 7404
rect 18946 7370 18955 7404
rect 18903 7332 18955 7370
rect 18903 7298 18912 7332
rect 18946 7298 18955 7332
rect 18903 7260 18955 7298
rect 18903 7226 18912 7260
rect 18946 7226 18955 7260
rect 18903 7188 18955 7226
rect 18903 7154 18912 7188
rect 18946 7154 18955 7188
rect 18903 7116 18955 7154
rect 18903 7099 18912 7116
rect 18946 7099 18955 7116
rect 18903 7044 18955 7047
rect 18903 7035 18912 7044
rect 18946 7035 18955 7044
rect 18903 6972 18955 6983
rect 18992 7908 19038 8038
rect 18992 7874 18998 7908
rect 19032 7874 19038 7908
rect 18992 7836 19038 7874
rect 18992 7802 18998 7836
rect 19032 7802 19038 7836
rect 18992 7764 19038 7802
rect 18992 7730 18998 7764
rect 19032 7730 19038 7764
rect 18992 7692 19038 7730
rect 18992 7658 18998 7692
rect 19032 7658 19038 7692
rect 18992 7620 19038 7658
rect 18992 7586 18998 7620
rect 19032 7586 19038 7620
rect 18992 7548 19038 7586
rect 18992 7514 18998 7548
rect 19032 7514 19038 7548
rect 18992 7476 19038 7514
rect 18992 7442 18998 7476
rect 19032 7442 19038 7476
rect 18992 7404 19038 7442
rect 18992 7370 18998 7404
rect 19032 7370 19038 7404
rect 18992 7332 19038 7370
rect 18992 7298 18998 7332
rect 19032 7298 19038 7332
rect 18992 7260 19038 7298
rect 18992 7226 18998 7260
rect 19032 7226 19038 7260
rect 18992 7188 19038 7226
rect 18992 7154 18998 7188
rect 19032 7154 19038 7188
rect 18992 7116 19038 7154
rect 18992 7082 18998 7116
rect 19032 7082 19038 7116
rect 18992 7044 19038 7082
rect 18992 7010 18998 7044
rect 19032 7010 19038 7044
rect 18992 6972 19038 7010
rect 19075 7908 19127 7942
rect 19075 7874 19084 7908
rect 19118 7874 19127 7908
rect 19075 7836 19127 7874
rect 19075 7802 19084 7836
rect 19118 7802 19127 7836
rect 19075 7764 19127 7802
rect 19075 7730 19084 7764
rect 19118 7730 19127 7764
rect 19075 7692 19127 7730
rect 19075 7658 19084 7692
rect 19118 7658 19127 7692
rect 19075 7620 19127 7658
rect 19075 7586 19084 7620
rect 19118 7586 19127 7620
rect 19075 7548 19127 7586
rect 19075 7514 19084 7548
rect 19118 7514 19127 7548
rect 19075 7476 19127 7514
rect 19075 7442 19084 7476
rect 19118 7442 19127 7476
rect 19075 7404 19127 7442
rect 19075 7370 19084 7404
rect 19118 7370 19127 7404
rect 19075 7332 19127 7370
rect 19075 7298 19084 7332
rect 19118 7298 19127 7332
rect 19075 7260 19127 7298
rect 19075 7226 19084 7260
rect 19118 7226 19127 7260
rect 19075 7188 19127 7226
rect 19075 7154 19084 7188
rect 19118 7154 19127 7188
rect 19075 7116 19127 7154
rect 19075 7099 19084 7116
rect 19118 7099 19127 7116
rect 19075 7044 19127 7047
rect 19075 7035 19084 7044
rect 19118 7035 19127 7044
rect 19075 6972 19127 6983
rect 19164 7908 19210 8038
rect 19164 7874 19170 7908
rect 19204 7874 19210 7908
rect 19164 7836 19210 7874
rect 19164 7802 19170 7836
rect 19204 7802 19210 7836
rect 19164 7764 19210 7802
rect 19164 7730 19170 7764
rect 19204 7730 19210 7764
rect 19164 7692 19210 7730
rect 19164 7658 19170 7692
rect 19204 7658 19210 7692
rect 19164 7620 19210 7658
rect 19164 7586 19170 7620
rect 19204 7586 19210 7620
rect 19164 7548 19210 7586
rect 19164 7514 19170 7548
rect 19204 7514 19210 7548
rect 19164 7476 19210 7514
rect 19164 7442 19170 7476
rect 19204 7442 19210 7476
rect 19164 7404 19210 7442
rect 19164 7370 19170 7404
rect 19204 7370 19210 7404
rect 19164 7332 19210 7370
rect 19164 7298 19170 7332
rect 19204 7298 19210 7332
rect 19164 7260 19210 7298
rect 19164 7226 19170 7260
rect 19204 7226 19210 7260
rect 19164 7188 19210 7226
rect 19164 7154 19170 7188
rect 19204 7154 19210 7188
rect 19164 7116 19210 7154
rect 19164 7082 19170 7116
rect 19204 7082 19210 7116
rect 19164 7044 19210 7082
rect 19164 7010 19170 7044
rect 19204 7010 19210 7044
rect 19164 6972 19210 7010
rect 19247 7908 19299 7942
rect 19247 7874 19256 7908
rect 19290 7874 19299 7908
rect 19247 7836 19299 7874
rect 19247 7802 19256 7836
rect 19290 7802 19299 7836
rect 19247 7764 19299 7802
rect 19247 7730 19256 7764
rect 19290 7730 19299 7764
rect 19247 7692 19299 7730
rect 19247 7658 19256 7692
rect 19290 7658 19299 7692
rect 19247 7620 19299 7658
rect 19247 7586 19256 7620
rect 19290 7586 19299 7620
rect 19247 7548 19299 7586
rect 19247 7514 19256 7548
rect 19290 7514 19299 7548
rect 19247 7476 19299 7514
rect 19247 7442 19256 7476
rect 19290 7442 19299 7476
rect 19247 7404 19299 7442
rect 19247 7370 19256 7404
rect 19290 7370 19299 7404
rect 19247 7332 19299 7370
rect 19247 7298 19256 7332
rect 19290 7298 19299 7332
rect 19247 7260 19299 7298
rect 19247 7226 19256 7260
rect 19290 7226 19299 7260
rect 19247 7188 19299 7226
rect 19247 7154 19256 7188
rect 19290 7154 19299 7188
rect 19247 7116 19299 7154
rect 19247 7099 19256 7116
rect 19290 7099 19299 7116
rect 19247 7044 19299 7047
rect 19247 7035 19256 7044
rect 19290 7035 19299 7044
rect 19247 6972 19299 6983
rect 19336 7908 19382 8038
rect 19336 7874 19342 7908
rect 19376 7874 19382 7908
rect 19336 7836 19382 7874
rect 19336 7802 19342 7836
rect 19376 7802 19382 7836
rect 19336 7764 19382 7802
rect 19336 7730 19342 7764
rect 19376 7730 19382 7764
rect 19336 7692 19382 7730
rect 19336 7658 19342 7692
rect 19376 7658 19382 7692
rect 19336 7620 19382 7658
rect 19336 7586 19342 7620
rect 19376 7586 19382 7620
rect 19336 7548 19382 7586
rect 19336 7514 19342 7548
rect 19376 7514 19382 7548
rect 19336 7476 19382 7514
rect 19336 7442 19342 7476
rect 19376 7442 19382 7476
rect 19336 7404 19382 7442
rect 19336 7370 19342 7404
rect 19376 7370 19382 7404
rect 19336 7332 19382 7370
rect 19336 7298 19342 7332
rect 19376 7298 19382 7332
rect 19336 7260 19382 7298
rect 19336 7226 19342 7260
rect 19376 7226 19382 7260
rect 19336 7188 19382 7226
rect 19336 7154 19342 7188
rect 19376 7154 19382 7188
rect 19336 7116 19382 7154
rect 19336 7082 19342 7116
rect 19376 7082 19382 7116
rect 19336 7044 19382 7082
rect 19336 7010 19342 7044
rect 19376 7010 19382 7044
rect 19336 6972 19382 7010
rect 19419 7908 19471 7942
rect 19419 7874 19428 7908
rect 19462 7874 19471 7908
rect 19419 7836 19471 7874
rect 19419 7802 19428 7836
rect 19462 7802 19471 7836
rect 19419 7764 19471 7802
rect 19419 7730 19428 7764
rect 19462 7730 19471 7764
rect 19419 7692 19471 7730
rect 19419 7658 19428 7692
rect 19462 7658 19471 7692
rect 19419 7620 19471 7658
rect 19419 7586 19428 7620
rect 19462 7586 19471 7620
rect 19419 7548 19471 7586
rect 19419 7514 19428 7548
rect 19462 7514 19471 7548
rect 19419 7476 19471 7514
rect 19419 7442 19428 7476
rect 19462 7442 19471 7476
rect 19419 7404 19471 7442
rect 19419 7370 19428 7404
rect 19462 7370 19471 7404
rect 19419 7332 19471 7370
rect 19419 7298 19428 7332
rect 19462 7298 19471 7332
rect 19419 7260 19471 7298
rect 19419 7226 19428 7260
rect 19462 7226 19471 7260
rect 19419 7188 19471 7226
rect 19419 7154 19428 7188
rect 19462 7154 19471 7188
rect 19419 7116 19471 7154
rect 19419 7099 19428 7116
rect 19462 7099 19471 7116
rect 19419 7044 19471 7047
rect 19419 7035 19428 7044
rect 19462 7035 19471 7044
rect 19419 6972 19471 6983
rect 19508 7908 19554 8038
rect 19508 7874 19514 7908
rect 19548 7874 19554 7908
rect 19508 7836 19554 7874
rect 19508 7802 19514 7836
rect 19548 7802 19554 7836
rect 19508 7764 19554 7802
rect 19508 7730 19514 7764
rect 19548 7730 19554 7764
rect 19508 7692 19554 7730
rect 19508 7658 19514 7692
rect 19548 7658 19554 7692
rect 19508 7620 19554 7658
rect 19508 7586 19514 7620
rect 19548 7586 19554 7620
rect 19508 7548 19554 7586
rect 19508 7514 19514 7548
rect 19548 7514 19554 7548
rect 19508 7476 19554 7514
rect 19508 7442 19514 7476
rect 19548 7442 19554 7476
rect 19508 7404 19554 7442
rect 19508 7370 19514 7404
rect 19548 7370 19554 7404
rect 19508 7332 19554 7370
rect 19508 7298 19514 7332
rect 19548 7298 19554 7332
rect 19508 7260 19554 7298
rect 19508 7226 19514 7260
rect 19548 7226 19554 7260
rect 19508 7188 19554 7226
rect 19508 7154 19514 7188
rect 19548 7154 19554 7188
rect 19508 7116 19554 7154
rect 19508 7082 19514 7116
rect 19548 7082 19554 7116
rect 19508 7044 19554 7082
rect 19508 7010 19514 7044
rect 19548 7010 19554 7044
rect 19508 6972 19554 7010
rect 19591 7908 19643 7942
rect 19591 7874 19600 7908
rect 19634 7874 19643 7908
rect 19591 7836 19643 7874
rect 19591 7802 19600 7836
rect 19634 7802 19643 7836
rect 19591 7764 19643 7802
rect 19591 7730 19600 7764
rect 19634 7730 19643 7764
rect 19591 7692 19643 7730
rect 19591 7658 19600 7692
rect 19634 7658 19643 7692
rect 19591 7620 19643 7658
rect 19591 7586 19600 7620
rect 19634 7586 19643 7620
rect 19591 7548 19643 7586
rect 19591 7514 19600 7548
rect 19634 7514 19643 7548
rect 19591 7476 19643 7514
rect 19591 7442 19600 7476
rect 19634 7442 19643 7476
rect 19591 7404 19643 7442
rect 19591 7370 19600 7404
rect 19634 7370 19643 7404
rect 19591 7332 19643 7370
rect 19591 7298 19600 7332
rect 19634 7298 19643 7332
rect 19591 7260 19643 7298
rect 19591 7226 19600 7260
rect 19634 7226 19643 7260
rect 19591 7188 19643 7226
rect 19591 7154 19600 7188
rect 19634 7154 19643 7188
rect 19591 7116 19643 7154
rect 19591 7099 19600 7116
rect 19634 7099 19643 7116
rect 19591 7044 19643 7047
rect 19591 7035 19600 7044
rect 19634 7035 19643 7044
rect 19591 6972 19643 6983
rect 19680 7908 19726 8038
rect 19680 7874 19686 7908
rect 19720 7874 19726 7908
rect 19680 7836 19726 7874
rect 19680 7802 19686 7836
rect 19720 7802 19726 7836
rect 19680 7764 19726 7802
rect 19680 7730 19686 7764
rect 19720 7730 19726 7764
rect 19680 7692 19726 7730
rect 19680 7658 19686 7692
rect 19720 7658 19726 7692
rect 19680 7620 19726 7658
rect 19680 7586 19686 7620
rect 19720 7586 19726 7620
rect 19680 7548 19726 7586
rect 19680 7514 19686 7548
rect 19720 7514 19726 7548
rect 19680 7476 19726 7514
rect 19680 7442 19686 7476
rect 19720 7442 19726 7476
rect 19680 7404 19726 7442
rect 19680 7370 19686 7404
rect 19720 7370 19726 7404
rect 19680 7332 19726 7370
rect 19680 7298 19686 7332
rect 19720 7298 19726 7332
rect 19680 7260 19726 7298
rect 19680 7226 19686 7260
rect 19720 7226 19726 7260
rect 19680 7188 19726 7226
rect 19680 7154 19686 7188
rect 19720 7154 19726 7188
rect 19680 7116 19726 7154
rect 19680 7082 19686 7116
rect 19720 7082 19726 7116
rect 19680 7044 19726 7082
rect 19680 7010 19686 7044
rect 19720 7010 19726 7044
rect 19680 6972 19726 7010
rect 19763 7908 19815 7942
rect 19763 7874 19772 7908
rect 19806 7874 19815 7908
rect 19763 7836 19815 7874
rect 19763 7802 19772 7836
rect 19806 7802 19815 7836
rect 19763 7764 19815 7802
rect 19763 7730 19772 7764
rect 19806 7730 19815 7764
rect 19763 7692 19815 7730
rect 19763 7658 19772 7692
rect 19806 7658 19815 7692
rect 19763 7620 19815 7658
rect 19763 7586 19772 7620
rect 19806 7586 19815 7620
rect 19763 7548 19815 7586
rect 19763 7514 19772 7548
rect 19806 7514 19815 7548
rect 19763 7476 19815 7514
rect 19763 7442 19772 7476
rect 19806 7442 19815 7476
rect 19763 7404 19815 7442
rect 19763 7370 19772 7404
rect 19806 7370 19815 7404
rect 19763 7332 19815 7370
rect 19763 7298 19772 7332
rect 19806 7298 19815 7332
rect 19763 7260 19815 7298
rect 19763 7226 19772 7260
rect 19806 7226 19815 7260
rect 19763 7188 19815 7226
rect 19763 7154 19772 7188
rect 19806 7154 19815 7188
rect 19763 7116 19815 7154
rect 19763 7099 19772 7116
rect 19806 7099 19815 7116
rect 19763 7044 19815 7047
rect 19763 7035 19772 7044
rect 19806 7035 19815 7044
rect 19763 6972 19815 6983
rect 19852 7908 19898 8038
rect 20024 7950 20070 8038
rect 19852 7874 19858 7908
rect 19892 7874 19898 7908
rect 19852 7836 19898 7874
rect 19852 7802 19858 7836
rect 19892 7802 19898 7836
rect 19852 7764 19898 7802
rect 19852 7730 19858 7764
rect 19892 7730 19898 7764
rect 19852 7692 19898 7730
rect 19852 7658 19858 7692
rect 19892 7658 19898 7692
rect 19852 7620 19898 7658
rect 19852 7586 19858 7620
rect 19892 7586 19898 7620
rect 19852 7548 19898 7586
rect 19852 7514 19858 7548
rect 19892 7514 19898 7548
rect 19852 7476 19898 7514
rect 19852 7442 19858 7476
rect 19892 7442 19898 7476
rect 19852 7404 19898 7442
rect 19852 7370 19858 7404
rect 19892 7370 19898 7404
rect 19852 7332 19898 7370
rect 19852 7298 19858 7332
rect 19892 7298 19898 7332
rect 19852 7260 19898 7298
rect 19852 7226 19858 7260
rect 19892 7226 19898 7260
rect 19852 7188 19898 7226
rect 19852 7154 19858 7188
rect 19892 7154 19898 7188
rect 19852 7116 19898 7154
rect 19852 7082 19858 7116
rect 19892 7082 19898 7116
rect 19852 7044 19898 7082
rect 19852 7010 19858 7044
rect 19892 7010 19898 7044
rect 19852 6972 19898 7010
rect 19935 7908 19987 7942
rect 19935 7874 19944 7908
rect 19978 7874 19987 7908
rect 19935 7836 19987 7874
rect 19935 7802 19944 7836
rect 19978 7802 19987 7836
rect 19935 7764 19987 7802
rect 19935 7730 19944 7764
rect 19978 7730 19987 7764
rect 19935 7692 19987 7730
rect 19935 7658 19944 7692
rect 19978 7658 19987 7692
rect 19935 7620 19987 7658
rect 19935 7586 19944 7620
rect 19978 7586 19987 7620
rect 19935 7548 19987 7586
rect 19935 7514 19944 7548
rect 19978 7514 19987 7548
rect 19935 7476 19987 7514
rect 19935 7442 19944 7476
rect 19978 7442 19987 7476
rect 19935 7404 19987 7442
rect 19935 7370 19944 7404
rect 19978 7370 19987 7404
rect 19935 7332 19987 7370
rect 19935 7298 19944 7332
rect 19978 7298 19987 7332
rect 19935 7260 19987 7298
rect 19935 7226 19944 7260
rect 19978 7226 19987 7260
rect 19935 7188 19987 7226
rect 19935 7154 19944 7188
rect 19978 7154 19987 7188
rect 19935 7116 19987 7154
rect 19935 7099 19944 7116
rect 19978 7099 19987 7116
rect 19935 7044 19987 7047
rect 19935 7035 19944 7044
rect 19978 7035 19987 7044
rect 19935 6972 19987 6983
rect 20024 7930 20198 7950
rect 20024 7908 20060 7930
rect 20024 7874 20030 7908
rect 20024 7836 20060 7874
rect 20024 7802 20030 7836
rect 20024 7764 20060 7802
rect 20024 7730 20030 7764
rect 20024 7692 20060 7730
rect 20024 7658 20030 7692
rect 20024 7620 20060 7658
rect 20024 7586 20030 7620
rect 20024 7548 20060 7586
rect 20024 7514 20030 7548
rect 20024 7476 20060 7514
rect 20024 7442 20030 7476
rect 20024 7404 20060 7442
rect 20024 7370 20030 7404
rect 20024 7332 20060 7370
rect 20024 7298 20030 7332
rect 20024 7260 20060 7298
rect 20024 7226 20030 7260
rect 20024 7188 20060 7226
rect 20024 7154 20030 7188
rect 20024 7116 20060 7154
rect 20024 7082 20030 7116
rect 20024 7044 20060 7082
rect 20024 7010 20030 7044
rect 20024 7000 20060 7010
rect 20180 7000 20198 7930
rect 20024 6990 20138 7000
rect 20178 6990 20198 7000
rect 20024 6972 20198 6990
rect 17498 6970 17658 6972
rect 20038 6970 20198 6972
rect 11801 6930 12147 6950
rect 11801 6896 11813 6930
rect 11847 6896 11885 6930
rect 11919 6896 11957 6930
rect 11991 6896 12029 6930
rect 12063 6896 12101 6930
rect 12135 6896 12147 6930
rect 11801 6884 12147 6896
rect 12367 6930 12713 6950
rect 12367 6896 12379 6930
rect 12413 6896 12451 6930
rect 12485 6896 12523 6930
rect 12557 6896 12595 6930
rect 12629 6896 12667 6930
rect 12701 6896 12713 6930
rect 12367 6884 12713 6896
rect 12933 6930 13279 6950
rect 12933 6896 12945 6930
rect 12979 6896 13017 6930
rect 13051 6896 13089 6930
rect 13123 6896 13161 6930
rect 13195 6896 13233 6930
rect 13267 6896 13279 6930
rect 12933 6884 13279 6896
rect 13499 6930 13845 6950
rect 13499 6896 13511 6930
rect 13545 6896 13583 6930
rect 13617 6896 13655 6930
rect 13689 6896 13727 6930
rect 13761 6896 13799 6930
rect 13833 6896 13845 6930
rect 13499 6884 13845 6896
rect 14065 6930 14411 6950
rect 14065 6896 14077 6930
rect 14111 6896 14149 6930
rect 14183 6896 14221 6930
rect 14255 6896 14293 6930
rect 14327 6896 14365 6930
rect 14399 6896 14411 6930
rect 14065 6884 14411 6896
rect 14631 6930 14977 6950
rect 14631 6896 14643 6930
rect 14677 6896 14715 6930
rect 14749 6896 14787 6930
rect 14821 6896 14859 6930
rect 14893 6896 14931 6930
rect 14965 6896 14977 6930
rect 14631 6884 14977 6896
rect 15197 6930 15543 6950
rect 15197 6896 15209 6930
rect 15243 6896 15281 6930
rect 15315 6896 15353 6930
rect 15387 6896 15425 6930
rect 15459 6896 15497 6930
rect 15531 6896 15543 6930
rect 15197 6884 15543 6896
rect 16134 6931 17168 6943
rect 16134 6897 16218 6931
rect 16252 6897 16290 6931
rect 16324 6897 16362 6931
rect 16396 6897 16562 6931
rect 16596 6897 16634 6931
rect 16668 6897 16706 6931
rect 16740 6897 16906 6931
rect 16940 6897 16978 6931
rect 17012 6897 17050 6931
rect 17084 6897 17168 6931
rect 11662 6838 11720 6850
rect 11662 6804 11674 6838
rect 11708 6804 11720 6838
rect 11662 6766 11720 6804
rect 11662 6732 11674 6766
rect 11708 6732 11720 6766
rect 11662 6694 11720 6732
rect 11662 6660 11674 6694
rect 11708 6660 11720 6694
rect 11662 6622 11720 6660
rect 11662 6588 11674 6622
rect 11708 6588 11720 6622
rect 11662 6550 11720 6588
rect 11662 6516 11674 6550
rect 11708 6516 11720 6550
rect 11662 6478 11720 6516
rect 11662 6444 11674 6478
rect 11708 6444 11720 6478
rect 11662 6406 11720 6444
rect 11662 6372 11674 6406
rect 11708 6372 11720 6406
rect 11662 6334 11720 6372
rect 11662 6300 11674 6334
rect 11708 6300 11720 6334
rect 11662 6262 11720 6300
rect 11662 6228 11674 6262
rect 11708 6228 11720 6262
rect 11662 6190 11720 6228
rect 11662 6156 11674 6190
rect 11708 6156 11720 6190
rect 11662 6118 11720 6156
rect 11662 6084 11674 6118
rect 11708 6084 11720 6118
rect 11662 6046 11720 6084
rect 11662 6012 11674 6046
rect 11708 6012 11720 6046
rect 11662 5974 11720 6012
rect 11662 5940 11674 5974
rect 11708 5940 11720 5974
rect 11662 5902 11720 5940
rect 11662 5868 11674 5902
rect 11708 5868 11720 5902
rect 11662 5470 11720 5868
rect 11776 6844 11828 6850
rect 11776 6780 11828 6792
rect 11776 6716 11828 6728
rect 11776 6660 11785 6664
rect 11819 6660 11828 6664
rect 11776 6652 11828 6660
rect 11776 6588 11785 6600
rect 11819 6588 11828 6600
rect 11776 6524 11785 6536
rect 11819 6524 11828 6536
rect 11776 6460 11785 6472
rect 11819 6460 11828 6472
rect 11776 6406 11828 6408
rect 11776 6396 11785 6406
rect 11819 6396 11828 6406
rect 11776 6334 11828 6344
rect 11776 6332 11785 6334
rect 11819 6332 11828 6334
rect 11776 6268 11828 6280
rect 11776 6204 11828 6216
rect 11776 6140 11828 6152
rect 11776 6084 11785 6088
rect 11819 6084 11828 6088
rect 11776 6076 11828 6084
rect 11776 6012 11785 6024
rect 11819 6012 11828 6024
rect 11776 5948 11785 5960
rect 11819 5948 11828 5960
rect 11776 5868 11785 5896
rect 11819 5868 11828 5896
rect 11776 5856 11828 5868
rect 11862 6838 11914 6850
rect 11862 6810 11871 6838
rect 11905 6810 11914 6838
rect 11862 6746 11871 6758
rect 11905 6746 11914 6758
rect 11862 6682 11871 6694
rect 11905 6682 11914 6694
rect 11862 6622 11914 6630
rect 11862 6618 11871 6622
rect 11905 6618 11914 6622
rect 11862 6554 11914 6566
rect 11862 6490 11914 6502
rect 11862 6426 11914 6438
rect 11862 6372 11871 6374
rect 11905 6372 11914 6374
rect 11862 6362 11914 6372
rect 11862 6300 11871 6310
rect 11905 6300 11914 6310
rect 11862 6298 11914 6300
rect 11862 6234 11871 6246
rect 11905 6234 11914 6246
rect 11862 6170 11871 6182
rect 11905 6170 11914 6182
rect 11862 6106 11871 6118
rect 11905 6106 11914 6118
rect 11862 6046 11914 6054
rect 11862 6042 11871 6046
rect 11905 6042 11914 6046
rect 11862 5978 11914 5990
rect 11862 5914 11914 5926
rect 11862 5856 11914 5862
rect 11948 6844 12000 6850
rect 11948 6780 12000 6792
rect 11948 6716 12000 6728
rect 11948 6660 11957 6664
rect 11991 6660 12000 6664
rect 11948 6652 12000 6660
rect 11948 6588 11957 6600
rect 11991 6588 12000 6600
rect 11948 6524 11957 6536
rect 11991 6524 12000 6536
rect 11948 6460 11957 6472
rect 11991 6460 12000 6472
rect 11948 6406 12000 6408
rect 11948 6396 11957 6406
rect 11991 6396 12000 6406
rect 11948 6334 12000 6344
rect 11948 6332 11957 6334
rect 11991 6332 12000 6334
rect 11948 6268 12000 6280
rect 11948 6204 12000 6216
rect 11948 6140 12000 6152
rect 11948 6084 11957 6088
rect 11991 6084 12000 6088
rect 11948 6076 12000 6084
rect 11948 6012 11957 6024
rect 11991 6012 12000 6024
rect 11948 5948 11957 5960
rect 11991 5948 12000 5960
rect 11948 5868 11957 5896
rect 11991 5868 12000 5896
rect 11948 5856 12000 5868
rect 12034 6838 12086 6850
rect 12034 6810 12043 6838
rect 12077 6810 12086 6838
rect 12034 6746 12043 6758
rect 12077 6746 12086 6758
rect 12034 6682 12043 6694
rect 12077 6682 12086 6694
rect 12034 6622 12086 6630
rect 12034 6618 12043 6622
rect 12077 6618 12086 6622
rect 12034 6554 12086 6566
rect 12034 6490 12086 6502
rect 12034 6426 12086 6438
rect 12034 6372 12043 6374
rect 12077 6372 12086 6374
rect 12034 6362 12086 6372
rect 12034 6300 12043 6310
rect 12077 6300 12086 6310
rect 12034 6298 12086 6300
rect 12034 6234 12043 6246
rect 12077 6234 12086 6246
rect 12034 6170 12043 6182
rect 12077 6170 12086 6182
rect 12034 6106 12043 6118
rect 12077 6106 12086 6118
rect 12034 6046 12086 6054
rect 12034 6042 12043 6046
rect 12077 6042 12086 6046
rect 12034 5978 12086 5990
rect 12034 5914 12086 5926
rect 12034 5856 12086 5862
rect 12120 6844 12172 6850
rect 12120 6780 12172 6792
rect 12120 6716 12172 6728
rect 12120 6660 12129 6664
rect 12163 6660 12172 6664
rect 12120 6652 12172 6660
rect 12120 6588 12129 6600
rect 12163 6588 12172 6600
rect 12120 6524 12129 6536
rect 12163 6524 12172 6536
rect 12120 6460 12129 6472
rect 12163 6460 12172 6472
rect 12120 6406 12172 6408
rect 12120 6396 12129 6406
rect 12163 6396 12172 6406
rect 12120 6334 12172 6344
rect 12120 6332 12129 6334
rect 12163 6332 12172 6334
rect 12120 6268 12172 6280
rect 12120 6204 12172 6216
rect 12120 6140 12172 6152
rect 12120 6084 12129 6088
rect 12163 6084 12172 6088
rect 12120 6076 12172 6084
rect 12120 6012 12129 6024
rect 12163 6012 12172 6024
rect 12120 5948 12129 5960
rect 12163 5948 12172 5960
rect 12120 5868 12129 5896
rect 12163 5868 12172 5896
rect 12120 5856 12172 5868
rect 12228 6838 12286 6850
rect 12228 6804 12240 6838
rect 12274 6804 12286 6838
rect 12228 6766 12286 6804
rect 12228 6732 12240 6766
rect 12274 6732 12286 6766
rect 12228 6694 12286 6732
rect 12228 6660 12240 6694
rect 12274 6660 12286 6694
rect 12228 6622 12286 6660
rect 12228 6588 12240 6622
rect 12274 6588 12286 6622
rect 12228 6550 12286 6588
rect 12228 6516 12240 6550
rect 12274 6516 12286 6550
rect 12228 6478 12286 6516
rect 12228 6444 12240 6478
rect 12274 6444 12286 6478
rect 12228 6406 12286 6444
rect 12228 6372 12240 6406
rect 12274 6372 12286 6406
rect 12228 6334 12286 6372
rect 12228 6300 12240 6334
rect 12274 6300 12286 6334
rect 12228 6262 12286 6300
rect 12228 6228 12240 6262
rect 12274 6228 12286 6262
rect 12228 6190 12286 6228
rect 12228 6156 12240 6190
rect 12274 6156 12286 6190
rect 12228 6118 12286 6156
rect 12228 6084 12240 6118
rect 12274 6084 12286 6118
rect 12228 6046 12286 6084
rect 12228 6012 12240 6046
rect 12274 6012 12286 6046
rect 12228 5974 12286 6012
rect 12228 5940 12240 5974
rect 12274 5940 12286 5974
rect 12228 5902 12286 5940
rect 12228 5868 12240 5902
rect 12274 5868 12286 5902
rect 11801 5810 12147 5822
rect 11801 5776 11813 5810
rect 11847 5776 11885 5810
rect 11919 5776 11957 5810
rect 11991 5776 12029 5810
rect 12063 5776 12101 5810
rect 12135 5776 12147 5810
rect 11801 5756 12147 5776
rect 11840 5590 11880 5756
rect 11920 5590 11960 5756
rect 12000 5590 12040 5756
rect 12080 5590 12120 5756
rect 11840 5570 12120 5590
rect 11840 5510 11860 5570
rect 12100 5510 12120 5570
rect 12228 5470 12286 5868
rect 12342 6844 12394 6850
rect 12342 6780 12394 6792
rect 12342 6716 12394 6728
rect 12342 6660 12351 6664
rect 12385 6660 12394 6664
rect 12342 6652 12394 6660
rect 12342 6588 12351 6600
rect 12385 6588 12394 6600
rect 12342 6524 12351 6536
rect 12385 6524 12394 6536
rect 12342 6460 12351 6472
rect 12385 6460 12394 6472
rect 12342 6406 12394 6408
rect 12342 6396 12351 6406
rect 12385 6396 12394 6406
rect 12342 6334 12394 6344
rect 12342 6332 12351 6334
rect 12385 6332 12394 6334
rect 12342 6268 12394 6280
rect 12342 6204 12394 6216
rect 12342 6140 12394 6152
rect 12342 6084 12351 6088
rect 12385 6084 12394 6088
rect 12342 6076 12394 6084
rect 12342 6012 12351 6024
rect 12385 6012 12394 6024
rect 12342 5948 12351 5960
rect 12385 5948 12394 5960
rect 12342 5868 12351 5896
rect 12385 5868 12394 5896
rect 12342 5856 12394 5868
rect 12428 6838 12480 6850
rect 12428 6810 12437 6838
rect 12471 6810 12480 6838
rect 12428 6746 12437 6758
rect 12471 6746 12480 6758
rect 12428 6682 12437 6694
rect 12471 6682 12480 6694
rect 12428 6622 12480 6630
rect 12428 6618 12437 6622
rect 12471 6618 12480 6622
rect 12428 6554 12480 6566
rect 12428 6490 12480 6502
rect 12428 6426 12480 6438
rect 12428 6372 12437 6374
rect 12471 6372 12480 6374
rect 12428 6362 12480 6372
rect 12428 6300 12437 6310
rect 12471 6300 12480 6310
rect 12428 6298 12480 6300
rect 12428 6234 12437 6246
rect 12471 6234 12480 6246
rect 12428 6170 12437 6182
rect 12471 6170 12480 6182
rect 12428 6106 12437 6118
rect 12471 6106 12480 6118
rect 12428 6046 12480 6054
rect 12428 6042 12437 6046
rect 12471 6042 12480 6046
rect 12428 5978 12480 5990
rect 12428 5914 12480 5926
rect 12428 5856 12480 5862
rect 12514 6844 12566 6850
rect 12514 6780 12566 6792
rect 12514 6716 12566 6728
rect 12514 6660 12523 6664
rect 12557 6660 12566 6664
rect 12514 6652 12566 6660
rect 12514 6588 12523 6600
rect 12557 6588 12566 6600
rect 12514 6524 12523 6536
rect 12557 6524 12566 6536
rect 12514 6460 12523 6472
rect 12557 6460 12566 6472
rect 12514 6406 12566 6408
rect 12514 6396 12523 6406
rect 12557 6396 12566 6406
rect 12514 6334 12566 6344
rect 12514 6332 12523 6334
rect 12557 6332 12566 6334
rect 12514 6268 12566 6280
rect 12514 6204 12566 6216
rect 12514 6140 12566 6152
rect 12514 6084 12523 6088
rect 12557 6084 12566 6088
rect 12514 6076 12566 6084
rect 12514 6012 12523 6024
rect 12557 6012 12566 6024
rect 12514 5948 12523 5960
rect 12557 5948 12566 5960
rect 12514 5868 12523 5896
rect 12557 5868 12566 5896
rect 12514 5856 12566 5868
rect 12600 6838 12652 6850
rect 12600 6810 12609 6838
rect 12643 6810 12652 6838
rect 12600 6746 12609 6758
rect 12643 6746 12652 6758
rect 12600 6682 12609 6694
rect 12643 6682 12652 6694
rect 12600 6622 12652 6630
rect 12600 6618 12609 6622
rect 12643 6618 12652 6622
rect 12600 6554 12652 6566
rect 12600 6490 12652 6502
rect 12600 6426 12652 6438
rect 12600 6372 12609 6374
rect 12643 6372 12652 6374
rect 12600 6362 12652 6372
rect 12600 6300 12609 6310
rect 12643 6300 12652 6310
rect 12600 6298 12652 6300
rect 12600 6234 12609 6246
rect 12643 6234 12652 6246
rect 12600 6170 12609 6182
rect 12643 6170 12652 6182
rect 12600 6106 12609 6118
rect 12643 6106 12652 6118
rect 12600 6046 12652 6054
rect 12600 6042 12609 6046
rect 12643 6042 12652 6046
rect 12600 5978 12652 5990
rect 12600 5914 12652 5926
rect 12600 5856 12652 5862
rect 12686 6844 12738 6850
rect 12686 6780 12738 6792
rect 12686 6716 12738 6728
rect 12686 6660 12695 6664
rect 12729 6660 12738 6664
rect 12686 6652 12738 6660
rect 12686 6588 12695 6600
rect 12729 6588 12738 6600
rect 12686 6524 12695 6536
rect 12729 6524 12738 6536
rect 12686 6460 12695 6472
rect 12729 6460 12738 6472
rect 12686 6406 12738 6408
rect 12686 6396 12695 6406
rect 12729 6396 12738 6406
rect 12686 6334 12738 6344
rect 12686 6332 12695 6334
rect 12729 6332 12738 6334
rect 12686 6268 12738 6280
rect 12686 6204 12738 6216
rect 12686 6140 12738 6152
rect 12686 6084 12695 6088
rect 12729 6084 12738 6088
rect 12686 6076 12738 6084
rect 12686 6012 12695 6024
rect 12729 6012 12738 6024
rect 12686 5948 12695 5960
rect 12729 5948 12738 5960
rect 12686 5868 12695 5896
rect 12729 5868 12738 5896
rect 12686 5856 12738 5868
rect 12794 6838 12852 6850
rect 12794 6804 12806 6838
rect 12840 6804 12852 6838
rect 12794 6766 12852 6804
rect 12794 6732 12806 6766
rect 12840 6732 12852 6766
rect 12794 6694 12852 6732
rect 12794 6660 12806 6694
rect 12840 6660 12852 6694
rect 12794 6622 12852 6660
rect 12794 6588 12806 6622
rect 12840 6588 12852 6622
rect 12794 6550 12852 6588
rect 12794 6516 12806 6550
rect 12840 6516 12852 6550
rect 12794 6478 12852 6516
rect 12794 6444 12806 6478
rect 12840 6444 12852 6478
rect 12794 6406 12852 6444
rect 12794 6372 12806 6406
rect 12840 6372 12852 6406
rect 12794 6334 12852 6372
rect 12794 6300 12806 6334
rect 12840 6300 12852 6334
rect 12794 6262 12852 6300
rect 12794 6228 12806 6262
rect 12840 6228 12852 6262
rect 12794 6190 12852 6228
rect 12794 6156 12806 6190
rect 12840 6156 12852 6190
rect 12794 6118 12852 6156
rect 12794 6084 12806 6118
rect 12840 6084 12852 6118
rect 12794 6046 12852 6084
rect 12794 6012 12806 6046
rect 12840 6012 12852 6046
rect 12794 5974 12852 6012
rect 12794 5940 12806 5974
rect 12840 5940 12852 5974
rect 12794 5902 12852 5940
rect 12794 5868 12806 5902
rect 12840 5868 12852 5902
rect 12367 5810 12713 5822
rect 12367 5776 12379 5810
rect 12413 5776 12451 5810
rect 12485 5776 12523 5810
rect 12557 5776 12595 5810
rect 12629 5776 12667 5810
rect 12701 5776 12713 5810
rect 12367 5756 12713 5776
rect 12400 5590 12440 5756
rect 12480 5590 12520 5756
rect 12560 5590 12600 5756
rect 12640 5590 12680 5756
rect 12400 5570 12680 5590
rect 12400 5510 12420 5570
rect 12660 5510 12680 5570
rect 12794 5470 12852 5868
rect 12908 6844 12960 6850
rect 12908 6780 12960 6792
rect 12908 6716 12960 6728
rect 12908 6660 12917 6664
rect 12951 6660 12960 6664
rect 12908 6652 12960 6660
rect 12908 6588 12917 6600
rect 12951 6588 12960 6600
rect 12908 6524 12917 6536
rect 12951 6524 12960 6536
rect 12908 6460 12917 6472
rect 12951 6460 12960 6472
rect 12908 6406 12960 6408
rect 12908 6396 12917 6406
rect 12951 6396 12960 6406
rect 12908 6334 12960 6344
rect 12908 6332 12917 6334
rect 12951 6332 12960 6334
rect 12908 6268 12960 6280
rect 12908 6204 12960 6216
rect 12908 6140 12960 6152
rect 12908 6084 12917 6088
rect 12951 6084 12960 6088
rect 12908 6076 12960 6084
rect 12908 6012 12917 6024
rect 12951 6012 12960 6024
rect 12908 5948 12917 5960
rect 12951 5948 12960 5960
rect 12908 5868 12917 5896
rect 12951 5868 12960 5896
rect 12908 5856 12960 5868
rect 12994 6838 13046 6850
rect 12994 6810 13003 6838
rect 13037 6810 13046 6838
rect 12994 6746 13003 6758
rect 13037 6746 13046 6758
rect 12994 6682 13003 6694
rect 13037 6682 13046 6694
rect 12994 6622 13046 6630
rect 12994 6618 13003 6622
rect 13037 6618 13046 6622
rect 12994 6554 13046 6566
rect 12994 6490 13046 6502
rect 12994 6426 13046 6438
rect 12994 6372 13003 6374
rect 13037 6372 13046 6374
rect 12994 6362 13046 6372
rect 12994 6300 13003 6310
rect 13037 6300 13046 6310
rect 12994 6298 13046 6300
rect 12994 6234 13003 6246
rect 13037 6234 13046 6246
rect 12994 6170 13003 6182
rect 13037 6170 13046 6182
rect 12994 6106 13003 6118
rect 13037 6106 13046 6118
rect 12994 6046 13046 6054
rect 12994 6042 13003 6046
rect 13037 6042 13046 6046
rect 12994 5978 13046 5990
rect 12994 5914 13046 5926
rect 12994 5856 13046 5862
rect 13080 6844 13132 6850
rect 13080 6780 13132 6792
rect 13080 6716 13132 6728
rect 13080 6660 13089 6664
rect 13123 6660 13132 6664
rect 13080 6652 13132 6660
rect 13080 6588 13089 6600
rect 13123 6588 13132 6600
rect 13080 6524 13089 6536
rect 13123 6524 13132 6536
rect 13080 6460 13089 6472
rect 13123 6460 13132 6472
rect 13080 6406 13132 6408
rect 13080 6396 13089 6406
rect 13123 6396 13132 6406
rect 13080 6334 13132 6344
rect 13080 6332 13089 6334
rect 13123 6332 13132 6334
rect 13080 6268 13132 6280
rect 13080 6204 13132 6216
rect 13080 6140 13132 6152
rect 13080 6084 13089 6088
rect 13123 6084 13132 6088
rect 13080 6076 13132 6084
rect 13080 6012 13089 6024
rect 13123 6012 13132 6024
rect 13080 5948 13089 5960
rect 13123 5948 13132 5960
rect 13080 5868 13089 5896
rect 13123 5868 13132 5896
rect 13080 5856 13132 5868
rect 13166 6838 13218 6850
rect 13166 6810 13175 6838
rect 13209 6810 13218 6838
rect 13166 6746 13175 6758
rect 13209 6746 13218 6758
rect 13166 6682 13175 6694
rect 13209 6682 13218 6694
rect 13166 6622 13218 6630
rect 13166 6618 13175 6622
rect 13209 6618 13218 6622
rect 13166 6554 13218 6566
rect 13166 6490 13218 6502
rect 13166 6426 13218 6438
rect 13166 6372 13175 6374
rect 13209 6372 13218 6374
rect 13166 6362 13218 6372
rect 13166 6300 13175 6310
rect 13209 6300 13218 6310
rect 13166 6298 13218 6300
rect 13166 6234 13175 6246
rect 13209 6234 13218 6246
rect 13166 6170 13175 6182
rect 13209 6170 13218 6182
rect 13166 6106 13175 6118
rect 13209 6106 13218 6118
rect 13166 6046 13218 6054
rect 13166 6042 13175 6046
rect 13209 6042 13218 6046
rect 13166 5978 13218 5990
rect 13166 5914 13218 5926
rect 13166 5856 13218 5862
rect 13252 6844 13304 6850
rect 13252 6780 13304 6792
rect 13252 6716 13304 6728
rect 13252 6660 13261 6664
rect 13295 6660 13304 6664
rect 13252 6652 13304 6660
rect 13252 6588 13261 6600
rect 13295 6588 13304 6600
rect 13252 6524 13261 6536
rect 13295 6524 13304 6536
rect 13252 6460 13261 6472
rect 13295 6460 13304 6472
rect 13252 6406 13304 6408
rect 13252 6396 13261 6406
rect 13295 6396 13304 6406
rect 13252 6334 13304 6344
rect 13252 6332 13261 6334
rect 13295 6332 13304 6334
rect 13252 6268 13304 6280
rect 13252 6204 13304 6216
rect 13252 6140 13304 6152
rect 13252 6084 13261 6088
rect 13295 6084 13304 6088
rect 13252 6076 13304 6084
rect 13252 6012 13261 6024
rect 13295 6012 13304 6024
rect 13252 5948 13261 5960
rect 13295 5948 13304 5960
rect 13252 5868 13261 5896
rect 13295 5868 13304 5896
rect 13252 5856 13304 5868
rect 13360 6838 13418 6850
rect 13360 6804 13372 6838
rect 13406 6804 13418 6838
rect 13360 6766 13418 6804
rect 13360 6732 13372 6766
rect 13406 6732 13418 6766
rect 13360 6694 13418 6732
rect 13360 6660 13372 6694
rect 13406 6660 13418 6694
rect 13360 6622 13418 6660
rect 13360 6588 13372 6622
rect 13406 6588 13418 6622
rect 13360 6550 13418 6588
rect 13360 6516 13372 6550
rect 13406 6516 13418 6550
rect 13360 6478 13418 6516
rect 13360 6444 13372 6478
rect 13406 6444 13418 6478
rect 13360 6406 13418 6444
rect 13360 6372 13372 6406
rect 13406 6372 13418 6406
rect 13360 6334 13418 6372
rect 13360 6300 13372 6334
rect 13406 6300 13418 6334
rect 13360 6262 13418 6300
rect 13360 6228 13372 6262
rect 13406 6228 13418 6262
rect 13360 6190 13418 6228
rect 13360 6156 13372 6190
rect 13406 6156 13418 6190
rect 13360 6118 13418 6156
rect 13360 6084 13372 6118
rect 13406 6084 13418 6118
rect 13360 6046 13418 6084
rect 13360 6012 13372 6046
rect 13406 6012 13418 6046
rect 13360 5974 13418 6012
rect 13360 5940 13372 5974
rect 13406 5940 13418 5974
rect 13360 5902 13418 5940
rect 13360 5868 13372 5902
rect 13406 5868 13418 5902
rect 12933 5810 13279 5822
rect 12933 5776 12945 5810
rect 12979 5776 13017 5810
rect 13051 5776 13089 5810
rect 13123 5776 13161 5810
rect 13195 5776 13233 5810
rect 13267 5776 13279 5810
rect 12933 5756 13279 5776
rect 12960 5590 13000 5756
rect 13040 5590 13080 5756
rect 13120 5590 13160 5756
rect 13200 5590 13240 5756
rect 12960 5570 13240 5590
rect 12960 5510 12980 5570
rect 13220 5510 13240 5570
rect 13360 5470 13418 5868
rect 13474 6844 13526 6850
rect 13474 6780 13526 6792
rect 13474 6716 13526 6728
rect 13474 6660 13483 6664
rect 13517 6660 13526 6664
rect 13474 6652 13526 6660
rect 13474 6588 13483 6600
rect 13517 6588 13526 6600
rect 13474 6524 13483 6536
rect 13517 6524 13526 6536
rect 13474 6460 13483 6472
rect 13517 6460 13526 6472
rect 13474 6406 13526 6408
rect 13474 6396 13483 6406
rect 13517 6396 13526 6406
rect 13474 6334 13526 6344
rect 13474 6332 13483 6334
rect 13517 6332 13526 6334
rect 13474 6268 13526 6280
rect 13474 6204 13526 6216
rect 13474 6140 13526 6152
rect 13474 6084 13483 6088
rect 13517 6084 13526 6088
rect 13474 6076 13526 6084
rect 13474 6012 13483 6024
rect 13517 6012 13526 6024
rect 13474 5948 13483 5960
rect 13517 5948 13526 5960
rect 13474 5868 13483 5896
rect 13517 5868 13526 5896
rect 13474 5856 13526 5868
rect 13560 6838 13612 6850
rect 13560 6810 13569 6838
rect 13603 6810 13612 6838
rect 13560 6746 13569 6758
rect 13603 6746 13612 6758
rect 13560 6682 13569 6694
rect 13603 6682 13612 6694
rect 13560 6622 13612 6630
rect 13560 6618 13569 6622
rect 13603 6618 13612 6622
rect 13560 6554 13612 6566
rect 13560 6490 13612 6502
rect 13560 6426 13612 6438
rect 13560 6372 13569 6374
rect 13603 6372 13612 6374
rect 13560 6362 13612 6372
rect 13560 6300 13569 6310
rect 13603 6300 13612 6310
rect 13560 6298 13612 6300
rect 13560 6234 13569 6246
rect 13603 6234 13612 6246
rect 13560 6170 13569 6182
rect 13603 6170 13612 6182
rect 13560 6106 13569 6118
rect 13603 6106 13612 6118
rect 13560 6046 13612 6054
rect 13560 6042 13569 6046
rect 13603 6042 13612 6046
rect 13560 5978 13612 5990
rect 13560 5914 13612 5926
rect 13560 5856 13612 5862
rect 13646 6844 13698 6850
rect 13646 6780 13698 6792
rect 13646 6716 13698 6728
rect 13646 6660 13655 6664
rect 13689 6660 13698 6664
rect 13646 6652 13698 6660
rect 13646 6588 13655 6600
rect 13689 6588 13698 6600
rect 13646 6524 13655 6536
rect 13689 6524 13698 6536
rect 13646 6460 13655 6472
rect 13689 6460 13698 6472
rect 13646 6406 13698 6408
rect 13646 6396 13655 6406
rect 13689 6396 13698 6406
rect 13646 6334 13698 6344
rect 13646 6332 13655 6334
rect 13689 6332 13698 6334
rect 13646 6268 13698 6280
rect 13646 6204 13698 6216
rect 13646 6140 13698 6152
rect 13646 6084 13655 6088
rect 13689 6084 13698 6088
rect 13646 6076 13698 6084
rect 13646 6012 13655 6024
rect 13689 6012 13698 6024
rect 13646 5948 13655 5960
rect 13689 5948 13698 5960
rect 13646 5868 13655 5896
rect 13689 5868 13698 5896
rect 13646 5856 13698 5868
rect 13732 6838 13784 6850
rect 13732 6810 13741 6838
rect 13775 6810 13784 6838
rect 13732 6746 13741 6758
rect 13775 6746 13784 6758
rect 13732 6682 13741 6694
rect 13775 6682 13784 6694
rect 13732 6622 13784 6630
rect 13732 6618 13741 6622
rect 13775 6618 13784 6622
rect 13732 6554 13784 6566
rect 13732 6490 13784 6502
rect 13732 6426 13784 6438
rect 13732 6372 13741 6374
rect 13775 6372 13784 6374
rect 13732 6362 13784 6372
rect 13732 6300 13741 6310
rect 13775 6300 13784 6310
rect 13732 6298 13784 6300
rect 13732 6234 13741 6246
rect 13775 6234 13784 6246
rect 13732 6170 13741 6182
rect 13775 6170 13784 6182
rect 13732 6106 13741 6118
rect 13775 6106 13784 6118
rect 13732 6046 13784 6054
rect 13732 6042 13741 6046
rect 13775 6042 13784 6046
rect 13732 5978 13784 5990
rect 13732 5914 13784 5926
rect 13732 5856 13784 5862
rect 13818 6844 13870 6850
rect 13818 6780 13870 6792
rect 13818 6716 13870 6728
rect 13818 6660 13827 6664
rect 13861 6660 13870 6664
rect 13818 6652 13870 6660
rect 13818 6588 13827 6600
rect 13861 6588 13870 6600
rect 13818 6524 13827 6536
rect 13861 6524 13870 6536
rect 13818 6460 13827 6472
rect 13861 6460 13870 6472
rect 13818 6406 13870 6408
rect 13818 6396 13827 6406
rect 13861 6396 13870 6406
rect 13818 6334 13870 6344
rect 13818 6332 13827 6334
rect 13861 6332 13870 6334
rect 13818 6268 13870 6280
rect 13818 6204 13870 6216
rect 13818 6140 13870 6152
rect 13818 6084 13827 6088
rect 13861 6084 13870 6088
rect 13818 6076 13870 6084
rect 13818 6012 13827 6024
rect 13861 6012 13870 6024
rect 13818 5948 13827 5960
rect 13861 5948 13870 5960
rect 13818 5868 13827 5896
rect 13861 5868 13870 5896
rect 13818 5856 13870 5868
rect 13926 6838 13984 6850
rect 13926 6804 13938 6838
rect 13972 6804 13984 6838
rect 13926 6766 13984 6804
rect 13926 6732 13938 6766
rect 13972 6732 13984 6766
rect 13926 6694 13984 6732
rect 13926 6660 13938 6694
rect 13972 6660 13984 6694
rect 13926 6622 13984 6660
rect 13926 6588 13938 6622
rect 13972 6588 13984 6622
rect 13926 6550 13984 6588
rect 13926 6516 13938 6550
rect 13972 6516 13984 6550
rect 13926 6478 13984 6516
rect 13926 6444 13938 6478
rect 13972 6444 13984 6478
rect 13926 6406 13984 6444
rect 13926 6372 13938 6406
rect 13972 6372 13984 6406
rect 13926 6334 13984 6372
rect 13926 6300 13938 6334
rect 13972 6300 13984 6334
rect 13926 6262 13984 6300
rect 13926 6228 13938 6262
rect 13972 6228 13984 6262
rect 13926 6190 13984 6228
rect 13926 6156 13938 6190
rect 13972 6156 13984 6190
rect 13926 6118 13984 6156
rect 13926 6084 13938 6118
rect 13972 6084 13984 6118
rect 13926 6046 13984 6084
rect 13926 6012 13938 6046
rect 13972 6012 13984 6046
rect 13926 5974 13984 6012
rect 13926 5940 13938 5974
rect 13972 5940 13984 5974
rect 13926 5902 13984 5940
rect 13926 5868 13938 5902
rect 13972 5868 13984 5902
rect 13499 5810 13845 5822
rect 13499 5776 13511 5810
rect 13545 5776 13583 5810
rect 13617 5776 13655 5810
rect 13689 5776 13727 5810
rect 13761 5776 13799 5810
rect 13833 5776 13845 5810
rect 13499 5756 13845 5776
rect 13540 5590 13580 5756
rect 13620 5590 13660 5756
rect 13700 5590 13740 5756
rect 13780 5590 13820 5756
rect 13540 5570 13820 5590
rect 13540 5510 13560 5570
rect 13800 5510 13820 5570
rect 13926 5470 13984 5868
rect 14040 6844 14092 6850
rect 14040 6780 14092 6792
rect 14040 6716 14092 6728
rect 14040 6660 14049 6664
rect 14083 6660 14092 6664
rect 14040 6652 14092 6660
rect 14040 6588 14049 6600
rect 14083 6588 14092 6600
rect 14040 6524 14049 6536
rect 14083 6524 14092 6536
rect 14040 6460 14049 6472
rect 14083 6460 14092 6472
rect 14040 6406 14092 6408
rect 14040 6396 14049 6406
rect 14083 6396 14092 6406
rect 14040 6334 14092 6344
rect 14040 6332 14049 6334
rect 14083 6332 14092 6334
rect 14040 6268 14092 6280
rect 14040 6204 14092 6216
rect 14040 6140 14092 6152
rect 14040 6084 14049 6088
rect 14083 6084 14092 6088
rect 14040 6076 14092 6084
rect 14040 6012 14049 6024
rect 14083 6012 14092 6024
rect 14040 5948 14049 5960
rect 14083 5948 14092 5960
rect 14040 5868 14049 5896
rect 14083 5868 14092 5896
rect 14040 5856 14092 5868
rect 14126 6838 14178 6850
rect 14126 6810 14135 6838
rect 14169 6810 14178 6838
rect 14126 6746 14135 6758
rect 14169 6746 14178 6758
rect 14126 6682 14135 6694
rect 14169 6682 14178 6694
rect 14126 6622 14178 6630
rect 14126 6618 14135 6622
rect 14169 6618 14178 6622
rect 14126 6554 14178 6566
rect 14126 6490 14178 6502
rect 14126 6426 14178 6438
rect 14126 6372 14135 6374
rect 14169 6372 14178 6374
rect 14126 6362 14178 6372
rect 14126 6300 14135 6310
rect 14169 6300 14178 6310
rect 14126 6298 14178 6300
rect 14126 6234 14135 6246
rect 14169 6234 14178 6246
rect 14126 6170 14135 6182
rect 14169 6170 14178 6182
rect 14126 6106 14135 6118
rect 14169 6106 14178 6118
rect 14126 6046 14178 6054
rect 14126 6042 14135 6046
rect 14169 6042 14178 6046
rect 14126 5978 14178 5990
rect 14126 5914 14178 5926
rect 14126 5856 14178 5862
rect 14212 6844 14264 6850
rect 14212 6780 14264 6792
rect 14212 6716 14264 6728
rect 14212 6660 14221 6664
rect 14255 6660 14264 6664
rect 14212 6652 14264 6660
rect 14212 6588 14221 6600
rect 14255 6588 14264 6600
rect 14212 6524 14221 6536
rect 14255 6524 14264 6536
rect 14212 6460 14221 6472
rect 14255 6460 14264 6472
rect 14212 6406 14264 6408
rect 14212 6396 14221 6406
rect 14255 6396 14264 6406
rect 14212 6334 14264 6344
rect 14212 6332 14221 6334
rect 14255 6332 14264 6334
rect 14212 6268 14264 6280
rect 14212 6204 14264 6216
rect 14212 6140 14264 6152
rect 14212 6084 14221 6088
rect 14255 6084 14264 6088
rect 14212 6076 14264 6084
rect 14212 6012 14221 6024
rect 14255 6012 14264 6024
rect 14212 5948 14221 5960
rect 14255 5948 14264 5960
rect 14212 5868 14221 5896
rect 14255 5868 14264 5896
rect 14212 5856 14264 5868
rect 14298 6838 14350 6850
rect 14298 6810 14307 6838
rect 14341 6810 14350 6838
rect 14298 6746 14307 6758
rect 14341 6746 14350 6758
rect 14298 6682 14307 6694
rect 14341 6682 14350 6694
rect 14298 6622 14350 6630
rect 14298 6618 14307 6622
rect 14341 6618 14350 6622
rect 14298 6554 14350 6566
rect 14298 6490 14350 6502
rect 14298 6426 14350 6438
rect 14298 6372 14307 6374
rect 14341 6372 14350 6374
rect 14298 6362 14350 6372
rect 14298 6300 14307 6310
rect 14341 6300 14350 6310
rect 14298 6298 14350 6300
rect 14298 6234 14307 6246
rect 14341 6234 14350 6246
rect 14298 6170 14307 6182
rect 14341 6170 14350 6182
rect 14298 6106 14307 6118
rect 14341 6106 14350 6118
rect 14298 6046 14350 6054
rect 14298 6042 14307 6046
rect 14341 6042 14350 6046
rect 14298 5978 14350 5990
rect 14298 5914 14350 5926
rect 14298 5856 14350 5862
rect 14384 6844 14436 6850
rect 14384 6780 14436 6792
rect 14384 6716 14436 6728
rect 14384 6660 14393 6664
rect 14427 6660 14436 6664
rect 14384 6652 14436 6660
rect 14384 6588 14393 6600
rect 14427 6588 14436 6600
rect 14384 6524 14393 6536
rect 14427 6524 14436 6536
rect 14384 6460 14393 6472
rect 14427 6460 14436 6472
rect 14384 6406 14436 6408
rect 14384 6396 14393 6406
rect 14427 6396 14436 6406
rect 14384 6334 14436 6344
rect 14384 6332 14393 6334
rect 14427 6332 14436 6334
rect 14384 6268 14436 6280
rect 14384 6204 14436 6216
rect 14384 6140 14436 6152
rect 14384 6084 14393 6088
rect 14427 6084 14436 6088
rect 14384 6076 14436 6084
rect 14384 6012 14393 6024
rect 14427 6012 14436 6024
rect 14384 5948 14393 5960
rect 14427 5948 14436 5960
rect 14384 5868 14393 5896
rect 14427 5868 14436 5896
rect 14384 5856 14436 5868
rect 14492 6838 14550 6850
rect 14492 6804 14504 6838
rect 14538 6804 14550 6838
rect 14492 6766 14550 6804
rect 14492 6732 14504 6766
rect 14538 6732 14550 6766
rect 14492 6694 14550 6732
rect 14492 6660 14504 6694
rect 14538 6660 14550 6694
rect 14492 6622 14550 6660
rect 14492 6588 14504 6622
rect 14538 6588 14550 6622
rect 14492 6550 14550 6588
rect 14492 6516 14504 6550
rect 14538 6516 14550 6550
rect 14492 6478 14550 6516
rect 14492 6444 14504 6478
rect 14538 6444 14550 6478
rect 14492 6406 14550 6444
rect 14492 6372 14504 6406
rect 14538 6372 14550 6406
rect 14492 6334 14550 6372
rect 14492 6300 14504 6334
rect 14538 6300 14550 6334
rect 14492 6262 14550 6300
rect 14492 6228 14504 6262
rect 14538 6228 14550 6262
rect 14492 6190 14550 6228
rect 14492 6156 14504 6190
rect 14538 6156 14550 6190
rect 14492 6118 14550 6156
rect 14492 6084 14504 6118
rect 14538 6084 14550 6118
rect 14492 6046 14550 6084
rect 14492 6012 14504 6046
rect 14538 6012 14550 6046
rect 14492 5974 14550 6012
rect 14492 5940 14504 5974
rect 14538 5940 14550 5974
rect 14492 5902 14550 5940
rect 14492 5868 14504 5902
rect 14538 5868 14550 5902
rect 14065 5810 14411 5822
rect 14065 5776 14077 5810
rect 14111 5776 14149 5810
rect 14183 5776 14221 5810
rect 14255 5776 14293 5810
rect 14327 5776 14365 5810
rect 14399 5776 14411 5810
rect 14065 5756 14411 5776
rect 14100 5590 14140 5756
rect 14180 5590 14220 5756
rect 14260 5590 14300 5756
rect 14340 5590 14380 5756
rect 14100 5570 14380 5590
rect 14100 5510 14120 5570
rect 14360 5510 14380 5570
rect 14492 5470 14550 5868
rect 14606 6844 14658 6850
rect 14606 6780 14658 6792
rect 14606 6716 14658 6728
rect 14606 6660 14615 6664
rect 14649 6660 14658 6664
rect 14606 6652 14658 6660
rect 14606 6588 14615 6600
rect 14649 6588 14658 6600
rect 14606 6524 14615 6536
rect 14649 6524 14658 6536
rect 14606 6460 14615 6472
rect 14649 6460 14658 6472
rect 14606 6406 14658 6408
rect 14606 6396 14615 6406
rect 14649 6396 14658 6406
rect 14606 6334 14658 6344
rect 14606 6332 14615 6334
rect 14649 6332 14658 6334
rect 14606 6268 14658 6280
rect 14606 6204 14658 6216
rect 14606 6140 14658 6152
rect 14606 6084 14615 6088
rect 14649 6084 14658 6088
rect 14606 6076 14658 6084
rect 14606 6012 14615 6024
rect 14649 6012 14658 6024
rect 14606 5948 14615 5960
rect 14649 5948 14658 5960
rect 14606 5868 14615 5896
rect 14649 5868 14658 5896
rect 14606 5856 14658 5868
rect 14692 6838 14744 6850
rect 14692 6810 14701 6838
rect 14735 6810 14744 6838
rect 14692 6746 14701 6758
rect 14735 6746 14744 6758
rect 14692 6682 14701 6694
rect 14735 6682 14744 6694
rect 14692 6622 14744 6630
rect 14692 6618 14701 6622
rect 14735 6618 14744 6622
rect 14692 6554 14744 6566
rect 14692 6490 14744 6502
rect 14692 6426 14744 6438
rect 14692 6372 14701 6374
rect 14735 6372 14744 6374
rect 14692 6362 14744 6372
rect 14692 6300 14701 6310
rect 14735 6300 14744 6310
rect 14692 6298 14744 6300
rect 14692 6234 14701 6246
rect 14735 6234 14744 6246
rect 14692 6170 14701 6182
rect 14735 6170 14744 6182
rect 14692 6106 14701 6118
rect 14735 6106 14744 6118
rect 14692 6046 14744 6054
rect 14692 6042 14701 6046
rect 14735 6042 14744 6046
rect 14692 5978 14744 5990
rect 14692 5914 14744 5926
rect 14692 5856 14744 5862
rect 14778 6844 14830 6850
rect 14778 6780 14830 6792
rect 14778 6716 14830 6728
rect 14778 6660 14787 6664
rect 14821 6660 14830 6664
rect 14778 6652 14830 6660
rect 14778 6588 14787 6600
rect 14821 6588 14830 6600
rect 14778 6524 14787 6536
rect 14821 6524 14830 6536
rect 14778 6460 14787 6472
rect 14821 6460 14830 6472
rect 14778 6406 14830 6408
rect 14778 6396 14787 6406
rect 14821 6396 14830 6406
rect 14778 6334 14830 6344
rect 14778 6332 14787 6334
rect 14821 6332 14830 6334
rect 14778 6268 14830 6280
rect 14778 6204 14830 6216
rect 14778 6140 14830 6152
rect 14778 6084 14787 6088
rect 14821 6084 14830 6088
rect 14778 6076 14830 6084
rect 14778 6012 14787 6024
rect 14821 6012 14830 6024
rect 14778 5948 14787 5960
rect 14821 5948 14830 5960
rect 14778 5868 14787 5896
rect 14821 5868 14830 5896
rect 14778 5856 14830 5868
rect 14864 6838 14916 6850
rect 14864 6810 14873 6838
rect 14907 6810 14916 6838
rect 14864 6746 14873 6758
rect 14907 6746 14916 6758
rect 14864 6682 14873 6694
rect 14907 6682 14916 6694
rect 14864 6622 14916 6630
rect 14864 6618 14873 6622
rect 14907 6618 14916 6622
rect 14864 6554 14916 6566
rect 14864 6490 14916 6502
rect 14864 6426 14916 6438
rect 14864 6372 14873 6374
rect 14907 6372 14916 6374
rect 14864 6362 14916 6372
rect 14864 6300 14873 6310
rect 14907 6300 14916 6310
rect 14864 6298 14916 6300
rect 14864 6234 14873 6246
rect 14907 6234 14916 6246
rect 14864 6170 14873 6182
rect 14907 6170 14916 6182
rect 14864 6106 14873 6118
rect 14907 6106 14916 6118
rect 14864 6046 14916 6054
rect 14864 6042 14873 6046
rect 14907 6042 14916 6046
rect 14864 5978 14916 5990
rect 14864 5914 14916 5926
rect 14864 5856 14916 5862
rect 14950 6844 15002 6850
rect 14950 6780 15002 6792
rect 14950 6716 15002 6728
rect 14950 6660 14959 6664
rect 14993 6660 15002 6664
rect 14950 6652 15002 6660
rect 14950 6588 14959 6600
rect 14993 6588 15002 6600
rect 14950 6524 14959 6536
rect 14993 6524 15002 6536
rect 14950 6460 14959 6472
rect 14993 6460 15002 6472
rect 14950 6406 15002 6408
rect 14950 6396 14959 6406
rect 14993 6396 15002 6406
rect 14950 6334 15002 6344
rect 14950 6332 14959 6334
rect 14993 6332 15002 6334
rect 14950 6268 15002 6280
rect 14950 6204 15002 6216
rect 14950 6140 15002 6152
rect 14950 6084 14959 6088
rect 14993 6084 15002 6088
rect 14950 6076 15002 6084
rect 14950 6012 14959 6024
rect 14993 6012 15002 6024
rect 14950 5948 14959 5960
rect 14993 5948 15002 5960
rect 14950 5868 14959 5896
rect 14993 5868 15002 5896
rect 14950 5856 15002 5868
rect 15058 6838 15116 6850
rect 15058 6804 15070 6838
rect 15104 6804 15116 6838
rect 15058 6766 15116 6804
rect 15058 6732 15070 6766
rect 15104 6732 15116 6766
rect 15058 6694 15116 6732
rect 15058 6660 15070 6694
rect 15104 6660 15116 6694
rect 15058 6622 15116 6660
rect 15058 6588 15070 6622
rect 15104 6588 15116 6622
rect 15058 6550 15116 6588
rect 15058 6516 15070 6550
rect 15104 6516 15116 6550
rect 15058 6478 15116 6516
rect 15058 6444 15070 6478
rect 15104 6444 15116 6478
rect 15058 6406 15116 6444
rect 15058 6372 15070 6406
rect 15104 6372 15116 6406
rect 15058 6334 15116 6372
rect 15058 6300 15070 6334
rect 15104 6300 15116 6334
rect 15058 6262 15116 6300
rect 15058 6228 15070 6262
rect 15104 6228 15116 6262
rect 15058 6190 15116 6228
rect 15058 6156 15070 6190
rect 15104 6156 15116 6190
rect 15058 6118 15116 6156
rect 15058 6084 15070 6118
rect 15104 6084 15116 6118
rect 15058 6046 15116 6084
rect 15058 6012 15070 6046
rect 15104 6012 15116 6046
rect 15058 5974 15116 6012
rect 15058 5940 15070 5974
rect 15104 5940 15116 5974
rect 15058 5902 15116 5940
rect 15058 5868 15070 5902
rect 15104 5868 15116 5902
rect 14631 5810 14977 5822
rect 14631 5776 14643 5810
rect 14677 5776 14715 5810
rect 14749 5776 14787 5810
rect 14821 5776 14859 5810
rect 14893 5776 14931 5810
rect 14965 5776 14977 5810
rect 14631 5756 14977 5776
rect 14680 5590 14720 5756
rect 14760 5590 14800 5756
rect 14840 5590 14880 5756
rect 14920 5590 14960 5756
rect 14680 5570 14960 5590
rect 14680 5510 14700 5570
rect 14940 5510 14960 5570
rect 15058 5470 15116 5868
rect 15172 6844 15224 6850
rect 15172 6780 15224 6792
rect 15172 6716 15224 6728
rect 15172 6660 15181 6664
rect 15215 6660 15224 6664
rect 15172 6652 15224 6660
rect 15172 6588 15181 6600
rect 15215 6588 15224 6600
rect 15172 6524 15181 6536
rect 15215 6524 15224 6536
rect 15172 6460 15181 6472
rect 15215 6460 15224 6472
rect 15172 6406 15224 6408
rect 15172 6396 15181 6406
rect 15215 6396 15224 6406
rect 15172 6334 15224 6344
rect 15172 6332 15181 6334
rect 15215 6332 15224 6334
rect 15172 6268 15224 6280
rect 15172 6204 15224 6216
rect 15172 6140 15224 6152
rect 15172 6084 15181 6088
rect 15215 6084 15224 6088
rect 15172 6076 15224 6084
rect 15172 6012 15181 6024
rect 15215 6012 15224 6024
rect 15172 5948 15181 5960
rect 15215 5948 15224 5960
rect 15172 5868 15181 5896
rect 15215 5868 15224 5896
rect 15172 5856 15224 5868
rect 15258 6838 15310 6850
rect 15258 6810 15267 6838
rect 15301 6810 15310 6838
rect 15258 6746 15267 6758
rect 15301 6746 15310 6758
rect 15258 6682 15267 6694
rect 15301 6682 15310 6694
rect 15258 6622 15310 6630
rect 15258 6618 15267 6622
rect 15301 6618 15310 6622
rect 15258 6554 15310 6566
rect 15258 6490 15310 6502
rect 15258 6426 15310 6438
rect 15258 6372 15267 6374
rect 15301 6372 15310 6374
rect 15258 6362 15310 6372
rect 15258 6300 15267 6310
rect 15301 6300 15310 6310
rect 15258 6298 15310 6300
rect 15258 6234 15267 6246
rect 15301 6234 15310 6246
rect 15258 6170 15267 6182
rect 15301 6170 15310 6182
rect 15258 6106 15267 6118
rect 15301 6106 15310 6118
rect 15258 6046 15310 6054
rect 15258 6042 15267 6046
rect 15301 6042 15310 6046
rect 15258 5978 15310 5990
rect 15258 5914 15310 5926
rect 15258 5856 15310 5862
rect 15344 6844 15396 6850
rect 15344 6780 15396 6792
rect 15344 6716 15396 6728
rect 15344 6660 15353 6664
rect 15387 6660 15396 6664
rect 15344 6652 15396 6660
rect 15344 6588 15353 6600
rect 15387 6588 15396 6600
rect 15344 6524 15353 6536
rect 15387 6524 15396 6536
rect 15344 6460 15353 6472
rect 15387 6460 15396 6472
rect 15344 6406 15396 6408
rect 15344 6396 15353 6406
rect 15387 6396 15396 6406
rect 15344 6334 15396 6344
rect 15344 6332 15353 6334
rect 15387 6332 15396 6334
rect 15344 6268 15396 6280
rect 15344 6204 15396 6216
rect 15344 6140 15396 6152
rect 15344 6084 15353 6088
rect 15387 6084 15396 6088
rect 15344 6076 15396 6084
rect 15344 6012 15353 6024
rect 15387 6012 15396 6024
rect 15344 5948 15353 5960
rect 15387 5948 15396 5960
rect 15344 5868 15353 5896
rect 15387 5868 15396 5896
rect 15344 5856 15396 5868
rect 15430 6838 15482 6850
rect 15430 6810 15439 6838
rect 15473 6810 15482 6838
rect 15430 6746 15439 6758
rect 15473 6746 15482 6758
rect 15430 6682 15439 6694
rect 15473 6682 15482 6694
rect 15430 6622 15482 6630
rect 15430 6618 15439 6622
rect 15473 6618 15482 6622
rect 15430 6554 15482 6566
rect 15430 6490 15482 6502
rect 15430 6426 15482 6438
rect 15430 6372 15439 6374
rect 15473 6372 15482 6374
rect 15430 6362 15482 6372
rect 15430 6300 15439 6310
rect 15473 6300 15482 6310
rect 15430 6298 15482 6300
rect 15430 6234 15439 6246
rect 15473 6234 15482 6246
rect 15430 6170 15439 6182
rect 15473 6170 15482 6182
rect 15430 6106 15439 6118
rect 15473 6106 15482 6118
rect 15430 6046 15482 6054
rect 15430 6042 15439 6046
rect 15473 6042 15482 6046
rect 15430 5978 15482 5990
rect 15430 5914 15482 5926
rect 15430 5856 15482 5862
rect 15516 6844 15568 6850
rect 15516 6780 15568 6792
rect 15516 6716 15568 6728
rect 15516 6660 15525 6664
rect 15559 6660 15568 6664
rect 15516 6652 15568 6660
rect 15516 6588 15525 6600
rect 15559 6588 15568 6600
rect 15516 6524 15525 6536
rect 15559 6524 15568 6536
rect 15516 6460 15525 6472
rect 15559 6460 15568 6472
rect 15516 6406 15568 6408
rect 15516 6396 15525 6406
rect 15559 6396 15568 6406
rect 15516 6334 15568 6344
rect 15516 6332 15525 6334
rect 15559 6332 15568 6334
rect 15516 6268 15568 6280
rect 15516 6204 15568 6216
rect 15516 6140 15568 6152
rect 15516 6084 15525 6088
rect 15559 6084 15568 6088
rect 15516 6076 15568 6084
rect 15516 6012 15525 6024
rect 15559 6012 15568 6024
rect 15516 5948 15525 5960
rect 15559 5948 15568 5960
rect 15516 5868 15525 5896
rect 15559 5868 15568 5896
rect 15516 5856 15568 5868
rect 15624 6838 15682 6850
rect 16134 6840 17168 6897
rect 17667 6908 20012 6920
rect 17667 6874 17686 6908
rect 17720 6874 17758 6908
rect 17792 6874 17830 6908
rect 17864 6874 17902 6908
rect 17936 6874 18030 6908
rect 18064 6874 18102 6908
rect 18136 6874 18174 6908
rect 18208 6874 18246 6908
rect 18280 6874 18374 6908
rect 18408 6874 18446 6908
rect 18480 6874 18518 6908
rect 18552 6874 18590 6908
rect 18624 6874 18718 6908
rect 18752 6874 18790 6908
rect 18824 6874 18862 6908
rect 18896 6874 18934 6908
rect 18968 6874 19062 6908
rect 19096 6874 19134 6908
rect 19168 6874 19206 6908
rect 19240 6874 19278 6908
rect 19312 6874 19406 6908
rect 19440 6874 19478 6908
rect 19512 6874 19550 6908
rect 19584 6874 19622 6908
rect 19656 6874 19750 6908
rect 19784 6874 19822 6908
rect 19856 6874 19894 6908
rect 19928 6874 19966 6908
rect 20000 6874 20012 6908
rect 15624 6804 15636 6838
rect 15670 6804 15682 6838
rect 15624 6766 15682 6804
rect 15624 6732 15636 6766
rect 15670 6732 15682 6766
rect 16130 6810 17180 6840
rect 16130 6750 16140 6810
rect 17130 6780 17180 6810
rect 17667 6820 20012 6874
rect 17130 6750 17140 6780
rect 16130 6740 17140 6750
rect 15624 6694 15682 6732
rect 17667 6710 17680 6820
rect 20000 6710 20012 6820
rect 17667 6704 20012 6710
rect 15624 6660 15636 6694
rect 15670 6660 15682 6694
rect 15624 6622 15682 6660
rect 15624 6588 15636 6622
rect 15670 6588 15682 6622
rect 15624 6550 15682 6588
rect 15624 6516 15636 6550
rect 15670 6516 15682 6550
rect 15624 6478 15682 6516
rect 17650 6500 20000 6510
rect 17650 6486 17660 6500
rect 15624 6444 15636 6478
rect 15670 6444 15682 6478
rect 15624 6406 15682 6444
rect 15624 6372 15636 6406
rect 15670 6372 15682 6406
rect 15624 6334 15682 6372
rect 15624 6300 15636 6334
rect 15670 6300 15682 6334
rect 16130 6410 17180 6420
rect 16130 6350 16140 6410
rect 17170 6350 17180 6410
rect 16130 6320 17180 6350
rect 17649 6390 17660 6486
rect 19980 6390 20000 6500
rect 17649 6380 20000 6390
rect 15624 6262 15682 6300
rect 15624 6228 15636 6262
rect 15670 6228 15682 6262
rect 15624 6190 15682 6228
rect 16134 6263 17168 6320
rect 17649 6316 19994 6380
rect 17649 6282 17668 6316
rect 17702 6282 17740 6316
rect 17774 6282 17812 6316
rect 17846 6282 17884 6316
rect 17918 6282 18012 6316
rect 18046 6282 18084 6316
rect 18118 6282 18156 6316
rect 18190 6282 18228 6316
rect 18262 6282 18356 6316
rect 18390 6282 18428 6316
rect 18462 6282 18500 6316
rect 18534 6282 18572 6316
rect 18606 6282 18700 6316
rect 18734 6282 18772 6316
rect 18806 6282 18844 6316
rect 18878 6282 18916 6316
rect 18950 6282 19044 6316
rect 19078 6282 19116 6316
rect 19150 6282 19188 6316
rect 19222 6282 19260 6316
rect 19294 6282 19388 6316
rect 19422 6282 19460 6316
rect 19494 6282 19532 6316
rect 19566 6282 19604 6316
rect 19638 6282 19732 6316
rect 19766 6282 19804 6316
rect 19838 6282 19876 6316
rect 19910 6282 19948 6316
rect 19982 6282 19994 6316
rect 17649 6270 19994 6282
rect 16134 6229 16218 6263
rect 16252 6229 16290 6263
rect 16324 6229 16362 6263
rect 16396 6229 16562 6263
rect 16596 6229 16634 6263
rect 16668 6229 16706 6263
rect 16740 6229 16906 6263
rect 16940 6229 16978 6263
rect 17012 6229 17050 6263
rect 17084 6229 17168 6263
rect 16134 6217 17168 6229
rect 17480 6218 17640 6220
rect 20020 6218 20180 6220
rect 17480 6200 17644 6218
rect 15624 6156 15636 6190
rect 15670 6156 15682 6190
rect 15970 6180 16040 6190
rect 16109 6180 16161 6183
rect 15970 6171 16161 6180
rect 15970 6170 16118 6171
rect 15624 6118 15682 6156
rect 15624 6084 15636 6118
rect 15670 6084 15682 6118
rect 15624 6046 15682 6084
rect 15624 6012 15636 6046
rect 15670 6012 15682 6046
rect 15624 5974 15682 6012
rect 15624 5940 15636 5974
rect 15670 5940 15682 5974
rect 15624 5902 15682 5940
rect 15624 5868 15636 5902
rect 15670 5868 15682 5902
rect 15197 5810 15543 5822
rect 15197 5776 15209 5810
rect 15243 5776 15281 5810
rect 15315 5776 15353 5810
rect 15387 5776 15425 5810
rect 15459 5776 15497 5810
rect 15531 5776 15543 5810
rect 15197 5756 15543 5776
rect 15240 5590 15280 5756
rect 15320 5590 15360 5756
rect 15400 5590 15440 5756
rect 15480 5590 15520 5756
rect 15240 5570 15520 5590
rect 15240 5510 15260 5570
rect 15500 5510 15520 5570
rect 15624 5470 15682 5868
rect 15950 6160 16118 6170
rect 11640 5460 15700 5470
rect 11640 5380 11650 5460
rect 15690 5380 15700 5460
rect 11640 5370 15700 5380
rect 15950 5050 15960 6160
rect 16100 6137 16118 6160
rect 16152 6137 16161 6171
rect 16100 6099 16161 6137
rect 16100 6065 16118 6099
rect 16152 6065 16161 6099
rect 16100 6027 16161 6065
rect 16100 5993 16118 6027
rect 16152 5993 16161 6027
rect 16100 5955 16161 5993
rect 16100 5921 16118 5955
rect 16152 5921 16161 5955
rect 16100 5883 16161 5921
rect 16100 5849 16118 5883
rect 16152 5849 16161 5883
rect 16100 5811 16161 5849
rect 16100 5777 16118 5811
rect 16152 5777 16161 5811
rect 16100 5739 16161 5777
rect 16100 5705 16118 5739
rect 16152 5705 16161 5739
rect 16100 5667 16161 5705
rect 16100 5633 16118 5667
rect 16152 5633 16161 5667
rect 16100 5595 16161 5633
rect 16100 5561 16118 5595
rect 16152 5561 16161 5595
rect 16100 5523 16161 5561
rect 16100 5489 16118 5523
rect 16152 5489 16161 5523
rect 16100 5451 16161 5489
rect 16100 5417 16118 5451
rect 16152 5417 16161 5451
rect 16100 5379 16161 5417
rect 16100 5345 16118 5379
rect 16152 5345 16161 5379
rect 16100 5307 16161 5345
rect 16100 5273 16118 5307
rect 16152 5273 16161 5307
rect 16100 5235 16161 5273
rect 16100 5201 16118 5235
rect 16152 5201 16161 5235
rect 16100 5099 16161 5201
rect 16195 6171 16247 6183
rect 16195 6137 16204 6171
rect 16238 6137 16247 6171
rect 16195 6111 16247 6137
rect 16195 6031 16247 6059
rect 16195 5955 16247 5979
rect 16195 5951 16204 5955
rect 16238 5951 16247 5955
rect 16195 5883 16247 5899
rect 16195 5871 16204 5883
rect 16238 5871 16247 5883
rect 16195 5811 16247 5819
rect 16195 5791 16204 5811
rect 16238 5791 16247 5811
rect 16195 5711 16204 5739
rect 16238 5711 16247 5739
rect 16195 5633 16204 5659
rect 16238 5633 16247 5659
rect 16195 5631 16247 5633
rect 16195 5561 16204 5579
rect 16238 5561 16247 5579
rect 16195 5551 16247 5561
rect 16195 5489 16204 5499
rect 16238 5489 16247 5499
rect 16195 5471 16247 5489
rect 16195 5417 16204 5419
rect 16238 5417 16247 5419
rect 16195 5391 16247 5417
rect 16195 5311 16247 5339
rect 16195 5235 16247 5259
rect 16195 5201 16204 5235
rect 16238 5201 16247 5235
rect 16195 5189 16247 5201
rect 16281 6171 16333 6183
rect 16281 6137 16290 6171
rect 16324 6137 16333 6171
rect 16281 6099 16333 6137
rect 16281 6065 16290 6099
rect 16324 6065 16333 6099
rect 16281 6027 16333 6065
rect 16281 5993 16290 6027
rect 16324 5993 16333 6027
rect 16281 5955 16333 5993
rect 16281 5921 16290 5955
rect 16324 5921 16333 5955
rect 16281 5883 16333 5921
rect 16281 5849 16290 5883
rect 16324 5849 16333 5883
rect 16281 5811 16333 5849
rect 16281 5777 16290 5811
rect 16324 5777 16333 5811
rect 16281 5739 16333 5777
rect 16281 5705 16290 5739
rect 16324 5705 16333 5739
rect 16281 5667 16333 5705
rect 16281 5633 16290 5667
rect 16324 5633 16333 5667
rect 16281 5595 16333 5633
rect 16281 5561 16290 5595
rect 16324 5561 16333 5595
rect 16281 5523 16333 5561
rect 16281 5489 16290 5523
rect 16324 5489 16333 5523
rect 16281 5451 16333 5489
rect 16281 5417 16290 5451
rect 16324 5417 16333 5451
rect 16281 5379 16333 5417
rect 16281 5345 16290 5379
rect 16324 5345 16333 5379
rect 16281 5307 16333 5345
rect 16281 5273 16290 5307
rect 16324 5273 16333 5307
rect 16281 5235 16333 5273
rect 16281 5201 16290 5235
rect 16324 5201 16333 5235
rect 16281 5099 16333 5201
rect 16367 6171 16419 6183
rect 16367 6137 16376 6171
rect 16410 6137 16419 6171
rect 16367 6111 16419 6137
rect 16367 6031 16419 6059
rect 16367 5955 16419 5979
rect 16367 5951 16376 5955
rect 16410 5951 16419 5955
rect 16367 5883 16419 5899
rect 16367 5871 16376 5883
rect 16410 5871 16419 5883
rect 16367 5811 16419 5819
rect 16367 5791 16376 5811
rect 16410 5791 16419 5811
rect 16367 5711 16376 5739
rect 16410 5711 16419 5739
rect 16367 5633 16376 5659
rect 16410 5633 16419 5659
rect 16367 5631 16419 5633
rect 16367 5561 16376 5579
rect 16410 5561 16419 5579
rect 16367 5551 16419 5561
rect 16367 5489 16376 5499
rect 16410 5489 16419 5499
rect 16367 5471 16419 5489
rect 16367 5417 16376 5419
rect 16410 5417 16419 5419
rect 16367 5391 16419 5417
rect 16367 5311 16419 5339
rect 16367 5235 16419 5259
rect 16367 5201 16376 5235
rect 16410 5201 16419 5235
rect 16367 5189 16419 5201
rect 16453 6171 16505 6183
rect 16453 6137 16462 6171
rect 16496 6137 16505 6171
rect 16453 6099 16505 6137
rect 16453 6065 16462 6099
rect 16496 6065 16505 6099
rect 16453 6027 16505 6065
rect 16453 5993 16462 6027
rect 16496 5993 16505 6027
rect 16453 5955 16505 5993
rect 16453 5921 16462 5955
rect 16496 5921 16505 5955
rect 16453 5883 16505 5921
rect 16453 5849 16462 5883
rect 16496 5849 16505 5883
rect 16453 5811 16505 5849
rect 16453 5777 16462 5811
rect 16496 5777 16505 5811
rect 16453 5739 16505 5777
rect 16453 5705 16462 5739
rect 16496 5705 16505 5739
rect 16453 5667 16505 5705
rect 16453 5633 16462 5667
rect 16496 5633 16505 5667
rect 16453 5595 16505 5633
rect 16453 5561 16462 5595
rect 16496 5561 16505 5595
rect 16453 5523 16505 5561
rect 16453 5489 16462 5523
rect 16496 5489 16505 5523
rect 16453 5451 16505 5489
rect 16453 5417 16462 5451
rect 16496 5417 16505 5451
rect 16453 5379 16505 5417
rect 16453 5345 16462 5379
rect 16496 5345 16505 5379
rect 16453 5307 16505 5345
rect 16453 5273 16462 5307
rect 16496 5273 16505 5307
rect 16453 5235 16505 5273
rect 16453 5201 16462 5235
rect 16496 5201 16505 5235
rect 16453 5099 16505 5201
rect 16539 6171 16591 6183
rect 16539 6137 16548 6171
rect 16582 6137 16591 6171
rect 16539 6111 16591 6137
rect 16539 6031 16591 6059
rect 16539 5955 16591 5979
rect 16539 5951 16548 5955
rect 16582 5951 16591 5955
rect 16539 5883 16591 5899
rect 16539 5871 16548 5883
rect 16582 5871 16591 5883
rect 16539 5811 16591 5819
rect 16539 5791 16548 5811
rect 16582 5791 16591 5811
rect 16539 5711 16548 5739
rect 16582 5711 16591 5739
rect 16539 5633 16548 5659
rect 16582 5633 16591 5659
rect 16539 5631 16591 5633
rect 16539 5561 16548 5579
rect 16582 5561 16591 5579
rect 16539 5551 16591 5561
rect 16539 5489 16548 5499
rect 16582 5489 16591 5499
rect 16539 5471 16591 5489
rect 16539 5417 16548 5419
rect 16582 5417 16591 5419
rect 16539 5391 16591 5417
rect 16539 5311 16591 5339
rect 16539 5235 16591 5259
rect 16539 5201 16548 5235
rect 16582 5201 16591 5235
rect 16539 5189 16591 5201
rect 16625 6171 16677 6183
rect 16625 6137 16634 6171
rect 16668 6137 16677 6171
rect 16625 6099 16677 6137
rect 16625 6065 16634 6099
rect 16668 6065 16677 6099
rect 16625 6027 16677 6065
rect 16625 5993 16634 6027
rect 16668 5993 16677 6027
rect 16625 5955 16677 5993
rect 16625 5921 16634 5955
rect 16668 5921 16677 5955
rect 16625 5883 16677 5921
rect 16625 5849 16634 5883
rect 16668 5849 16677 5883
rect 16625 5811 16677 5849
rect 16625 5777 16634 5811
rect 16668 5777 16677 5811
rect 16625 5739 16677 5777
rect 16625 5705 16634 5739
rect 16668 5705 16677 5739
rect 16625 5667 16677 5705
rect 16625 5633 16634 5667
rect 16668 5633 16677 5667
rect 16625 5595 16677 5633
rect 16625 5561 16634 5595
rect 16668 5561 16677 5595
rect 16625 5523 16677 5561
rect 16625 5489 16634 5523
rect 16668 5489 16677 5523
rect 16625 5451 16677 5489
rect 16625 5417 16634 5451
rect 16668 5417 16677 5451
rect 16625 5379 16677 5417
rect 16625 5345 16634 5379
rect 16668 5345 16677 5379
rect 16625 5307 16677 5345
rect 16625 5273 16634 5307
rect 16668 5273 16677 5307
rect 16625 5235 16677 5273
rect 16625 5201 16634 5235
rect 16668 5201 16677 5235
rect 16625 5099 16677 5201
rect 16711 6171 16763 6183
rect 16711 6137 16720 6171
rect 16754 6137 16763 6171
rect 16711 6111 16763 6137
rect 16711 6031 16763 6059
rect 16711 5955 16763 5979
rect 16711 5951 16720 5955
rect 16754 5951 16763 5955
rect 16711 5883 16763 5899
rect 16711 5871 16720 5883
rect 16754 5871 16763 5883
rect 16711 5811 16763 5819
rect 16711 5791 16720 5811
rect 16754 5791 16763 5811
rect 16711 5711 16720 5739
rect 16754 5711 16763 5739
rect 16711 5633 16720 5659
rect 16754 5633 16763 5659
rect 16711 5631 16763 5633
rect 16711 5561 16720 5579
rect 16754 5561 16763 5579
rect 16711 5551 16763 5561
rect 16711 5489 16720 5499
rect 16754 5489 16763 5499
rect 16711 5471 16763 5489
rect 16711 5417 16720 5419
rect 16754 5417 16763 5419
rect 16711 5391 16763 5417
rect 16711 5311 16763 5339
rect 16711 5235 16763 5259
rect 16711 5201 16720 5235
rect 16754 5201 16763 5235
rect 16711 5189 16763 5201
rect 16797 6171 16849 6183
rect 16797 6137 16806 6171
rect 16840 6137 16849 6171
rect 16797 6099 16849 6137
rect 16797 6065 16806 6099
rect 16840 6065 16849 6099
rect 16797 6027 16849 6065
rect 16797 5993 16806 6027
rect 16840 5993 16849 6027
rect 16797 5955 16849 5993
rect 16797 5921 16806 5955
rect 16840 5921 16849 5955
rect 16797 5883 16849 5921
rect 16797 5849 16806 5883
rect 16840 5849 16849 5883
rect 16797 5811 16849 5849
rect 16797 5777 16806 5811
rect 16840 5777 16849 5811
rect 16797 5739 16849 5777
rect 16797 5705 16806 5739
rect 16840 5705 16849 5739
rect 16797 5667 16849 5705
rect 16797 5633 16806 5667
rect 16840 5633 16849 5667
rect 16797 5595 16849 5633
rect 16797 5561 16806 5595
rect 16840 5561 16849 5595
rect 16797 5523 16849 5561
rect 16797 5489 16806 5523
rect 16840 5489 16849 5523
rect 16797 5451 16849 5489
rect 16797 5417 16806 5451
rect 16840 5417 16849 5451
rect 16797 5379 16849 5417
rect 16797 5345 16806 5379
rect 16840 5345 16849 5379
rect 16797 5307 16849 5345
rect 16797 5273 16806 5307
rect 16840 5273 16849 5307
rect 16797 5235 16849 5273
rect 16797 5201 16806 5235
rect 16840 5201 16849 5235
rect 16797 5099 16849 5201
rect 16883 6171 16935 6183
rect 16883 6137 16892 6171
rect 16926 6137 16935 6171
rect 16883 6111 16935 6137
rect 16883 6031 16935 6059
rect 16883 5955 16935 5979
rect 16883 5951 16892 5955
rect 16926 5951 16935 5955
rect 16883 5883 16935 5899
rect 16883 5871 16892 5883
rect 16926 5871 16935 5883
rect 16883 5811 16935 5819
rect 16883 5791 16892 5811
rect 16926 5791 16935 5811
rect 16883 5711 16892 5739
rect 16926 5711 16935 5739
rect 16883 5633 16892 5659
rect 16926 5633 16935 5659
rect 16883 5631 16935 5633
rect 16883 5561 16892 5579
rect 16926 5561 16935 5579
rect 16883 5551 16935 5561
rect 16883 5489 16892 5499
rect 16926 5489 16935 5499
rect 16883 5471 16935 5489
rect 16883 5417 16892 5419
rect 16926 5417 16935 5419
rect 16883 5391 16935 5417
rect 16883 5311 16935 5339
rect 16883 5235 16935 5259
rect 16883 5201 16892 5235
rect 16926 5201 16935 5235
rect 16883 5189 16935 5201
rect 16969 6171 17021 6183
rect 16969 6137 16978 6171
rect 17012 6137 17021 6171
rect 16969 6099 17021 6137
rect 16969 6065 16978 6099
rect 17012 6065 17021 6099
rect 16969 6027 17021 6065
rect 16969 5993 16978 6027
rect 17012 5993 17021 6027
rect 16969 5955 17021 5993
rect 16969 5921 16978 5955
rect 17012 5921 17021 5955
rect 16969 5883 17021 5921
rect 16969 5849 16978 5883
rect 17012 5849 17021 5883
rect 16969 5811 17021 5849
rect 16969 5777 16978 5811
rect 17012 5777 17021 5811
rect 16969 5739 17021 5777
rect 16969 5705 16978 5739
rect 17012 5705 17021 5739
rect 16969 5667 17021 5705
rect 16969 5633 16978 5667
rect 17012 5633 17021 5667
rect 16969 5595 17021 5633
rect 16969 5561 16978 5595
rect 17012 5561 17021 5595
rect 16969 5523 17021 5561
rect 16969 5489 16978 5523
rect 17012 5489 17021 5523
rect 16969 5451 17021 5489
rect 16969 5417 16978 5451
rect 17012 5417 17021 5451
rect 16969 5379 17021 5417
rect 16969 5345 16978 5379
rect 17012 5345 17021 5379
rect 16969 5307 17021 5345
rect 16969 5273 16978 5307
rect 17012 5273 17021 5307
rect 16969 5235 17021 5273
rect 16969 5201 16978 5235
rect 17012 5201 17021 5235
rect 16969 5099 17021 5201
rect 17055 6171 17107 6183
rect 17055 6137 17064 6171
rect 17098 6137 17107 6171
rect 17055 6111 17107 6137
rect 17055 6031 17107 6059
rect 17055 5955 17107 5979
rect 17055 5951 17064 5955
rect 17098 5951 17107 5955
rect 17055 5883 17107 5899
rect 17055 5871 17064 5883
rect 17098 5871 17107 5883
rect 17055 5811 17107 5819
rect 17055 5791 17064 5811
rect 17098 5791 17107 5811
rect 17055 5711 17064 5739
rect 17098 5711 17107 5739
rect 17055 5633 17064 5659
rect 17098 5633 17107 5659
rect 17055 5631 17107 5633
rect 17055 5561 17064 5579
rect 17098 5561 17107 5579
rect 17055 5551 17107 5561
rect 17055 5489 17064 5499
rect 17098 5489 17107 5499
rect 17055 5471 17107 5489
rect 17055 5417 17064 5419
rect 17098 5417 17107 5419
rect 17055 5391 17107 5417
rect 17055 5311 17107 5339
rect 17055 5235 17107 5259
rect 17055 5201 17064 5235
rect 17098 5201 17107 5235
rect 17055 5189 17107 5201
rect 17141 6180 17193 6183
rect 17260 6180 17330 6190
rect 17141 6171 17330 6180
rect 17141 6137 17150 6171
rect 17184 6154 17330 6171
rect 17184 6137 17280 6154
rect 17141 6120 17280 6137
rect 17314 6120 17330 6154
rect 17141 6099 17330 6120
rect 17141 6065 17150 6099
rect 17184 6074 17330 6099
rect 17184 6065 17280 6074
rect 17141 6040 17280 6065
rect 17314 6040 17330 6074
rect 17141 6027 17330 6040
rect 17141 5993 17150 6027
rect 17184 5994 17330 6027
rect 17184 5993 17280 5994
rect 17141 5960 17280 5993
rect 17314 5960 17330 5994
rect 17141 5955 17330 5960
rect 17141 5921 17150 5955
rect 17184 5921 17330 5955
rect 17141 5914 17330 5921
rect 17141 5883 17280 5914
rect 17141 5849 17150 5883
rect 17184 5880 17280 5883
rect 17314 5880 17330 5914
rect 17184 5849 17330 5880
rect 17141 5834 17330 5849
rect 17141 5811 17280 5834
rect 17141 5777 17150 5811
rect 17184 5800 17280 5811
rect 17314 5800 17330 5834
rect 17184 5777 17330 5800
rect 17141 5754 17330 5777
rect 17141 5739 17280 5754
rect 17141 5705 17150 5739
rect 17184 5720 17280 5739
rect 17314 5720 17330 5754
rect 17184 5705 17330 5720
rect 17141 5674 17330 5705
rect 17141 5667 17280 5674
rect 17141 5633 17150 5667
rect 17184 5640 17280 5667
rect 17314 5640 17330 5674
rect 17184 5633 17330 5640
rect 17141 5595 17330 5633
rect 17141 5561 17150 5595
rect 17184 5594 17330 5595
rect 17184 5561 17280 5594
rect 17141 5560 17280 5561
rect 17314 5560 17330 5594
rect 17141 5523 17330 5560
rect 17141 5489 17150 5523
rect 17184 5514 17330 5523
rect 17184 5489 17280 5514
rect 17141 5480 17280 5489
rect 17314 5480 17330 5514
rect 17141 5451 17330 5480
rect 17141 5417 17150 5451
rect 17184 5434 17330 5451
rect 17184 5417 17280 5434
rect 17141 5400 17280 5417
rect 17314 5400 17330 5434
rect 17141 5379 17330 5400
rect 17141 5345 17150 5379
rect 17184 5354 17330 5379
rect 17184 5345 17280 5354
rect 17141 5320 17280 5345
rect 17314 5320 17330 5354
rect 17141 5307 17330 5320
rect 17141 5273 17150 5307
rect 17184 5274 17330 5307
rect 17184 5273 17280 5274
rect 17141 5240 17280 5273
rect 17314 5240 17330 5274
rect 17480 5260 17500 6200
rect 17540 6180 17644 6200
rect 17540 6146 17604 6180
rect 17638 6146 17644 6180
rect 17540 6108 17644 6146
rect 17540 6074 17604 6108
rect 17638 6074 17644 6108
rect 17540 6036 17644 6074
rect 17540 6002 17604 6036
rect 17638 6002 17644 6036
rect 17540 5964 17644 6002
rect 17540 5930 17604 5964
rect 17638 5930 17644 5964
rect 17540 5892 17644 5930
rect 17540 5858 17604 5892
rect 17638 5858 17644 5892
rect 17540 5820 17644 5858
rect 17540 5786 17604 5820
rect 17638 5786 17644 5820
rect 17540 5748 17644 5786
rect 17540 5714 17604 5748
rect 17638 5714 17644 5748
rect 17540 5676 17644 5714
rect 17540 5642 17604 5676
rect 17638 5642 17644 5676
rect 17540 5604 17644 5642
rect 17540 5570 17604 5604
rect 17638 5570 17644 5604
rect 17540 5532 17644 5570
rect 17540 5498 17604 5532
rect 17638 5498 17644 5532
rect 17540 5460 17644 5498
rect 17540 5426 17604 5460
rect 17638 5426 17644 5460
rect 17540 5388 17644 5426
rect 17540 5354 17604 5388
rect 17638 5354 17644 5388
rect 17540 5316 17644 5354
rect 17540 5282 17604 5316
rect 17638 5282 17644 5316
rect 17540 5260 17644 5282
rect 17480 5240 17644 5260
rect 17681 6207 17733 6218
rect 17681 6146 17690 6155
rect 17724 6146 17733 6155
rect 17681 6143 17733 6146
rect 17681 6074 17690 6091
rect 17724 6074 17733 6091
rect 17681 6036 17733 6074
rect 17681 6002 17690 6036
rect 17724 6002 17733 6036
rect 17681 5964 17733 6002
rect 17681 5930 17690 5964
rect 17724 5930 17733 5964
rect 17681 5892 17733 5930
rect 17681 5858 17690 5892
rect 17724 5858 17733 5892
rect 17681 5820 17733 5858
rect 17681 5786 17690 5820
rect 17724 5786 17733 5820
rect 17681 5748 17733 5786
rect 17681 5714 17690 5748
rect 17724 5714 17733 5748
rect 17681 5676 17733 5714
rect 17681 5642 17690 5676
rect 17724 5642 17733 5676
rect 17681 5604 17733 5642
rect 17681 5570 17690 5604
rect 17724 5570 17733 5604
rect 17681 5532 17733 5570
rect 17681 5498 17690 5532
rect 17724 5498 17733 5532
rect 17681 5460 17733 5498
rect 17681 5426 17690 5460
rect 17724 5426 17733 5460
rect 17681 5388 17733 5426
rect 17681 5354 17690 5388
rect 17724 5354 17733 5388
rect 17681 5316 17733 5354
rect 17681 5282 17690 5316
rect 17724 5282 17733 5316
rect 17681 5248 17733 5282
rect 17770 6180 17816 6218
rect 17770 6146 17776 6180
rect 17810 6146 17816 6180
rect 17770 6108 17816 6146
rect 17770 6074 17776 6108
rect 17810 6074 17816 6108
rect 17770 6036 17816 6074
rect 17770 6002 17776 6036
rect 17810 6002 17816 6036
rect 17770 5964 17816 6002
rect 17770 5930 17776 5964
rect 17810 5930 17816 5964
rect 17770 5892 17816 5930
rect 17770 5858 17776 5892
rect 17810 5858 17816 5892
rect 17770 5820 17816 5858
rect 17770 5786 17776 5820
rect 17810 5786 17816 5820
rect 17770 5748 17816 5786
rect 17770 5714 17776 5748
rect 17810 5714 17816 5748
rect 17770 5676 17816 5714
rect 17770 5642 17776 5676
rect 17810 5642 17816 5676
rect 17770 5604 17816 5642
rect 17770 5570 17776 5604
rect 17810 5570 17816 5604
rect 17770 5532 17816 5570
rect 17770 5498 17776 5532
rect 17810 5498 17816 5532
rect 17770 5460 17816 5498
rect 17770 5426 17776 5460
rect 17810 5426 17816 5460
rect 17770 5388 17816 5426
rect 17770 5354 17776 5388
rect 17810 5354 17816 5388
rect 17770 5316 17816 5354
rect 17770 5282 17776 5316
rect 17810 5282 17816 5316
rect 17141 5235 17330 5240
rect 17141 5201 17150 5235
rect 17184 5201 17330 5235
rect 17141 5194 17330 5201
rect 17141 5160 17280 5194
rect 17314 5160 17330 5194
rect 17141 5099 17330 5160
rect 17598 5152 17644 5240
rect 17770 5152 17816 5282
rect 17853 6207 17905 6218
rect 17853 6146 17862 6155
rect 17896 6146 17905 6155
rect 17853 6143 17905 6146
rect 17853 6074 17862 6091
rect 17896 6074 17905 6091
rect 17853 6036 17905 6074
rect 17853 6002 17862 6036
rect 17896 6002 17905 6036
rect 17853 5964 17905 6002
rect 17853 5930 17862 5964
rect 17896 5930 17905 5964
rect 17853 5892 17905 5930
rect 17853 5858 17862 5892
rect 17896 5858 17905 5892
rect 17853 5820 17905 5858
rect 17853 5786 17862 5820
rect 17896 5786 17905 5820
rect 17853 5748 17905 5786
rect 17853 5714 17862 5748
rect 17896 5714 17905 5748
rect 17853 5676 17905 5714
rect 17853 5642 17862 5676
rect 17896 5642 17905 5676
rect 17853 5604 17905 5642
rect 17853 5570 17862 5604
rect 17896 5570 17905 5604
rect 17853 5532 17905 5570
rect 17853 5498 17862 5532
rect 17896 5498 17905 5532
rect 17853 5460 17905 5498
rect 17853 5426 17862 5460
rect 17896 5426 17905 5460
rect 17853 5388 17905 5426
rect 17853 5354 17862 5388
rect 17896 5354 17905 5388
rect 17853 5316 17905 5354
rect 17853 5282 17862 5316
rect 17896 5282 17905 5316
rect 17853 5248 17905 5282
rect 17942 6180 17988 6218
rect 17942 6146 17948 6180
rect 17982 6146 17988 6180
rect 17942 6108 17988 6146
rect 17942 6074 17948 6108
rect 17982 6074 17988 6108
rect 17942 6036 17988 6074
rect 17942 6002 17948 6036
rect 17982 6002 17988 6036
rect 17942 5964 17988 6002
rect 17942 5930 17948 5964
rect 17982 5930 17988 5964
rect 17942 5892 17988 5930
rect 17942 5858 17948 5892
rect 17982 5858 17988 5892
rect 17942 5820 17988 5858
rect 17942 5786 17948 5820
rect 17982 5786 17988 5820
rect 17942 5748 17988 5786
rect 17942 5714 17948 5748
rect 17982 5714 17988 5748
rect 17942 5676 17988 5714
rect 17942 5642 17948 5676
rect 17982 5642 17988 5676
rect 17942 5604 17988 5642
rect 17942 5570 17948 5604
rect 17982 5570 17988 5604
rect 17942 5532 17988 5570
rect 17942 5498 17948 5532
rect 17982 5498 17988 5532
rect 17942 5460 17988 5498
rect 17942 5426 17948 5460
rect 17982 5426 17988 5460
rect 17942 5388 17988 5426
rect 17942 5354 17948 5388
rect 17982 5354 17988 5388
rect 17942 5316 17988 5354
rect 17942 5282 17948 5316
rect 17982 5282 17988 5316
rect 17942 5152 17988 5282
rect 18025 6207 18077 6218
rect 18025 6146 18034 6155
rect 18068 6146 18077 6155
rect 18025 6143 18077 6146
rect 18025 6074 18034 6091
rect 18068 6074 18077 6091
rect 18025 6036 18077 6074
rect 18025 6002 18034 6036
rect 18068 6002 18077 6036
rect 18025 5964 18077 6002
rect 18025 5930 18034 5964
rect 18068 5930 18077 5964
rect 18025 5892 18077 5930
rect 18025 5858 18034 5892
rect 18068 5858 18077 5892
rect 18025 5820 18077 5858
rect 18025 5786 18034 5820
rect 18068 5786 18077 5820
rect 18025 5748 18077 5786
rect 18025 5714 18034 5748
rect 18068 5714 18077 5748
rect 18025 5676 18077 5714
rect 18025 5642 18034 5676
rect 18068 5642 18077 5676
rect 18025 5604 18077 5642
rect 18025 5570 18034 5604
rect 18068 5570 18077 5604
rect 18025 5532 18077 5570
rect 18025 5498 18034 5532
rect 18068 5498 18077 5532
rect 18025 5460 18077 5498
rect 18025 5426 18034 5460
rect 18068 5426 18077 5460
rect 18025 5388 18077 5426
rect 18025 5354 18034 5388
rect 18068 5354 18077 5388
rect 18025 5316 18077 5354
rect 18025 5282 18034 5316
rect 18068 5282 18077 5316
rect 18025 5248 18077 5282
rect 18114 6180 18160 6218
rect 18114 6146 18120 6180
rect 18154 6146 18160 6180
rect 18114 6108 18160 6146
rect 18114 6074 18120 6108
rect 18154 6074 18160 6108
rect 18114 6036 18160 6074
rect 18114 6002 18120 6036
rect 18154 6002 18160 6036
rect 18114 5964 18160 6002
rect 18114 5930 18120 5964
rect 18154 5930 18160 5964
rect 18114 5892 18160 5930
rect 18114 5858 18120 5892
rect 18154 5858 18160 5892
rect 18114 5820 18160 5858
rect 18114 5786 18120 5820
rect 18154 5786 18160 5820
rect 18114 5748 18160 5786
rect 18114 5714 18120 5748
rect 18154 5714 18160 5748
rect 18114 5676 18160 5714
rect 18114 5642 18120 5676
rect 18154 5642 18160 5676
rect 18114 5604 18160 5642
rect 18114 5570 18120 5604
rect 18154 5570 18160 5604
rect 18114 5532 18160 5570
rect 18114 5498 18120 5532
rect 18154 5498 18160 5532
rect 18114 5460 18160 5498
rect 18114 5426 18120 5460
rect 18154 5426 18160 5460
rect 18114 5388 18160 5426
rect 18114 5354 18120 5388
rect 18154 5354 18160 5388
rect 18114 5316 18160 5354
rect 18114 5282 18120 5316
rect 18154 5282 18160 5316
rect 18114 5152 18160 5282
rect 18197 6207 18249 6218
rect 18197 6146 18206 6155
rect 18240 6146 18249 6155
rect 18197 6143 18249 6146
rect 18197 6074 18206 6091
rect 18240 6074 18249 6091
rect 18197 6036 18249 6074
rect 18197 6002 18206 6036
rect 18240 6002 18249 6036
rect 18197 5964 18249 6002
rect 18197 5930 18206 5964
rect 18240 5930 18249 5964
rect 18197 5892 18249 5930
rect 18197 5858 18206 5892
rect 18240 5858 18249 5892
rect 18197 5820 18249 5858
rect 18197 5786 18206 5820
rect 18240 5786 18249 5820
rect 18197 5748 18249 5786
rect 18197 5714 18206 5748
rect 18240 5714 18249 5748
rect 18197 5676 18249 5714
rect 18197 5642 18206 5676
rect 18240 5642 18249 5676
rect 18197 5604 18249 5642
rect 18197 5570 18206 5604
rect 18240 5570 18249 5604
rect 18197 5532 18249 5570
rect 18197 5498 18206 5532
rect 18240 5498 18249 5532
rect 18197 5460 18249 5498
rect 18197 5426 18206 5460
rect 18240 5426 18249 5460
rect 18197 5388 18249 5426
rect 18197 5354 18206 5388
rect 18240 5354 18249 5388
rect 18197 5316 18249 5354
rect 18197 5282 18206 5316
rect 18240 5282 18249 5316
rect 18197 5248 18249 5282
rect 18286 6180 18332 6218
rect 18286 6146 18292 6180
rect 18326 6146 18332 6180
rect 18286 6108 18332 6146
rect 18286 6074 18292 6108
rect 18326 6074 18332 6108
rect 18286 6036 18332 6074
rect 18286 6002 18292 6036
rect 18326 6002 18332 6036
rect 18286 5964 18332 6002
rect 18286 5930 18292 5964
rect 18326 5930 18332 5964
rect 18286 5892 18332 5930
rect 18286 5858 18292 5892
rect 18326 5858 18332 5892
rect 18286 5820 18332 5858
rect 18286 5786 18292 5820
rect 18326 5786 18332 5820
rect 18286 5748 18332 5786
rect 18286 5714 18292 5748
rect 18326 5714 18332 5748
rect 18286 5676 18332 5714
rect 18286 5642 18292 5676
rect 18326 5642 18332 5676
rect 18286 5604 18332 5642
rect 18286 5570 18292 5604
rect 18326 5570 18332 5604
rect 18286 5532 18332 5570
rect 18286 5498 18292 5532
rect 18326 5498 18332 5532
rect 18286 5460 18332 5498
rect 18286 5426 18292 5460
rect 18326 5426 18332 5460
rect 18286 5388 18332 5426
rect 18286 5354 18292 5388
rect 18326 5354 18332 5388
rect 18286 5316 18332 5354
rect 18286 5282 18292 5316
rect 18326 5282 18332 5316
rect 18286 5152 18332 5282
rect 18369 6207 18421 6218
rect 18369 6146 18378 6155
rect 18412 6146 18421 6155
rect 18369 6143 18421 6146
rect 18369 6074 18378 6091
rect 18412 6074 18421 6091
rect 18369 6036 18421 6074
rect 18369 6002 18378 6036
rect 18412 6002 18421 6036
rect 18369 5964 18421 6002
rect 18369 5930 18378 5964
rect 18412 5930 18421 5964
rect 18369 5892 18421 5930
rect 18369 5858 18378 5892
rect 18412 5858 18421 5892
rect 18369 5820 18421 5858
rect 18369 5786 18378 5820
rect 18412 5786 18421 5820
rect 18369 5748 18421 5786
rect 18369 5714 18378 5748
rect 18412 5714 18421 5748
rect 18369 5676 18421 5714
rect 18369 5642 18378 5676
rect 18412 5642 18421 5676
rect 18369 5604 18421 5642
rect 18369 5570 18378 5604
rect 18412 5570 18421 5604
rect 18369 5532 18421 5570
rect 18369 5498 18378 5532
rect 18412 5498 18421 5532
rect 18369 5460 18421 5498
rect 18369 5426 18378 5460
rect 18412 5426 18421 5460
rect 18369 5388 18421 5426
rect 18369 5354 18378 5388
rect 18412 5354 18421 5388
rect 18369 5316 18421 5354
rect 18369 5282 18378 5316
rect 18412 5282 18421 5316
rect 18369 5248 18421 5282
rect 18458 6180 18504 6218
rect 18458 6146 18464 6180
rect 18498 6146 18504 6180
rect 18458 6108 18504 6146
rect 18458 6074 18464 6108
rect 18498 6074 18504 6108
rect 18458 6036 18504 6074
rect 18458 6002 18464 6036
rect 18498 6002 18504 6036
rect 18458 5964 18504 6002
rect 18458 5930 18464 5964
rect 18498 5930 18504 5964
rect 18458 5892 18504 5930
rect 18458 5858 18464 5892
rect 18498 5858 18504 5892
rect 18458 5820 18504 5858
rect 18458 5786 18464 5820
rect 18498 5786 18504 5820
rect 18458 5748 18504 5786
rect 18458 5714 18464 5748
rect 18498 5714 18504 5748
rect 18458 5676 18504 5714
rect 18458 5642 18464 5676
rect 18498 5642 18504 5676
rect 18458 5604 18504 5642
rect 18458 5570 18464 5604
rect 18498 5570 18504 5604
rect 18458 5532 18504 5570
rect 18458 5498 18464 5532
rect 18498 5498 18504 5532
rect 18458 5460 18504 5498
rect 18458 5426 18464 5460
rect 18498 5426 18504 5460
rect 18458 5388 18504 5426
rect 18458 5354 18464 5388
rect 18498 5354 18504 5388
rect 18458 5316 18504 5354
rect 18458 5282 18464 5316
rect 18498 5282 18504 5316
rect 18458 5152 18504 5282
rect 18541 6207 18593 6218
rect 18541 6146 18550 6155
rect 18584 6146 18593 6155
rect 18541 6143 18593 6146
rect 18541 6074 18550 6091
rect 18584 6074 18593 6091
rect 18541 6036 18593 6074
rect 18541 6002 18550 6036
rect 18584 6002 18593 6036
rect 18541 5964 18593 6002
rect 18541 5930 18550 5964
rect 18584 5930 18593 5964
rect 18541 5892 18593 5930
rect 18541 5858 18550 5892
rect 18584 5858 18593 5892
rect 18541 5820 18593 5858
rect 18541 5786 18550 5820
rect 18584 5786 18593 5820
rect 18541 5748 18593 5786
rect 18541 5714 18550 5748
rect 18584 5714 18593 5748
rect 18541 5676 18593 5714
rect 18541 5642 18550 5676
rect 18584 5642 18593 5676
rect 18541 5604 18593 5642
rect 18541 5570 18550 5604
rect 18584 5570 18593 5604
rect 18541 5532 18593 5570
rect 18541 5498 18550 5532
rect 18584 5498 18593 5532
rect 18541 5460 18593 5498
rect 18541 5426 18550 5460
rect 18584 5426 18593 5460
rect 18541 5388 18593 5426
rect 18541 5354 18550 5388
rect 18584 5354 18593 5388
rect 18541 5316 18593 5354
rect 18541 5282 18550 5316
rect 18584 5282 18593 5316
rect 18541 5248 18593 5282
rect 18630 6180 18676 6218
rect 18630 6146 18636 6180
rect 18670 6146 18676 6180
rect 18630 6108 18676 6146
rect 18630 6074 18636 6108
rect 18670 6074 18676 6108
rect 18630 6036 18676 6074
rect 18630 6002 18636 6036
rect 18670 6002 18676 6036
rect 18630 5964 18676 6002
rect 18630 5930 18636 5964
rect 18670 5930 18676 5964
rect 18630 5892 18676 5930
rect 18630 5858 18636 5892
rect 18670 5858 18676 5892
rect 18630 5820 18676 5858
rect 18630 5786 18636 5820
rect 18670 5786 18676 5820
rect 18630 5748 18676 5786
rect 18630 5714 18636 5748
rect 18670 5714 18676 5748
rect 18630 5676 18676 5714
rect 18630 5642 18636 5676
rect 18670 5642 18676 5676
rect 18630 5604 18676 5642
rect 18630 5570 18636 5604
rect 18670 5570 18676 5604
rect 18630 5532 18676 5570
rect 18630 5498 18636 5532
rect 18670 5498 18676 5532
rect 18630 5460 18676 5498
rect 18630 5426 18636 5460
rect 18670 5426 18676 5460
rect 18630 5388 18676 5426
rect 18630 5354 18636 5388
rect 18670 5354 18676 5388
rect 18630 5316 18676 5354
rect 18630 5282 18636 5316
rect 18670 5282 18676 5316
rect 18630 5152 18676 5282
rect 18713 6207 18765 6218
rect 18713 6146 18722 6155
rect 18756 6146 18765 6155
rect 18713 6143 18765 6146
rect 18713 6074 18722 6091
rect 18756 6074 18765 6091
rect 18713 6036 18765 6074
rect 18713 6002 18722 6036
rect 18756 6002 18765 6036
rect 18713 5964 18765 6002
rect 18713 5930 18722 5964
rect 18756 5930 18765 5964
rect 18713 5892 18765 5930
rect 18713 5858 18722 5892
rect 18756 5858 18765 5892
rect 18713 5820 18765 5858
rect 18713 5786 18722 5820
rect 18756 5786 18765 5820
rect 18713 5748 18765 5786
rect 18713 5714 18722 5748
rect 18756 5714 18765 5748
rect 18713 5676 18765 5714
rect 18713 5642 18722 5676
rect 18756 5642 18765 5676
rect 18713 5604 18765 5642
rect 18713 5570 18722 5604
rect 18756 5570 18765 5604
rect 18713 5532 18765 5570
rect 18713 5498 18722 5532
rect 18756 5498 18765 5532
rect 18713 5460 18765 5498
rect 18713 5426 18722 5460
rect 18756 5426 18765 5460
rect 18713 5388 18765 5426
rect 18713 5354 18722 5388
rect 18756 5354 18765 5388
rect 18713 5316 18765 5354
rect 18713 5282 18722 5316
rect 18756 5282 18765 5316
rect 18713 5248 18765 5282
rect 18802 6180 18848 6218
rect 18802 6146 18808 6180
rect 18842 6146 18848 6180
rect 18802 6108 18848 6146
rect 18802 6074 18808 6108
rect 18842 6074 18848 6108
rect 18802 6036 18848 6074
rect 18802 6002 18808 6036
rect 18842 6002 18848 6036
rect 18802 5964 18848 6002
rect 18802 5930 18808 5964
rect 18842 5930 18848 5964
rect 18802 5892 18848 5930
rect 18802 5858 18808 5892
rect 18842 5858 18848 5892
rect 18802 5820 18848 5858
rect 18802 5786 18808 5820
rect 18842 5786 18848 5820
rect 18802 5748 18848 5786
rect 18802 5714 18808 5748
rect 18842 5714 18848 5748
rect 18802 5676 18848 5714
rect 18802 5642 18808 5676
rect 18842 5642 18848 5676
rect 18802 5604 18848 5642
rect 18802 5570 18808 5604
rect 18842 5570 18848 5604
rect 18802 5532 18848 5570
rect 18802 5498 18808 5532
rect 18842 5498 18848 5532
rect 18802 5460 18848 5498
rect 18802 5426 18808 5460
rect 18842 5426 18848 5460
rect 18802 5388 18848 5426
rect 18802 5354 18808 5388
rect 18842 5354 18848 5388
rect 18802 5316 18848 5354
rect 18802 5282 18808 5316
rect 18842 5282 18848 5316
rect 18802 5152 18848 5282
rect 18885 6207 18937 6218
rect 18885 6146 18894 6155
rect 18928 6146 18937 6155
rect 18885 6143 18937 6146
rect 18885 6074 18894 6091
rect 18928 6074 18937 6091
rect 18885 6036 18937 6074
rect 18885 6002 18894 6036
rect 18928 6002 18937 6036
rect 18885 5964 18937 6002
rect 18885 5930 18894 5964
rect 18928 5930 18937 5964
rect 18885 5892 18937 5930
rect 18885 5858 18894 5892
rect 18928 5858 18937 5892
rect 18885 5820 18937 5858
rect 18885 5786 18894 5820
rect 18928 5786 18937 5820
rect 18885 5748 18937 5786
rect 18885 5714 18894 5748
rect 18928 5714 18937 5748
rect 18885 5676 18937 5714
rect 18885 5642 18894 5676
rect 18928 5642 18937 5676
rect 18885 5604 18937 5642
rect 18885 5570 18894 5604
rect 18928 5570 18937 5604
rect 18885 5532 18937 5570
rect 18885 5498 18894 5532
rect 18928 5498 18937 5532
rect 18885 5460 18937 5498
rect 18885 5426 18894 5460
rect 18928 5426 18937 5460
rect 18885 5388 18937 5426
rect 18885 5354 18894 5388
rect 18928 5354 18937 5388
rect 18885 5316 18937 5354
rect 18885 5282 18894 5316
rect 18928 5282 18937 5316
rect 18885 5248 18937 5282
rect 18974 6180 19020 6218
rect 18974 6146 18980 6180
rect 19014 6146 19020 6180
rect 18974 6108 19020 6146
rect 18974 6074 18980 6108
rect 19014 6074 19020 6108
rect 18974 6036 19020 6074
rect 18974 6002 18980 6036
rect 19014 6002 19020 6036
rect 18974 5964 19020 6002
rect 18974 5930 18980 5964
rect 19014 5930 19020 5964
rect 18974 5892 19020 5930
rect 18974 5858 18980 5892
rect 19014 5858 19020 5892
rect 18974 5820 19020 5858
rect 18974 5786 18980 5820
rect 19014 5786 19020 5820
rect 18974 5748 19020 5786
rect 18974 5714 18980 5748
rect 19014 5714 19020 5748
rect 18974 5676 19020 5714
rect 18974 5642 18980 5676
rect 19014 5642 19020 5676
rect 18974 5604 19020 5642
rect 18974 5570 18980 5604
rect 19014 5570 19020 5604
rect 18974 5532 19020 5570
rect 18974 5498 18980 5532
rect 19014 5498 19020 5532
rect 18974 5460 19020 5498
rect 18974 5426 18980 5460
rect 19014 5426 19020 5460
rect 18974 5388 19020 5426
rect 18974 5354 18980 5388
rect 19014 5354 19020 5388
rect 18974 5316 19020 5354
rect 18974 5282 18980 5316
rect 19014 5282 19020 5316
rect 18974 5152 19020 5282
rect 19057 6207 19109 6218
rect 19057 6146 19066 6155
rect 19100 6146 19109 6155
rect 19057 6143 19109 6146
rect 19057 6074 19066 6091
rect 19100 6074 19109 6091
rect 19057 6036 19109 6074
rect 19057 6002 19066 6036
rect 19100 6002 19109 6036
rect 19057 5964 19109 6002
rect 19057 5930 19066 5964
rect 19100 5930 19109 5964
rect 19057 5892 19109 5930
rect 19057 5858 19066 5892
rect 19100 5858 19109 5892
rect 19057 5820 19109 5858
rect 19057 5786 19066 5820
rect 19100 5786 19109 5820
rect 19057 5748 19109 5786
rect 19057 5714 19066 5748
rect 19100 5714 19109 5748
rect 19057 5676 19109 5714
rect 19057 5642 19066 5676
rect 19100 5642 19109 5676
rect 19057 5604 19109 5642
rect 19057 5570 19066 5604
rect 19100 5570 19109 5604
rect 19057 5532 19109 5570
rect 19057 5498 19066 5532
rect 19100 5498 19109 5532
rect 19057 5460 19109 5498
rect 19057 5426 19066 5460
rect 19100 5426 19109 5460
rect 19057 5388 19109 5426
rect 19057 5354 19066 5388
rect 19100 5354 19109 5388
rect 19057 5316 19109 5354
rect 19057 5282 19066 5316
rect 19100 5282 19109 5316
rect 19057 5248 19109 5282
rect 19146 6180 19192 6218
rect 19146 6146 19152 6180
rect 19186 6146 19192 6180
rect 19146 6108 19192 6146
rect 19146 6074 19152 6108
rect 19186 6074 19192 6108
rect 19146 6036 19192 6074
rect 19146 6002 19152 6036
rect 19186 6002 19192 6036
rect 19146 5964 19192 6002
rect 19146 5930 19152 5964
rect 19186 5930 19192 5964
rect 19146 5892 19192 5930
rect 19146 5858 19152 5892
rect 19186 5858 19192 5892
rect 19146 5820 19192 5858
rect 19146 5786 19152 5820
rect 19186 5786 19192 5820
rect 19146 5748 19192 5786
rect 19146 5714 19152 5748
rect 19186 5714 19192 5748
rect 19146 5676 19192 5714
rect 19146 5642 19152 5676
rect 19186 5642 19192 5676
rect 19146 5604 19192 5642
rect 19146 5570 19152 5604
rect 19186 5570 19192 5604
rect 19146 5532 19192 5570
rect 19146 5498 19152 5532
rect 19186 5498 19192 5532
rect 19146 5460 19192 5498
rect 19146 5426 19152 5460
rect 19186 5426 19192 5460
rect 19146 5388 19192 5426
rect 19146 5354 19152 5388
rect 19186 5354 19192 5388
rect 19146 5316 19192 5354
rect 19146 5282 19152 5316
rect 19186 5282 19192 5316
rect 19146 5152 19192 5282
rect 19229 6207 19281 6218
rect 19229 6146 19238 6155
rect 19272 6146 19281 6155
rect 19229 6143 19281 6146
rect 19229 6074 19238 6091
rect 19272 6074 19281 6091
rect 19229 6036 19281 6074
rect 19229 6002 19238 6036
rect 19272 6002 19281 6036
rect 19229 5964 19281 6002
rect 19229 5930 19238 5964
rect 19272 5930 19281 5964
rect 19229 5892 19281 5930
rect 19229 5858 19238 5892
rect 19272 5858 19281 5892
rect 19229 5820 19281 5858
rect 19229 5786 19238 5820
rect 19272 5786 19281 5820
rect 19229 5748 19281 5786
rect 19229 5714 19238 5748
rect 19272 5714 19281 5748
rect 19229 5676 19281 5714
rect 19229 5642 19238 5676
rect 19272 5642 19281 5676
rect 19229 5604 19281 5642
rect 19229 5570 19238 5604
rect 19272 5570 19281 5604
rect 19229 5532 19281 5570
rect 19229 5498 19238 5532
rect 19272 5498 19281 5532
rect 19229 5460 19281 5498
rect 19229 5426 19238 5460
rect 19272 5426 19281 5460
rect 19229 5388 19281 5426
rect 19229 5354 19238 5388
rect 19272 5354 19281 5388
rect 19229 5316 19281 5354
rect 19229 5282 19238 5316
rect 19272 5282 19281 5316
rect 19229 5248 19281 5282
rect 19318 6180 19364 6218
rect 19318 6146 19324 6180
rect 19358 6146 19364 6180
rect 19318 6108 19364 6146
rect 19318 6074 19324 6108
rect 19358 6074 19364 6108
rect 19318 6036 19364 6074
rect 19318 6002 19324 6036
rect 19358 6002 19364 6036
rect 19318 5964 19364 6002
rect 19318 5930 19324 5964
rect 19358 5930 19364 5964
rect 19318 5892 19364 5930
rect 19318 5858 19324 5892
rect 19358 5858 19364 5892
rect 19318 5820 19364 5858
rect 19318 5786 19324 5820
rect 19358 5786 19364 5820
rect 19318 5748 19364 5786
rect 19318 5714 19324 5748
rect 19358 5714 19364 5748
rect 19318 5676 19364 5714
rect 19318 5642 19324 5676
rect 19358 5642 19364 5676
rect 19318 5604 19364 5642
rect 19318 5570 19324 5604
rect 19358 5570 19364 5604
rect 19318 5532 19364 5570
rect 19318 5498 19324 5532
rect 19358 5498 19364 5532
rect 19318 5460 19364 5498
rect 19318 5426 19324 5460
rect 19358 5426 19364 5460
rect 19318 5388 19364 5426
rect 19318 5354 19324 5388
rect 19358 5354 19364 5388
rect 19318 5316 19364 5354
rect 19318 5282 19324 5316
rect 19358 5282 19364 5316
rect 19318 5152 19364 5282
rect 19401 6207 19453 6218
rect 19401 6146 19410 6155
rect 19444 6146 19453 6155
rect 19401 6143 19453 6146
rect 19401 6074 19410 6091
rect 19444 6074 19453 6091
rect 19401 6036 19453 6074
rect 19401 6002 19410 6036
rect 19444 6002 19453 6036
rect 19401 5964 19453 6002
rect 19401 5930 19410 5964
rect 19444 5930 19453 5964
rect 19401 5892 19453 5930
rect 19401 5858 19410 5892
rect 19444 5858 19453 5892
rect 19401 5820 19453 5858
rect 19401 5786 19410 5820
rect 19444 5786 19453 5820
rect 19401 5748 19453 5786
rect 19401 5714 19410 5748
rect 19444 5714 19453 5748
rect 19401 5676 19453 5714
rect 19401 5642 19410 5676
rect 19444 5642 19453 5676
rect 19401 5604 19453 5642
rect 19401 5570 19410 5604
rect 19444 5570 19453 5604
rect 19401 5532 19453 5570
rect 19401 5498 19410 5532
rect 19444 5498 19453 5532
rect 19401 5460 19453 5498
rect 19401 5426 19410 5460
rect 19444 5426 19453 5460
rect 19401 5388 19453 5426
rect 19401 5354 19410 5388
rect 19444 5354 19453 5388
rect 19401 5316 19453 5354
rect 19401 5282 19410 5316
rect 19444 5282 19453 5316
rect 19401 5248 19453 5282
rect 19490 6180 19536 6218
rect 19490 6146 19496 6180
rect 19530 6146 19536 6180
rect 19490 6108 19536 6146
rect 19490 6074 19496 6108
rect 19530 6074 19536 6108
rect 19490 6036 19536 6074
rect 19490 6002 19496 6036
rect 19530 6002 19536 6036
rect 19490 5964 19536 6002
rect 19490 5930 19496 5964
rect 19530 5930 19536 5964
rect 19490 5892 19536 5930
rect 19490 5858 19496 5892
rect 19530 5858 19536 5892
rect 19490 5820 19536 5858
rect 19490 5786 19496 5820
rect 19530 5786 19536 5820
rect 19490 5748 19536 5786
rect 19490 5714 19496 5748
rect 19530 5714 19536 5748
rect 19490 5676 19536 5714
rect 19490 5642 19496 5676
rect 19530 5642 19536 5676
rect 19490 5604 19536 5642
rect 19490 5570 19496 5604
rect 19530 5570 19536 5604
rect 19490 5532 19536 5570
rect 19490 5498 19496 5532
rect 19530 5498 19536 5532
rect 19490 5460 19536 5498
rect 19490 5426 19496 5460
rect 19530 5426 19536 5460
rect 19490 5388 19536 5426
rect 19490 5354 19496 5388
rect 19530 5354 19536 5388
rect 19490 5316 19536 5354
rect 19490 5282 19496 5316
rect 19530 5282 19536 5316
rect 19490 5152 19536 5282
rect 19573 6207 19625 6218
rect 19573 6146 19582 6155
rect 19616 6146 19625 6155
rect 19573 6143 19625 6146
rect 19573 6074 19582 6091
rect 19616 6074 19625 6091
rect 19573 6036 19625 6074
rect 19573 6002 19582 6036
rect 19616 6002 19625 6036
rect 19573 5964 19625 6002
rect 19573 5930 19582 5964
rect 19616 5930 19625 5964
rect 19573 5892 19625 5930
rect 19573 5858 19582 5892
rect 19616 5858 19625 5892
rect 19573 5820 19625 5858
rect 19573 5786 19582 5820
rect 19616 5786 19625 5820
rect 19573 5748 19625 5786
rect 19573 5714 19582 5748
rect 19616 5714 19625 5748
rect 19573 5676 19625 5714
rect 19573 5642 19582 5676
rect 19616 5642 19625 5676
rect 19573 5604 19625 5642
rect 19573 5570 19582 5604
rect 19616 5570 19625 5604
rect 19573 5532 19625 5570
rect 19573 5498 19582 5532
rect 19616 5498 19625 5532
rect 19573 5460 19625 5498
rect 19573 5426 19582 5460
rect 19616 5426 19625 5460
rect 19573 5388 19625 5426
rect 19573 5354 19582 5388
rect 19616 5354 19625 5388
rect 19573 5316 19625 5354
rect 19573 5282 19582 5316
rect 19616 5282 19625 5316
rect 19573 5248 19625 5282
rect 19662 6180 19708 6218
rect 19662 6146 19668 6180
rect 19702 6146 19708 6180
rect 19662 6108 19708 6146
rect 19662 6074 19668 6108
rect 19702 6074 19708 6108
rect 19662 6036 19708 6074
rect 19662 6002 19668 6036
rect 19702 6002 19708 6036
rect 19662 5964 19708 6002
rect 19662 5930 19668 5964
rect 19702 5930 19708 5964
rect 19662 5892 19708 5930
rect 19662 5858 19668 5892
rect 19702 5858 19708 5892
rect 19662 5820 19708 5858
rect 19662 5786 19668 5820
rect 19702 5786 19708 5820
rect 19662 5748 19708 5786
rect 19662 5714 19668 5748
rect 19702 5714 19708 5748
rect 19662 5676 19708 5714
rect 19662 5642 19668 5676
rect 19702 5642 19708 5676
rect 19662 5604 19708 5642
rect 19662 5570 19668 5604
rect 19702 5570 19708 5604
rect 19662 5532 19708 5570
rect 19662 5498 19668 5532
rect 19702 5498 19708 5532
rect 19662 5460 19708 5498
rect 19662 5426 19668 5460
rect 19702 5426 19708 5460
rect 19662 5388 19708 5426
rect 19662 5354 19668 5388
rect 19702 5354 19708 5388
rect 19662 5316 19708 5354
rect 19662 5282 19668 5316
rect 19702 5282 19708 5316
rect 19662 5152 19708 5282
rect 19745 6207 19797 6218
rect 19745 6146 19754 6155
rect 19788 6146 19797 6155
rect 19745 6143 19797 6146
rect 19745 6074 19754 6091
rect 19788 6074 19797 6091
rect 19745 6036 19797 6074
rect 19745 6002 19754 6036
rect 19788 6002 19797 6036
rect 19745 5964 19797 6002
rect 19745 5930 19754 5964
rect 19788 5930 19797 5964
rect 19745 5892 19797 5930
rect 19745 5858 19754 5892
rect 19788 5858 19797 5892
rect 19745 5820 19797 5858
rect 19745 5786 19754 5820
rect 19788 5786 19797 5820
rect 19745 5748 19797 5786
rect 19745 5714 19754 5748
rect 19788 5714 19797 5748
rect 19745 5676 19797 5714
rect 19745 5642 19754 5676
rect 19788 5642 19797 5676
rect 19745 5604 19797 5642
rect 19745 5570 19754 5604
rect 19788 5570 19797 5604
rect 19745 5532 19797 5570
rect 19745 5498 19754 5532
rect 19788 5498 19797 5532
rect 19745 5460 19797 5498
rect 19745 5426 19754 5460
rect 19788 5426 19797 5460
rect 19745 5388 19797 5426
rect 19745 5354 19754 5388
rect 19788 5354 19797 5388
rect 19745 5316 19797 5354
rect 19745 5282 19754 5316
rect 19788 5282 19797 5316
rect 19745 5248 19797 5282
rect 19834 6180 19880 6218
rect 19834 6146 19840 6180
rect 19874 6146 19880 6180
rect 19834 6108 19880 6146
rect 19834 6074 19840 6108
rect 19874 6074 19880 6108
rect 19834 6036 19880 6074
rect 19834 6002 19840 6036
rect 19874 6002 19880 6036
rect 19834 5964 19880 6002
rect 19834 5930 19840 5964
rect 19874 5930 19880 5964
rect 19834 5892 19880 5930
rect 19834 5858 19840 5892
rect 19874 5858 19880 5892
rect 19834 5820 19880 5858
rect 19834 5786 19840 5820
rect 19874 5786 19880 5820
rect 19834 5748 19880 5786
rect 19834 5714 19840 5748
rect 19874 5714 19880 5748
rect 19834 5676 19880 5714
rect 19834 5642 19840 5676
rect 19874 5642 19880 5676
rect 19834 5604 19880 5642
rect 19834 5570 19840 5604
rect 19874 5570 19880 5604
rect 19834 5532 19880 5570
rect 19834 5498 19840 5532
rect 19874 5498 19880 5532
rect 19834 5460 19880 5498
rect 19834 5426 19840 5460
rect 19874 5426 19880 5460
rect 19834 5388 19880 5426
rect 19834 5354 19840 5388
rect 19874 5354 19880 5388
rect 19834 5316 19880 5354
rect 19834 5282 19840 5316
rect 19874 5282 19880 5316
rect 19834 5152 19880 5282
rect 19917 6207 19969 6218
rect 19917 6146 19926 6155
rect 19960 6146 19969 6155
rect 19917 6143 19969 6146
rect 19917 6074 19926 6091
rect 19960 6074 19969 6091
rect 19917 6036 19969 6074
rect 19917 6002 19926 6036
rect 19960 6002 19969 6036
rect 19917 5964 19969 6002
rect 19917 5930 19926 5964
rect 19960 5930 19969 5964
rect 19917 5892 19969 5930
rect 19917 5858 19926 5892
rect 19960 5858 19969 5892
rect 19917 5820 19969 5858
rect 19917 5786 19926 5820
rect 19960 5786 19969 5820
rect 19917 5748 19969 5786
rect 19917 5714 19926 5748
rect 19960 5714 19969 5748
rect 19917 5676 19969 5714
rect 19917 5642 19926 5676
rect 19960 5642 19969 5676
rect 19917 5604 19969 5642
rect 19917 5570 19926 5604
rect 19960 5570 19969 5604
rect 19917 5532 19969 5570
rect 19917 5498 19926 5532
rect 19960 5498 19969 5532
rect 19917 5460 19969 5498
rect 19917 5426 19926 5460
rect 19960 5426 19969 5460
rect 19917 5388 19969 5426
rect 19917 5354 19926 5388
rect 19960 5354 19969 5388
rect 19917 5316 19969 5354
rect 19917 5282 19926 5316
rect 19960 5282 19969 5316
rect 19917 5248 19969 5282
rect 20006 6200 20180 6218
rect 20006 6190 20120 6200
rect 20160 6190 20180 6200
rect 20006 6180 20060 6190
rect 20006 6146 20012 6180
rect 20046 6146 20060 6180
rect 20006 6108 20060 6146
rect 20006 6074 20012 6108
rect 20046 6074 20060 6108
rect 20006 6036 20060 6074
rect 20006 6002 20012 6036
rect 20046 6002 20060 6036
rect 20006 5964 20060 6002
rect 20006 5930 20012 5964
rect 20046 5930 20060 5964
rect 20006 5892 20060 5930
rect 20006 5858 20012 5892
rect 20046 5858 20060 5892
rect 20006 5820 20060 5858
rect 20006 5786 20012 5820
rect 20046 5786 20060 5820
rect 20006 5748 20060 5786
rect 20006 5714 20012 5748
rect 20046 5714 20060 5748
rect 20006 5676 20060 5714
rect 20006 5642 20012 5676
rect 20046 5642 20060 5676
rect 20006 5604 20060 5642
rect 20006 5570 20012 5604
rect 20046 5570 20060 5604
rect 20006 5532 20060 5570
rect 20006 5498 20012 5532
rect 20046 5498 20060 5532
rect 20006 5460 20060 5498
rect 20006 5426 20012 5460
rect 20046 5426 20060 5460
rect 20006 5388 20060 5426
rect 20006 5354 20012 5388
rect 20046 5354 20060 5388
rect 20006 5316 20060 5354
rect 20006 5282 20012 5316
rect 20046 5282 20060 5316
rect 20006 5260 20060 5282
rect 20006 5240 20180 5260
rect 20006 5152 20052 5240
rect 17598 5140 20052 5152
rect 16100 5084 17330 5099
rect 16114 5050 16160 5084
rect 16194 5050 16240 5084
rect 16274 5050 16320 5084
rect 16354 5050 16400 5084
rect 16434 5050 16480 5084
rect 16514 5050 16560 5084
rect 16594 5050 16640 5084
rect 16674 5050 16720 5084
rect 16754 5050 16800 5084
rect 16834 5050 16880 5084
rect 16914 5050 16960 5084
rect 16994 5050 17040 5084
rect 17074 5050 17120 5084
rect 17154 5050 17330 5084
rect 15950 5040 17330 5050
rect 15970 5030 17330 5040
rect 17380 5100 17620 5140
rect 20040 5100 20230 5140
rect 15980 5010 16100 5030
rect 16550 4818 17319 5030
rect 17380 5000 17420 5100
rect 20140 5000 20230 5100
rect 17380 4960 20230 5000
rect 16550 4811 20116 4818
rect 16550 4802 16638 4811
rect 16550 4768 16635 4802
rect 16550 4765 16638 4768
rect 16550 4713 16557 4765
rect 16609 4759 16638 4765
rect 16690 4759 16702 4811
rect 16754 4759 16766 4811
rect 16818 4759 16830 4811
rect 16882 4802 16894 4811
rect 16946 4802 16958 4811
rect 17010 4802 17022 4811
rect 17074 4802 17086 4811
rect 17138 4802 17150 4811
rect 17202 4802 17214 4811
rect 16885 4768 16894 4802
rect 16957 4768 16958 4802
rect 17138 4768 17139 4802
rect 17202 4768 17211 4802
rect 16882 4759 16894 4768
rect 16946 4759 16958 4768
rect 17010 4759 17022 4768
rect 17074 4759 17086 4768
rect 17138 4759 17150 4768
rect 17202 4759 17214 4768
rect 17266 4759 17278 4811
rect 17330 4802 17492 4811
rect 17330 4768 17355 4802
rect 17389 4768 17427 4802
rect 17461 4768 17492 4802
rect 17330 4759 17492 4768
rect 17544 4759 17556 4811
rect 17608 4759 17620 4811
rect 17672 4802 17684 4811
rect 17736 4802 17748 4811
rect 17800 4802 17812 4811
rect 17864 4802 17876 4811
rect 17928 4802 17940 4811
rect 17992 4802 18004 4811
rect 17677 4768 17684 4802
rect 17928 4768 17931 4802
rect 17992 4768 18003 4802
rect 17672 4759 17684 4768
rect 17736 4759 17748 4768
rect 17800 4759 17812 4768
rect 17864 4759 17876 4768
rect 17928 4759 17940 4768
rect 17992 4759 18004 4768
rect 18056 4759 18068 4811
rect 18120 4759 18132 4811
rect 18184 4802 18488 4811
rect 18184 4768 18485 4802
rect 18184 4765 18488 4768
rect 18184 4759 18207 4765
rect 16609 4752 18207 4759
rect 16609 4713 16616 4752
rect 16550 4701 16566 4713
rect 16600 4701 16616 4713
rect 16550 4649 16557 4701
rect 16609 4649 16616 4701
rect 16550 4637 16566 4649
rect 16600 4637 16616 4649
rect 16550 4585 16557 4637
rect 16609 4585 16616 4637
rect 16550 4573 16566 4585
rect 16600 4573 16616 4585
rect 16550 4521 16557 4573
rect 16609 4521 16616 4573
rect 16550 4519 16616 4521
rect 16550 4509 16566 4519
rect 16600 4509 16616 4519
rect 16550 4457 16557 4509
rect 16609 4457 16616 4509
rect 16550 4447 16616 4457
rect 16550 4445 16566 4447
rect 16600 4445 16616 4447
rect 16550 4393 16557 4445
rect 16609 4393 16616 4445
rect 16550 4381 16616 4393
rect 16550 4329 16557 4381
rect 16609 4329 16616 4381
rect 16550 4317 16616 4329
rect 16550 4265 16557 4317
rect 16609 4265 16616 4317
rect 16550 4253 16616 4265
rect 16550 4201 16557 4253
rect 16609 4201 16616 4253
rect 16550 4197 16566 4201
rect 16600 4197 16616 4201
rect 16550 4189 16616 4197
rect 16550 4137 16557 4189
rect 16609 4137 16616 4189
rect 16550 4125 16566 4137
rect 16600 4125 16616 4137
rect 16550 4087 16616 4125
rect 16550 4053 16566 4087
rect 16600 4053 16616 4087
rect 16550 4015 16616 4053
rect 16550 3981 16566 4015
rect 16600 3981 16616 4015
rect 16550 3943 16616 3981
rect 16550 3931 16566 3943
rect 16600 3931 16616 3943
rect 16550 3879 16557 3931
rect 16609 3879 16616 3931
rect 16550 3871 16616 3879
rect 16550 3867 16566 3871
rect 16600 3867 16616 3871
rect 16550 3815 16557 3867
rect 16609 3815 16616 3867
rect 16550 3803 16616 3815
rect 16550 3751 16557 3803
rect 16609 3751 16616 3803
rect 16550 3739 16616 3751
rect 16550 3687 16557 3739
rect 16609 3687 16616 3739
rect 16550 3675 16616 3687
rect 16550 3623 16557 3675
rect 16609 3623 16616 3675
rect 16550 3621 16566 3623
rect 16600 3621 16616 3623
rect 16550 3611 16616 3621
rect 16550 3559 16557 3611
rect 16609 3559 16616 3611
rect 16550 3549 16566 3559
rect 16600 3549 16616 3559
rect 16550 3547 16616 3549
rect 16550 3495 16557 3547
rect 16609 3495 16616 3547
rect 16550 3483 16566 3495
rect 16600 3483 16616 3495
rect 16550 3431 16557 3483
rect 16609 3431 16616 3483
rect 16550 3419 16566 3431
rect 16600 3419 16616 3431
rect 16550 3367 16557 3419
rect 16609 3367 16616 3419
rect 16550 3355 16566 3367
rect 16600 3355 16616 3367
rect 16550 3303 16557 3355
rect 16609 3316 16616 3355
rect 16649 4066 16677 4724
rect 16705 4094 16733 4752
rect 16761 4066 16789 4724
rect 16817 4094 16845 4752
rect 16873 4066 16901 4724
rect 16929 4094 16957 4752
rect 16985 4066 17013 4724
rect 17041 4094 17069 4752
rect 17097 4066 17125 4724
rect 17153 4094 17181 4752
rect 17209 4066 17237 4724
rect 17265 4094 17293 4752
rect 17321 4066 17349 4724
rect 17381 4718 17435 4724
rect 17381 4666 17382 4718
rect 17434 4666 17435 4718
rect 17381 4654 17435 4666
rect 17381 4602 17382 4654
rect 17434 4602 17435 4654
rect 17381 4590 17435 4602
rect 17381 4538 17382 4590
rect 17434 4538 17435 4590
rect 17381 4526 17435 4538
rect 17381 4474 17382 4526
rect 17434 4474 17435 4526
rect 17381 4462 17435 4474
rect 17381 4410 17382 4462
rect 17434 4410 17435 4462
rect 17381 4398 17435 4410
rect 17381 4346 17382 4398
rect 17434 4346 17435 4398
rect 17381 4334 17435 4346
rect 17381 4282 17382 4334
rect 17434 4282 17435 4334
rect 17381 4270 17435 4282
rect 17381 4218 17382 4270
rect 17434 4218 17435 4270
rect 17381 4206 17435 4218
rect 17381 4154 17382 4206
rect 17434 4154 17435 4206
rect 17381 4142 17435 4154
rect 17381 4090 17382 4142
rect 17434 4090 17435 4142
rect 17381 4066 17435 4090
rect 17467 4066 17495 4724
rect 17523 4094 17551 4752
rect 17579 4066 17607 4724
rect 17635 4094 17663 4752
rect 17691 4066 17719 4724
rect 17747 4094 17775 4752
rect 17803 4066 17831 4724
rect 17859 4094 17887 4752
rect 17915 4066 17943 4724
rect 17971 4094 17999 4752
rect 18027 4066 18055 4724
rect 18083 4094 18111 4752
rect 18139 4066 18167 4724
rect 16649 4060 18167 4066
rect 16649 4008 16655 4060
rect 16707 4008 16719 4060
rect 16771 4008 16783 4060
rect 16835 4008 16847 4060
rect 16899 4008 16911 4060
rect 16963 4008 16975 4060
rect 17027 4008 17039 4060
rect 17091 4008 17103 4060
rect 17155 4008 17167 4060
rect 17219 4008 17231 4060
rect 17283 4008 17295 4060
rect 17347 4008 17469 4060
rect 17521 4008 17533 4060
rect 17585 4008 17597 4060
rect 17649 4008 17661 4060
rect 17713 4008 17725 4060
rect 17777 4008 17789 4060
rect 17841 4008 17853 4060
rect 17905 4008 17917 4060
rect 17969 4008 17981 4060
rect 18033 4008 18045 4060
rect 18097 4008 18109 4060
rect 18161 4008 18167 4060
rect 16649 4002 18167 4008
rect 16649 3344 16677 4002
rect 16705 3316 16733 3974
rect 16761 3344 16789 4002
rect 16817 3316 16845 3974
rect 16873 3344 16901 4002
rect 16929 3316 16957 3974
rect 16985 3344 17013 4002
rect 17041 3316 17069 3974
rect 17097 3344 17125 4002
rect 17153 3316 17181 3974
rect 17209 3344 17237 4002
rect 17265 3316 17293 3974
rect 17321 3344 17349 4002
rect 17381 3978 17435 4002
rect 17381 3926 17382 3978
rect 17434 3926 17435 3978
rect 17381 3914 17435 3926
rect 17381 3862 17382 3914
rect 17434 3862 17435 3914
rect 17381 3850 17435 3862
rect 17381 3798 17382 3850
rect 17434 3798 17435 3850
rect 17381 3786 17435 3798
rect 17381 3734 17382 3786
rect 17434 3734 17435 3786
rect 17381 3722 17435 3734
rect 17381 3670 17382 3722
rect 17434 3670 17435 3722
rect 17381 3658 17435 3670
rect 17381 3606 17382 3658
rect 17434 3606 17435 3658
rect 17381 3594 17435 3606
rect 17381 3542 17382 3594
rect 17434 3542 17435 3594
rect 17381 3530 17435 3542
rect 17381 3478 17382 3530
rect 17434 3478 17435 3530
rect 17381 3466 17435 3478
rect 17381 3414 17382 3466
rect 17434 3414 17435 3466
rect 17381 3402 17435 3414
rect 17381 3350 17382 3402
rect 17434 3350 17435 3402
rect 17381 3344 17435 3350
rect 17467 3344 17495 4002
rect 17523 3316 17551 3974
rect 17579 3344 17607 4002
rect 17635 3316 17663 3974
rect 17691 3344 17719 4002
rect 17747 3316 17775 3974
rect 17803 3344 17831 4002
rect 17859 3316 17887 3974
rect 17915 3344 17943 4002
rect 17971 3316 17999 3974
rect 18027 3344 18055 4002
rect 18083 3316 18111 3974
rect 18139 3344 18167 4002
rect 18200 4713 18207 4752
rect 18259 4713 18407 4765
rect 18459 4759 18488 4765
rect 18540 4759 18552 4811
rect 18604 4759 18616 4811
rect 18668 4759 18680 4811
rect 18732 4802 18744 4811
rect 18796 4802 18808 4811
rect 18860 4802 18872 4811
rect 18924 4802 18936 4811
rect 18988 4802 19000 4811
rect 19052 4802 19064 4811
rect 18735 4768 18744 4802
rect 18807 4768 18808 4802
rect 18988 4768 18989 4802
rect 19052 4768 19061 4802
rect 18732 4759 18744 4768
rect 18796 4759 18808 4768
rect 18860 4759 18872 4768
rect 18924 4759 18936 4768
rect 18988 4759 19000 4768
rect 19052 4759 19064 4768
rect 19116 4759 19128 4811
rect 19180 4802 19342 4811
rect 19180 4768 19205 4802
rect 19239 4768 19277 4802
rect 19311 4768 19342 4802
rect 19180 4759 19342 4768
rect 19394 4759 19406 4811
rect 19458 4759 19470 4811
rect 19522 4802 19534 4811
rect 19586 4802 19598 4811
rect 19650 4802 19662 4811
rect 19714 4802 19726 4811
rect 19778 4802 19790 4811
rect 19842 4802 19854 4811
rect 19527 4768 19534 4802
rect 19778 4768 19781 4802
rect 19842 4768 19853 4802
rect 19522 4759 19534 4768
rect 19586 4759 19598 4768
rect 19650 4759 19662 4768
rect 19714 4759 19726 4768
rect 19778 4759 19790 4768
rect 19842 4759 19854 4768
rect 19906 4759 19918 4811
rect 19970 4759 19982 4811
rect 20034 4765 20116 4811
rect 20034 4759 20057 4765
rect 18459 4752 20057 4759
rect 18459 4713 18466 4752
rect 18200 4701 18216 4713
rect 18250 4701 18416 4713
rect 18450 4701 18466 4713
rect 18200 4649 18207 4701
rect 18259 4649 18407 4701
rect 18459 4649 18466 4701
rect 18200 4637 18216 4649
rect 18250 4637 18416 4649
rect 18450 4637 18466 4649
rect 18200 4585 18207 4637
rect 18259 4585 18407 4637
rect 18459 4585 18466 4637
rect 18200 4573 18216 4585
rect 18250 4573 18416 4585
rect 18450 4573 18466 4585
rect 18200 4521 18207 4573
rect 18259 4521 18407 4573
rect 18459 4521 18466 4573
rect 18200 4519 18466 4521
rect 18200 4509 18216 4519
rect 18250 4509 18416 4519
rect 18450 4509 18466 4519
rect 18200 4457 18207 4509
rect 18259 4457 18407 4509
rect 18459 4457 18466 4509
rect 18200 4447 18466 4457
rect 18200 4445 18216 4447
rect 18250 4445 18416 4447
rect 18450 4445 18466 4447
rect 18200 4393 18207 4445
rect 18259 4393 18407 4445
rect 18459 4393 18466 4445
rect 18200 4381 18466 4393
rect 18200 4329 18207 4381
rect 18259 4329 18407 4381
rect 18459 4329 18466 4381
rect 18200 4317 18466 4329
rect 18200 4265 18207 4317
rect 18259 4265 18407 4317
rect 18459 4265 18466 4317
rect 18200 4253 18466 4265
rect 18200 4201 18207 4253
rect 18259 4201 18407 4253
rect 18459 4201 18466 4253
rect 18200 4197 18216 4201
rect 18250 4197 18416 4201
rect 18450 4197 18466 4201
rect 18200 4189 18466 4197
rect 18200 4137 18207 4189
rect 18259 4137 18407 4189
rect 18459 4137 18466 4189
rect 18200 4125 18216 4137
rect 18250 4125 18416 4137
rect 18450 4125 18466 4137
rect 18200 4087 18466 4125
rect 18200 4053 18216 4087
rect 18250 4053 18416 4087
rect 18450 4053 18466 4087
rect 18200 4015 18466 4053
rect 18200 3981 18216 4015
rect 18250 3981 18416 4015
rect 18450 3981 18466 4015
rect 18200 3943 18466 3981
rect 18200 3931 18216 3943
rect 18250 3931 18416 3943
rect 18450 3931 18466 3943
rect 18200 3879 18207 3931
rect 18259 3879 18407 3931
rect 18459 3879 18466 3931
rect 18200 3871 18466 3879
rect 18200 3867 18216 3871
rect 18250 3867 18416 3871
rect 18450 3867 18466 3871
rect 18200 3815 18207 3867
rect 18259 3815 18407 3867
rect 18459 3815 18466 3867
rect 18200 3803 18466 3815
rect 18200 3751 18207 3803
rect 18259 3751 18407 3803
rect 18459 3751 18466 3803
rect 18200 3739 18466 3751
rect 18200 3687 18207 3739
rect 18259 3687 18407 3739
rect 18459 3687 18466 3739
rect 18200 3675 18466 3687
rect 18200 3623 18207 3675
rect 18259 3623 18407 3675
rect 18459 3623 18466 3675
rect 18200 3621 18216 3623
rect 18250 3621 18416 3623
rect 18450 3621 18466 3623
rect 18200 3611 18466 3621
rect 18200 3559 18207 3611
rect 18259 3559 18407 3611
rect 18459 3559 18466 3611
rect 18200 3549 18216 3559
rect 18250 3549 18416 3559
rect 18450 3549 18466 3559
rect 18200 3547 18466 3549
rect 18200 3495 18207 3547
rect 18259 3495 18407 3547
rect 18459 3495 18466 3547
rect 18200 3483 18216 3495
rect 18250 3483 18416 3495
rect 18450 3483 18466 3495
rect 18200 3431 18207 3483
rect 18259 3431 18407 3483
rect 18459 3431 18466 3483
rect 18200 3419 18216 3431
rect 18250 3419 18416 3431
rect 18450 3419 18466 3431
rect 18200 3367 18207 3419
rect 18259 3367 18407 3419
rect 18459 3367 18466 3419
rect 18200 3355 18216 3367
rect 18250 3355 18416 3367
rect 18450 3355 18466 3367
rect 18200 3316 18207 3355
rect 16609 3309 18207 3316
rect 16609 3303 16638 3309
rect 16550 3300 16638 3303
rect 16550 3266 16635 3300
rect 16550 3257 16638 3266
rect 16690 3257 16702 3309
rect 16754 3257 16766 3309
rect 16818 3257 16830 3309
rect 16882 3300 16894 3309
rect 16946 3300 16958 3309
rect 17010 3300 17022 3309
rect 17074 3300 17086 3309
rect 17138 3300 17150 3309
rect 17202 3300 17214 3309
rect 16885 3266 16894 3300
rect 16957 3266 16958 3300
rect 17138 3266 17139 3300
rect 17202 3266 17211 3300
rect 16882 3257 16894 3266
rect 16946 3257 16958 3266
rect 17010 3257 17022 3266
rect 17074 3257 17086 3266
rect 17138 3257 17150 3266
rect 17202 3257 17214 3266
rect 17266 3257 17278 3309
rect 17330 3300 17492 3309
rect 17330 3266 17355 3300
rect 17389 3266 17427 3300
rect 17461 3266 17492 3300
rect 17330 3257 17492 3266
rect 17544 3257 17556 3309
rect 17608 3257 17620 3309
rect 17672 3300 17684 3309
rect 17736 3300 17748 3309
rect 17800 3300 17812 3309
rect 17864 3300 17876 3309
rect 17928 3300 17940 3309
rect 17992 3300 18004 3309
rect 17677 3266 17684 3300
rect 17928 3266 17931 3300
rect 17992 3266 18003 3300
rect 17672 3257 17684 3266
rect 17736 3257 17748 3266
rect 17800 3257 17812 3266
rect 17864 3257 17876 3266
rect 17928 3257 17940 3266
rect 17992 3257 18004 3266
rect 18056 3257 18068 3309
rect 18120 3257 18132 3309
rect 18184 3303 18207 3309
rect 18259 3303 18407 3355
rect 18459 3316 18466 3355
rect 18499 4066 18527 4724
rect 18555 4094 18583 4752
rect 18611 4066 18639 4724
rect 18667 4094 18695 4752
rect 18723 4066 18751 4724
rect 18779 4094 18807 4752
rect 18835 4066 18863 4724
rect 18891 4094 18919 4752
rect 18947 4066 18975 4724
rect 19003 4094 19031 4752
rect 19059 4066 19087 4724
rect 19115 4094 19143 4752
rect 19171 4066 19199 4724
rect 19231 4718 19285 4724
rect 19231 4666 19232 4718
rect 19284 4666 19285 4718
rect 19231 4654 19285 4666
rect 19231 4602 19232 4654
rect 19284 4602 19285 4654
rect 19231 4590 19285 4602
rect 19231 4538 19232 4590
rect 19284 4538 19285 4590
rect 19231 4526 19285 4538
rect 19231 4474 19232 4526
rect 19284 4474 19285 4526
rect 19231 4462 19285 4474
rect 19231 4410 19232 4462
rect 19284 4410 19285 4462
rect 19231 4398 19285 4410
rect 19231 4346 19232 4398
rect 19284 4346 19285 4398
rect 19231 4334 19285 4346
rect 19231 4282 19232 4334
rect 19284 4282 19285 4334
rect 19231 4270 19285 4282
rect 19231 4218 19232 4270
rect 19284 4218 19285 4270
rect 19231 4206 19285 4218
rect 19231 4154 19232 4206
rect 19284 4154 19285 4206
rect 19231 4142 19285 4154
rect 19231 4090 19232 4142
rect 19284 4090 19285 4142
rect 19231 4066 19285 4090
rect 19317 4066 19345 4724
rect 19373 4094 19401 4752
rect 19429 4066 19457 4724
rect 19485 4094 19513 4752
rect 19541 4066 19569 4724
rect 19597 4094 19625 4752
rect 19653 4066 19681 4724
rect 19709 4094 19737 4752
rect 19765 4066 19793 4724
rect 19821 4094 19849 4752
rect 19877 4066 19905 4724
rect 19933 4094 19961 4752
rect 19989 4066 20017 4724
rect 18499 4060 20017 4066
rect 18499 4008 18505 4060
rect 18557 4008 18569 4060
rect 18621 4008 18633 4060
rect 18685 4008 18697 4060
rect 18749 4008 18761 4060
rect 18813 4008 18825 4060
rect 18877 4008 18889 4060
rect 18941 4008 18953 4060
rect 19005 4008 19017 4060
rect 19069 4008 19081 4060
rect 19133 4008 19145 4060
rect 19197 4008 19319 4060
rect 19371 4008 19383 4060
rect 19435 4008 19447 4060
rect 19499 4008 19511 4060
rect 19563 4008 19575 4060
rect 19627 4008 19639 4060
rect 19691 4008 19703 4060
rect 19755 4008 19767 4060
rect 19819 4008 19831 4060
rect 19883 4008 19895 4060
rect 19947 4008 19959 4060
rect 20011 4008 20017 4060
rect 18499 4002 20017 4008
rect 18499 3344 18527 4002
rect 18555 3316 18583 3974
rect 18611 3344 18639 4002
rect 18667 3316 18695 3974
rect 18723 3344 18751 4002
rect 18779 3316 18807 3974
rect 18835 3344 18863 4002
rect 18891 3316 18919 3974
rect 18947 3344 18975 4002
rect 19003 3316 19031 3974
rect 19059 3344 19087 4002
rect 19115 3316 19143 3974
rect 19171 3344 19199 4002
rect 19231 3978 19285 4002
rect 19231 3926 19232 3978
rect 19284 3926 19285 3978
rect 19231 3914 19285 3926
rect 19231 3862 19232 3914
rect 19284 3862 19285 3914
rect 19231 3850 19285 3862
rect 19231 3798 19232 3850
rect 19284 3798 19285 3850
rect 19231 3786 19285 3798
rect 19231 3734 19232 3786
rect 19284 3734 19285 3786
rect 19231 3722 19285 3734
rect 19231 3670 19232 3722
rect 19284 3670 19285 3722
rect 19231 3658 19285 3670
rect 19231 3606 19232 3658
rect 19284 3606 19285 3658
rect 19231 3594 19285 3606
rect 19231 3542 19232 3594
rect 19284 3542 19285 3594
rect 19231 3530 19285 3542
rect 19231 3478 19232 3530
rect 19284 3478 19285 3530
rect 19231 3466 19285 3478
rect 19231 3414 19232 3466
rect 19284 3414 19285 3466
rect 19231 3402 19285 3414
rect 19231 3350 19232 3402
rect 19284 3350 19285 3402
rect 19231 3344 19285 3350
rect 19317 3344 19345 4002
rect 19373 3316 19401 3974
rect 19429 3344 19457 4002
rect 19485 3316 19513 3974
rect 19541 3344 19569 4002
rect 19597 3316 19625 3974
rect 19653 3344 19681 4002
rect 19709 3316 19737 3974
rect 19765 3344 19793 4002
rect 19821 3316 19849 3974
rect 19877 3344 19905 4002
rect 19933 3316 19961 3974
rect 19989 3344 20017 4002
rect 20050 4713 20057 4752
rect 20109 4713 20116 4765
rect 20050 4701 20066 4713
rect 20100 4701 20116 4713
rect 20050 4649 20057 4701
rect 20109 4649 20116 4701
rect 20050 4637 20066 4649
rect 20100 4637 20116 4649
rect 20050 4585 20057 4637
rect 20109 4585 20116 4637
rect 20050 4573 20066 4585
rect 20100 4573 20116 4585
rect 20050 4521 20057 4573
rect 20109 4521 20116 4573
rect 20050 4519 20116 4521
rect 20050 4509 20066 4519
rect 20100 4509 20116 4519
rect 20050 4457 20057 4509
rect 20109 4457 20116 4509
rect 20050 4447 20116 4457
rect 20050 4445 20066 4447
rect 20100 4445 20116 4447
rect 20050 4393 20057 4445
rect 20109 4393 20116 4445
rect 20050 4381 20116 4393
rect 20050 4329 20057 4381
rect 20109 4329 20116 4381
rect 20050 4317 20116 4329
rect 20050 4265 20057 4317
rect 20109 4265 20116 4317
rect 20050 4253 20116 4265
rect 20050 4201 20057 4253
rect 20109 4201 20116 4253
rect 20050 4197 20066 4201
rect 20100 4197 20116 4201
rect 20050 4189 20116 4197
rect 20050 4137 20057 4189
rect 20109 4137 20116 4189
rect 20050 4125 20066 4137
rect 20100 4125 20116 4137
rect 20050 4087 20116 4125
rect 20050 4053 20066 4087
rect 20100 4053 20116 4087
rect 20050 4015 20116 4053
rect 20050 3981 20066 4015
rect 20100 3981 20116 4015
rect 20050 3943 20116 3981
rect 20050 3931 20066 3943
rect 20100 3931 20116 3943
rect 20050 3879 20057 3931
rect 20109 3879 20116 3931
rect 20050 3871 20116 3879
rect 20050 3867 20066 3871
rect 20100 3867 20116 3871
rect 20050 3815 20057 3867
rect 20109 3815 20116 3867
rect 20050 3803 20116 3815
rect 20050 3751 20057 3803
rect 20109 3751 20116 3803
rect 20050 3739 20116 3751
rect 20050 3687 20057 3739
rect 20109 3687 20116 3739
rect 20050 3675 20116 3687
rect 20050 3623 20057 3675
rect 20109 3623 20116 3675
rect 20050 3621 20066 3623
rect 20100 3621 20116 3623
rect 20050 3611 20116 3621
rect 20050 3559 20057 3611
rect 20109 3559 20116 3611
rect 20050 3549 20066 3559
rect 20100 3549 20116 3559
rect 20050 3547 20116 3549
rect 20050 3495 20057 3547
rect 20109 3495 20116 3547
rect 20050 3483 20066 3495
rect 20100 3483 20116 3495
rect 20050 3431 20057 3483
rect 20109 3431 20116 3483
rect 20050 3419 20066 3431
rect 20100 3419 20116 3431
rect 20050 3367 20057 3419
rect 20109 3367 20116 3419
rect 20050 3355 20066 3367
rect 20100 3355 20116 3367
rect 20050 3316 20057 3355
rect 18459 3309 20057 3316
rect 18459 3303 18488 3309
rect 18184 3300 18488 3303
rect 18184 3266 18485 3300
rect 18184 3257 18488 3266
rect 18540 3257 18552 3309
rect 18604 3257 18616 3309
rect 18668 3257 18680 3309
rect 18732 3300 18744 3309
rect 18796 3300 18808 3309
rect 18860 3300 18872 3309
rect 18924 3300 18936 3309
rect 18988 3300 19000 3309
rect 19052 3300 19064 3309
rect 18735 3266 18744 3300
rect 18807 3266 18808 3300
rect 18988 3266 18989 3300
rect 19052 3266 19061 3300
rect 18732 3257 18744 3266
rect 18796 3257 18808 3266
rect 18860 3257 18872 3266
rect 18924 3257 18936 3266
rect 18988 3257 19000 3266
rect 19052 3257 19064 3266
rect 19116 3257 19128 3309
rect 19180 3300 19342 3309
rect 19180 3266 19205 3300
rect 19239 3266 19277 3300
rect 19311 3266 19342 3300
rect 19180 3257 19342 3266
rect 19394 3257 19406 3309
rect 19458 3257 19470 3309
rect 19522 3300 19534 3309
rect 19586 3300 19598 3309
rect 19650 3300 19662 3309
rect 19714 3300 19726 3309
rect 19778 3300 19790 3309
rect 19842 3300 19854 3309
rect 19527 3266 19534 3300
rect 19778 3266 19781 3300
rect 19842 3266 19853 3300
rect 19522 3257 19534 3266
rect 19586 3257 19598 3266
rect 19650 3257 19662 3266
rect 19714 3257 19726 3266
rect 19778 3257 19790 3266
rect 19842 3257 19854 3266
rect 19906 3257 19918 3309
rect 19970 3257 19982 3309
rect 20034 3303 20057 3309
rect 20109 3303 20116 3355
rect 20034 3257 20116 3303
rect 16550 3250 20116 3257
<< via1 >>
rect 16638 9852 16690 9861
rect 16638 9818 16669 9852
rect 16669 9818 16690 9852
rect 16557 9785 16609 9815
rect 16638 9809 16690 9818
rect 16702 9852 16754 9861
rect 16702 9818 16707 9852
rect 16707 9818 16741 9852
rect 16741 9818 16754 9852
rect 16702 9809 16754 9818
rect 16766 9852 16818 9861
rect 16766 9818 16779 9852
rect 16779 9818 16813 9852
rect 16813 9818 16818 9852
rect 16766 9809 16818 9818
rect 16830 9852 16882 9861
rect 16894 9852 16946 9861
rect 16958 9852 17010 9861
rect 17022 9852 17074 9861
rect 17086 9852 17138 9861
rect 17150 9852 17202 9861
rect 17214 9852 17266 9861
rect 16830 9818 16851 9852
rect 16851 9818 16882 9852
rect 16894 9818 16923 9852
rect 16923 9818 16946 9852
rect 16958 9818 16995 9852
rect 16995 9818 17010 9852
rect 17022 9818 17029 9852
rect 17029 9818 17067 9852
rect 17067 9818 17074 9852
rect 17086 9818 17101 9852
rect 17101 9818 17138 9852
rect 17150 9818 17173 9852
rect 17173 9818 17202 9852
rect 17214 9818 17245 9852
rect 17245 9818 17266 9852
rect 16830 9809 16882 9818
rect 16894 9809 16946 9818
rect 16958 9809 17010 9818
rect 17022 9809 17074 9818
rect 17086 9809 17138 9818
rect 17150 9809 17202 9818
rect 17214 9809 17266 9818
rect 17278 9852 17330 9861
rect 17492 9852 17544 9861
rect 17278 9818 17283 9852
rect 17283 9818 17317 9852
rect 17317 9818 17330 9852
rect 17492 9818 17499 9852
rect 17499 9818 17533 9852
rect 17533 9818 17544 9852
rect 17278 9809 17330 9818
rect 17492 9809 17544 9818
rect 17556 9852 17608 9861
rect 17556 9818 17571 9852
rect 17571 9818 17605 9852
rect 17605 9818 17608 9852
rect 17556 9809 17608 9818
rect 17620 9852 17672 9861
rect 17684 9852 17736 9861
rect 17748 9852 17800 9861
rect 17812 9852 17864 9861
rect 17876 9852 17928 9861
rect 17940 9852 17992 9861
rect 18004 9852 18056 9861
rect 17620 9818 17643 9852
rect 17643 9818 17672 9852
rect 17684 9818 17715 9852
rect 17715 9818 17736 9852
rect 17748 9818 17749 9852
rect 17749 9818 17787 9852
rect 17787 9818 17800 9852
rect 17812 9818 17821 9852
rect 17821 9818 17859 9852
rect 17859 9818 17864 9852
rect 17876 9818 17893 9852
rect 17893 9818 17928 9852
rect 17940 9818 17965 9852
rect 17965 9818 17992 9852
rect 18004 9818 18037 9852
rect 18037 9818 18056 9852
rect 17620 9809 17672 9818
rect 17684 9809 17736 9818
rect 17748 9809 17800 9818
rect 17812 9809 17864 9818
rect 17876 9809 17928 9818
rect 17940 9809 17992 9818
rect 18004 9809 18056 9818
rect 18068 9852 18120 9861
rect 18068 9818 18075 9852
rect 18075 9818 18109 9852
rect 18109 9818 18120 9852
rect 18068 9809 18120 9818
rect 18132 9852 18184 9861
rect 18488 9852 18540 9861
rect 18132 9818 18147 9852
rect 18147 9818 18181 9852
rect 18181 9818 18184 9852
rect 18488 9818 18519 9852
rect 18519 9818 18540 9852
rect 18132 9809 18184 9818
rect 16557 9763 16566 9785
rect 16566 9763 16600 9785
rect 16600 9763 16609 9785
rect 16557 9713 16609 9751
rect 16557 9699 16566 9713
rect 16566 9699 16600 9713
rect 16600 9699 16609 9713
rect 16557 9679 16566 9687
rect 16566 9679 16600 9687
rect 16600 9679 16609 9687
rect 16557 9641 16609 9679
rect 16557 9635 16566 9641
rect 16566 9635 16600 9641
rect 16600 9635 16609 9641
rect 16557 9607 16566 9623
rect 16566 9607 16600 9623
rect 16600 9607 16609 9623
rect 16557 9571 16609 9607
rect 16557 9535 16566 9559
rect 16566 9535 16600 9559
rect 16600 9535 16609 9559
rect 16557 9507 16609 9535
rect 16557 9463 16566 9495
rect 16566 9463 16600 9495
rect 16600 9463 16609 9495
rect 16557 9443 16609 9463
rect 16557 9425 16609 9431
rect 16557 9391 16566 9425
rect 16566 9391 16600 9425
rect 16600 9391 16609 9425
rect 16557 9379 16609 9391
rect 16557 9353 16609 9367
rect 16557 9319 16566 9353
rect 16566 9319 16600 9353
rect 16600 9319 16609 9353
rect 16557 9315 16609 9319
rect 16557 9281 16609 9303
rect 16557 9251 16566 9281
rect 16566 9251 16600 9281
rect 16600 9251 16609 9281
rect 16557 9209 16609 9239
rect 16557 9187 16566 9209
rect 16566 9187 16600 9209
rect 16600 9187 16609 9209
rect 16557 8959 16566 8981
rect 16566 8959 16600 8981
rect 16600 8959 16609 8981
rect 16557 8929 16609 8959
rect 16557 8887 16566 8917
rect 16566 8887 16600 8917
rect 16600 8887 16609 8917
rect 16557 8865 16609 8887
rect 16557 8849 16609 8853
rect 16557 8815 16566 8849
rect 16566 8815 16600 8849
rect 16600 8815 16609 8849
rect 16557 8801 16609 8815
rect 16557 8777 16609 8789
rect 16557 8743 16566 8777
rect 16566 8743 16600 8777
rect 16600 8743 16609 8777
rect 16557 8737 16609 8743
rect 16557 8705 16609 8725
rect 16557 8673 16566 8705
rect 16566 8673 16600 8705
rect 16600 8673 16609 8705
rect 16557 8633 16609 8661
rect 16557 8609 16566 8633
rect 16566 8609 16600 8633
rect 16600 8609 16609 8633
rect 16557 8561 16609 8597
rect 16557 8545 16566 8561
rect 16566 8545 16600 8561
rect 16600 8545 16609 8561
rect 16557 8527 16566 8533
rect 16566 8527 16600 8533
rect 16600 8527 16609 8533
rect 16557 8489 16609 8527
rect 16557 8481 16566 8489
rect 16566 8481 16600 8489
rect 16600 8481 16609 8489
rect 16557 8455 16566 8469
rect 16566 8455 16600 8469
rect 16600 8455 16609 8469
rect 16557 8417 16609 8455
rect 16557 8383 16566 8405
rect 16566 8383 16600 8405
rect 16600 8383 16609 8405
rect 16557 8353 16609 8383
rect 17382 9716 17434 9768
rect 17382 9652 17434 9704
rect 17382 9588 17434 9640
rect 17382 9524 17434 9576
rect 17382 9460 17434 9512
rect 17382 9396 17434 9448
rect 17382 9332 17434 9384
rect 17382 9268 17434 9320
rect 17382 9204 17434 9256
rect 17382 9140 17434 9192
rect 16655 9058 16707 9110
rect 16719 9058 16771 9110
rect 16783 9058 16835 9110
rect 16847 9058 16899 9110
rect 16911 9058 16963 9110
rect 16975 9058 17027 9110
rect 17039 9058 17091 9110
rect 17103 9058 17155 9110
rect 17167 9058 17219 9110
rect 17231 9058 17283 9110
rect 17295 9058 17347 9110
rect 17469 9058 17521 9110
rect 17533 9058 17585 9110
rect 17597 9058 17649 9110
rect 17661 9058 17713 9110
rect 17725 9058 17777 9110
rect 17789 9058 17841 9110
rect 17853 9058 17905 9110
rect 17917 9058 17969 9110
rect 17981 9058 18033 9110
rect 18045 9058 18097 9110
rect 18109 9058 18161 9110
rect 17382 8976 17434 9028
rect 17382 8912 17434 8964
rect 17382 8848 17434 8900
rect 17382 8784 17434 8836
rect 17382 8720 17434 8772
rect 17382 8656 17434 8708
rect 17382 8592 17434 8644
rect 17382 8528 17434 8580
rect 17382 8464 17434 8516
rect 17382 8400 17434 8452
rect 18207 9785 18259 9815
rect 18207 9763 18216 9785
rect 18216 9763 18250 9785
rect 18250 9763 18259 9785
rect 18407 9785 18459 9815
rect 18488 9809 18540 9818
rect 18552 9852 18604 9861
rect 18552 9818 18557 9852
rect 18557 9818 18591 9852
rect 18591 9818 18604 9852
rect 18552 9809 18604 9818
rect 18616 9852 18668 9861
rect 18616 9818 18629 9852
rect 18629 9818 18663 9852
rect 18663 9818 18668 9852
rect 18616 9809 18668 9818
rect 18680 9852 18732 9861
rect 18744 9852 18796 9861
rect 18808 9852 18860 9861
rect 18872 9852 18924 9861
rect 18936 9852 18988 9861
rect 19000 9852 19052 9861
rect 19064 9852 19116 9861
rect 18680 9818 18701 9852
rect 18701 9818 18732 9852
rect 18744 9818 18773 9852
rect 18773 9818 18796 9852
rect 18808 9818 18845 9852
rect 18845 9818 18860 9852
rect 18872 9818 18879 9852
rect 18879 9818 18917 9852
rect 18917 9818 18924 9852
rect 18936 9818 18951 9852
rect 18951 9818 18988 9852
rect 19000 9818 19023 9852
rect 19023 9818 19052 9852
rect 19064 9818 19095 9852
rect 19095 9818 19116 9852
rect 18680 9809 18732 9818
rect 18744 9809 18796 9818
rect 18808 9809 18860 9818
rect 18872 9809 18924 9818
rect 18936 9809 18988 9818
rect 19000 9809 19052 9818
rect 19064 9809 19116 9818
rect 19128 9852 19180 9861
rect 19342 9852 19394 9861
rect 19128 9818 19133 9852
rect 19133 9818 19167 9852
rect 19167 9818 19180 9852
rect 19342 9818 19349 9852
rect 19349 9818 19383 9852
rect 19383 9818 19394 9852
rect 19128 9809 19180 9818
rect 19342 9809 19394 9818
rect 19406 9852 19458 9861
rect 19406 9818 19421 9852
rect 19421 9818 19455 9852
rect 19455 9818 19458 9852
rect 19406 9809 19458 9818
rect 19470 9852 19522 9861
rect 19534 9852 19586 9861
rect 19598 9852 19650 9861
rect 19662 9852 19714 9861
rect 19726 9852 19778 9861
rect 19790 9852 19842 9861
rect 19854 9852 19906 9861
rect 19470 9818 19493 9852
rect 19493 9818 19522 9852
rect 19534 9818 19565 9852
rect 19565 9818 19586 9852
rect 19598 9818 19599 9852
rect 19599 9818 19637 9852
rect 19637 9818 19650 9852
rect 19662 9818 19671 9852
rect 19671 9818 19709 9852
rect 19709 9818 19714 9852
rect 19726 9818 19743 9852
rect 19743 9818 19778 9852
rect 19790 9818 19815 9852
rect 19815 9818 19842 9852
rect 19854 9818 19887 9852
rect 19887 9818 19906 9852
rect 19470 9809 19522 9818
rect 19534 9809 19586 9818
rect 19598 9809 19650 9818
rect 19662 9809 19714 9818
rect 19726 9809 19778 9818
rect 19790 9809 19842 9818
rect 19854 9809 19906 9818
rect 19918 9852 19970 9861
rect 19918 9818 19925 9852
rect 19925 9818 19959 9852
rect 19959 9818 19970 9852
rect 19918 9809 19970 9818
rect 19982 9852 20034 9861
rect 19982 9818 19997 9852
rect 19997 9818 20031 9852
rect 20031 9818 20034 9852
rect 19982 9809 20034 9818
rect 18407 9763 18416 9785
rect 18416 9763 18450 9785
rect 18450 9763 18459 9785
rect 18207 9713 18259 9751
rect 18207 9699 18216 9713
rect 18216 9699 18250 9713
rect 18250 9699 18259 9713
rect 18407 9713 18459 9751
rect 18407 9699 18416 9713
rect 18416 9699 18450 9713
rect 18450 9699 18459 9713
rect 18207 9679 18216 9687
rect 18216 9679 18250 9687
rect 18250 9679 18259 9687
rect 18207 9641 18259 9679
rect 18207 9635 18216 9641
rect 18216 9635 18250 9641
rect 18250 9635 18259 9641
rect 18407 9679 18416 9687
rect 18416 9679 18450 9687
rect 18450 9679 18459 9687
rect 18407 9641 18459 9679
rect 18407 9635 18416 9641
rect 18416 9635 18450 9641
rect 18450 9635 18459 9641
rect 18207 9607 18216 9623
rect 18216 9607 18250 9623
rect 18250 9607 18259 9623
rect 18207 9571 18259 9607
rect 18407 9607 18416 9623
rect 18416 9607 18450 9623
rect 18450 9607 18459 9623
rect 18407 9571 18459 9607
rect 18207 9535 18216 9559
rect 18216 9535 18250 9559
rect 18250 9535 18259 9559
rect 18207 9507 18259 9535
rect 18407 9535 18416 9559
rect 18416 9535 18450 9559
rect 18450 9535 18459 9559
rect 18407 9507 18459 9535
rect 18207 9463 18216 9495
rect 18216 9463 18250 9495
rect 18250 9463 18259 9495
rect 18207 9443 18259 9463
rect 18407 9463 18416 9495
rect 18416 9463 18450 9495
rect 18450 9463 18459 9495
rect 18407 9443 18459 9463
rect 18207 9425 18259 9431
rect 18207 9391 18216 9425
rect 18216 9391 18250 9425
rect 18250 9391 18259 9425
rect 18207 9379 18259 9391
rect 18407 9425 18459 9431
rect 18407 9391 18416 9425
rect 18416 9391 18450 9425
rect 18450 9391 18459 9425
rect 18407 9379 18459 9391
rect 18207 9353 18259 9367
rect 18207 9319 18216 9353
rect 18216 9319 18250 9353
rect 18250 9319 18259 9353
rect 18207 9315 18259 9319
rect 18407 9353 18459 9367
rect 18407 9319 18416 9353
rect 18416 9319 18450 9353
rect 18450 9319 18459 9353
rect 18407 9315 18459 9319
rect 18207 9281 18259 9303
rect 18207 9251 18216 9281
rect 18216 9251 18250 9281
rect 18250 9251 18259 9281
rect 18407 9281 18459 9303
rect 18407 9251 18416 9281
rect 18416 9251 18450 9281
rect 18450 9251 18459 9281
rect 18207 9209 18259 9239
rect 18207 9187 18216 9209
rect 18216 9187 18250 9209
rect 18250 9187 18259 9209
rect 18407 9209 18459 9239
rect 18407 9187 18416 9209
rect 18416 9187 18450 9209
rect 18450 9187 18459 9209
rect 18207 8959 18216 8981
rect 18216 8959 18250 8981
rect 18250 8959 18259 8981
rect 18207 8929 18259 8959
rect 18407 8959 18416 8981
rect 18416 8959 18450 8981
rect 18450 8959 18459 8981
rect 18407 8929 18459 8959
rect 18207 8887 18216 8917
rect 18216 8887 18250 8917
rect 18250 8887 18259 8917
rect 18207 8865 18259 8887
rect 18407 8887 18416 8917
rect 18416 8887 18450 8917
rect 18450 8887 18459 8917
rect 18407 8865 18459 8887
rect 18207 8849 18259 8853
rect 18207 8815 18216 8849
rect 18216 8815 18250 8849
rect 18250 8815 18259 8849
rect 18207 8801 18259 8815
rect 18407 8849 18459 8853
rect 18407 8815 18416 8849
rect 18416 8815 18450 8849
rect 18450 8815 18459 8849
rect 18407 8801 18459 8815
rect 18207 8777 18259 8789
rect 18207 8743 18216 8777
rect 18216 8743 18250 8777
rect 18250 8743 18259 8777
rect 18207 8737 18259 8743
rect 18407 8777 18459 8789
rect 18407 8743 18416 8777
rect 18416 8743 18450 8777
rect 18450 8743 18459 8777
rect 18407 8737 18459 8743
rect 18207 8705 18259 8725
rect 18207 8673 18216 8705
rect 18216 8673 18250 8705
rect 18250 8673 18259 8705
rect 18407 8705 18459 8725
rect 18407 8673 18416 8705
rect 18416 8673 18450 8705
rect 18450 8673 18459 8705
rect 18207 8633 18259 8661
rect 18207 8609 18216 8633
rect 18216 8609 18250 8633
rect 18250 8609 18259 8633
rect 18407 8633 18459 8661
rect 18407 8609 18416 8633
rect 18416 8609 18450 8633
rect 18450 8609 18459 8633
rect 18207 8561 18259 8597
rect 18207 8545 18216 8561
rect 18216 8545 18250 8561
rect 18250 8545 18259 8561
rect 18407 8561 18459 8597
rect 18407 8545 18416 8561
rect 18416 8545 18450 8561
rect 18450 8545 18459 8561
rect 18207 8527 18216 8533
rect 18216 8527 18250 8533
rect 18250 8527 18259 8533
rect 18207 8489 18259 8527
rect 18207 8481 18216 8489
rect 18216 8481 18250 8489
rect 18250 8481 18259 8489
rect 18407 8527 18416 8533
rect 18416 8527 18450 8533
rect 18450 8527 18459 8533
rect 18407 8489 18459 8527
rect 18407 8481 18416 8489
rect 18416 8481 18450 8489
rect 18450 8481 18459 8489
rect 18207 8455 18216 8469
rect 18216 8455 18250 8469
rect 18250 8455 18259 8469
rect 18207 8417 18259 8455
rect 18407 8455 18416 8469
rect 18416 8455 18450 8469
rect 18450 8455 18459 8469
rect 18407 8417 18459 8455
rect 18207 8383 18216 8405
rect 18216 8383 18250 8405
rect 18250 8383 18259 8405
rect 16638 8350 16690 8359
rect 16638 8316 16669 8350
rect 16669 8316 16690 8350
rect 16638 8307 16690 8316
rect 16702 8350 16754 8359
rect 16702 8316 16707 8350
rect 16707 8316 16741 8350
rect 16741 8316 16754 8350
rect 16702 8307 16754 8316
rect 16766 8350 16818 8359
rect 16766 8316 16779 8350
rect 16779 8316 16813 8350
rect 16813 8316 16818 8350
rect 16766 8307 16818 8316
rect 16830 8350 16882 8359
rect 16894 8350 16946 8359
rect 16958 8350 17010 8359
rect 17022 8350 17074 8359
rect 17086 8350 17138 8359
rect 17150 8350 17202 8359
rect 17214 8350 17266 8359
rect 16830 8316 16851 8350
rect 16851 8316 16882 8350
rect 16894 8316 16923 8350
rect 16923 8316 16946 8350
rect 16958 8316 16995 8350
rect 16995 8316 17010 8350
rect 17022 8316 17029 8350
rect 17029 8316 17067 8350
rect 17067 8316 17074 8350
rect 17086 8316 17101 8350
rect 17101 8316 17138 8350
rect 17150 8316 17173 8350
rect 17173 8316 17202 8350
rect 17214 8316 17245 8350
rect 17245 8316 17266 8350
rect 16830 8307 16882 8316
rect 16894 8307 16946 8316
rect 16958 8307 17010 8316
rect 17022 8307 17074 8316
rect 17086 8307 17138 8316
rect 17150 8307 17202 8316
rect 17214 8307 17266 8316
rect 17278 8350 17330 8359
rect 17492 8350 17544 8359
rect 17278 8316 17283 8350
rect 17283 8316 17317 8350
rect 17317 8316 17330 8350
rect 17492 8316 17499 8350
rect 17499 8316 17533 8350
rect 17533 8316 17544 8350
rect 17278 8307 17330 8316
rect 17492 8307 17544 8316
rect 17556 8350 17608 8359
rect 17556 8316 17571 8350
rect 17571 8316 17605 8350
rect 17605 8316 17608 8350
rect 17556 8307 17608 8316
rect 17620 8350 17672 8359
rect 17684 8350 17736 8359
rect 17748 8350 17800 8359
rect 17812 8350 17864 8359
rect 17876 8350 17928 8359
rect 17940 8350 17992 8359
rect 18004 8350 18056 8359
rect 17620 8316 17643 8350
rect 17643 8316 17672 8350
rect 17684 8316 17715 8350
rect 17715 8316 17736 8350
rect 17748 8316 17749 8350
rect 17749 8316 17787 8350
rect 17787 8316 17800 8350
rect 17812 8316 17821 8350
rect 17821 8316 17859 8350
rect 17859 8316 17864 8350
rect 17876 8316 17893 8350
rect 17893 8316 17928 8350
rect 17940 8316 17965 8350
rect 17965 8316 17992 8350
rect 18004 8316 18037 8350
rect 18037 8316 18056 8350
rect 17620 8307 17672 8316
rect 17684 8307 17736 8316
rect 17748 8307 17800 8316
rect 17812 8307 17864 8316
rect 17876 8307 17928 8316
rect 17940 8307 17992 8316
rect 18004 8307 18056 8316
rect 18068 8350 18120 8359
rect 18068 8316 18075 8350
rect 18075 8316 18109 8350
rect 18109 8316 18120 8350
rect 18068 8307 18120 8316
rect 18132 8350 18184 8359
rect 18207 8353 18259 8383
rect 18407 8383 18416 8405
rect 18416 8383 18450 8405
rect 18450 8383 18459 8405
rect 18407 8353 18459 8383
rect 19232 9716 19284 9768
rect 19232 9652 19284 9704
rect 19232 9588 19284 9640
rect 19232 9524 19284 9576
rect 19232 9460 19284 9512
rect 19232 9396 19284 9448
rect 19232 9332 19284 9384
rect 19232 9268 19284 9320
rect 19232 9204 19284 9256
rect 19232 9140 19284 9192
rect 18505 9058 18557 9110
rect 18569 9058 18621 9110
rect 18633 9058 18685 9110
rect 18697 9058 18749 9110
rect 18761 9058 18813 9110
rect 18825 9058 18877 9110
rect 18889 9058 18941 9110
rect 18953 9058 19005 9110
rect 19017 9058 19069 9110
rect 19081 9058 19133 9110
rect 19145 9058 19197 9110
rect 19319 9058 19371 9110
rect 19383 9058 19435 9110
rect 19447 9058 19499 9110
rect 19511 9058 19563 9110
rect 19575 9058 19627 9110
rect 19639 9058 19691 9110
rect 19703 9058 19755 9110
rect 19767 9058 19819 9110
rect 19831 9058 19883 9110
rect 19895 9058 19947 9110
rect 19959 9058 20011 9110
rect 19232 8976 19284 9028
rect 19232 8912 19284 8964
rect 19232 8848 19284 8900
rect 19232 8784 19284 8836
rect 19232 8720 19284 8772
rect 19232 8656 19284 8708
rect 19232 8592 19284 8644
rect 19232 8528 19284 8580
rect 19232 8464 19284 8516
rect 19232 8400 19284 8452
rect 20057 9785 20109 9815
rect 20057 9763 20066 9785
rect 20066 9763 20100 9785
rect 20100 9763 20109 9785
rect 20057 9713 20109 9751
rect 20057 9699 20066 9713
rect 20066 9699 20100 9713
rect 20100 9699 20109 9713
rect 20057 9679 20066 9687
rect 20066 9679 20100 9687
rect 20100 9679 20109 9687
rect 20057 9641 20109 9679
rect 20057 9635 20066 9641
rect 20066 9635 20100 9641
rect 20100 9635 20109 9641
rect 20057 9607 20066 9623
rect 20066 9607 20100 9623
rect 20100 9607 20109 9623
rect 20057 9571 20109 9607
rect 20057 9535 20066 9559
rect 20066 9535 20100 9559
rect 20100 9535 20109 9559
rect 20057 9507 20109 9535
rect 20057 9463 20066 9495
rect 20066 9463 20100 9495
rect 20100 9463 20109 9495
rect 20057 9443 20109 9463
rect 20057 9425 20109 9431
rect 20057 9391 20066 9425
rect 20066 9391 20100 9425
rect 20100 9391 20109 9425
rect 20057 9379 20109 9391
rect 20057 9353 20109 9367
rect 20057 9319 20066 9353
rect 20066 9319 20100 9353
rect 20100 9319 20109 9353
rect 20057 9315 20109 9319
rect 20057 9281 20109 9303
rect 20057 9251 20066 9281
rect 20066 9251 20100 9281
rect 20100 9251 20109 9281
rect 20057 9209 20109 9239
rect 20057 9187 20066 9209
rect 20066 9187 20100 9209
rect 20100 9187 20109 9209
rect 20057 8959 20066 8981
rect 20066 8959 20100 8981
rect 20100 8959 20109 8981
rect 20057 8929 20109 8959
rect 20057 8887 20066 8917
rect 20066 8887 20100 8917
rect 20100 8887 20109 8917
rect 20057 8865 20109 8887
rect 20057 8849 20109 8853
rect 20057 8815 20066 8849
rect 20066 8815 20100 8849
rect 20100 8815 20109 8849
rect 20057 8801 20109 8815
rect 20057 8777 20109 8789
rect 20057 8743 20066 8777
rect 20066 8743 20100 8777
rect 20100 8743 20109 8777
rect 20057 8737 20109 8743
rect 20057 8705 20109 8725
rect 20057 8673 20066 8705
rect 20066 8673 20100 8705
rect 20100 8673 20109 8705
rect 20057 8633 20109 8661
rect 20057 8609 20066 8633
rect 20066 8609 20100 8633
rect 20100 8609 20109 8633
rect 20057 8561 20109 8597
rect 20057 8545 20066 8561
rect 20066 8545 20100 8561
rect 20100 8545 20109 8561
rect 20057 8527 20066 8533
rect 20066 8527 20100 8533
rect 20100 8527 20109 8533
rect 20057 8489 20109 8527
rect 20057 8481 20066 8489
rect 20066 8481 20100 8489
rect 20100 8481 20109 8489
rect 20057 8455 20066 8469
rect 20066 8455 20100 8469
rect 20100 8455 20109 8469
rect 20057 8417 20109 8455
rect 20057 8383 20066 8405
rect 20066 8383 20100 8405
rect 20100 8383 20109 8405
rect 18488 8350 18540 8359
rect 18132 8316 18147 8350
rect 18147 8316 18181 8350
rect 18181 8316 18184 8350
rect 18488 8316 18519 8350
rect 18519 8316 18540 8350
rect 18132 8307 18184 8316
rect 18488 8307 18540 8316
rect 18552 8350 18604 8359
rect 18552 8316 18557 8350
rect 18557 8316 18591 8350
rect 18591 8316 18604 8350
rect 18552 8307 18604 8316
rect 18616 8350 18668 8359
rect 18616 8316 18629 8350
rect 18629 8316 18663 8350
rect 18663 8316 18668 8350
rect 18616 8307 18668 8316
rect 18680 8350 18732 8359
rect 18744 8350 18796 8359
rect 18808 8350 18860 8359
rect 18872 8350 18924 8359
rect 18936 8350 18988 8359
rect 19000 8350 19052 8359
rect 19064 8350 19116 8359
rect 18680 8316 18701 8350
rect 18701 8316 18732 8350
rect 18744 8316 18773 8350
rect 18773 8316 18796 8350
rect 18808 8316 18845 8350
rect 18845 8316 18860 8350
rect 18872 8316 18879 8350
rect 18879 8316 18917 8350
rect 18917 8316 18924 8350
rect 18936 8316 18951 8350
rect 18951 8316 18988 8350
rect 19000 8316 19023 8350
rect 19023 8316 19052 8350
rect 19064 8316 19095 8350
rect 19095 8316 19116 8350
rect 18680 8307 18732 8316
rect 18744 8307 18796 8316
rect 18808 8307 18860 8316
rect 18872 8307 18924 8316
rect 18936 8307 18988 8316
rect 19000 8307 19052 8316
rect 19064 8307 19116 8316
rect 19128 8350 19180 8359
rect 19342 8350 19394 8359
rect 19128 8316 19133 8350
rect 19133 8316 19167 8350
rect 19167 8316 19180 8350
rect 19342 8316 19349 8350
rect 19349 8316 19383 8350
rect 19383 8316 19394 8350
rect 19128 8307 19180 8316
rect 19342 8307 19394 8316
rect 19406 8350 19458 8359
rect 19406 8316 19421 8350
rect 19421 8316 19455 8350
rect 19455 8316 19458 8350
rect 19406 8307 19458 8316
rect 19470 8350 19522 8359
rect 19534 8350 19586 8359
rect 19598 8350 19650 8359
rect 19662 8350 19714 8359
rect 19726 8350 19778 8359
rect 19790 8350 19842 8359
rect 19854 8350 19906 8359
rect 19470 8316 19493 8350
rect 19493 8316 19522 8350
rect 19534 8316 19565 8350
rect 19565 8316 19586 8350
rect 19598 8316 19599 8350
rect 19599 8316 19637 8350
rect 19637 8316 19650 8350
rect 19662 8316 19671 8350
rect 19671 8316 19709 8350
rect 19709 8316 19714 8350
rect 19726 8316 19743 8350
rect 19743 8316 19778 8350
rect 19790 8316 19815 8350
rect 19815 8316 19842 8350
rect 19854 8316 19887 8350
rect 19887 8316 19906 8350
rect 19470 8307 19522 8316
rect 19534 8307 19586 8316
rect 19598 8307 19650 8316
rect 19662 8307 19714 8316
rect 19726 8307 19778 8316
rect 19790 8307 19842 8316
rect 19854 8307 19906 8316
rect 19918 8350 19970 8359
rect 19918 8316 19925 8350
rect 19925 8316 19959 8350
rect 19959 8316 19970 8350
rect 19918 8307 19970 8316
rect 19982 8350 20034 8359
rect 20057 8353 20109 8383
rect 19982 8316 19997 8350
rect 19997 8316 20031 8350
rect 20031 8316 20034 8350
rect 19982 8307 20034 8316
rect 16510 8120 17260 8220
rect 15960 8000 16060 8110
rect 15960 7966 15990 8000
rect 15990 7966 16024 8000
rect 16024 7966 16060 8000
rect 15960 7920 16060 7966
rect 15960 7886 15990 7920
rect 15990 7886 16024 7920
rect 16024 7886 16060 7920
rect 15960 7840 16060 7886
rect 15960 7806 15990 7840
rect 15990 7806 16024 7840
rect 16024 7806 16060 7840
rect 15960 7760 16060 7806
rect 15960 7726 15990 7760
rect 15990 7726 16024 7760
rect 16024 7726 16060 7760
rect 15960 7680 16060 7726
rect 15960 7646 15990 7680
rect 15990 7646 16024 7680
rect 16024 7646 16060 7680
rect 15960 7600 16060 7646
rect 15960 7566 15990 7600
rect 15990 7566 16024 7600
rect 16024 7566 16060 7600
rect 15960 7520 16060 7566
rect 15960 7486 15990 7520
rect 15990 7486 16024 7520
rect 16024 7486 16060 7520
rect 15960 7440 16060 7486
rect 15960 7406 15990 7440
rect 15990 7406 16024 7440
rect 16024 7406 16060 7440
rect 15960 7360 16060 7406
rect 15960 7326 15990 7360
rect 15990 7326 16024 7360
rect 16024 7326 16060 7360
rect 15960 7280 16060 7326
rect 15960 7246 15990 7280
rect 15990 7246 16024 7280
rect 16024 7246 16060 7280
rect 15960 7200 16060 7246
rect 15960 7166 15990 7200
rect 15990 7166 16024 7200
rect 16024 7166 16060 7200
rect 15960 7120 16060 7166
rect 15960 7086 15990 7120
rect 15990 7086 16024 7120
rect 16024 7086 16060 7120
rect 15960 7040 16060 7086
rect 15960 7006 15990 7040
rect 15990 7006 16024 7040
rect 16024 7006 16060 7040
rect 15960 7000 16060 7006
rect 16195 7887 16247 7901
rect 16195 7853 16204 7887
rect 16204 7853 16238 7887
rect 16238 7853 16247 7887
rect 16195 7849 16247 7853
rect 16195 7815 16247 7821
rect 16195 7781 16204 7815
rect 16204 7781 16238 7815
rect 16238 7781 16247 7815
rect 16195 7769 16247 7781
rect 16195 7709 16204 7741
rect 16204 7709 16238 7741
rect 16238 7709 16247 7741
rect 16195 7689 16247 7709
rect 16195 7637 16204 7661
rect 16204 7637 16238 7661
rect 16238 7637 16247 7661
rect 16195 7609 16247 7637
rect 16195 7565 16204 7581
rect 16204 7565 16238 7581
rect 16238 7565 16247 7581
rect 16195 7529 16247 7565
rect 16195 7493 16204 7501
rect 16204 7493 16238 7501
rect 16238 7493 16247 7501
rect 16195 7455 16247 7493
rect 16195 7449 16204 7455
rect 16204 7449 16238 7455
rect 16238 7449 16247 7455
rect 16195 7383 16247 7421
rect 16195 7369 16204 7383
rect 16204 7369 16238 7383
rect 16238 7369 16247 7383
rect 16195 7311 16247 7341
rect 16195 7289 16204 7311
rect 16204 7289 16238 7311
rect 16238 7289 16247 7311
rect 16195 7239 16247 7261
rect 16195 7209 16204 7239
rect 16204 7209 16238 7239
rect 16238 7209 16247 7239
rect 16195 7167 16247 7181
rect 16195 7133 16204 7167
rect 16204 7133 16238 7167
rect 16238 7133 16247 7167
rect 16195 7129 16247 7133
rect 16195 7095 16247 7101
rect 16195 7061 16204 7095
rect 16204 7061 16238 7095
rect 16238 7061 16247 7095
rect 16195 7049 16247 7061
rect 16367 7887 16419 7901
rect 16367 7853 16376 7887
rect 16376 7853 16410 7887
rect 16410 7853 16419 7887
rect 16367 7849 16419 7853
rect 16367 7815 16419 7821
rect 16367 7781 16376 7815
rect 16376 7781 16410 7815
rect 16410 7781 16419 7815
rect 16367 7769 16419 7781
rect 16367 7709 16376 7741
rect 16376 7709 16410 7741
rect 16410 7709 16419 7741
rect 16367 7689 16419 7709
rect 16367 7637 16376 7661
rect 16376 7637 16410 7661
rect 16410 7637 16419 7661
rect 16367 7609 16419 7637
rect 16367 7565 16376 7581
rect 16376 7565 16410 7581
rect 16410 7565 16419 7581
rect 16367 7529 16419 7565
rect 16367 7493 16376 7501
rect 16376 7493 16410 7501
rect 16410 7493 16419 7501
rect 16367 7455 16419 7493
rect 16367 7449 16376 7455
rect 16376 7449 16410 7455
rect 16410 7449 16419 7455
rect 16367 7383 16419 7421
rect 16367 7369 16376 7383
rect 16376 7369 16410 7383
rect 16410 7369 16419 7383
rect 16367 7311 16419 7341
rect 16367 7289 16376 7311
rect 16376 7289 16410 7311
rect 16410 7289 16419 7311
rect 16367 7239 16419 7261
rect 16367 7209 16376 7239
rect 16376 7209 16410 7239
rect 16410 7209 16419 7239
rect 16367 7167 16419 7181
rect 16367 7133 16376 7167
rect 16376 7133 16410 7167
rect 16410 7133 16419 7167
rect 16367 7129 16419 7133
rect 16367 7095 16419 7101
rect 16367 7061 16376 7095
rect 16376 7061 16410 7095
rect 16410 7061 16419 7095
rect 16367 7049 16419 7061
rect 16539 7887 16591 7901
rect 16539 7853 16548 7887
rect 16548 7853 16582 7887
rect 16582 7853 16591 7887
rect 16539 7849 16591 7853
rect 16539 7815 16591 7821
rect 16539 7781 16548 7815
rect 16548 7781 16582 7815
rect 16582 7781 16591 7815
rect 16539 7769 16591 7781
rect 16539 7709 16548 7741
rect 16548 7709 16582 7741
rect 16582 7709 16591 7741
rect 16539 7689 16591 7709
rect 16539 7637 16548 7661
rect 16548 7637 16582 7661
rect 16582 7637 16591 7661
rect 16539 7609 16591 7637
rect 16539 7565 16548 7581
rect 16548 7565 16582 7581
rect 16582 7565 16591 7581
rect 16539 7529 16591 7565
rect 16539 7493 16548 7501
rect 16548 7493 16582 7501
rect 16582 7493 16591 7501
rect 16539 7455 16591 7493
rect 16539 7449 16548 7455
rect 16548 7449 16582 7455
rect 16582 7449 16591 7455
rect 16539 7383 16591 7421
rect 16539 7369 16548 7383
rect 16548 7369 16582 7383
rect 16582 7369 16591 7383
rect 16539 7311 16591 7341
rect 16539 7289 16548 7311
rect 16548 7289 16582 7311
rect 16582 7289 16591 7311
rect 16539 7239 16591 7261
rect 16539 7209 16548 7239
rect 16548 7209 16582 7239
rect 16582 7209 16591 7239
rect 16539 7167 16591 7181
rect 16539 7133 16548 7167
rect 16548 7133 16582 7167
rect 16582 7133 16591 7167
rect 16539 7129 16591 7133
rect 16539 7095 16591 7101
rect 16539 7061 16548 7095
rect 16548 7061 16582 7095
rect 16582 7061 16591 7095
rect 16539 7049 16591 7061
rect 16711 7887 16763 7901
rect 16711 7853 16720 7887
rect 16720 7853 16754 7887
rect 16754 7853 16763 7887
rect 16711 7849 16763 7853
rect 16711 7815 16763 7821
rect 16711 7781 16720 7815
rect 16720 7781 16754 7815
rect 16754 7781 16763 7815
rect 16711 7769 16763 7781
rect 16711 7709 16720 7741
rect 16720 7709 16754 7741
rect 16754 7709 16763 7741
rect 16711 7689 16763 7709
rect 16711 7637 16720 7661
rect 16720 7637 16754 7661
rect 16754 7637 16763 7661
rect 16711 7609 16763 7637
rect 16711 7565 16720 7581
rect 16720 7565 16754 7581
rect 16754 7565 16763 7581
rect 16711 7529 16763 7565
rect 16711 7493 16720 7501
rect 16720 7493 16754 7501
rect 16754 7493 16763 7501
rect 16711 7455 16763 7493
rect 16711 7449 16720 7455
rect 16720 7449 16754 7455
rect 16754 7449 16763 7455
rect 16711 7383 16763 7421
rect 16711 7369 16720 7383
rect 16720 7369 16754 7383
rect 16754 7369 16763 7383
rect 16711 7311 16763 7341
rect 16711 7289 16720 7311
rect 16720 7289 16754 7311
rect 16754 7289 16763 7311
rect 16711 7239 16763 7261
rect 16711 7209 16720 7239
rect 16720 7209 16754 7239
rect 16754 7209 16763 7239
rect 16711 7167 16763 7181
rect 16711 7133 16720 7167
rect 16720 7133 16754 7167
rect 16754 7133 16763 7167
rect 16711 7129 16763 7133
rect 16711 7095 16763 7101
rect 16711 7061 16720 7095
rect 16720 7061 16754 7095
rect 16754 7061 16763 7095
rect 16711 7049 16763 7061
rect 16883 7887 16935 7901
rect 16883 7853 16892 7887
rect 16892 7853 16926 7887
rect 16926 7853 16935 7887
rect 16883 7849 16935 7853
rect 16883 7815 16935 7821
rect 16883 7781 16892 7815
rect 16892 7781 16926 7815
rect 16926 7781 16935 7815
rect 16883 7769 16935 7781
rect 16883 7709 16892 7741
rect 16892 7709 16926 7741
rect 16926 7709 16935 7741
rect 16883 7689 16935 7709
rect 16883 7637 16892 7661
rect 16892 7637 16926 7661
rect 16926 7637 16935 7661
rect 16883 7609 16935 7637
rect 16883 7565 16892 7581
rect 16892 7565 16926 7581
rect 16926 7565 16935 7581
rect 16883 7529 16935 7565
rect 16883 7493 16892 7501
rect 16892 7493 16926 7501
rect 16926 7493 16935 7501
rect 16883 7455 16935 7493
rect 16883 7449 16892 7455
rect 16892 7449 16926 7455
rect 16926 7449 16935 7455
rect 16883 7383 16935 7421
rect 16883 7369 16892 7383
rect 16892 7369 16926 7383
rect 16926 7369 16935 7383
rect 16883 7311 16935 7341
rect 16883 7289 16892 7311
rect 16892 7289 16926 7311
rect 16926 7289 16935 7311
rect 16883 7239 16935 7261
rect 16883 7209 16892 7239
rect 16892 7209 16926 7239
rect 16926 7209 16935 7239
rect 16883 7167 16935 7181
rect 16883 7133 16892 7167
rect 16892 7133 16926 7167
rect 16926 7133 16935 7167
rect 16883 7129 16935 7133
rect 16883 7095 16935 7101
rect 16883 7061 16892 7095
rect 16892 7061 16926 7095
rect 16926 7061 16935 7095
rect 16883 7049 16935 7061
rect 17420 8090 20140 8180
rect 17420 8080 17638 8090
rect 17638 8080 20058 8090
rect 20058 8080 20140 8090
rect 17055 7887 17107 7901
rect 17055 7853 17064 7887
rect 17064 7853 17098 7887
rect 17098 7853 17107 7887
rect 17055 7849 17107 7853
rect 17055 7815 17107 7821
rect 17055 7781 17064 7815
rect 17064 7781 17098 7815
rect 17098 7781 17107 7815
rect 17055 7769 17107 7781
rect 17055 7709 17064 7741
rect 17064 7709 17098 7741
rect 17098 7709 17107 7741
rect 17055 7689 17107 7709
rect 17055 7637 17064 7661
rect 17064 7637 17098 7661
rect 17098 7637 17107 7661
rect 17055 7609 17107 7637
rect 17055 7565 17064 7581
rect 17064 7565 17098 7581
rect 17098 7565 17107 7581
rect 17055 7529 17107 7565
rect 17055 7493 17064 7501
rect 17064 7493 17098 7501
rect 17098 7493 17107 7501
rect 17055 7455 17107 7493
rect 17055 7449 17064 7455
rect 17064 7449 17098 7455
rect 17098 7449 17107 7455
rect 17055 7383 17107 7421
rect 17055 7369 17064 7383
rect 17064 7369 17098 7383
rect 17098 7369 17107 7383
rect 17055 7311 17107 7341
rect 17055 7289 17064 7311
rect 17064 7289 17098 7311
rect 17098 7289 17107 7311
rect 17055 7239 17107 7261
rect 17055 7209 17064 7239
rect 17064 7209 17098 7239
rect 17098 7209 17107 7239
rect 17055 7167 17107 7181
rect 17055 7133 17064 7167
rect 17064 7133 17098 7167
rect 17098 7133 17107 7167
rect 17055 7129 17107 7133
rect 17055 7095 17107 7101
rect 17055 7061 17064 7095
rect 17064 7061 17098 7095
rect 17098 7061 17107 7095
rect 17055 7049 17107 7061
rect 17699 7082 17708 7099
rect 17708 7082 17742 7099
rect 17742 7082 17751 7099
rect 17699 7047 17751 7082
rect 17699 7010 17708 7035
rect 17708 7010 17742 7035
rect 17742 7010 17751 7035
rect 17699 6983 17751 7010
rect 17871 7082 17880 7099
rect 17880 7082 17914 7099
rect 17914 7082 17923 7099
rect 17871 7047 17923 7082
rect 17871 7010 17880 7035
rect 17880 7010 17914 7035
rect 17914 7010 17923 7035
rect 17871 6983 17923 7010
rect 18043 7082 18052 7099
rect 18052 7082 18086 7099
rect 18086 7082 18095 7099
rect 18043 7047 18095 7082
rect 18043 7010 18052 7035
rect 18052 7010 18086 7035
rect 18086 7010 18095 7035
rect 18043 6983 18095 7010
rect 18215 7082 18224 7099
rect 18224 7082 18258 7099
rect 18258 7082 18267 7099
rect 18215 7047 18267 7082
rect 18215 7010 18224 7035
rect 18224 7010 18258 7035
rect 18258 7010 18267 7035
rect 18215 6983 18267 7010
rect 18387 7082 18396 7099
rect 18396 7082 18430 7099
rect 18430 7082 18439 7099
rect 18387 7047 18439 7082
rect 18387 7010 18396 7035
rect 18396 7010 18430 7035
rect 18430 7010 18439 7035
rect 18387 6983 18439 7010
rect 18559 7082 18568 7099
rect 18568 7082 18602 7099
rect 18602 7082 18611 7099
rect 18559 7047 18611 7082
rect 18559 7010 18568 7035
rect 18568 7010 18602 7035
rect 18602 7010 18611 7035
rect 18559 6983 18611 7010
rect 18731 7082 18740 7099
rect 18740 7082 18774 7099
rect 18774 7082 18783 7099
rect 18731 7047 18783 7082
rect 18731 7010 18740 7035
rect 18740 7010 18774 7035
rect 18774 7010 18783 7035
rect 18731 6983 18783 7010
rect 18903 7082 18912 7099
rect 18912 7082 18946 7099
rect 18946 7082 18955 7099
rect 18903 7047 18955 7082
rect 18903 7010 18912 7035
rect 18912 7010 18946 7035
rect 18946 7010 18955 7035
rect 18903 6983 18955 7010
rect 19075 7082 19084 7099
rect 19084 7082 19118 7099
rect 19118 7082 19127 7099
rect 19075 7047 19127 7082
rect 19075 7010 19084 7035
rect 19084 7010 19118 7035
rect 19118 7010 19127 7035
rect 19075 6983 19127 7010
rect 19247 7082 19256 7099
rect 19256 7082 19290 7099
rect 19290 7082 19299 7099
rect 19247 7047 19299 7082
rect 19247 7010 19256 7035
rect 19256 7010 19290 7035
rect 19290 7010 19299 7035
rect 19247 6983 19299 7010
rect 19419 7082 19428 7099
rect 19428 7082 19462 7099
rect 19462 7082 19471 7099
rect 19419 7047 19471 7082
rect 19419 7010 19428 7035
rect 19428 7010 19462 7035
rect 19462 7010 19471 7035
rect 19419 6983 19471 7010
rect 19591 7082 19600 7099
rect 19600 7082 19634 7099
rect 19634 7082 19643 7099
rect 19591 7047 19643 7082
rect 19591 7010 19600 7035
rect 19600 7010 19634 7035
rect 19634 7010 19643 7035
rect 19591 6983 19643 7010
rect 19763 7082 19772 7099
rect 19772 7082 19806 7099
rect 19806 7082 19815 7099
rect 19763 7047 19815 7082
rect 19763 7010 19772 7035
rect 19772 7010 19806 7035
rect 19806 7010 19815 7035
rect 19763 6983 19815 7010
rect 19935 7082 19944 7099
rect 19944 7082 19978 7099
rect 19978 7082 19987 7099
rect 19935 7047 19987 7082
rect 19935 7010 19944 7035
rect 19944 7010 19978 7035
rect 19978 7010 19987 7035
rect 19935 6983 19987 7010
rect 20060 7908 20138 7930
rect 20060 7874 20064 7908
rect 20064 7874 20138 7908
rect 20060 7836 20138 7874
rect 20060 7802 20064 7836
rect 20064 7802 20138 7836
rect 20060 7764 20138 7802
rect 20060 7730 20064 7764
rect 20064 7730 20138 7764
rect 20060 7692 20138 7730
rect 20060 7658 20064 7692
rect 20064 7658 20138 7692
rect 20060 7620 20138 7658
rect 20060 7586 20064 7620
rect 20064 7586 20138 7620
rect 20060 7548 20138 7586
rect 20060 7514 20064 7548
rect 20064 7514 20138 7548
rect 20060 7476 20138 7514
rect 20060 7442 20064 7476
rect 20064 7442 20138 7476
rect 20060 7404 20138 7442
rect 20060 7370 20064 7404
rect 20064 7370 20138 7404
rect 20060 7332 20138 7370
rect 20060 7298 20064 7332
rect 20064 7298 20138 7332
rect 20060 7260 20138 7298
rect 20060 7226 20064 7260
rect 20064 7226 20138 7260
rect 20060 7188 20138 7226
rect 20060 7154 20064 7188
rect 20064 7154 20138 7188
rect 20060 7116 20138 7154
rect 20060 7082 20064 7116
rect 20064 7082 20138 7116
rect 20060 7044 20138 7082
rect 20060 7010 20064 7044
rect 20064 7010 20138 7044
rect 20060 7000 20138 7010
rect 20138 7000 20178 7930
rect 20178 7000 20180 7930
rect 11776 6838 11828 6844
rect 11776 6804 11785 6838
rect 11785 6804 11819 6838
rect 11819 6804 11828 6838
rect 11776 6792 11828 6804
rect 11776 6766 11828 6780
rect 11776 6732 11785 6766
rect 11785 6732 11819 6766
rect 11819 6732 11828 6766
rect 11776 6728 11828 6732
rect 11776 6694 11828 6716
rect 11776 6664 11785 6694
rect 11785 6664 11819 6694
rect 11819 6664 11828 6694
rect 11776 6622 11828 6652
rect 11776 6600 11785 6622
rect 11785 6600 11819 6622
rect 11819 6600 11828 6622
rect 11776 6550 11828 6588
rect 11776 6536 11785 6550
rect 11785 6536 11819 6550
rect 11819 6536 11828 6550
rect 11776 6516 11785 6524
rect 11785 6516 11819 6524
rect 11819 6516 11828 6524
rect 11776 6478 11828 6516
rect 11776 6472 11785 6478
rect 11785 6472 11819 6478
rect 11819 6472 11828 6478
rect 11776 6444 11785 6460
rect 11785 6444 11819 6460
rect 11819 6444 11828 6460
rect 11776 6408 11828 6444
rect 11776 6372 11785 6396
rect 11785 6372 11819 6396
rect 11819 6372 11828 6396
rect 11776 6344 11828 6372
rect 11776 6300 11785 6332
rect 11785 6300 11819 6332
rect 11819 6300 11828 6332
rect 11776 6280 11828 6300
rect 11776 6262 11828 6268
rect 11776 6228 11785 6262
rect 11785 6228 11819 6262
rect 11819 6228 11828 6262
rect 11776 6216 11828 6228
rect 11776 6190 11828 6204
rect 11776 6156 11785 6190
rect 11785 6156 11819 6190
rect 11819 6156 11828 6190
rect 11776 6152 11828 6156
rect 11776 6118 11828 6140
rect 11776 6088 11785 6118
rect 11785 6088 11819 6118
rect 11819 6088 11828 6118
rect 11776 6046 11828 6076
rect 11776 6024 11785 6046
rect 11785 6024 11819 6046
rect 11819 6024 11828 6046
rect 11776 5974 11828 6012
rect 11776 5960 11785 5974
rect 11785 5960 11819 5974
rect 11819 5960 11828 5974
rect 11776 5940 11785 5948
rect 11785 5940 11819 5948
rect 11819 5940 11828 5948
rect 11776 5902 11828 5940
rect 11776 5896 11785 5902
rect 11785 5896 11819 5902
rect 11819 5896 11828 5902
rect 11862 6804 11871 6810
rect 11871 6804 11905 6810
rect 11905 6804 11914 6810
rect 11862 6766 11914 6804
rect 11862 6758 11871 6766
rect 11871 6758 11905 6766
rect 11905 6758 11914 6766
rect 11862 6732 11871 6746
rect 11871 6732 11905 6746
rect 11905 6732 11914 6746
rect 11862 6694 11914 6732
rect 11862 6660 11871 6682
rect 11871 6660 11905 6682
rect 11905 6660 11914 6682
rect 11862 6630 11914 6660
rect 11862 6588 11871 6618
rect 11871 6588 11905 6618
rect 11905 6588 11914 6618
rect 11862 6566 11914 6588
rect 11862 6550 11914 6554
rect 11862 6516 11871 6550
rect 11871 6516 11905 6550
rect 11905 6516 11914 6550
rect 11862 6502 11914 6516
rect 11862 6478 11914 6490
rect 11862 6444 11871 6478
rect 11871 6444 11905 6478
rect 11905 6444 11914 6478
rect 11862 6438 11914 6444
rect 11862 6406 11914 6426
rect 11862 6374 11871 6406
rect 11871 6374 11905 6406
rect 11905 6374 11914 6406
rect 11862 6334 11914 6362
rect 11862 6310 11871 6334
rect 11871 6310 11905 6334
rect 11905 6310 11914 6334
rect 11862 6262 11914 6298
rect 11862 6246 11871 6262
rect 11871 6246 11905 6262
rect 11905 6246 11914 6262
rect 11862 6228 11871 6234
rect 11871 6228 11905 6234
rect 11905 6228 11914 6234
rect 11862 6190 11914 6228
rect 11862 6182 11871 6190
rect 11871 6182 11905 6190
rect 11905 6182 11914 6190
rect 11862 6156 11871 6170
rect 11871 6156 11905 6170
rect 11905 6156 11914 6170
rect 11862 6118 11914 6156
rect 11862 6084 11871 6106
rect 11871 6084 11905 6106
rect 11905 6084 11914 6106
rect 11862 6054 11914 6084
rect 11862 6012 11871 6042
rect 11871 6012 11905 6042
rect 11905 6012 11914 6042
rect 11862 5990 11914 6012
rect 11862 5974 11914 5978
rect 11862 5940 11871 5974
rect 11871 5940 11905 5974
rect 11905 5940 11914 5974
rect 11862 5926 11914 5940
rect 11862 5902 11914 5914
rect 11862 5868 11871 5902
rect 11871 5868 11905 5902
rect 11905 5868 11914 5902
rect 11862 5862 11914 5868
rect 11948 6838 12000 6844
rect 11948 6804 11957 6838
rect 11957 6804 11991 6838
rect 11991 6804 12000 6838
rect 11948 6792 12000 6804
rect 11948 6766 12000 6780
rect 11948 6732 11957 6766
rect 11957 6732 11991 6766
rect 11991 6732 12000 6766
rect 11948 6728 12000 6732
rect 11948 6694 12000 6716
rect 11948 6664 11957 6694
rect 11957 6664 11991 6694
rect 11991 6664 12000 6694
rect 11948 6622 12000 6652
rect 11948 6600 11957 6622
rect 11957 6600 11991 6622
rect 11991 6600 12000 6622
rect 11948 6550 12000 6588
rect 11948 6536 11957 6550
rect 11957 6536 11991 6550
rect 11991 6536 12000 6550
rect 11948 6516 11957 6524
rect 11957 6516 11991 6524
rect 11991 6516 12000 6524
rect 11948 6478 12000 6516
rect 11948 6472 11957 6478
rect 11957 6472 11991 6478
rect 11991 6472 12000 6478
rect 11948 6444 11957 6460
rect 11957 6444 11991 6460
rect 11991 6444 12000 6460
rect 11948 6408 12000 6444
rect 11948 6372 11957 6396
rect 11957 6372 11991 6396
rect 11991 6372 12000 6396
rect 11948 6344 12000 6372
rect 11948 6300 11957 6332
rect 11957 6300 11991 6332
rect 11991 6300 12000 6332
rect 11948 6280 12000 6300
rect 11948 6262 12000 6268
rect 11948 6228 11957 6262
rect 11957 6228 11991 6262
rect 11991 6228 12000 6262
rect 11948 6216 12000 6228
rect 11948 6190 12000 6204
rect 11948 6156 11957 6190
rect 11957 6156 11991 6190
rect 11991 6156 12000 6190
rect 11948 6152 12000 6156
rect 11948 6118 12000 6140
rect 11948 6088 11957 6118
rect 11957 6088 11991 6118
rect 11991 6088 12000 6118
rect 11948 6046 12000 6076
rect 11948 6024 11957 6046
rect 11957 6024 11991 6046
rect 11991 6024 12000 6046
rect 11948 5974 12000 6012
rect 11948 5960 11957 5974
rect 11957 5960 11991 5974
rect 11991 5960 12000 5974
rect 11948 5940 11957 5948
rect 11957 5940 11991 5948
rect 11991 5940 12000 5948
rect 11948 5902 12000 5940
rect 11948 5896 11957 5902
rect 11957 5896 11991 5902
rect 11991 5896 12000 5902
rect 12034 6804 12043 6810
rect 12043 6804 12077 6810
rect 12077 6804 12086 6810
rect 12034 6766 12086 6804
rect 12034 6758 12043 6766
rect 12043 6758 12077 6766
rect 12077 6758 12086 6766
rect 12034 6732 12043 6746
rect 12043 6732 12077 6746
rect 12077 6732 12086 6746
rect 12034 6694 12086 6732
rect 12034 6660 12043 6682
rect 12043 6660 12077 6682
rect 12077 6660 12086 6682
rect 12034 6630 12086 6660
rect 12034 6588 12043 6618
rect 12043 6588 12077 6618
rect 12077 6588 12086 6618
rect 12034 6566 12086 6588
rect 12034 6550 12086 6554
rect 12034 6516 12043 6550
rect 12043 6516 12077 6550
rect 12077 6516 12086 6550
rect 12034 6502 12086 6516
rect 12034 6478 12086 6490
rect 12034 6444 12043 6478
rect 12043 6444 12077 6478
rect 12077 6444 12086 6478
rect 12034 6438 12086 6444
rect 12034 6406 12086 6426
rect 12034 6374 12043 6406
rect 12043 6374 12077 6406
rect 12077 6374 12086 6406
rect 12034 6334 12086 6362
rect 12034 6310 12043 6334
rect 12043 6310 12077 6334
rect 12077 6310 12086 6334
rect 12034 6262 12086 6298
rect 12034 6246 12043 6262
rect 12043 6246 12077 6262
rect 12077 6246 12086 6262
rect 12034 6228 12043 6234
rect 12043 6228 12077 6234
rect 12077 6228 12086 6234
rect 12034 6190 12086 6228
rect 12034 6182 12043 6190
rect 12043 6182 12077 6190
rect 12077 6182 12086 6190
rect 12034 6156 12043 6170
rect 12043 6156 12077 6170
rect 12077 6156 12086 6170
rect 12034 6118 12086 6156
rect 12034 6084 12043 6106
rect 12043 6084 12077 6106
rect 12077 6084 12086 6106
rect 12034 6054 12086 6084
rect 12034 6012 12043 6042
rect 12043 6012 12077 6042
rect 12077 6012 12086 6042
rect 12034 5990 12086 6012
rect 12034 5974 12086 5978
rect 12034 5940 12043 5974
rect 12043 5940 12077 5974
rect 12077 5940 12086 5974
rect 12034 5926 12086 5940
rect 12034 5902 12086 5914
rect 12034 5868 12043 5902
rect 12043 5868 12077 5902
rect 12077 5868 12086 5902
rect 12034 5862 12086 5868
rect 12120 6838 12172 6844
rect 12120 6804 12129 6838
rect 12129 6804 12163 6838
rect 12163 6804 12172 6838
rect 12120 6792 12172 6804
rect 12120 6766 12172 6780
rect 12120 6732 12129 6766
rect 12129 6732 12163 6766
rect 12163 6732 12172 6766
rect 12120 6728 12172 6732
rect 12120 6694 12172 6716
rect 12120 6664 12129 6694
rect 12129 6664 12163 6694
rect 12163 6664 12172 6694
rect 12120 6622 12172 6652
rect 12120 6600 12129 6622
rect 12129 6600 12163 6622
rect 12163 6600 12172 6622
rect 12120 6550 12172 6588
rect 12120 6536 12129 6550
rect 12129 6536 12163 6550
rect 12163 6536 12172 6550
rect 12120 6516 12129 6524
rect 12129 6516 12163 6524
rect 12163 6516 12172 6524
rect 12120 6478 12172 6516
rect 12120 6472 12129 6478
rect 12129 6472 12163 6478
rect 12163 6472 12172 6478
rect 12120 6444 12129 6460
rect 12129 6444 12163 6460
rect 12163 6444 12172 6460
rect 12120 6408 12172 6444
rect 12120 6372 12129 6396
rect 12129 6372 12163 6396
rect 12163 6372 12172 6396
rect 12120 6344 12172 6372
rect 12120 6300 12129 6332
rect 12129 6300 12163 6332
rect 12163 6300 12172 6332
rect 12120 6280 12172 6300
rect 12120 6262 12172 6268
rect 12120 6228 12129 6262
rect 12129 6228 12163 6262
rect 12163 6228 12172 6262
rect 12120 6216 12172 6228
rect 12120 6190 12172 6204
rect 12120 6156 12129 6190
rect 12129 6156 12163 6190
rect 12163 6156 12172 6190
rect 12120 6152 12172 6156
rect 12120 6118 12172 6140
rect 12120 6088 12129 6118
rect 12129 6088 12163 6118
rect 12163 6088 12172 6118
rect 12120 6046 12172 6076
rect 12120 6024 12129 6046
rect 12129 6024 12163 6046
rect 12163 6024 12172 6046
rect 12120 5974 12172 6012
rect 12120 5960 12129 5974
rect 12129 5960 12163 5974
rect 12163 5960 12172 5974
rect 12120 5940 12129 5948
rect 12129 5940 12163 5948
rect 12163 5940 12172 5948
rect 12120 5902 12172 5940
rect 12120 5896 12129 5902
rect 12129 5896 12163 5902
rect 12163 5896 12172 5902
rect 11860 5510 12100 5570
rect 12342 6838 12394 6844
rect 12342 6804 12351 6838
rect 12351 6804 12385 6838
rect 12385 6804 12394 6838
rect 12342 6792 12394 6804
rect 12342 6766 12394 6780
rect 12342 6732 12351 6766
rect 12351 6732 12385 6766
rect 12385 6732 12394 6766
rect 12342 6728 12394 6732
rect 12342 6694 12394 6716
rect 12342 6664 12351 6694
rect 12351 6664 12385 6694
rect 12385 6664 12394 6694
rect 12342 6622 12394 6652
rect 12342 6600 12351 6622
rect 12351 6600 12385 6622
rect 12385 6600 12394 6622
rect 12342 6550 12394 6588
rect 12342 6536 12351 6550
rect 12351 6536 12385 6550
rect 12385 6536 12394 6550
rect 12342 6516 12351 6524
rect 12351 6516 12385 6524
rect 12385 6516 12394 6524
rect 12342 6478 12394 6516
rect 12342 6472 12351 6478
rect 12351 6472 12385 6478
rect 12385 6472 12394 6478
rect 12342 6444 12351 6460
rect 12351 6444 12385 6460
rect 12385 6444 12394 6460
rect 12342 6408 12394 6444
rect 12342 6372 12351 6396
rect 12351 6372 12385 6396
rect 12385 6372 12394 6396
rect 12342 6344 12394 6372
rect 12342 6300 12351 6332
rect 12351 6300 12385 6332
rect 12385 6300 12394 6332
rect 12342 6280 12394 6300
rect 12342 6262 12394 6268
rect 12342 6228 12351 6262
rect 12351 6228 12385 6262
rect 12385 6228 12394 6262
rect 12342 6216 12394 6228
rect 12342 6190 12394 6204
rect 12342 6156 12351 6190
rect 12351 6156 12385 6190
rect 12385 6156 12394 6190
rect 12342 6152 12394 6156
rect 12342 6118 12394 6140
rect 12342 6088 12351 6118
rect 12351 6088 12385 6118
rect 12385 6088 12394 6118
rect 12342 6046 12394 6076
rect 12342 6024 12351 6046
rect 12351 6024 12385 6046
rect 12385 6024 12394 6046
rect 12342 5974 12394 6012
rect 12342 5960 12351 5974
rect 12351 5960 12385 5974
rect 12385 5960 12394 5974
rect 12342 5940 12351 5948
rect 12351 5940 12385 5948
rect 12385 5940 12394 5948
rect 12342 5902 12394 5940
rect 12342 5896 12351 5902
rect 12351 5896 12385 5902
rect 12385 5896 12394 5902
rect 12428 6804 12437 6810
rect 12437 6804 12471 6810
rect 12471 6804 12480 6810
rect 12428 6766 12480 6804
rect 12428 6758 12437 6766
rect 12437 6758 12471 6766
rect 12471 6758 12480 6766
rect 12428 6732 12437 6746
rect 12437 6732 12471 6746
rect 12471 6732 12480 6746
rect 12428 6694 12480 6732
rect 12428 6660 12437 6682
rect 12437 6660 12471 6682
rect 12471 6660 12480 6682
rect 12428 6630 12480 6660
rect 12428 6588 12437 6618
rect 12437 6588 12471 6618
rect 12471 6588 12480 6618
rect 12428 6566 12480 6588
rect 12428 6550 12480 6554
rect 12428 6516 12437 6550
rect 12437 6516 12471 6550
rect 12471 6516 12480 6550
rect 12428 6502 12480 6516
rect 12428 6478 12480 6490
rect 12428 6444 12437 6478
rect 12437 6444 12471 6478
rect 12471 6444 12480 6478
rect 12428 6438 12480 6444
rect 12428 6406 12480 6426
rect 12428 6374 12437 6406
rect 12437 6374 12471 6406
rect 12471 6374 12480 6406
rect 12428 6334 12480 6362
rect 12428 6310 12437 6334
rect 12437 6310 12471 6334
rect 12471 6310 12480 6334
rect 12428 6262 12480 6298
rect 12428 6246 12437 6262
rect 12437 6246 12471 6262
rect 12471 6246 12480 6262
rect 12428 6228 12437 6234
rect 12437 6228 12471 6234
rect 12471 6228 12480 6234
rect 12428 6190 12480 6228
rect 12428 6182 12437 6190
rect 12437 6182 12471 6190
rect 12471 6182 12480 6190
rect 12428 6156 12437 6170
rect 12437 6156 12471 6170
rect 12471 6156 12480 6170
rect 12428 6118 12480 6156
rect 12428 6084 12437 6106
rect 12437 6084 12471 6106
rect 12471 6084 12480 6106
rect 12428 6054 12480 6084
rect 12428 6012 12437 6042
rect 12437 6012 12471 6042
rect 12471 6012 12480 6042
rect 12428 5990 12480 6012
rect 12428 5974 12480 5978
rect 12428 5940 12437 5974
rect 12437 5940 12471 5974
rect 12471 5940 12480 5974
rect 12428 5926 12480 5940
rect 12428 5902 12480 5914
rect 12428 5868 12437 5902
rect 12437 5868 12471 5902
rect 12471 5868 12480 5902
rect 12428 5862 12480 5868
rect 12514 6838 12566 6844
rect 12514 6804 12523 6838
rect 12523 6804 12557 6838
rect 12557 6804 12566 6838
rect 12514 6792 12566 6804
rect 12514 6766 12566 6780
rect 12514 6732 12523 6766
rect 12523 6732 12557 6766
rect 12557 6732 12566 6766
rect 12514 6728 12566 6732
rect 12514 6694 12566 6716
rect 12514 6664 12523 6694
rect 12523 6664 12557 6694
rect 12557 6664 12566 6694
rect 12514 6622 12566 6652
rect 12514 6600 12523 6622
rect 12523 6600 12557 6622
rect 12557 6600 12566 6622
rect 12514 6550 12566 6588
rect 12514 6536 12523 6550
rect 12523 6536 12557 6550
rect 12557 6536 12566 6550
rect 12514 6516 12523 6524
rect 12523 6516 12557 6524
rect 12557 6516 12566 6524
rect 12514 6478 12566 6516
rect 12514 6472 12523 6478
rect 12523 6472 12557 6478
rect 12557 6472 12566 6478
rect 12514 6444 12523 6460
rect 12523 6444 12557 6460
rect 12557 6444 12566 6460
rect 12514 6408 12566 6444
rect 12514 6372 12523 6396
rect 12523 6372 12557 6396
rect 12557 6372 12566 6396
rect 12514 6344 12566 6372
rect 12514 6300 12523 6332
rect 12523 6300 12557 6332
rect 12557 6300 12566 6332
rect 12514 6280 12566 6300
rect 12514 6262 12566 6268
rect 12514 6228 12523 6262
rect 12523 6228 12557 6262
rect 12557 6228 12566 6262
rect 12514 6216 12566 6228
rect 12514 6190 12566 6204
rect 12514 6156 12523 6190
rect 12523 6156 12557 6190
rect 12557 6156 12566 6190
rect 12514 6152 12566 6156
rect 12514 6118 12566 6140
rect 12514 6088 12523 6118
rect 12523 6088 12557 6118
rect 12557 6088 12566 6118
rect 12514 6046 12566 6076
rect 12514 6024 12523 6046
rect 12523 6024 12557 6046
rect 12557 6024 12566 6046
rect 12514 5974 12566 6012
rect 12514 5960 12523 5974
rect 12523 5960 12557 5974
rect 12557 5960 12566 5974
rect 12514 5940 12523 5948
rect 12523 5940 12557 5948
rect 12557 5940 12566 5948
rect 12514 5902 12566 5940
rect 12514 5896 12523 5902
rect 12523 5896 12557 5902
rect 12557 5896 12566 5902
rect 12600 6804 12609 6810
rect 12609 6804 12643 6810
rect 12643 6804 12652 6810
rect 12600 6766 12652 6804
rect 12600 6758 12609 6766
rect 12609 6758 12643 6766
rect 12643 6758 12652 6766
rect 12600 6732 12609 6746
rect 12609 6732 12643 6746
rect 12643 6732 12652 6746
rect 12600 6694 12652 6732
rect 12600 6660 12609 6682
rect 12609 6660 12643 6682
rect 12643 6660 12652 6682
rect 12600 6630 12652 6660
rect 12600 6588 12609 6618
rect 12609 6588 12643 6618
rect 12643 6588 12652 6618
rect 12600 6566 12652 6588
rect 12600 6550 12652 6554
rect 12600 6516 12609 6550
rect 12609 6516 12643 6550
rect 12643 6516 12652 6550
rect 12600 6502 12652 6516
rect 12600 6478 12652 6490
rect 12600 6444 12609 6478
rect 12609 6444 12643 6478
rect 12643 6444 12652 6478
rect 12600 6438 12652 6444
rect 12600 6406 12652 6426
rect 12600 6374 12609 6406
rect 12609 6374 12643 6406
rect 12643 6374 12652 6406
rect 12600 6334 12652 6362
rect 12600 6310 12609 6334
rect 12609 6310 12643 6334
rect 12643 6310 12652 6334
rect 12600 6262 12652 6298
rect 12600 6246 12609 6262
rect 12609 6246 12643 6262
rect 12643 6246 12652 6262
rect 12600 6228 12609 6234
rect 12609 6228 12643 6234
rect 12643 6228 12652 6234
rect 12600 6190 12652 6228
rect 12600 6182 12609 6190
rect 12609 6182 12643 6190
rect 12643 6182 12652 6190
rect 12600 6156 12609 6170
rect 12609 6156 12643 6170
rect 12643 6156 12652 6170
rect 12600 6118 12652 6156
rect 12600 6084 12609 6106
rect 12609 6084 12643 6106
rect 12643 6084 12652 6106
rect 12600 6054 12652 6084
rect 12600 6012 12609 6042
rect 12609 6012 12643 6042
rect 12643 6012 12652 6042
rect 12600 5990 12652 6012
rect 12600 5974 12652 5978
rect 12600 5940 12609 5974
rect 12609 5940 12643 5974
rect 12643 5940 12652 5974
rect 12600 5926 12652 5940
rect 12600 5902 12652 5914
rect 12600 5868 12609 5902
rect 12609 5868 12643 5902
rect 12643 5868 12652 5902
rect 12600 5862 12652 5868
rect 12686 6838 12738 6844
rect 12686 6804 12695 6838
rect 12695 6804 12729 6838
rect 12729 6804 12738 6838
rect 12686 6792 12738 6804
rect 12686 6766 12738 6780
rect 12686 6732 12695 6766
rect 12695 6732 12729 6766
rect 12729 6732 12738 6766
rect 12686 6728 12738 6732
rect 12686 6694 12738 6716
rect 12686 6664 12695 6694
rect 12695 6664 12729 6694
rect 12729 6664 12738 6694
rect 12686 6622 12738 6652
rect 12686 6600 12695 6622
rect 12695 6600 12729 6622
rect 12729 6600 12738 6622
rect 12686 6550 12738 6588
rect 12686 6536 12695 6550
rect 12695 6536 12729 6550
rect 12729 6536 12738 6550
rect 12686 6516 12695 6524
rect 12695 6516 12729 6524
rect 12729 6516 12738 6524
rect 12686 6478 12738 6516
rect 12686 6472 12695 6478
rect 12695 6472 12729 6478
rect 12729 6472 12738 6478
rect 12686 6444 12695 6460
rect 12695 6444 12729 6460
rect 12729 6444 12738 6460
rect 12686 6408 12738 6444
rect 12686 6372 12695 6396
rect 12695 6372 12729 6396
rect 12729 6372 12738 6396
rect 12686 6344 12738 6372
rect 12686 6300 12695 6332
rect 12695 6300 12729 6332
rect 12729 6300 12738 6332
rect 12686 6280 12738 6300
rect 12686 6262 12738 6268
rect 12686 6228 12695 6262
rect 12695 6228 12729 6262
rect 12729 6228 12738 6262
rect 12686 6216 12738 6228
rect 12686 6190 12738 6204
rect 12686 6156 12695 6190
rect 12695 6156 12729 6190
rect 12729 6156 12738 6190
rect 12686 6152 12738 6156
rect 12686 6118 12738 6140
rect 12686 6088 12695 6118
rect 12695 6088 12729 6118
rect 12729 6088 12738 6118
rect 12686 6046 12738 6076
rect 12686 6024 12695 6046
rect 12695 6024 12729 6046
rect 12729 6024 12738 6046
rect 12686 5974 12738 6012
rect 12686 5960 12695 5974
rect 12695 5960 12729 5974
rect 12729 5960 12738 5974
rect 12686 5940 12695 5948
rect 12695 5940 12729 5948
rect 12729 5940 12738 5948
rect 12686 5902 12738 5940
rect 12686 5896 12695 5902
rect 12695 5896 12729 5902
rect 12729 5896 12738 5902
rect 12420 5510 12660 5570
rect 12908 6838 12960 6844
rect 12908 6804 12917 6838
rect 12917 6804 12951 6838
rect 12951 6804 12960 6838
rect 12908 6792 12960 6804
rect 12908 6766 12960 6780
rect 12908 6732 12917 6766
rect 12917 6732 12951 6766
rect 12951 6732 12960 6766
rect 12908 6728 12960 6732
rect 12908 6694 12960 6716
rect 12908 6664 12917 6694
rect 12917 6664 12951 6694
rect 12951 6664 12960 6694
rect 12908 6622 12960 6652
rect 12908 6600 12917 6622
rect 12917 6600 12951 6622
rect 12951 6600 12960 6622
rect 12908 6550 12960 6588
rect 12908 6536 12917 6550
rect 12917 6536 12951 6550
rect 12951 6536 12960 6550
rect 12908 6516 12917 6524
rect 12917 6516 12951 6524
rect 12951 6516 12960 6524
rect 12908 6478 12960 6516
rect 12908 6472 12917 6478
rect 12917 6472 12951 6478
rect 12951 6472 12960 6478
rect 12908 6444 12917 6460
rect 12917 6444 12951 6460
rect 12951 6444 12960 6460
rect 12908 6408 12960 6444
rect 12908 6372 12917 6396
rect 12917 6372 12951 6396
rect 12951 6372 12960 6396
rect 12908 6344 12960 6372
rect 12908 6300 12917 6332
rect 12917 6300 12951 6332
rect 12951 6300 12960 6332
rect 12908 6280 12960 6300
rect 12908 6262 12960 6268
rect 12908 6228 12917 6262
rect 12917 6228 12951 6262
rect 12951 6228 12960 6262
rect 12908 6216 12960 6228
rect 12908 6190 12960 6204
rect 12908 6156 12917 6190
rect 12917 6156 12951 6190
rect 12951 6156 12960 6190
rect 12908 6152 12960 6156
rect 12908 6118 12960 6140
rect 12908 6088 12917 6118
rect 12917 6088 12951 6118
rect 12951 6088 12960 6118
rect 12908 6046 12960 6076
rect 12908 6024 12917 6046
rect 12917 6024 12951 6046
rect 12951 6024 12960 6046
rect 12908 5974 12960 6012
rect 12908 5960 12917 5974
rect 12917 5960 12951 5974
rect 12951 5960 12960 5974
rect 12908 5940 12917 5948
rect 12917 5940 12951 5948
rect 12951 5940 12960 5948
rect 12908 5902 12960 5940
rect 12908 5896 12917 5902
rect 12917 5896 12951 5902
rect 12951 5896 12960 5902
rect 12994 6804 13003 6810
rect 13003 6804 13037 6810
rect 13037 6804 13046 6810
rect 12994 6766 13046 6804
rect 12994 6758 13003 6766
rect 13003 6758 13037 6766
rect 13037 6758 13046 6766
rect 12994 6732 13003 6746
rect 13003 6732 13037 6746
rect 13037 6732 13046 6746
rect 12994 6694 13046 6732
rect 12994 6660 13003 6682
rect 13003 6660 13037 6682
rect 13037 6660 13046 6682
rect 12994 6630 13046 6660
rect 12994 6588 13003 6618
rect 13003 6588 13037 6618
rect 13037 6588 13046 6618
rect 12994 6566 13046 6588
rect 12994 6550 13046 6554
rect 12994 6516 13003 6550
rect 13003 6516 13037 6550
rect 13037 6516 13046 6550
rect 12994 6502 13046 6516
rect 12994 6478 13046 6490
rect 12994 6444 13003 6478
rect 13003 6444 13037 6478
rect 13037 6444 13046 6478
rect 12994 6438 13046 6444
rect 12994 6406 13046 6426
rect 12994 6374 13003 6406
rect 13003 6374 13037 6406
rect 13037 6374 13046 6406
rect 12994 6334 13046 6362
rect 12994 6310 13003 6334
rect 13003 6310 13037 6334
rect 13037 6310 13046 6334
rect 12994 6262 13046 6298
rect 12994 6246 13003 6262
rect 13003 6246 13037 6262
rect 13037 6246 13046 6262
rect 12994 6228 13003 6234
rect 13003 6228 13037 6234
rect 13037 6228 13046 6234
rect 12994 6190 13046 6228
rect 12994 6182 13003 6190
rect 13003 6182 13037 6190
rect 13037 6182 13046 6190
rect 12994 6156 13003 6170
rect 13003 6156 13037 6170
rect 13037 6156 13046 6170
rect 12994 6118 13046 6156
rect 12994 6084 13003 6106
rect 13003 6084 13037 6106
rect 13037 6084 13046 6106
rect 12994 6054 13046 6084
rect 12994 6012 13003 6042
rect 13003 6012 13037 6042
rect 13037 6012 13046 6042
rect 12994 5990 13046 6012
rect 12994 5974 13046 5978
rect 12994 5940 13003 5974
rect 13003 5940 13037 5974
rect 13037 5940 13046 5974
rect 12994 5926 13046 5940
rect 12994 5902 13046 5914
rect 12994 5868 13003 5902
rect 13003 5868 13037 5902
rect 13037 5868 13046 5902
rect 12994 5862 13046 5868
rect 13080 6838 13132 6844
rect 13080 6804 13089 6838
rect 13089 6804 13123 6838
rect 13123 6804 13132 6838
rect 13080 6792 13132 6804
rect 13080 6766 13132 6780
rect 13080 6732 13089 6766
rect 13089 6732 13123 6766
rect 13123 6732 13132 6766
rect 13080 6728 13132 6732
rect 13080 6694 13132 6716
rect 13080 6664 13089 6694
rect 13089 6664 13123 6694
rect 13123 6664 13132 6694
rect 13080 6622 13132 6652
rect 13080 6600 13089 6622
rect 13089 6600 13123 6622
rect 13123 6600 13132 6622
rect 13080 6550 13132 6588
rect 13080 6536 13089 6550
rect 13089 6536 13123 6550
rect 13123 6536 13132 6550
rect 13080 6516 13089 6524
rect 13089 6516 13123 6524
rect 13123 6516 13132 6524
rect 13080 6478 13132 6516
rect 13080 6472 13089 6478
rect 13089 6472 13123 6478
rect 13123 6472 13132 6478
rect 13080 6444 13089 6460
rect 13089 6444 13123 6460
rect 13123 6444 13132 6460
rect 13080 6408 13132 6444
rect 13080 6372 13089 6396
rect 13089 6372 13123 6396
rect 13123 6372 13132 6396
rect 13080 6344 13132 6372
rect 13080 6300 13089 6332
rect 13089 6300 13123 6332
rect 13123 6300 13132 6332
rect 13080 6280 13132 6300
rect 13080 6262 13132 6268
rect 13080 6228 13089 6262
rect 13089 6228 13123 6262
rect 13123 6228 13132 6262
rect 13080 6216 13132 6228
rect 13080 6190 13132 6204
rect 13080 6156 13089 6190
rect 13089 6156 13123 6190
rect 13123 6156 13132 6190
rect 13080 6152 13132 6156
rect 13080 6118 13132 6140
rect 13080 6088 13089 6118
rect 13089 6088 13123 6118
rect 13123 6088 13132 6118
rect 13080 6046 13132 6076
rect 13080 6024 13089 6046
rect 13089 6024 13123 6046
rect 13123 6024 13132 6046
rect 13080 5974 13132 6012
rect 13080 5960 13089 5974
rect 13089 5960 13123 5974
rect 13123 5960 13132 5974
rect 13080 5940 13089 5948
rect 13089 5940 13123 5948
rect 13123 5940 13132 5948
rect 13080 5902 13132 5940
rect 13080 5896 13089 5902
rect 13089 5896 13123 5902
rect 13123 5896 13132 5902
rect 13166 6804 13175 6810
rect 13175 6804 13209 6810
rect 13209 6804 13218 6810
rect 13166 6766 13218 6804
rect 13166 6758 13175 6766
rect 13175 6758 13209 6766
rect 13209 6758 13218 6766
rect 13166 6732 13175 6746
rect 13175 6732 13209 6746
rect 13209 6732 13218 6746
rect 13166 6694 13218 6732
rect 13166 6660 13175 6682
rect 13175 6660 13209 6682
rect 13209 6660 13218 6682
rect 13166 6630 13218 6660
rect 13166 6588 13175 6618
rect 13175 6588 13209 6618
rect 13209 6588 13218 6618
rect 13166 6566 13218 6588
rect 13166 6550 13218 6554
rect 13166 6516 13175 6550
rect 13175 6516 13209 6550
rect 13209 6516 13218 6550
rect 13166 6502 13218 6516
rect 13166 6478 13218 6490
rect 13166 6444 13175 6478
rect 13175 6444 13209 6478
rect 13209 6444 13218 6478
rect 13166 6438 13218 6444
rect 13166 6406 13218 6426
rect 13166 6374 13175 6406
rect 13175 6374 13209 6406
rect 13209 6374 13218 6406
rect 13166 6334 13218 6362
rect 13166 6310 13175 6334
rect 13175 6310 13209 6334
rect 13209 6310 13218 6334
rect 13166 6262 13218 6298
rect 13166 6246 13175 6262
rect 13175 6246 13209 6262
rect 13209 6246 13218 6262
rect 13166 6228 13175 6234
rect 13175 6228 13209 6234
rect 13209 6228 13218 6234
rect 13166 6190 13218 6228
rect 13166 6182 13175 6190
rect 13175 6182 13209 6190
rect 13209 6182 13218 6190
rect 13166 6156 13175 6170
rect 13175 6156 13209 6170
rect 13209 6156 13218 6170
rect 13166 6118 13218 6156
rect 13166 6084 13175 6106
rect 13175 6084 13209 6106
rect 13209 6084 13218 6106
rect 13166 6054 13218 6084
rect 13166 6012 13175 6042
rect 13175 6012 13209 6042
rect 13209 6012 13218 6042
rect 13166 5990 13218 6012
rect 13166 5974 13218 5978
rect 13166 5940 13175 5974
rect 13175 5940 13209 5974
rect 13209 5940 13218 5974
rect 13166 5926 13218 5940
rect 13166 5902 13218 5914
rect 13166 5868 13175 5902
rect 13175 5868 13209 5902
rect 13209 5868 13218 5902
rect 13166 5862 13218 5868
rect 13252 6838 13304 6844
rect 13252 6804 13261 6838
rect 13261 6804 13295 6838
rect 13295 6804 13304 6838
rect 13252 6792 13304 6804
rect 13252 6766 13304 6780
rect 13252 6732 13261 6766
rect 13261 6732 13295 6766
rect 13295 6732 13304 6766
rect 13252 6728 13304 6732
rect 13252 6694 13304 6716
rect 13252 6664 13261 6694
rect 13261 6664 13295 6694
rect 13295 6664 13304 6694
rect 13252 6622 13304 6652
rect 13252 6600 13261 6622
rect 13261 6600 13295 6622
rect 13295 6600 13304 6622
rect 13252 6550 13304 6588
rect 13252 6536 13261 6550
rect 13261 6536 13295 6550
rect 13295 6536 13304 6550
rect 13252 6516 13261 6524
rect 13261 6516 13295 6524
rect 13295 6516 13304 6524
rect 13252 6478 13304 6516
rect 13252 6472 13261 6478
rect 13261 6472 13295 6478
rect 13295 6472 13304 6478
rect 13252 6444 13261 6460
rect 13261 6444 13295 6460
rect 13295 6444 13304 6460
rect 13252 6408 13304 6444
rect 13252 6372 13261 6396
rect 13261 6372 13295 6396
rect 13295 6372 13304 6396
rect 13252 6344 13304 6372
rect 13252 6300 13261 6332
rect 13261 6300 13295 6332
rect 13295 6300 13304 6332
rect 13252 6280 13304 6300
rect 13252 6262 13304 6268
rect 13252 6228 13261 6262
rect 13261 6228 13295 6262
rect 13295 6228 13304 6262
rect 13252 6216 13304 6228
rect 13252 6190 13304 6204
rect 13252 6156 13261 6190
rect 13261 6156 13295 6190
rect 13295 6156 13304 6190
rect 13252 6152 13304 6156
rect 13252 6118 13304 6140
rect 13252 6088 13261 6118
rect 13261 6088 13295 6118
rect 13295 6088 13304 6118
rect 13252 6046 13304 6076
rect 13252 6024 13261 6046
rect 13261 6024 13295 6046
rect 13295 6024 13304 6046
rect 13252 5974 13304 6012
rect 13252 5960 13261 5974
rect 13261 5960 13295 5974
rect 13295 5960 13304 5974
rect 13252 5940 13261 5948
rect 13261 5940 13295 5948
rect 13295 5940 13304 5948
rect 13252 5902 13304 5940
rect 13252 5896 13261 5902
rect 13261 5896 13295 5902
rect 13295 5896 13304 5902
rect 12980 5510 13220 5570
rect 13474 6838 13526 6844
rect 13474 6804 13483 6838
rect 13483 6804 13517 6838
rect 13517 6804 13526 6838
rect 13474 6792 13526 6804
rect 13474 6766 13526 6780
rect 13474 6732 13483 6766
rect 13483 6732 13517 6766
rect 13517 6732 13526 6766
rect 13474 6728 13526 6732
rect 13474 6694 13526 6716
rect 13474 6664 13483 6694
rect 13483 6664 13517 6694
rect 13517 6664 13526 6694
rect 13474 6622 13526 6652
rect 13474 6600 13483 6622
rect 13483 6600 13517 6622
rect 13517 6600 13526 6622
rect 13474 6550 13526 6588
rect 13474 6536 13483 6550
rect 13483 6536 13517 6550
rect 13517 6536 13526 6550
rect 13474 6516 13483 6524
rect 13483 6516 13517 6524
rect 13517 6516 13526 6524
rect 13474 6478 13526 6516
rect 13474 6472 13483 6478
rect 13483 6472 13517 6478
rect 13517 6472 13526 6478
rect 13474 6444 13483 6460
rect 13483 6444 13517 6460
rect 13517 6444 13526 6460
rect 13474 6408 13526 6444
rect 13474 6372 13483 6396
rect 13483 6372 13517 6396
rect 13517 6372 13526 6396
rect 13474 6344 13526 6372
rect 13474 6300 13483 6332
rect 13483 6300 13517 6332
rect 13517 6300 13526 6332
rect 13474 6280 13526 6300
rect 13474 6262 13526 6268
rect 13474 6228 13483 6262
rect 13483 6228 13517 6262
rect 13517 6228 13526 6262
rect 13474 6216 13526 6228
rect 13474 6190 13526 6204
rect 13474 6156 13483 6190
rect 13483 6156 13517 6190
rect 13517 6156 13526 6190
rect 13474 6152 13526 6156
rect 13474 6118 13526 6140
rect 13474 6088 13483 6118
rect 13483 6088 13517 6118
rect 13517 6088 13526 6118
rect 13474 6046 13526 6076
rect 13474 6024 13483 6046
rect 13483 6024 13517 6046
rect 13517 6024 13526 6046
rect 13474 5974 13526 6012
rect 13474 5960 13483 5974
rect 13483 5960 13517 5974
rect 13517 5960 13526 5974
rect 13474 5940 13483 5948
rect 13483 5940 13517 5948
rect 13517 5940 13526 5948
rect 13474 5902 13526 5940
rect 13474 5896 13483 5902
rect 13483 5896 13517 5902
rect 13517 5896 13526 5902
rect 13560 6804 13569 6810
rect 13569 6804 13603 6810
rect 13603 6804 13612 6810
rect 13560 6766 13612 6804
rect 13560 6758 13569 6766
rect 13569 6758 13603 6766
rect 13603 6758 13612 6766
rect 13560 6732 13569 6746
rect 13569 6732 13603 6746
rect 13603 6732 13612 6746
rect 13560 6694 13612 6732
rect 13560 6660 13569 6682
rect 13569 6660 13603 6682
rect 13603 6660 13612 6682
rect 13560 6630 13612 6660
rect 13560 6588 13569 6618
rect 13569 6588 13603 6618
rect 13603 6588 13612 6618
rect 13560 6566 13612 6588
rect 13560 6550 13612 6554
rect 13560 6516 13569 6550
rect 13569 6516 13603 6550
rect 13603 6516 13612 6550
rect 13560 6502 13612 6516
rect 13560 6478 13612 6490
rect 13560 6444 13569 6478
rect 13569 6444 13603 6478
rect 13603 6444 13612 6478
rect 13560 6438 13612 6444
rect 13560 6406 13612 6426
rect 13560 6374 13569 6406
rect 13569 6374 13603 6406
rect 13603 6374 13612 6406
rect 13560 6334 13612 6362
rect 13560 6310 13569 6334
rect 13569 6310 13603 6334
rect 13603 6310 13612 6334
rect 13560 6262 13612 6298
rect 13560 6246 13569 6262
rect 13569 6246 13603 6262
rect 13603 6246 13612 6262
rect 13560 6228 13569 6234
rect 13569 6228 13603 6234
rect 13603 6228 13612 6234
rect 13560 6190 13612 6228
rect 13560 6182 13569 6190
rect 13569 6182 13603 6190
rect 13603 6182 13612 6190
rect 13560 6156 13569 6170
rect 13569 6156 13603 6170
rect 13603 6156 13612 6170
rect 13560 6118 13612 6156
rect 13560 6084 13569 6106
rect 13569 6084 13603 6106
rect 13603 6084 13612 6106
rect 13560 6054 13612 6084
rect 13560 6012 13569 6042
rect 13569 6012 13603 6042
rect 13603 6012 13612 6042
rect 13560 5990 13612 6012
rect 13560 5974 13612 5978
rect 13560 5940 13569 5974
rect 13569 5940 13603 5974
rect 13603 5940 13612 5974
rect 13560 5926 13612 5940
rect 13560 5902 13612 5914
rect 13560 5868 13569 5902
rect 13569 5868 13603 5902
rect 13603 5868 13612 5902
rect 13560 5862 13612 5868
rect 13646 6838 13698 6844
rect 13646 6804 13655 6838
rect 13655 6804 13689 6838
rect 13689 6804 13698 6838
rect 13646 6792 13698 6804
rect 13646 6766 13698 6780
rect 13646 6732 13655 6766
rect 13655 6732 13689 6766
rect 13689 6732 13698 6766
rect 13646 6728 13698 6732
rect 13646 6694 13698 6716
rect 13646 6664 13655 6694
rect 13655 6664 13689 6694
rect 13689 6664 13698 6694
rect 13646 6622 13698 6652
rect 13646 6600 13655 6622
rect 13655 6600 13689 6622
rect 13689 6600 13698 6622
rect 13646 6550 13698 6588
rect 13646 6536 13655 6550
rect 13655 6536 13689 6550
rect 13689 6536 13698 6550
rect 13646 6516 13655 6524
rect 13655 6516 13689 6524
rect 13689 6516 13698 6524
rect 13646 6478 13698 6516
rect 13646 6472 13655 6478
rect 13655 6472 13689 6478
rect 13689 6472 13698 6478
rect 13646 6444 13655 6460
rect 13655 6444 13689 6460
rect 13689 6444 13698 6460
rect 13646 6408 13698 6444
rect 13646 6372 13655 6396
rect 13655 6372 13689 6396
rect 13689 6372 13698 6396
rect 13646 6344 13698 6372
rect 13646 6300 13655 6332
rect 13655 6300 13689 6332
rect 13689 6300 13698 6332
rect 13646 6280 13698 6300
rect 13646 6262 13698 6268
rect 13646 6228 13655 6262
rect 13655 6228 13689 6262
rect 13689 6228 13698 6262
rect 13646 6216 13698 6228
rect 13646 6190 13698 6204
rect 13646 6156 13655 6190
rect 13655 6156 13689 6190
rect 13689 6156 13698 6190
rect 13646 6152 13698 6156
rect 13646 6118 13698 6140
rect 13646 6088 13655 6118
rect 13655 6088 13689 6118
rect 13689 6088 13698 6118
rect 13646 6046 13698 6076
rect 13646 6024 13655 6046
rect 13655 6024 13689 6046
rect 13689 6024 13698 6046
rect 13646 5974 13698 6012
rect 13646 5960 13655 5974
rect 13655 5960 13689 5974
rect 13689 5960 13698 5974
rect 13646 5940 13655 5948
rect 13655 5940 13689 5948
rect 13689 5940 13698 5948
rect 13646 5902 13698 5940
rect 13646 5896 13655 5902
rect 13655 5896 13689 5902
rect 13689 5896 13698 5902
rect 13732 6804 13741 6810
rect 13741 6804 13775 6810
rect 13775 6804 13784 6810
rect 13732 6766 13784 6804
rect 13732 6758 13741 6766
rect 13741 6758 13775 6766
rect 13775 6758 13784 6766
rect 13732 6732 13741 6746
rect 13741 6732 13775 6746
rect 13775 6732 13784 6746
rect 13732 6694 13784 6732
rect 13732 6660 13741 6682
rect 13741 6660 13775 6682
rect 13775 6660 13784 6682
rect 13732 6630 13784 6660
rect 13732 6588 13741 6618
rect 13741 6588 13775 6618
rect 13775 6588 13784 6618
rect 13732 6566 13784 6588
rect 13732 6550 13784 6554
rect 13732 6516 13741 6550
rect 13741 6516 13775 6550
rect 13775 6516 13784 6550
rect 13732 6502 13784 6516
rect 13732 6478 13784 6490
rect 13732 6444 13741 6478
rect 13741 6444 13775 6478
rect 13775 6444 13784 6478
rect 13732 6438 13784 6444
rect 13732 6406 13784 6426
rect 13732 6374 13741 6406
rect 13741 6374 13775 6406
rect 13775 6374 13784 6406
rect 13732 6334 13784 6362
rect 13732 6310 13741 6334
rect 13741 6310 13775 6334
rect 13775 6310 13784 6334
rect 13732 6262 13784 6298
rect 13732 6246 13741 6262
rect 13741 6246 13775 6262
rect 13775 6246 13784 6262
rect 13732 6228 13741 6234
rect 13741 6228 13775 6234
rect 13775 6228 13784 6234
rect 13732 6190 13784 6228
rect 13732 6182 13741 6190
rect 13741 6182 13775 6190
rect 13775 6182 13784 6190
rect 13732 6156 13741 6170
rect 13741 6156 13775 6170
rect 13775 6156 13784 6170
rect 13732 6118 13784 6156
rect 13732 6084 13741 6106
rect 13741 6084 13775 6106
rect 13775 6084 13784 6106
rect 13732 6054 13784 6084
rect 13732 6012 13741 6042
rect 13741 6012 13775 6042
rect 13775 6012 13784 6042
rect 13732 5990 13784 6012
rect 13732 5974 13784 5978
rect 13732 5940 13741 5974
rect 13741 5940 13775 5974
rect 13775 5940 13784 5974
rect 13732 5926 13784 5940
rect 13732 5902 13784 5914
rect 13732 5868 13741 5902
rect 13741 5868 13775 5902
rect 13775 5868 13784 5902
rect 13732 5862 13784 5868
rect 13818 6838 13870 6844
rect 13818 6804 13827 6838
rect 13827 6804 13861 6838
rect 13861 6804 13870 6838
rect 13818 6792 13870 6804
rect 13818 6766 13870 6780
rect 13818 6732 13827 6766
rect 13827 6732 13861 6766
rect 13861 6732 13870 6766
rect 13818 6728 13870 6732
rect 13818 6694 13870 6716
rect 13818 6664 13827 6694
rect 13827 6664 13861 6694
rect 13861 6664 13870 6694
rect 13818 6622 13870 6652
rect 13818 6600 13827 6622
rect 13827 6600 13861 6622
rect 13861 6600 13870 6622
rect 13818 6550 13870 6588
rect 13818 6536 13827 6550
rect 13827 6536 13861 6550
rect 13861 6536 13870 6550
rect 13818 6516 13827 6524
rect 13827 6516 13861 6524
rect 13861 6516 13870 6524
rect 13818 6478 13870 6516
rect 13818 6472 13827 6478
rect 13827 6472 13861 6478
rect 13861 6472 13870 6478
rect 13818 6444 13827 6460
rect 13827 6444 13861 6460
rect 13861 6444 13870 6460
rect 13818 6408 13870 6444
rect 13818 6372 13827 6396
rect 13827 6372 13861 6396
rect 13861 6372 13870 6396
rect 13818 6344 13870 6372
rect 13818 6300 13827 6332
rect 13827 6300 13861 6332
rect 13861 6300 13870 6332
rect 13818 6280 13870 6300
rect 13818 6262 13870 6268
rect 13818 6228 13827 6262
rect 13827 6228 13861 6262
rect 13861 6228 13870 6262
rect 13818 6216 13870 6228
rect 13818 6190 13870 6204
rect 13818 6156 13827 6190
rect 13827 6156 13861 6190
rect 13861 6156 13870 6190
rect 13818 6152 13870 6156
rect 13818 6118 13870 6140
rect 13818 6088 13827 6118
rect 13827 6088 13861 6118
rect 13861 6088 13870 6118
rect 13818 6046 13870 6076
rect 13818 6024 13827 6046
rect 13827 6024 13861 6046
rect 13861 6024 13870 6046
rect 13818 5974 13870 6012
rect 13818 5960 13827 5974
rect 13827 5960 13861 5974
rect 13861 5960 13870 5974
rect 13818 5940 13827 5948
rect 13827 5940 13861 5948
rect 13861 5940 13870 5948
rect 13818 5902 13870 5940
rect 13818 5896 13827 5902
rect 13827 5896 13861 5902
rect 13861 5896 13870 5902
rect 13560 5510 13800 5570
rect 14040 6838 14092 6844
rect 14040 6804 14049 6838
rect 14049 6804 14083 6838
rect 14083 6804 14092 6838
rect 14040 6792 14092 6804
rect 14040 6766 14092 6780
rect 14040 6732 14049 6766
rect 14049 6732 14083 6766
rect 14083 6732 14092 6766
rect 14040 6728 14092 6732
rect 14040 6694 14092 6716
rect 14040 6664 14049 6694
rect 14049 6664 14083 6694
rect 14083 6664 14092 6694
rect 14040 6622 14092 6652
rect 14040 6600 14049 6622
rect 14049 6600 14083 6622
rect 14083 6600 14092 6622
rect 14040 6550 14092 6588
rect 14040 6536 14049 6550
rect 14049 6536 14083 6550
rect 14083 6536 14092 6550
rect 14040 6516 14049 6524
rect 14049 6516 14083 6524
rect 14083 6516 14092 6524
rect 14040 6478 14092 6516
rect 14040 6472 14049 6478
rect 14049 6472 14083 6478
rect 14083 6472 14092 6478
rect 14040 6444 14049 6460
rect 14049 6444 14083 6460
rect 14083 6444 14092 6460
rect 14040 6408 14092 6444
rect 14040 6372 14049 6396
rect 14049 6372 14083 6396
rect 14083 6372 14092 6396
rect 14040 6344 14092 6372
rect 14040 6300 14049 6332
rect 14049 6300 14083 6332
rect 14083 6300 14092 6332
rect 14040 6280 14092 6300
rect 14040 6262 14092 6268
rect 14040 6228 14049 6262
rect 14049 6228 14083 6262
rect 14083 6228 14092 6262
rect 14040 6216 14092 6228
rect 14040 6190 14092 6204
rect 14040 6156 14049 6190
rect 14049 6156 14083 6190
rect 14083 6156 14092 6190
rect 14040 6152 14092 6156
rect 14040 6118 14092 6140
rect 14040 6088 14049 6118
rect 14049 6088 14083 6118
rect 14083 6088 14092 6118
rect 14040 6046 14092 6076
rect 14040 6024 14049 6046
rect 14049 6024 14083 6046
rect 14083 6024 14092 6046
rect 14040 5974 14092 6012
rect 14040 5960 14049 5974
rect 14049 5960 14083 5974
rect 14083 5960 14092 5974
rect 14040 5940 14049 5948
rect 14049 5940 14083 5948
rect 14083 5940 14092 5948
rect 14040 5902 14092 5940
rect 14040 5896 14049 5902
rect 14049 5896 14083 5902
rect 14083 5896 14092 5902
rect 14126 6804 14135 6810
rect 14135 6804 14169 6810
rect 14169 6804 14178 6810
rect 14126 6766 14178 6804
rect 14126 6758 14135 6766
rect 14135 6758 14169 6766
rect 14169 6758 14178 6766
rect 14126 6732 14135 6746
rect 14135 6732 14169 6746
rect 14169 6732 14178 6746
rect 14126 6694 14178 6732
rect 14126 6660 14135 6682
rect 14135 6660 14169 6682
rect 14169 6660 14178 6682
rect 14126 6630 14178 6660
rect 14126 6588 14135 6618
rect 14135 6588 14169 6618
rect 14169 6588 14178 6618
rect 14126 6566 14178 6588
rect 14126 6550 14178 6554
rect 14126 6516 14135 6550
rect 14135 6516 14169 6550
rect 14169 6516 14178 6550
rect 14126 6502 14178 6516
rect 14126 6478 14178 6490
rect 14126 6444 14135 6478
rect 14135 6444 14169 6478
rect 14169 6444 14178 6478
rect 14126 6438 14178 6444
rect 14126 6406 14178 6426
rect 14126 6374 14135 6406
rect 14135 6374 14169 6406
rect 14169 6374 14178 6406
rect 14126 6334 14178 6362
rect 14126 6310 14135 6334
rect 14135 6310 14169 6334
rect 14169 6310 14178 6334
rect 14126 6262 14178 6298
rect 14126 6246 14135 6262
rect 14135 6246 14169 6262
rect 14169 6246 14178 6262
rect 14126 6228 14135 6234
rect 14135 6228 14169 6234
rect 14169 6228 14178 6234
rect 14126 6190 14178 6228
rect 14126 6182 14135 6190
rect 14135 6182 14169 6190
rect 14169 6182 14178 6190
rect 14126 6156 14135 6170
rect 14135 6156 14169 6170
rect 14169 6156 14178 6170
rect 14126 6118 14178 6156
rect 14126 6084 14135 6106
rect 14135 6084 14169 6106
rect 14169 6084 14178 6106
rect 14126 6054 14178 6084
rect 14126 6012 14135 6042
rect 14135 6012 14169 6042
rect 14169 6012 14178 6042
rect 14126 5990 14178 6012
rect 14126 5974 14178 5978
rect 14126 5940 14135 5974
rect 14135 5940 14169 5974
rect 14169 5940 14178 5974
rect 14126 5926 14178 5940
rect 14126 5902 14178 5914
rect 14126 5868 14135 5902
rect 14135 5868 14169 5902
rect 14169 5868 14178 5902
rect 14126 5862 14178 5868
rect 14212 6838 14264 6844
rect 14212 6804 14221 6838
rect 14221 6804 14255 6838
rect 14255 6804 14264 6838
rect 14212 6792 14264 6804
rect 14212 6766 14264 6780
rect 14212 6732 14221 6766
rect 14221 6732 14255 6766
rect 14255 6732 14264 6766
rect 14212 6728 14264 6732
rect 14212 6694 14264 6716
rect 14212 6664 14221 6694
rect 14221 6664 14255 6694
rect 14255 6664 14264 6694
rect 14212 6622 14264 6652
rect 14212 6600 14221 6622
rect 14221 6600 14255 6622
rect 14255 6600 14264 6622
rect 14212 6550 14264 6588
rect 14212 6536 14221 6550
rect 14221 6536 14255 6550
rect 14255 6536 14264 6550
rect 14212 6516 14221 6524
rect 14221 6516 14255 6524
rect 14255 6516 14264 6524
rect 14212 6478 14264 6516
rect 14212 6472 14221 6478
rect 14221 6472 14255 6478
rect 14255 6472 14264 6478
rect 14212 6444 14221 6460
rect 14221 6444 14255 6460
rect 14255 6444 14264 6460
rect 14212 6408 14264 6444
rect 14212 6372 14221 6396
rect 14221 6372 14255 6396
rect 14255 6372 14264 6396
rect 14212 6344 14264 6372
rect 14212 6300 14221 6332
rect 14221 6300 14255 6332
rect 14255 6300 14264 6332
rect 14212 6280 14264 6300
rect 14212 6262 14264 6268
rect 14212 6228 14221 6262
rect 14221 6228 14255 6262
rect 14255 6228 14264 6262
rect 14212 6216 14264 6228
rect 14212 6190 14264 6204
rect 14212 6156 14221 6190
rect 14221 6156 14255 6190
rect 14255 6156 14264 6190
rect 14212 6152 14264 6156
rect 14212 6118 14264 6140
rect 14212 6088 14221 6118
rect 14221 6088 14255 6118
rect 14255 6088 14264 6118
rect 14212 6046 14264 6076
rect 14212 6024 14221 6046
rect 14221 6024 14255 6046
rect 14255 6024 14264 6046
rect 14212 5974 14264 6012
rect 14212 5960 14221 5974
rect 14221 5960 14255 5974
rect 14255 5960 14264 5974
rect 14212 5940 14221 5948
rect 14221 5940 14255 5948
rect 14255 5940 14264 5948
rect 14212 5902 14264 5940
rect 14212 5896 14221 5902
rect 14221 5896 14255 5902
rect 14255 5896 14264 5902
rect 14298 6804 14307 6810
rect 14307 6804 14341 6810
rect 14341 6804 14350 6810
rect 14298 6766 14350 6804
rect 14298 6758 14307 6766
rect 14307 6758 14341 6766
rect 14341 6758 14350 6766
rect 14298 6732 14307 6746
rect 14307 6732 14341 6746
rect 14341 6732 14350 6746
rect 14298 6694 14350 6732
rect 14298 6660 14307 6682
rect 14307 6660 14341 6682
rect 14341 6660 14350 6682
rect 14298 6630 14350 6660
rect 14298 6588 14307 6618
rect 14307 6588 14341 6618
rect 14341 6588 14350 6618
rect 14298 6566 14350 6588
rect 14298 6550 14350 6554
rect 14298 6516 14307 6550
rect 14307 6516 14341 6550
rect 14341 6516 14350 6550
rect 14298 6502 14350 6516
rect 14298 6478 14350 6490
rect 14298 6444 14307 6478
rect 14307 6444 14341 6478
rect 14341 6444 14350 6478
rect 14298 6438 14350 6444
rect 14298 6406 14350 6426
rect 14298 6374 14307 6406
rect 14307 6374 14341 6406
rect 14341 6374 14350 6406
rect 14298 6334 14350 6362
rect 14298 6310 14307 6334
rect 14307 6310 14341 6334
rect 14341 6310 14350 6334
rect 14298 6262 14350 6298
rect 14298 6246 14307 6262
rect 14307 6246 14341 6262
rect 14341 6246 14350 6262
rect 14298 6228 14307 6234
rect 14307 6228 14341 6234
rect 14341 6228 14350 6234
rect 14298 6190 14350 6228
rect 14298 6182 14307 6190
rect 14307 6182 14341 6190
rect 14341 6182 14350 6190
rect 14298 6156 14307 6170
rect 14307 6156 14341 6170
rect 14341 6156 14350 6170
rect 14298 6118 14350 6156
rect 14298 6084 14307 6106
rect 14307 6084 14341 6106
rect 14341 6084 14350 6106
rect 14298 6054 14350 6084
rect 14298 6012 14307 6042
rect 14307 6012 14341 6042
rect 14341 6012 14350 6042
rect 14298 5990 14350 6012
rect 14298 5974 14350 5978
rect 14298 5940 14307 5974
rect 14307 5940 14341 5974
rect 14341 5940 14350 5974
rect 14298 5926 14350 5940
rect 14298 5902 14350 5914
rect 14298 5868 14307 5902
rect 14307 5868 14341 5902
rect 14341 5868 14350 5902
rect 14298 5862 14350 5868
rect 14384 6838 14436 6844
rect 14384 6804 14393 6838
rect 14393 6804 14427 6838
rect 14427 6804 14436 6838
rect 14384 6792 14436 6804
rect 14384 6766 14436 6780
rect 14384 6732 14393 6766
rect 14393 6732 14427 6766
rect 14427 6732 14436 6766
rect 14384 6728 14436 6732
rect 14384 6694 14436 6716
rect 14384 6664 14393 6694
rect 14393 6664 14427 6694
rect 14427 6664 14436 6694
rect 14384 6622 14436 6652
rect 14384 6600 14393 6622
rect 14393 6600 14427 6622
rect 14427 6600 14436 6622
rect 14384 6550 14436 6588
rect 14384 6536 14393 6550
rect 14393 6536 14427 6550
rect 14427 6536 14436 6550
rect 14384 6516 14393 6524
rect 14393 6516 14427 6524
rect 14427 6516 14436 6524
rect 14384 6478 14436 6516
rect 14384 6472 14393 6478
rect 14393 6472 14427 6478
rect 14427 6472 14436 6478
rect 14384 6444 14393 6460
rect 14393 6444 14427 6460
rect 14427 6444 14436 6460
rect 14384 6408 14436 6444
rect 14384 6372 14393 6396
rect 14393 6372 14427 6396
rect 14427 6372 14436 6396
rect 14384 6344 14436 6372
rect 14384 6300 14393 6332
rect 14393 6300 14427 6332
rect 14427 6300 14436 6332
rect 14384 6280 14436 6300
rect 14384 6262 14436 6268
rect 14384 6228 14393 6262
rect 14393 6228 14427 6262
rect 14427 6228 14436 6262
rect 14384 6216 14436 6228
rect 14384 6190 14436 6204
rect 14384 6156 14393 6190
rect 14393 6156 14427 6190
rect 14427 6156 14436 6190
rect 14384 6152 14436 6156
rect 14384 6118 14436 6140
rect 14384 6088 14393 6118
rect 14393 6088 14427 6118
rect 14427 6088 14436 6118
rect 14384 6046 14436 6076
rect 14384 6024 14393 6046
rect 14393 6024 14427 6046
rect 14427 6024 14436 6046
rect 14384 5974 14436 6012
rect 14384 5960 14393 5974
rect 14393 5960 14427 5974
rect 14427 5960 14436 5974
rect 14384 5940 14393 5948
rect 14393 5940 14427 5948
rect 14427 5940 14436 5948
rect 14384 5902 14436 5940
rect 14384 5896 14393 5902
rect 14393 5896 14427 5902
rect 14427 5896 14436 5902
rect 14120 5510 14360 5570
rect 14606 6838 14658 6844
rect 14606 6804 14615 6838
rect 14615 6804 14649 6838
rect 14649 6804 14658 6838
rect 14606 6792 14658 6804
rect 14606 6766 14658 6780
rect 14606 6732 14615 6766
rect 14615 6732 14649 6766
rect 14649 6732 14658 6766
rect 14606 6728 14658 6732
rect 14606 6694 14658 6716
rect 14606 6664 14615 6694
rect 14615 6664 14649 6694
rect 14649 6664 14658 6694
rect 14606 6622 14658 6652
rect 14606 6600 14615 6622
rect 14615 6600 14649 6622
rect 14649 6600 14658 6622
rect 14606 6550 14658 6588
rect 14606 6536 14615 6550
rect 14615 6536 14649 6550
rect 14649 6536 14658 6550
rect 14606 6516 14615 6524
rect 14615 6516 14649 6524
rect 14649 6516 14658 6524
rect 14606 6478 14658 6516
rect 14606 6472 14615 6478
rect 14615 6472 14649 6478
rect 14649 6472 14658 6478
rect 14606 6444 14615 6460
rect 14615 6444 14649 6460
rect 14649 6444 14658 6460
rect 14606 6408 14658 6444
rect 14606 6372 14615 6396
rect 14615 6372 14649 6396
rect 14649 6372 14658 6396
rect 14606 6344 14658 6372
rect 14606 6300 14615 6332
rect 14615 6300 14649 6332
rect 14649 6300 14658 6332
rect 14606 6280 14658 6300
rect 14606 6262 14658 6268
rect 14606 6228 14615 6262
rect 14615 6228 14649 6262
rect 14649 6228 14658 6262
rect 14606 6216 14658 6228
rect 14606 6190 14658 6204
rect 14606 6156 14615 6190
rect 14615 6156 14649 6190
rect 14649 6156 14658 6190
rect 14606 6152 14658 6156
rect 14606 6118 14658 6140
rect 14606 6088 14615 6118
rect 14615 6088 14649 6118
rect 14649 6088 14658 6118
rect 14606 6046 14658 6076
rect 14606 6024 14615 6046
rect 14615 6024 14649 6046
rect 14649 6024 14658 6046
rect 14606 5974 14658 6012
rect 14606 5960 14615 5974
rect 14615 5960 14649 5974
rect 14649 5960 14658 5974
rect 14606 5940 14615 5948
rect 14615 5940 14649 5948
rect 14649 5940 14658 5948
rect 14606 5902 14658 5940
rect 14606 5896 14615 5902
rect 14615 5896 14649 5902
rect 14649 5896 14658 5902
rect 14692 6804 14701 6810
rect 14701 6804 14735 6810
rect 14735 6804 14744 6810
rect 14692 6766 14744 6804
rect 14692 6758 14701 6766
rect 14701 6758 14735 6766
rect 14735 6758 14744 6766
rect 14692 6732 14701 6746
rect 14701 6732 14735 6746
rect 14735 6732 14744 6746
rect 14692 6694 14744 6732
rect 14692 6660 14701 6682
rect 14701 6660 14735 6682
rect 14735 6660 14744 6682
rect 14692 6630 14744 6660
rect 14692 6588 14701 6618
rect 14701 6588 14735 6618
rect 14735 6588 14744 6618
rect 14692 6566 14744 6588
rect 14692 6550 14744 6554
rect 14692 6516 14701 6550
rect 14701 6516 14735 6550
rect 14735 6516 14744 6550
rect 14692 6502 14744 6516
rect 14692 6478 14744 6490
rect 14692 6444 14701 6478
rect 14701 6444 14735 6478
rect 14735 6444 14744 6478
rect 14692 6438 14744 6444
rect 14692 6406 14744 6426
rect 14692 6374 14701 6406
rect 14701 6374 14735 6406
rect 14735 6374 14744 6406
rect 14692 6334 14744 6362
rect 14692 6310 14701 6334
rect 14701 6310 14735 6334
rect 14735 6310 14744 6334
rect 14692 6262 14744 6298
rect 14692 6246 14701 6262
rect 14701 6246 14735 6262
rect 14735 6246 14744 6262
rect 14692 6228 14701 6234
rect 14701 6228 14735 6234
rect 14735 6228 14744 6234
rect 14692 6190 14744 6228
rect 14692 6182 14701 6190
rect 14701 6182 14735 6190
rect 14735 6182 14744 6190
rect 14692 6156 14701 6170
rect 14701 6156 14735 6170
rect 14735 6156 14744 6170
rect 14692 6118 14744 6156
rect 14692 6084 14701 6106
rect 14701 6084 14735 6106
rect 14735 6084 14744 6106
rect 14692 6054 14744 6084
rect 14692 6012 14701 6042
rect 14701 6012 14735 6042
rect 14735 6012 14744 6042
rect 14692 5990 14744 6012
rect 14692 5974 14744 5978
rect 14692 5940 14701 5974
rect 14701 5940 14735 5974
rect 14735 5940 14744 5974
rect 14692 5926 14744 5940
rect 14692 5902 14744 5914
rect 14692 5868 14701 5902
rect 14701 5868 14735 5902
rect 14735 5868 14744 5902
rect 14692 5862 14744 5868
rect 14778 6838 14830 6844
rect 14778 6804 14787 6838
rect 14787 6804 14821 6838
rect 14821 6804 14830 6838
rect 14778 6792 14830 6804
rect 14778 6766 14830 6780
rect 14778 6732 14787 6766
rect 14787 6732 14821 6766
rect 14821 6732 14830 6766
rect 14778 6728 14830 6732
rect 14778 6694 14830 6716
rect 14778 6664 14787 6694
rect 14787 6664 14821 6694
rect 14821 6664 14830 6694
rect 14778 6622 14830 6652
rect 14778 6600 14787 6622
rect 14787 6600 14821 6622
rect 14821 6600 14830 6622
rect 14778 6550 14830 6588
rect 14778 6536 14787 6550
rect 14787 6536 14821 6550
rect 14821 6536 14830 6550
rect 14778 6516 14787 6524
rect 14787 6516 14821 6524
rect 14821 6516 14830 6524
rect 14778 6478 14830 6516
rect 14778 6472 14787 6478
rect 14787 6472 14821 6478
rect 14821 6472 14830 6478
rect 14778 6444 14787 6460
rect 14787 6444 14821 6460
rect 14821 6444 14830 6460
rect 14778 6408 14830 6444
rect 14778 6372 14787 6396
rect 14787 6372 14821 6396
rect 14821 6372 14830 6396
rect 14778 6344 14830 6372
rect 14778 6300 14787 6332
rect 14787 6300 14821 6332
rect 14821 6300 14830 6332
rect 14778 6280 14830 6300
rect 14778 6262 14830 6268
rect 14778 6228 14787 6262
rect 14787 6228 14821 6262
rect 14821 6228 14830 6262
rect 14778 6216 14830 6228
rect 14778 6190 14830 6204
rect 14778 6156 14787 6190
rect 14787 6156 14821 6190
rect 14821 6156 14830 6190
rect 14778 6152 14830 6156
rect 14778 6118 14830 6140
rect 14778 6088 14787 6118
rect 14787 6088 14821 6118
rect 14821 6088 14830 6118
rect 14778 6046 14830 6076
rect 14778 6024 14787 6046
rect 14787 6024 14821 6046
rect 14821 6024 14830 6046
rect 14778 5974 14830 6012
rect 14778 5960 14787 5974
rect 14787 5960 14821 5974
rect 14821 5960 14830 5974
rect 14778 5940 14787 5948
rect 14787 5940 14821 5948
rect 14821 5940 14830 5948
rect 14778 5902 14830 5940
rect 14778 5896 14787 5902
rect 14787 5896 14821 5902
rect 14821 5896 14830 5902
rect 14864 6804 14873 6810
rect 14873 6804 14907 6810
rect 14907 6804 14916 6810
rect 14864 6766 14916 6804
rect 14864 6758 14873 6766
rect 14873 6758 14907 6766
rect 14907 6758 14916 6766
rect 14864 6732 14873 6746
rect 14873 6732 14907 6746
rect 14907 6732 14916 6746
rect 14864 6694 14916 6732
rect 14864 6660 14873 6682
rect 14873 6660 14907 6682
rect 14907 6660 14916 6682
rect 14864 6630 14916 6660
rect 14864 6588 14873 6618
rect 14873 6588 14907 6618
rect 14907 6588 14916 6618
rect 14864 6566 14916 6588
rect 14864 6550 14916 6554
rect 14864 6516 14873 6550
rect 14873 6516 14907 6550
rect 14907 6516 14916 6550
rect 14864 6502 14916 6516
rect 14864 6478 14916 6490
rect 14864 6444 14873 6478
rect 14873 6444 14907 6478
rect 14907 6444 14916 6478
rect 14864 6438 14916 6444
rect 14864 6406 14916 6426
rect 14864 6374 14873 6406
rect 14873 6374 14907 6406
rect 14907 6374 14916 6406
rect 14864 6334 14916 6362
rect 14864 6310 14873 6334
rect 14873 6310 14907 6334
rect 14907 6310 14916 6334
rect 14864 6262 14916 6298
rect 14864 6246 14873 6262
rect 14873 6246 14907 6262
rect 14907 6246 14916 6262
rect 14864 6228 14873 6234
rect 14873 6228 14907 6234
rect 14907 6228 14916 6234
rect 14864 6190 14916 6228
rect 14864 6182 14873 6190
rect 14873 6182 14907 6190
rect 14907 6182 14916 6190
rect 14864 6156 14873 6170
rect 14873 6156 14907 6170
rect 14907 6156 14916 6170
rect 14864 6118 14916 6156
rect 14864 6084 14873 6106
rect 14873 6084 14907 6106
rect 14907 6084 14916 6106
rect 14864 6054 14916 6084
rect 14864 6012 14873 6042
rect 14873 6012 14907 6042
rect 14907 6012 14916 6042
rect 14864 5990 14916 6012
rect 14864 5974 14916 5978
rect 14864 5940 14873 5974
rect 14873 5940 14907 5974
rect 14907 5940 14916 5974
rect 14864 5926 14916 5940
rect 14864 5902 14916 5914
rect 14864 5868 14873 5902
rect 14873 5868 14907 5902
rect 14907 5868 14916 5902
rect 14864 5862 14916 5868
rect 14950 6838 15002 6844
rect 14950 6804 14959 6838
rect 14959 6804 14993 6838
rect 14993 6804 15002 6838
rect 14950 6792 15002 6804
rect 14950 6766 15002 6780
rect 14950 6732 14959 6766
rect 14959 6732 14993 6766
rect 14993 6732 15002 6766
rect 14950 6728 15002 6732
rect 14950 6694 15002 6716
rect 14950 6664 14959 6694
rect 14959 6664 14993 6694
rect 14993 6664 15002 6694
rect 14950 6622 15002 6652
rect 14950 6600 14959 6622
rect 14959 6600 14993 6622
rect 14993 6600 15002 6622
rect 14950 6550 15002 6588
rect 14950 6536 14959 6550
rect 14959 6536 14993 6550
rect 14993 6536 15002 6550
rect 14950 6516 14959 6524
rect 14959 6516 14993 6524
rect 14993 6516 15002 6524
rect 14950 6478 15002 6516
rect 14950 6472 14959 6478
rect 14959 6472 14993 6478
rect 14993 6472 15002 6478
rect 14950 6444 14959 6460
rect 14959 6444 14993 6460
rect 14993 6444 15002 6460
rect 14950 6408 15002 6444
rect 14950 6372 14959 6396
rect 14959 6372 14993 6396
rect 14993 6372 15002 6396
rect 14950 6344 15002 6372
rect 14950 6300 14959 6332
rect 14959 6300 14993 6332
rect 14993 6300 15002 6332
rect 14950 6280 15002 6300
rect 14950 6262 15002 6268
rect 14950 6228 14959 6262
rect 14959 6228 14993 6262
rect 14993 6228 15002 6262
rect 14950 6216 15002 6228
rect 14950 6190 15002 6204
rect 14950 6156 14959 6190
rect 14959 6156 14993 6190
rect 14993 6156 15002 6190
rect 14950 6152 15002 6156
rect 14950 6118 15002 6140
rect 14950 6088 14959 6118
rect 14959 6088 14993 6118
rect 14993 6088 15002 6118
rect 14950 6046 15002 6076
rect 14950 6024 14959 6046
rect 14959 6024 14993 6046
rect 14993 6024 15002 6046
rect 14950 5974 15002 6012
rect 14950 5960 14959 5974
rect 14959 5960 14993 5974
rect 14993 5960 15002 5974
rect 14950 5940 14959 5948
rect 14959 5940 14993 5948
rect 14993 5940 15002 5948
rect 14950 5902 15002 5940
rect 14950 5896 14959 5902
rect 14959 5896 14993 5902
rect 14993 5896 15002 5902
rect 14700 5510 14940 5570
rect 15172 6838 15224 6844
rect 15172 6804 15181 6838
rect 15181 6804 15215 6838
rect 15215 6804 15224 6838
rect 15172 6792 15224 6804
rect 15172 6766 15224 6780
rect 15172 6732 15181 6766
rect 15181 6732 15215 6766
rect 15215 6732 15224 6766
rect 15172 6728 15224 6732
rect 15172 6694 15224 6716
rect 15172 6664 15181 6694
rect 15181 6664 15215 6694
rect 15215 6664 15224 6694
rect 15172 6622 15224 6652
rect 15172 6600 15181 6622
rect 15181 6600 15215 6622
rect 15215 6600 15224 6622
rect 15172 6550 15224 6588
rect 15172 6536 15181 6550
rect 15181 6536 15215 6550
rect 15215 6536 15224 6550
rect 15172 6516 15181 6524
rect 15181 6516 15215 6524
rect 15215 6516 15224 6524
rect 15172 6478 15224 6516
rect 15172 6472 15181 6478
rect 15181 6472 15215 6478
rect 15215 6472 15224 6478
rect 15172 6444 15181 6460
rect 15181 6444 15215 6460
rect 15215 6444 15224 6460
rect 15172 6408 15224 6444
rect 15172 6372 15181 6396
rect 15181 6372 15215 6396
rect 15215 6372 15224 6396
rect 15172 6344 15224 6372
rect 15172 6300 15181 6332
rect 15181 6300 15215 6332
rect 15215 6300 15224 6332
rect 15172 6280 15224 6300
rect 15172 6262 15224 6268
rect 15172 6228 15181 6262
rect 15181 6228 15215 6262
rect 15215 6228 15224 6262
rect 15172 6216 15224 6228
rect 15172 6190 15224 6204
rect 15172 6156 15181 6190
rect 15181 6156 15215 6190
rect 15215 6156 15224 6190
rect 15172 6152 15224 6156
rect 15172 6118 15224 6140
rect 15172 6088 15181 6118
rect 15181 6088 15215 6118
rect 15215 6088 15224 6118
rect 15172 6046 15224 6076
rect 15172 6024 15181 6046
rect 15181 6024 15215 6046
rect 15215 6024 15224 6046
rect 15172 5974 15224 6012
rect 15172 5960 15181 5974
rect 15181 5960 15215 5974
rect 15215 5960 15224 5974
rect 15172 5940 15181 5948
rect 15181 5940 15215 5948
rect 15215 5940 15224 5948
rect 15172 5902 15224 5940
rect 15172 5896 15181 5902
rect 15181 5896 15215 5902
rect 15215 5896 15224 5902
rect 15258 6804 15267 6810
rect 15267 6804 15301 6810
rect 15301 6804 15310 6810
rect 15258 6766 15310 6804
rect 15258 6758 15267 6766
rect 15267 6758 15301 6766
rect 15301 6758 15310 6766
rect 15258 6732 15267 6746
rect 15267 6732 15301 6746
rect 15301 6732 15310 6746
rect 15258 6694 15310 6732
rect 15258 6660 15267 6682
rect 15267 6660 15301 6682
rect 15301 6660 15310 6682
rect 15258 6630 15310 6660
rect 15258 6588 15267 6618
rect 15267 6588 15301 6618
rect 15301 6588 15310 6618
rect 15258 6566 15310 6588
rect 15258 6550 15310 6554
rect 15258 6516 15267 6550
rect 15267 6516 15301 6550
rect 15301 6516 15310 6550
rect 15258 6502 15310 6516
rect 15258 6478 15310 6490
rect 15258 6444 15267 6478
rect 15267 6444 15301 6478
rect 15301 6444 15310 6478
rect 15258 6438 15310 6444
rect 15258 6406 15310 6426
rect 15258 6374 15267 6406
rect 15267 6374 15301 6406
rect 15301 6374 15310 6406
rect 15258 6334 15310 6362
rect 15258 6310 15267 6334
rect 15267 6310 15301 6334
rect 15301 6310 15310 6334
rect 15258 6262 15310 6298
rect 15258 6246 15267 6262
rect 15267 6246 15301 6262
rect 15301 6246 15310 6262
rect 15258 6228 15267 6234
rect 15267 6228 15301 6234
rect 15301 6228 15310 6234
rect 15258 6190 15310 6228
rect 15258 6182 15267 6190
rect 15267 6182 15301 6190
rect 15301 6182 15310 6190
rect 15258 6156 15267 6170
rect 15267 6156 15301 6170
rect 15301 6156 15310 6170
rect 15258 6118 15310 6156
rect 15258 6084 15267 6106
rect 15267 6084 15301 6106
rect 15301 6084 15310 6106
rect 15258 6054 15310 6084
rect 15258 6012 15267 6042
rect 15267 6012 15301 6042
rect 15301 6012 15310 6042
rect 15258 5990 15310 6012
rect 15258 5974 15310 5978
rect 15258 5940 15267 5974
rect 15267 5940 15301 5974
rect 15301 5940 15310 5974
rect 15258 5926 15310 5940
rect 15258 5902 15310 5914
rect 15258 5868 15267 5902
rect 15267 5868 15301 5902
rect 15301 5868 15310 5902
rect 15258 5862 15310 5868
rect 15344 6838 15396 6844
rect 15344 6804 15353 6838
rect 15353 6804 15387 6838
rect 15387 6804 15396 6838
rect 15344 6792 15396 6804
rect 15344 6766 15396 6780
rect 15344 6732 15353 6766
rect 15353 6732 15387 6766
rect 15387 6732 15396 6766
rect 15344 6728 15396 6732
rect 15344 6694 15396 6716
rect 15344 6664 15353 6694
rect 15353 6664 15387 6694
rect 15387 6664 15396 6694
rect 15344 6622 15396 6652
rect 15344 6600 15353 6622
rect 15353 6600 15387 6622
rect 15387 6600 15396 6622
rect 15344 6550 15396 6588
rect 15344 6536 15353 6550
rect 15353 6536 15387 6550
rect 15387 6536 15396 6550
rect 15344 6516 15353 6524
rect 15353 6516 15387 6524
rect 15387 6516 15396 6524
rect 15344 6478 15396 6516
rect 15344 6472 15353 6478
rect 15353 6472 15387 6478
rect 15387 6472 15396 6478
rect 15344 6444 15353 6460
rect 15353 6444 15387 6460
rect 15387 6444 15396 6460
rect 15344 6408 15396 6444
rect 15344 6372 15353 6396
rect 15353 6372 15387 6396
rect 15387 6372 15396 6396
rect 15344 6344 15396 6372
rect 15344 6300 15353 6332
rect 15353 6300 15387 6332
rect 15387 6300 15396 6332
rect 15344 6280 15396 6300
rect 15344 6262 15396 6268
rect 15344 6228 15353 6262
rect 15353 6228 15387 6262
rect 15387 6228 15396 6262
rect 15344 6216 15396 6228
rect 15344 6190 15396 6204
rect 15344 6156 15353 6190
rect 15353 6156 15387 6190
rect 15387 6156 15396 6190
rect 15344 6152 15396 6156
rect 15344 6118 15396 6140
rect 15344 6088 15353 6118
rect 15353 6088 15387 6118
rect 15387 6088 15396 6118
rect 15344 6046 15396 6076
rect 15344 6024 15353 6046
rect 15353 6024 15387 6046
rect 15387 6024 15396 6046
rect 15344 5974 15396 6012
rect 15344 5960 15353 5974
rect 15353 5960 15387 5974
rect 15387 5960 15396 5974
rect 15344 5940 15353 5948
rect 15353 5940 15387 5948
rect 15387 5940 15396 5948
rect 15344 5902 15396 5940
rect 15344 5896 15353 5902
rect 15353 5896 15387 5902
rect 15387 5896 15396 5902
rect 15430 6804 15439 6810
rect 15439 6804 15473 6810
rect 15473 6804 15482 6810
rect 15430 6766 15482 6804
rect 15430 6758 15439 6766
rect 15439 6758 15473 6766
rect 15473 6758 15482 6766
rect 15430 6732 15439 6746
rect 15439 6732 15473 6746
rect 15473 6732 15482 6746
rect 15430 6694 15482 6732
rect 15430 6660 15439 6682
rect 15439 6660 15473 6682
rect 15473 6660 15482 6682
rect 15430 6630 15482 6660
rect 15430 6588 15439 6618
rect 15439 6588 15473 6618
rect 15473 6588 15482 6618
rect 15430 6566 15482 6588
rect 15430 6550 15482 6554
rect 15430 6516 15439 6550
rect 15439 6516 15473 6550
rect 15473 6516 15482 6550
rect 15430 6502 15482 6516
rect 15430 6478 15482 6490
rect 15430 6444 15439 6478
rect 15439 6444 15473 6478
rect 15473 6444 15482 6478
rect 15430 6438 15482 6444
rect 15430 6406 15482 6426
rect 15430 6374 15439 6406
rect 15439 6374 15473 6406
rect 15473 6374 15482 6406
rect 15430 6334 15482 6362
rect 15430 6310 15439 6334
rect 15439 6310 15473 6334
rect 15473 6310 15482 6334
rect 15430 6262 15482 6298
rect 15430 6246 15439 6262
rect 15439 6246 15473 6262
rect 15473 6246 15482 6262
rect 15430 6228 15439 6234
rect 15439 6228 15473 6234
rect 15473 6228 15482 6234
rect 15430 6190 15482 6228
rect 15430 6182 15439 6190
rect 15439 6182 15473 6190
rect 15473 6182 15482 6190
rect 15430 6156 15439 6170
rect 15439 6156 15473 6170
rect 15473 6156 15482 6170
rect 15430 6118 15482 6156
rect 15430 6084 15439 6106
rect 15439 6084 15473 6106
rect 15473 6084 15482 6106
rect 15430 6054 15482 6084
rect 15430 6012 15439 6042
rect 15439 6012 15473 6042
rect 15473 6012 15482 6042
rect 15430 5990 15482 6012
rect 15430 5974 15482 5978
rect 15430 5940 15439 5974
rect 15439 5940 15473 5974
rect 15473 5940 15482 5974
rect 15430 5926 15482 5940
rect 15430 5902 15482 5914
rect 15430 5868 15439 5902
rect 15439 5868 15473 5902
rect 15473 5868 15482 5902
rect 15430 5862 15482 5868
rect 15516 6838 15568 6844
rect 15516 6804 15525 6838
rect 15525 6804 15559 6838
rect 15559 6804 15568 6838
rect 15516 6792 15568 6804
rect 15516 6766 15568 6780
rect 15516 6732 15525 6766
rect 15525 6732 15559 6766
rect 15559 6732 15568 6766
rect 15516 6728 15568 6732
rect 15516 6694 15568 6716
rect 15516 6664 15525 6694
rect 15525 6664 15559 6694
rect 15559 6664 15568 6694
rect 15516 6622 15568 6652
rect 15516 6600 15525 6622
rect 15525 6600 15559 6622
rect 15559 6600 15568 6622
rect 15516 6550 15568 6588
rect 15516 6536 15525 6550
rect 15525 6536 15559 6550
rect 15559 6536 15568 6550
rect 15516 6516 15525 6524
rect 15525 6516 15559 6524
rect 15559 6516 15568 6524
rect 15516 6478 15568 6516
rect 15516 6472 15525 6478
rect 15525 6472 15559 6478
rect 15559 6472 15568 6478
rect 15516 6444 15525 6460
rect 15525 6444 15559 6460
rect 15559 6444 15568 6460
rect 15516 6408 15568 6444
rect 15516 6372 15525 6396
rect 15525 6372 15559 6396
rect 15559 6372 15568 6396
rect 15516 6344 15568 6372
rect 15516 6300 15525 6332
rect 15525 6300 15559 6332
rect 15559 6300 15568 6332
rect 15516 6280 15568 6300
rect 15516 6262 15568 6268
rect 15516 6228 15525 6262
rect 15525 6228 15559 6262
rect 15559 6228 15568 6262
rect 15516 6216 15568 6228
rect 15516 6190 15568 6204
rect 15516 6156 15525 6190
rect 15525 6156 15559 6190
rect 15559 6156 15568 6190
rect 15516 6152 15568 6156
rect 15516 6118 15568 6140
rect 15516 6088 15525 6118
rect 15525 6088 15559 6118
rect 15559 6088 15568 6118
rect 15516 6046 15568 6076
rect 15516 6024 15525 6046
rect 15525 6024 15559 6046
rect 15559 6024 15568 6046
rect 15516 5974 15568 6012
rect 15516 5960 15525 5974
rect 15525 5960 15559 5974
rect 15559 5960 15568 5974
rect 15516 5940 15525 5948
rect 15525 5940 15559 5948
rect 15559 5940 15568 5948
rect 15516 5902 15568 5940
rect 15516 5896 15525 5902
rect 15525 5896 15559 5902
rect 15559 5896 15568 5902
rect 16140 6750 17130 6810
rect 17680 6710 20000 6820
rect 16140 6350 17170 6410
rect 17660 6390 19980 6500
rect 15260 5510 15500 5570
rect 11650 5380 15690 5460
rect 15960 6154 16100 6160
rect 15960 6120 15990 6154
rect 15990 6120 16024 6154
rect 16024 6120 16100 6154
rect 15960 6074 16100 6120
rect 15960 6040 15990 6074
rect 15990 6040 16024 6074
rect 16024 6040 16100 6074
rect 15960 5994 16100 6040
rect 15960 5960 15990 5994
rect 15990 5960 16024 5994
rect 16024 5960 16100 5994
rect 15960 5914 16100 5960
rect 15960 5880 15990 5914
rect 15990 5880 16024 5914
rect 16024 5880 16100 5914
rect 15960 5834 16100 5880
rect 15960 5800 15990 5834
rect 15990 5800 16024 5834
rect 16024 5800 16100 5834
rect 15960 5754 16100 5800
rect 15960 5720 15990 5754
rect 15990 5720 16024 5754
rect 16024 5720 16100 5754
rect 15960 5674 16100 5720
rect 15960 5640 15990 5674
rect 15990 5640 16024 5674
rect 16024 5640 16100 5674
rect 15960 5594 16100 5640
rect 15960 5560 15990 5594
rect 15990 5560 16024 5594
rect 16024 5560 16100 5594
rect 15960 5514 16100 5560
rect 15960 5480 15990 5514
rect 15990 5480 16024 5514
rect 16024 5480 16100 5514
rect 15960 5434 16100 5480
rect 15960 5400 15990 5434
rect 15990 5400 16024 5434
rect 16024 5400 16100 5434
rect 15960 5354 16100 5400
rect 15960 5320 15990 5354
rect 15990 5320 16024 5354
rect 16024 5320 16100 5354
rect 15960 5274 16100 5320
rect 15960 5240 15990 5274
rect 15990 5240 16024 5274
rect 16024 5240 16100 5274
rect 15960 5194 16100 5240
rect 15960 5160 15990 5194
rect 15990 5160 16024 5194
rect 16024 5160 16100 5194
rect 15960 5084 16100 5160
rect 16195 6099 16247 6111
rect 16195 6065 16204 6099
rect 16204 6065 16238 6099
rect 16238 6065 16247 6099
rect 16195 6059 16247 6065
rect 16195 6027 16247 6031
rect 16195 5993 16204 6027
rect 16204 5993 16238 6027
rect 16238 5993 16247 6027
rect 16195 5979 16247 5993
rect 16195 5921 16204 5951
rect 16204 5921 16238 5951
rect 16238 5921 16247 5951
rect 16195 5899 16247 5921
rect 16195 5849 16204 5871
rect 16204 5849 16238 5871
rect 16238 5849 16247 5871
rect 16195 5819 16247 5849
rect 16195 5777 16204 5791
rect 16204 5777 16238 5791
rect 16238 5777 16247 5791
rect 16195 5739 16247 5777
rect 16195 5705 16204 5711
rect 16204 5705 16238 5711
rect 16238 5705 16247 5711
rect 16195 5667 16247 5705
rect 16195 5659 16204 5667
rect 16204 5659 16238 5667
rect 16238 5659 16247 5667
rect 16195 5595 16247 5631
rect 16195 5579 16204 5595
rect 16204 5579 16238 5595
rect 16238 5579 16247 5595
rect 16195 5523 16247 5551
rect 16195 5499 16204 5523
rect 16204 5499 16238 5523
rect 16238 5499 16247 5523
rect 16195 5451 16247 5471
rect 16195 5419 16204 5451
rect 16204 5419 16238 5451
rect 16238 5419 16247 5451
rect 16195 5379 16247 5391
rect 16195 5345 16204 5379
rect 16204 5345 16238 5379
rect 16238 5345 16247 5379
rect 16195 5339 16247 5345
rect 16195 5307 16247 5311
rect 16195 5273 16204 5307
rect 16204 5273 16238 5307
rect 16238 5273 16247 5307
rect 16195 5259 16247 5273
rect 16367 6099 16419 6111
rect 16367 6065 16376 6099
rect 16376 6065 16410 6099
rect 16410 6065 16419 6099
rect 16367 6059 16419 6065
rect 16367 6027 16419 6031
rect 16367 5993 16376 6027
rect 16376 5993 16410 6027
rect 16410 5993 16419 6027
rect 16367 5979 16419 5993
rect 16367 5921 16376 5951
rect 16376 5921 16410 5951
rect 16410 5921 16419 5951
rect 16367 5899 16419 5921
rect 16367 5849 16376 5871
rect 16376 5849 16410 5871
rect 16410 5849 16419 5871
rect 16367 5819 16419 5849
rect 16367 5777 16376 5791
rect 16376 5777 16410 5791
rect 16410 5777 16419 5791
rect 16367 5739 16419 5777
rect 16367 5705 16376 5711
rect 16376 5705 16410 5711
rect 16410 5705 16419 5711
rect 16367 5667 16419 5705
rect 16367 5659 16376 5667
rect 16376 5659 16410 5667
rect 16410 5659 16419 5667
rect 16367 5595 16419 5631
rect 16367 5579 16376 5595
rect 16376 5579 16410 5595
rect 16410 5579 16419 5595
rect 16367 5523 16419 5551
rect 16367 5499 16376 5523
rect 16376 5499 16410 5523
rect 16410 5499 16419 5523
rect 16367 5451 16419 5471
rect 16367 5419 16376 5451
rect 16376 5419 16410 5451
rect 16410 5419 16419 5451
rect 16367 5379 16419 5391
rect 16367 5345 16376 5379
rect 16376 5345 16410 5379
rect 16410 5345 16419 5379
rect 16367 5339 16419 5345
rect 16367 5307 16419 5311
rect 16367 5273 16376 5307
rect 16376 5273 16410 5307
rect 16410 5273 16419 5307
rect 16367 5259 16419 5273
rect 16539 6099 16591 6111
rect 16539 6065 16548 6099
rect 16548 6065 16582 6099
rect 16582 6065 16591 6099
rect 16539 6059 16591 6065
rect 16539 6027 16591 6031
rect 16539 5993 16548 6027
rect 16548 5993 16582 6027
rect 16582 5993 16591 6027
rect 16539 5979 16591 5993
rect 16539 5921 16548 5951
rect 16548 5921 16582 5951
rect 16582 5921 16591 5951
rect 16539 5899 16591 5921
rect 16539 5849 16548 5871
rect 16548 5849 16582 5871
rect 16582 5849 16591 5871
rect 16539 5819 16591 5849
rect 16539 5777 16548 5791
rect 16548 5777 16582 5791
rect 16582 5777 16591 5791
rect 16539 5739 16591 5777
rect 16539 5705 16548 5711
rect 16548 5705 16582 5711
rect 16582 5705 16591 5711
rect 16539 5667 16591 5705
rect 16539 5659 16548 5667
rect 16548 5659 16582 5667
rect 16582 5659 16591 5667
rect 16539 5595 16591 5631
rect 16539 5579 16548 5595
rect 16548 5579 16582 5595
rect 16582 5579 16591 5595
rect 16539 5523 16591 5551
rect 16539 5499 16548 5523
rect 16548 5499 16582 5523
rect 16582 5499 16591 5523
rect 16539 5451 16591 5471
rect 16539 5419 16548 5451
rect 16548 5419 16582 5451
rect 16582 5419 16591 5451
rect 16539 5379 16591 5391
rect 16539 5345 16548 5379
rect 16548 5345 16582 5379
rect 16582 5345 16591 5379
rect 16539 5339 16591 5345
rect 16539 5307 16591 5311
rect 16539 5273 16548 5307
rect 16548 5273 16582 5307
rect 16582 5273 16591 5307
rect 16539 5259 16591 5273
rect 16711 6099 16763 6111
rect 16711 6065 16720 6099
rect 16720 6065 16754 6099
rect 16754 6065 16763 6099
rect 16711 6059 16763 6065
rect 16711 6027 16763 6031
rect 16711 5993 16720 6027
rect 16720 5993 16754 6027
rect 16754 5993 16763 6027
rect 16711 5979 16763 5993
rect 16711 5921 16720 5951
rect 16720 5921 16754 5951
rect 16754 5921 16763 5951
rect 16711 5899 16763 5921
rect 16711 5849 16720 5871
rect 16720 5849 16754 5871
rect 16754 5849 16763 5871
rect 16711 5819 16763 5849
rect 16711 5777 16720 5791
rect 16720 5777 16754 5791
rect 16754 5777 16763 5791
rect 16711 5739 16763 5777
rect 16711 5705 16720 5711
rect 16720 5705 16754 5711
rect 16754 5705 16763 5711
rect 16711 5667 16763 5705
rect 16711 5659 16720 5667
rect 16720 5659 16754 5667
rect 16754 5659 16763 5667
rect 16711 5595 16763 5631
rect 16711 5579 16720 5595
rect 16720 5579 16754 5595
rect 16754 5579 16763 5595
rect 16711 5523 16763 5551
rect 16711 5499 16720 5523
rect 16720 5499 16754 5523
rect 16754 5499 16763 5523
rect 16711 5451 16763 5471
rect 16711 5419 16720 5451
rect 16720 5419 16754 5451
rect 16754 5419 16763 5451
rect 16711 5379 16763 5391
rect 16711 5345 16720 5379
rect 16720 5345 16754 5379
rect 16754 5345 16763 5379
rect 16711 5339 16763 5345
rect 16711 5307 16763 5311
rect 16711 5273 16720 5307
rect 16720 5273 16754 5307
rect 16754 5273 16763 5307
rect 16711 5259 16763 5273
rect 16883 6099 16935 6111
rect 16883 6065 16892 6099
rect 16892 6065 16926 6099
rect 16926 6065 16935 6099
rect 16883 6059 16935 6065
rect 16883 6027 16935 6031
rect 16883 5993 16892 6027
rect 16892 5993 16926 6027
rect 16926 5993 16935 6027
rect 16883 5979 16935 5993
rect 16883 5921 16892 5951
rect 16892 5921 16926 5951
rect 16926 5921 16935 5951
rect 16883 5899 16935 5921
rect 16883 5849 16892 5871
rect 16892 5849 16926 5871
rect 16926 5849 16935 5871
rect 16883 5819 16935 5849
rect 16883 5777 16892 5791
rect 16892 5777 16926 5791
rect 16926 5777 16935 5791
rect 16883 5739 16935 5777
rect 16883 5705 16892 5711
rect 16892 5705 16926 5711
rect 16926 5705 16935 5711
rect 16883 5667 16935 5705
rect 16883 5659 16892 5667
rect 16892 5659 16926 5667
rect 16926 5659 16935 5667
rect 16883 5595 16935 5631
rect 16883 5579 16892 5595
rect 16892 5579 16926 5595
rect 16926 5579 16935 5595
rect 16883 5523 16935 5551
rect 16883 5499 16892 5523
rect 16892 5499 16926 5523
rect 16926 5499 16935 5523
rect 16883 5451 16935 5471
rect 16883 5419 16892 5451
rect 16892 5419 16926 5451
rect 16926 5419 16935 5451
rect 16883 5379 16935 5391
rect 16883 5345 16892 5379
rect 16892 5345 16926 5379
rect 16926 5345 16935 5379
rect 16883 5339 16935 5345
rect 16883 5307 16935 5311
rect 16883 5273 16892 5307
rect 16892 5273 16926 5307
rect 16926 5273 16935 5307
rect 16883 5259 16935 5273
rect 17055 6099 17107 6111
rect 17055 6065 17064 6099
rect 17064 6065 17098 6099
rect 17098 6065 17107 6099
rect 17055 6059 17107 6065
rect 17055 6027 17107 6031
rect 17055 5993 17064 6027
rect 17064 5993 17098 6027
rect 17098 5993 17107 6027
rect 17055 5979 17107 5993
rect 17055 5921 17064 5951
rect 17064 5921 17098 5951
rect 17098 5921 17107 5951
rect 17055 5899 17107 5921
rect 17055 5849 17064 5871
rect 17064 5849 17098 5871
rect 17098 5849 17107 5871
rect 17055 5819 17107 5849
rect 17055 5777 17064 5791
rect 17064 5777 17098 5791
rect 17098 5777 17107 5791
rect 17055 5739 17107 5777
rect 17055 5705 17064 5711
rect 17064 5705 17098 5711
rect 17098 5705 17107 5711
rect 17055 5667 17107 5705
rect 17055 5659 17064 5667
rect 17064 5659 17098 5667
rect 17098 5659 17107 5667
rect 17055 5595 17107 5631
rect 17055 5579 17064 5595
rect 17064 5579 17098 5595
rect 17098 5579 17107 5595
rect 17055 5523 17107 5551
rect 17055 5499 17064 5523
rect 17064 5499 17098 5523
rect 17098 5499 17107 5523
rect 17055 5451 17107 5471
rect 17055 5419 17064 5451
rect 17064 5419 17098 5451
rect 17098 5419 17107 5451
rect 17055 5379 17107 5391
rect 17055 5345 17064 5379
rect 17064 5345 17098 5379
rect 17098 5345 17107 5379
rect 17055 5339 17107 5345
rect 17055 5307 17107 5311
rect 17055 5273 17064 5307
rect 17064 5273 17098 5307
rect 17098 5273 17107 5307
rect 17055 5259 17107 5273
rect 17681 6180 17733 6207
rect 17681 6155 17690 6180
rect 17690 6155 17724 6180
rect 17724 6155 17733 6180
rect 17681 6108 17733 6143
rect 17681 6091 17690 6108
rect 17690 6091 17724 6108
rect 17724 6091 17733 6108
rect 17853 6180 17905 6207
rect 17853 6155 17862 6180
rect 17862 6155 17896 6180
rect 17896 6155 17905 6180
rect 17853 6108 17905 6143
rect 17853 6091 17862 6108
rect 17862 6091 17896 6108
rect 17896 6091 17905 6108
rect 18025 6180 18077 6207
rect 18025 6155 18034 6180
rect 18034 6155 18068 6180
rect 18068 6155 18077 6180
rect 18025 6108 18077 6143
rect 18025 6091 18034 6108
rect 18034 6091 18068 6108
rect 18068 6091 18077 6108
rect 18197 6180 18249 6207
rect 18197 6155 18206 6180
rect 18206 6155 18240 6180
rect 18240 6155 18249 6180
rect 18197 6108 18249 6143
rect 18197 6091 18206 6108
rect 18206 6091 18240 6108
rect 18240 6091 18249 6108
rect 18369 6180 18421 6207
rect 18369 6155 18378 6180
rect 18378 6155 18412 6180
rect 18412 6155 18421 6180
rect 18369 6108 18421 6143
rect 18369 6091 18378 6108
rect 18378 6091 18412 6108
rect 18412 6091 18421 6108
rect 18541 6180 18593 6207
rect 18541 6155 18550 6180
rect 18550 6155 18584 6180
rect 18584 6155 18593 6180
rect 18541 6108 18593 6143
rect 18541 6091 18550 6108
rect 18550 6091 18584 6108
rect 18584 6091 18593 6108
rect 18713 6180 18765 6207
rect 18713 6155 18722 6180
rect 18722 6155 18756 6180
rect 18756 6155 18765 6180
rect 18713 6108 18765 6143
rect 18713 6091 18722 6108
rect 18722 6091 18756 6108
rect 18756 6091 18765 6108
rect 18885 6180 18937 6207
rect 18885 6155 18894 6180
rect 18894 6155 18928 6180
rect 18928 6155 18937 6180
rect 18885 6108 18937 6143
rect 18885 6091 18894 6108
rect 18894 6091 18928 6108
rect 18928 6091 18937 6108
rect 19057 6180 19109 6207
rect 19057 6155 19066 6180
rect 19066 6155 19100 6180
rect 19100 6155 19109 6180
rect 19057 6108 19109 6143
rect 19057 6091 19066 6108
rect 19066 6091 19100 6108
rect 19100 6091 19109 6108
rect 19229 6180 19281 6207
rect 19229 6155 19238 6180
rect 19238 6155 19272 6180
rect 19272 6155 19281 6180
rect 19229 6108 19281 6143
rect 19229 6091 19238 6108
rect 19238 6091 19272 6108
rect 19272 6091 19281 6108
rect 19401 6180 19453 6207
rect 19401 6155 19410 6180
rect 19410 6155 19444 6180
rect 19444 6155 19453 6180
rect 19401 6108 19453 6143
rect 19401 6091 19410 6108
rect 19410 6091 19444 6108
rect 19444 6091 19453 6108
rect 19573 6180 19625 6207
rect 19573 6155 19582 6180
rect 19582 6155 19616 6180
rect 19616 6155 19625 6180
rect 19573 6108 19625 6143
rect 19573 6091 19582 6108
rect 19582 6091 19616 6108
rect 19616 6091 19625 6108
rect 19745 6180 19797 6207
rect 19745 6155 19754 6180
rect 19754 6155 19788 6180
rect 19788 6155 19797 6180
rect 19745 6108 19797 6143
rect 19745 6091 19754 6108
rect 19754 6091 19788 6108
rect 19788 6091 19797 6108
rect 19917 6180 19969 6207
rect 19917 6155 19926 6180
rect 19926 6155 19960 6180
rect 19960 6155 19969 6180
rect 19917 6108 19969 6143
rect 19917 6091 19926 6108
rect 19926 6091 19960 6108
rect 19960 6091 19969 6108
rect 20060 5260 20120 6190
rect 20120 5260 20160 6190
rect 20160 5260 20180 6190
rect 15960 5050 16080 5084
rect 16080 5050 16100 5084
rect 17420 5000 20140 5100
rect 16638 4802 16690 4811
rect 16638 4768 16669 4802
rect 16669 4768 16690 4802
rect 16557 4735 16609 4765
rect 16638 4759 16690 4768
rect 16702 4802 16754 4811
rect 16702 4768 16707 4802
rect 16707 4768 16741 4802
rect 16741 4768 16754 4802
rect 16702 4759 16754 4768
rect 16766 4802 16818 4811
rect 16766 4768 16779 4802
rect 16779 4768 16813 4802
rect 16813 4768 16818 4802
rect 16766 4759 16818 4768
rect 16830 4802 16882 4811
rect 16894 4802 16946 4811
rect 16958 4802 17010 4811
rect 17022 4802 17074 4811
rect 17086 4802 17138 4811
rect 17150 4802 17202 4811
rect 17214 4802 17266 4811
rect 16830 4768 16851 4802
rect 16851 4768 16882 4802
rect 16894 4768 16923 4802
rect 16923 4768 16946 4802
rect 16958 4768 16995 4802
rect 16995 4768 17010 4802
rect 17022 4768 17029 4802
rect 17029 4768 17067 4802
rect 17067 4768 17074 4802
rect 17086 4768 17101 4802
rect 17101 4768 17138 4802
rect 17150 4768 17173 4802
rect 17173 4768 17202 4802
rect 17214 4768 17245 4802
rect 17245 4768 17266 4802
rect 16830 4759 16882 4768
rect 16894 4759 16946 4768
rect 16958 4759 17010 4768
rect 17022 4759 17074 4768
rect 17086 4759 17138 4768
rect 17150 4759 17202 4768
rect 17214 4759 17266 4768
rect 17278 4802 17330 4811
rect 17492 4802 17544 4811
rect 17278 4768 17283 4802
rect 17283 4768 17317 4802
rect 17317 4768 17330 4802
rect 17492 4768 17499 4802
rect 17499 4768 17533 4802
rect 17533 4768 17544 4802
rect 17278 4759 17330 4768
rect 17492 4759 17544 4768
rect 17556 4802 17608 4811
rect 17556 4768 17571 4802
rect 17571 4768 17605 4802
rect 17605 4768 17608 4802
rect 17556 4759 17608 4768
rect 17620 4802 17672 4811
rect 17684 4802 17736 4811
rect 17748 4802 17800 4811
rect 17812 4802 17864 4811
rect 17876 4802 17928 4811
rect 17940 4802 17992 4811
rect 18004 4802 18056 4811
rect 17620 4768 17643 4802
rect 17643 4768 17672 4802
rect 17684 4768 17715 4802
rect 17715 4768 17736 4802
rect 17748 4768 17749 4802
rect 17749 4768 17787 4802
rect 17787 4768 17800 4802
rect 17812 4768 17821 4802
rect 17821 4768 17859 4802
rect 17859 4768 17864 4802
rect 17876 4768 17893 4802
rect 17893 4768 17928 4802
rect 17940 4768 17965 4802
rect 17965 4768 17992 4802
rect 18004 4768 18037 4802
rect 18037 4768 18056 4802
rect 17620 4759 17672 4768
rect 17684 4759 17736 4768
rect 17748 4759 17800 4768
rect 17812 4759 17864 4768
rect 17876 4759 17928 4768
rect 17940 4759 17992 4768
rect 18004 4759 18056 4768
rect 18068 4802 18120 4811
rect 18068 4768 18075 4802
rect 18075 4768 18109 4802
rect 18109 4768 18120 4802
rect 18068 4759 18120 4768
rect 18132 4802 18184 4811
rect 18488 4802 18540 4811
rect 18132 4768 18147 4802
rect 18147 4768 18181 4802
rect 18181 4768 18184 4802
rect 18488 4768 18519 4802
rect 18519 4768 18540 4802
rect 18132 4759 18184 4768
rect 16557 4713 16566 4735
rect 16566 4713 16600 4735
rect 16600 4713 16609 4735
rect 16557 4663 16609 4701
rect 16557 4649 16566 4663
rect 16566 4649 16600 4663
rect 16600 4649 16609 4663
rect 16557 4629 16566 4637
rect 16566 4629 16600 4637
rect 16600 4629 16609 4637
rect 16557 4591 16609 4629
rect 16557 4585 16566 4591
rect 16566 4585 16600 4591
rect 16600 4585 16609 4591
rect 16557 4557 16566 4573
rect 16566 4557 16600 4573
rect 16600 4557 16609 4573
rect 16557 4521 16609 4557
rect 16557 4485 16566 4509
rect 16566 4485 16600 4509
rect 16600 4485 16609 4509
rect 16557 4457 16609 4485
rect 16557 4413 16566 4445
rect 16566 4413 16600 4445
rect 16600 4413 16609 4445
rect 16557 4393 16609 4413
rect 16557 4375 16609 4381
rect 16557 4341 16566 4375
rect 16566 4341 16600 4375
rect 16600 4341 16609 4375
rect 16557 4329 16609 4341
rect 16557 4303 16609 4317
rect 16557 4269 16566 4303
rect 16566 4269 16600 4303
rect 16600 4269 16609 4303
rect 16557 4265 16609 4269
rect 16557 4231 16609 4253
rect 16557 4201 16566 4231
rect 16566 4201 16600 4231
rect 16600 4201 16609 4231
rect 16557 4159 16609 4189
rect 16557 4137 16566 4159
rect 16566 4137 16600 4159
rect 16600 4137 16609 4159
rect 16557 3909 16566 3931
rect 16566 3909 16600 3931
rect 16600 3909 16609 3931
rect 16557 3879 16609 3909
rect 16557 3837 16566 3867
rect 16566 3837 16600 3867
rect 16600 3837 16609 3867
rect 16557 3815 16609 3837
rect 16557 3799 16609 3803
rect 16557 3765 16566 3799
rect 16566 3765 16600 3799
rect 16600 3765 16609 3799
rect 16557 3751 16609 3765
rect 16557 3727 16609 3739
rect 16557 3693 16566 3727
rect 16566 3693 16600 3727
rect 16600 3693 16609 3727
rect 16557 3687 16609 3693
rect 16557 3655 16609 3675
rect 16557 3623 16566 3655
rect 16566 3623 16600 3655
rect 16600 3623 16609 3655
rect 16557 3583 16609 3611
rect 16557 3559 16566 3583
rect 16566 3559 16600 3583
rect 16600 3559 16609 3583
rect 16557 3511 16609 3547
rect 16557 3495 16566 3511
rect 16566 3495 16600 3511
rect 16600 3495 16609 3511
rect 16557 3477 16566 3483
rect 16566 3477 16600 3483
rect 16600 3477 16609 3483
rect 16557 3439 16609 3477
rect 16557 3431 16566 3439
rect 16566 3431 16600 3439
rect 16600 3431 16609 3439
rect 16557 3405 16566 3419
rect 16566 3405 16600 3419
rect 16600 3405 16609 3419
rect 16557 3367 16609 3405
rect 16557 3333 16566 3355
rect 16566 3333 16600 3355
rect 16600 3333 16609 3355
rect 16557 3303 16609 3333
rect 17382 4666 17434 4718
rect 17382 4602 17434 4654
rect 17382 4538 17434 4590
rect 17382 4474 17434 4526
rect 17382 4410 17434 4462
rect 17382 4346 17434 4398
rect 17382 4282 17434 4334
rect 17382 4218 17434 4270
rect 17382 4154 17434 4206
rect 17382 4090 17434 4142
rect 16655 4008 16707 4060
rect 16719 4008 16771 4060
rect 16783 4008 16835 4060
rect 16847 4008 16899 4060
rect 16911 4008 16963 4060
rect 16975 4008 17027 4060
rect 17039 4008 17091 4060
rect 17103 4008 17155 4060
rect 17167 4008 17219 4060
rect 17231 4008 17283 4060
rect 17295 4008 17347 4060
rect 17469 4008 17521 4060
rect 17533 4008 17585 4060
rect 17597 4008 17649 4060
rect 17661 4008 17713 4060
rect 17725 4008 17777 4060
rect 17789 4008 17841 4060
rect 17853 4008 17905 4060
rect 17917 4008 17969 4060
rect 17981 4008 18033 4060
rect 18045 4008 18097 4060
rect 18109 4008 18161 4060
rect 17382 3926 17434 3978
rect 17382 3862 17434 3914
rect 17382 3798 17434 3850
rect 17382 3734 17434 3786
rect 17382 3670 17434 3722
rect 17382 3606 17434 3658
rect 17382 3542 17434 3594
rect 17382 3478 17434 3530
rect 17382 3414 17434 3466
rect 17382 3350 17434 3402
rect 18207 4735 18259 4765
rect 18207 4713 18216 4735
rect 18216 4713 18250 4735
rect 18250 4713 18259 4735
rect 18407 4735 18459 4765
rect 18488 4759 18540 4768
rect 18552 4802 18604 4811
rect 18552 4768 18557 4802
rect 18557 4768 18591 4802
rect 18591 4768 18604 4802
rect 18552 4759 18604 4768
rect 18616 4802 18668 4811
rect 18616 4768 18629 4802
rect 18629 4768 18663 4802
rect 18663 4768 18668 4802
rect 18616 4759 18668 4768
rect 18680 4802 18732 4811
rect 18744 4802 18796 4811
rect 18808 4802 18860 4811
rect 18872 4802 18924 4811
rect 18936 4802 18988 4811
rect 19000 4802 19052 4811
rect 19064 4802 19116 4811
rect 18680 4768 18701 4802
rect 18701 4768 18732 4802
rect 18744 4768 18773 4802
rect 18773 4768 18796 4802
rect 18808 4768 18845 4802
rect 18845 4768 18860 4802
rect 18872 4768 18879 4802
rect 18879 4768 18917 4802
rect 18917 4768 18924 4802
rect 18936 4768 18951 4802
rect 18951 4768 18988 4802
rect 19000 4768 19023 4802
rect 19023 4768 19052 4802
rect 19064 4768 19095 4802
rect 19095 4768 19116 4802
rect 18680 4759 18732 4768
rect 18744 4759 18796 4768
rect 18808 4759 18860 4768
rect 18872 4759 18924 4768
rect 18936 4759 18988 4768
rect 19000 4759 19052 4768
rect 19064 4759 19116 4768
rect 19128 4802 19180 4811
rect 19342 4802 19394 4811
rect 19128 4768 19133 4802
rect 19133 4768 19167 4802
rect 19167 4768 19180 4802
rect 19342 4768 19349 4802
rect 19349 4768 19383 4802
rect 19383 4768 19394 4802
rect 19128 4759 19180 4768
rect 19342 4759 19394 4768
rect 19406 4802 19458 4811
rect 19406 4768 19421 4802
rect 19421 4768 19455 4802
rect 19455 4768 19458 4802
rect 19406 4759 19458 4768
rect 19470 4802 19522 4811
rect 19534 4802 19586 4811
rect 19598 4802 19650 4811
rect 19662 4802 19714 4811
rect 19726 4802 19778 4811
rect 19790 4802 19842 4811
rect 19854 4802 19906 4811
rect 19470 4768 19493 4802
rect 19493 4768 19522 4802
rect 19534 4768 19565 4802
rect 19565 4768 19586 4802
rect 19598 4768 19599 4802
rect 19599 4768 19637 4802
rect 19637 4768 19650 4802
rect 19662 4768 19671 4802
rect 19671 4768 19709 4802
rect 19709 4768 19714 4802
rect 19726 4768 19743 4802
rect 19743 4768 19778 4802
rect 19790 4768 19815 4802
rect 19815 4768 19842 4802
rect 19854 4768 19887 4802
rect 19887 4768 19906 4802
rect 19470 4759 19522 4768
rect 19534 4759 19586 4768
rect 19598 4759 19650 4768
rect 19662 4759 19714 4768
rect 19726 4759 19778 4768
rect 19790 4759 19842 4768
rect 19854 4759 19906 4768
rect 19918 4802 19970 4811
rect 19918 4768 19925 4802
rect 19925 4768 19959 4802
rect 19959 4768 19970 4802
rect 19918 4759 19970 4768
rect 19982 4802 20034 4811
rect 19982 4768 19997 4802
rect 19997 4768 20031 4802
rect 20031 4768 20034 4802
rect 19982 4759 20034 4768
rect 18407 4713 18416 4735
rect 18416 4713 18450 4735
rect 18450 4713 18459 4735
rect 18207 4663 18259 4701
rect 18207 4649 18216 4663
rect 18216 4649 18250 4663
rect 18250 4649 18259 4663
rect 18407 4663 18459 4701
rect 18407 4649 18416 4663
rect 18416 4649 18450 4663
rect 18450 4649 18459 4663
rect 18207 4629 18216 4637
rect 18216 4629 18250 4637
rect 18250 4629 18259 4637
rect 18207 4591 18259 4629
rect 18207 4585 18216 4591
rect 18216 4585 18250 4591
rect 18250 4585 18259 4591
rect 18407 4629 18416 4637
rect 18416 4629 18450 4637
rect 18450 4629 18459 4637
rect 18407 4591 18459 4629
rect 18407 4585 18416 4591
rect 18416 4585 18450 4591
rect 18450 4585 18459 4591
rect 18207 4557 18216 4573
rect 18216 4557 18250 4573
rect 18250 4557 18259 4573
rect 18207 4521 18259 4557
rect 18407 4557 18416 4573
rect 18416 4557 18450 4573
rect 18450 4557 18459 4573
rect 18407 4521 18459 4557
rect 18207 4485 18216 4509
rect 18216 4485 18250 4509
rect 18250 4485 18259 4509
rect 18207 4457 18259 4485
rect 18407 4485 18416 4509
rect 18416 4485 18450 4509
rect 18450 4485 18459 4509
rect 18407 4457 18459 4485
rect 18207 4413 18216 4445
rect 18216 4413 18250 4445
rect 18250 4413 18259 4445
rect 18207 4393 18259 4413
rect 18407 4413 18416 4445
rect 18416 4413 18450 4445
rect 18450 4413 18459 4445
rect 18407 4393 18459 4413
rect 18207 4375 18259 4381
rect 18207 4341 18216 4375
rect 18216 4341 18250 4375
rect 18250 4341 18259 4375
rect 18207 4329 18259 4341
rect 18407 4375 18459 4381
rect 18407 4341 18416 4375
rect 18416 4341 18450 4375
rect 18450 4341 18459 4375
rect 18407 4329 18459 4341
rect 18207 4303 18259 4317
rect 18207 4269 18216 4303
rect 18216 4269 18250 4303
rect 18250 4269 18259 4303
rect 18207 4265 18259 4269
rect 18407 4303 18459 4317
rect 18407 4269 18416 4303
rect 18416 4269 18450 4303
rect 18450 4269 18459 4303
rect 18407 4265 18459 4269
rect 18207 4231 18259 4253
rect 18207 4201 18216 4231
rect 18216 4201 18250 4231
rect 18250 4201 18259 4231
rect 18407 4231 18459 4253
rect 18407 4201 18416 4231
rect 18416 4201 18450 4231
rect 18450 4201 18459 4231
rect 18207 4159 18259 4189
rect 18207 4137 18216 4159
rect 18216 4137 18250 4159
rect 18250 4137 18259 4159
rect 18407 4159 18459 4189
rect 18407 4137 18416 4159
rect 18416 4137 18450 4159
rect 18450 4137 18459 4159
rect 18207 3909 18216 3931
rect 18216 3909 18250 3931
rect 18250 3909 18259 3931
rect 18207 3879 18259 3909
rect 18407 3909 18416 3931
rect 18416 3909 18450 3931
rect 18450 3909 18459 3931
rect 18407 3879 18459 3909
rect 18207 3837 18216 3867
rect 18216 3837 18250 3867
rect 18250 3837 18259 3867
rect 18207 3815 18259 3837
rect 18407 3837 18416 3867
rect 18416 3837 18450 3867
rect 18450 3837 18459 3867
rect 18407 3815 18459 3837
rect 18207 3799 18259 3803
rect 18207 3765 18216 3799
rect 18216 3765 18250 3799
rect 18250 3765 18259 3799
rect 18207 3751 18259 3765
rect 18407 3799 18459 3803
rect 18407 3765 18416 3799
rect 18416 3765 18450 3799
rect 18450 3765 18459 3799
rect 18407 3751 18459 3765
rect 18207 3727 18259 3739
rect 18207 3693 18216 3727
rect 18216 3693 18250 3727
rect 18250 3693 18259 3727
rect 18207 3687 18259 3693
rect 18407 3727 18459 3739
rect 18407 3693 18416 3727
rect 18416 3693 18450 3727
rect 18450 3693 18459 3727
rect 18407 3687 18459 3693
rect 18207 3655 18259 3675
rect 18207 3623 18216 3655
rect 18216 3623 18250 3655
rect 18250 3623 18259 3655
rect 18407 3655 18459 3675
rect 18407 3623 18416 3655
rect 18416 3623 18450 3655
rect 18450 3623 18459 3655
rect 18207 3583 18259 3611
rect 18207 3559 18216 3583
rect 18216 3559 18250 3583
rect 18250 3559 18259 3583
rect 18407 3583 18459 3611
rect 18407 3559 18416 3583
rect 18416 3559 18450 3583
rect 18450 3559 18459 3583
rect 18207 3511 18259 3547
rect 18207 3495 18216 3511
rect 18216 3495 18250 3511
rect 18250 3495 18259 3511
rect 18407 3511 18459 3547
rect 18407 3495 18416 3511
rect 18416 3495 18450 3511
rect 18450 3495 18459 3511
rect 18207 3477 18216 3483
rect 18216 3477 18250 3483
rect 18250 3477 18259 3483
rect 18207 3439 18259 3477
rect 18207 3431 18216 3439
rect 18216 3431 18250 3439
rect 18250 3431 18259 3439
rect 18407 3477 18416 3483
rect 18416 3477 18450 3483
rect 18450 3477 18459 3483
rect 18407 3439 18459 3477
rect 18407 3431 18416 3439
rect 18416 3431 18450 3439
rect 18450 3431 18459 3439
rect 18207 3405 18216 3419
rect 18216 3405 18250 3419
rect 18250 3405 18259 3419
rect 18207 3367 18259 3405
rect 18407 3405 18416 3419
rect 18416 3405 18450 3419
rect 18450 3405 18459 3419
rect 18407 3367 18459 3405
rect 18207 3333 18216 3355
rect 18216 3333 18250 3355
rect 18250 3333 18259 3355
rect 16638 3300 16690 3309
rect 16638 3266 16669 3300
rect 16669 3266 16690 3300
rect 16638 3257 16690 3266
rect 16702 3300 16754 3309
rect 16702 3266 16707 3300
rect 16707 3266 16741 3300
rect 16741 3266 16754 3300
rect 16702 3257 16754 3266
rect 16766 3300 16818 3309
rect 16766 3266 16779 3300
rect 16779 3266 16813 3300
rect 16813 3266 16818 3300
rect 16766 3257 16818 3266
rect 16830 3300 16882 3309
rect 16894 3300 16946 3309
rect 16958 3300 17010 3309
rect 17022 3300 17074 3309
rect 17086 3300 17138 3309
rect 17150 3300 17202 3309
rect 17214 3300 17266 3309
rect 16830 3266 16851 3300
rect 16851 3266 16882 3300
rect 16894 3266 16923 3300
rect 16923 3266 16946 3300
rect 16958 3266 16995 3300
rect 16995 3266 17010 3300
rect 17022 3266 17029 3300
rect 17029 3266 17067 3300
rect 17067 3266 17074 3300
rect 17086 3266 17101 3300
rect 17101 3266 17138 3300
rect 17150 3266 17173 3300
rect 17173 3266 17202 3300
rect 17214 3266 17245 3300
rect 17245 3266 17266 3300
rect 16830 3257 16882 3266
rect 16894 3257 16946 3266
rect 16958 3257 17010 3266
rect 17022 3257 17074 3266
rect 17086 3257 17138 3266
rect 17150 3257 17202 3266
rect 17214 3257 17266 3266
rect 17278 3300 17330 3309
rect 17492 3300 17544 3309
rect 17278 3266 17283 3300
rect 17283 3266 17317 3300
rect 17317 3266 17330 3300
rect 17492 3266 17499 3300
rect 17499 3266 17533 3300
rect 17533 3266 17544 3300
rect 17278 3257 17330 3266
rect 17492 3257 17544 3266
rect 17556 3300 17608 3309
rect 17556 3266 17571 3300
rect 17571 3266 17605 3300
rect 17605 3266 17608 3300
rect 17556 3257 17608 3266
rect 17620 3300 17672 3309
rect 17684 3300 17736 3309
rect 17748 3300 17800 3309
rect 17812 3300 17864 3309
rect 17876 3300 17928 3309
rect 17940 3300 17992 3309
rect 18004 3300 18056 3309
rect 17620 3266 17643 3300
rect 17643 3266 17672 3300
rect 17684 3266 17715 3300
rect 17715 3266 17736 3300
rect 17748 3266 17749 3300
rect 17749 3266 17787 3300
rect 17787 3266 17800 3300
rect 17812 3266 17821 3300
rect 17821 3266 17859 3300
rect 17859 3266 17864 3300
rect 17876 3266 17893 3300
rect 17893 3266 17928 3300
rect 17940 3266 17965 3300
rect 17965 3266 17992 3300
rect 18004 3266 18037 3300
rect 18037 3266 18056 3300
rect 17620 3257 17672 3266
rect 17684 3257 17736 3266
rect 17748 3257 17800 3266
rect 17812 3257 17864 3266
rect 17876 3257 17928 3266
rect 17940 3257 17992 3266
rect 18004 3257 18056 3266
rect 18068 3300 18120 3309
rect 18068 3266 18075 3300
rect 18075 3266 18109 3300
rect 18109 3266 18120 3300
rect 18068 3257 18120 3266
rect 18132 3300 18184 3309
rect 18207 3303 18259 3333
rect 18407 3333 18416 3355
rect 18416 3333 18450 3355
rect 18450 3333 18459 3355
rect 18407 3303 18459 3333
rect 19232 4666 19284 4718
rect 19232 4602 19284 4654
rect 19232 4538 19284 4590
rect 19232 4474 19284 4526
rect 19232 4410 19284 4462
rect 19232 4346 19284 4398
rect 19232 4282 19284 4334
rect 19232 4218 19284 4270
rect 19232 4154 19284 4206
rect 19232 4090 19284 4142
rect 18505 4008 18557 4060
rect 18569 4008 18621 4060
rect 18633 4008 18685 4060
rect 18697 4008 18749 4060
rect 18761 4008 18813 4060
rect 18825 4008 18877 4060
rect 18889 4008 18941 4060
rect 18953 4008 19005 4060
rect 19017 4008 19069 4060
rect 19081 4008 19133 4060
rect 19145 4008 19197 4060
rect 19319 4008 19371 4060
rect 19383 4008 19435 4060
rect 19447 4008 19499 4060
rect 19511 4008 19563 4060
rect 19575 4008 19627 4060
rect 19639 4008 19691 4060
rect 19703 4008 19755 4060
rect 19767 4008 19819 4060
rect 19831 4008 19883 4060
rect 19895 4008 19947 4060
rect 19959 4008 20011 4060
rect 19232 3926 19284 3978
rect 19232 3862 19284 3914
rect 19232 3798 19284 3850
rect 19232 3734 19284 3786
rect 19232 3670 19284 3722
rect 19232 3606 19284 3658
rect 19232 3542 19284 3594
rect 19232 3478 19284 3530
rect 19232 3414 19284 3466
rect 19232 3350 19284 3402
rect 20057 4735 20109 4765
rect 20057 4713 20066 4735
rect 20066 4713 20100 4735
rect 20100 4713 20109 4735
rect 20057 4663 20109 4701
rect 20057 4649 20066 4663
rect 20066 4649 20100 4663
rect 20100 4649 20109 4663
rect 20057 4629 20066 4637
rect 20066 4629 20100 4637
rect 20100 4629 20109 4637
rect 20057 4591 20109 4629
rect 20057 4585 20066 4591
rect 20066 4585 20100 4591
rect 20100 4585 20109 4591
rect 20057 4557 20066 4573
rect 20066 4557 20100 4573
rect 20100 4557 20109 4573
rect 20057 4521 20109 4557
rect 20057 4485 20066 4509
rect 20066 4485 20100 4509
rect 20100 4485 20109 4509
rect 20057 4457 20109 4485
rect 20057 4413 20066 4445
rect 20066 4413 20100 4445
rect 20100 4413 20109 4445
rect 20057 4393 20109 4413
rect 20057 4375 20109 4381
rect 20057 4341 20066 4375
rect 20066 4341 20100 4375
rect 20100 4341 20109 4375
rect 20057 4329 20109 4341
rect 20057 4303 20109 4317
rect 20057 4269 20066 4303
rect 20066 4269 20100 4303
rect 20100 4269 20109 4303
rect 20057 4265 20109 4269
rect 20057 4231 20109 4253
rect 20057 4201 20066 4231
rect 20066 4201 20100 4231
rect 20100 4201 20109 4231
rect 20057 4159 20109 4189
rect 20057 4137 20066 4159
rect 20066 4137 20100 4159
rect 20100 4137 20109 4159
rect 20057 3909 20066 3931
rect 20066 3909 20100 3931
rect 20100 3909 20109 3931
rect 20057 3879 20109 3909
rect 20057 3837 20066 3867
rect 20066 3837 20100 3867
rect 20100 3837 20109 3867
rect 20057 3815 20109 3837
rect 20057 3799 20109 3803
rect 20057 3765 20066 3799
rect 20066 3765 20100 3799
rect 20100 3765 20109 3799
rect 20057 3751 20109 3765
rect 20057 3727 20109 3739
rect 20057 3693 20066 3727
rect 20066 3693 20100 3727
rect 20100 3693 20109 3727
rect 20057 3687 20109 3693
rect 20057 3655 20109 3675
rect 20057 3623 20066 3655
rect 20066 3623 20100 3655
rect 20100 3623 20109 3655
rect 20057 3583 20109 3611
rect 20057 3559 20066 3583
rect 20066 3559 20100 3583
rect 20100 3559 20109 3583
rect 20057 3511 20109 3547
rect 20057 3495 20066 3511
rect 20066 3495 20100 3511
rect 20100 3495 20109 3511
rect 20057 3477 20066 3483
rect 20066 3477 20100 3483
rect 20100 3477 20109 3483
rect 20057 3439 20109 3477
rect 20057 3431 20066 3439
rect 20066 3431 20100 3439
rect 20100 3431 20109 3439
rect 20057 3405 20066 3419
rect 20066 3405 20100 3419
rect 20100 3405 20109 3419
rect 20057 3367 20109 3405
rect 20057 3333 20066 3355
rect 20066 3333 20100 3355
rect 20100 3333 20109 3355
rect 18488 3300 18540 3309
rect 18132 3266 18147 3300
rect 18147 3266 18181 3300
rect 18181 3266 18184 3300
rect 18488 3266 18519 3300
rect 18519 3266 18540 3300
rect 18132 3257 18184 3266
rect 18488 3257 18540 3266
rect 18552 3300 18604 3309
rect 18552 3266 18557 3300
rect 18557 3266 18591 3300
rect 18591 3266 18604 3300
rect 18552 3257 18604 3266
rect 18616 3300 18668 3309
rect 18616 3266 18629 3300
rect 18629 3266 18663 3300
rect 18663 3266 18668 3300
rect 18616 3257 18668 3266
rect 18680 3300 18732 3309
rect 18744 3300 18796 3309
rect 18808 3300 18860 3309
rect 18872 3300 18924 3309
rect 18936 3300 18988 3309
rect 19000 3300 19052 3309
rect 19064 3300 19116 3309
rect 18680 3266 18701 3300
rect 18701 3266 18732 3300
rect 18744 3266 18773 3300
rect 18773 3266 18796 3300
rect 18808 3266 18845 3300
rect 18845 3266 18860 3300
rect 18872 3266 18879 3300
rect 18879 3266 18917 3300
rect 18917 3266 18924 3300
rect 18936 3266 18951 3300
rect 18951 3266 18988 3300
rect 19000 3266 19023 3300
rect 19023 3266 19052 3300
rect 19064 3266 19095 3300
rect 19095 3266 19116 3300
rect 18680 3257 18732 3266
rect 18744 3257 18796 3266
rect 18808 3257 18860 3266
rect 18872 3257 18924 3266
rect 18936 3257 18988 3266
rect 19000 3257 19052 3266
rect 19064 3257 19116 3266
rect 19128 3300 19180 3309
rect 19342 3300 19394 3309
rect 19128 3266 19133 3300
rect 19133 3266 19167 3300
rect 19167 3266 19180 3300
rect 19342 3266 19349 3300
rect 19349 3266 19383 3300
rect 19383 3266 19394 3300
rect 19128 3257 19180 3266
rect 19342 3257 19394 3266
rect 19406 3300 19458 3309
rect 19406 3266 19421 3300
rect 19421 3266 19455 3300
rect 19455 3266 19458 3300
rect 19406 3257 19458 3266
rect 19470 3300 19522 3309
rect 19534 3300 19586 3309
rect 19598 3300 19650 3309
rect 19662 3300 19714 3309
rect 19726 3300 19778 3309
rect 19790 3300 19842 3309
rect 19854 3300 19906 3309
rect 19470 3266 19493 3300
rect 19493 3266 19522 3300
rect 19534 3266 19565 3300
rect 19565 3266 19586 3300
rect 19598 3266 19599 3300
rect 19599 3266 19637 3300
rect 19637 3266 19650 3300
rect 19662 3266 19671 3300
rect 19671 3266 19709 3300
rect 19709 3266 19714 3300
rect 19726 3266 19743 3300
rect 19743 3266 19778 3300
rect 19790 3266 19815 3300
rect 19815 3266 19842 3300
rect 19854 3266 19887 3300
rect 19887 3266 19906 3300
rect 19470 3257 19522 3266
rect 19534 3257 19586 3266
rect 19598 3257 19650 3266
rect 19662 3257 19714 3266
rect 19726 3257 19778 3266
rect 19790 3257 19842 3266
rect 19854 3257 19906 3266
rect 19918 3300 19970 3309
rect 19918 3266 19925 3300
rect 19925 3266 19959 3300
rect 19959 3266 19970 3300
rect 19918 3257 19970 3266
rect 19982 3300 20034 3309
rect 20057 3303 20109 3333
rect 19982 3266 19997 3300
rect 19997 3266 20031 3300
rect 20031 3266 20034 3300
rect 19982 3257 20034 3266
<< metal2 >>
rect 16550 9863 17353 9868
rect 16550 9861 16648 9863
rect 16704 9861 16728 9863
rect 16784 9861 16808 9863
rect 16864 9861 16888 9863
rect 16944 9861 16968 9863
rect 17024 9861 17048 9863
rect 17104 9861 17128 9863
rect 17184 9861 17208 9863
rect 17264 9861 17288 9863
rect 16550 9815 16638 9861
rect 15300 9300 16500 9800
rect 16200 8300 16500 9300
rect 16550 9764 16557 9815
rect 16609 9809 16638 9815
rect 16882 9809 16888 9861
rect 16946 9809 16958 9861
rect 17202 9809 17208 9861
rect 17266 9809 17278 9861
rect 16609 9807 16648 9809
rect 16704 9807 16728 9809
rect 16784 9807 16808 9809
rect 16864 9807 16888 9809
rect 16944 9807 16968 9809
rect 17024 9807 17048 9809
rect 17104 9807 17128 9809
rect 17184 9807 17208 9809
rect 17264 9807 17288 9809
rect 17344 9807 17353 9863
rect 16609 9802 17353 9807
rect 16609 9764 16616 9802
rect 17381 9774 17435 9868
rect 17463 9863 18266 9868
rect 17463 9807 17472 9863
rect 17528 9861 17552 9863
rect 17608 9861 17632 9863
rect 17688 9861 17712 9863
rect 17768 9861 17792 9863
rect 17848 9861 17872 9863
rect 17928 9861 17952 9863
rect 18008 9861 18032 9863
rect 18088 9861 18112 9863
rect 18168 9861 18266 9863
rect 17544 9809 17552 9861
rect 17608 9809 17620 9861
rect 17864 9809 17872 9861
rect 17928 9809 17940 9861
rect 18184 9860 18266 9861
rect 18400 9863 19203 9868
rect 18400 9861 18498 9863
rect 18554 9861 18578 9863
rect 18634 9861 18658 9863
rect 18714 9861 18738 9863
rect 18794 9861 18818 9863
rect 18874 9861 18898 9863
rect 18954 9861 18978 9863
rect 19034 9861 19058 9863
rect 19114 9861 19138 9863
rect 18400 9860 18488 9861
rect 18184 9815 18488 9860
rect 18184 9809 18207 9815
rect 17528 9807 17552 9809
rect 17608 9807 17632 9809
rect 17688 9807 17712 9809
rect 17768 9807 17792 9809
rect 17848 9807 17872 9809
rect 17928 9807 17952 9809
rect 18008 9807 18032 9809
rect 18088 9807 18112 9809
rect 18168 9807 18207 9809
rect 17463 9802 18207 9807
rect 16550 9708 16555 9764
rect 16611 9718 16616 9764
rect 16644 9768 18172 9774
rect 16644 9746 17382 9768
rect 16611 9708 17352 9718
rect 16550 9699 16557 9708
rect 16609 9699 17352 9708
rect 16550 9690 17352 9699
rect 17380 9716 17382 9746
rect 17434 9746 18172 9768
rect 18200 9764 18207 9802
rect 18259 9764 18407 9815
rect 18459 9809 18488 9815
rect 18732 9809 18738 9861
rect 18796 9809 18808 9861
rect 19052 9809 19058 9861
rect 19116 9809 19128 9861
rect 18459 9807 18498 9809
rect 18554 9807 18578 9809
rect 18634 9807 18658 9809
rect 18714 9807 18738 9809
rect 18794 9807 18818 9809
rect 18874 9807 18898 9809
rect 18954 9807 18978 9809
rect 19034 9807 19058 9809
rect 19114 9807 19138 9809
rect 19194 9807 19203 9863
rect 18459 9802 19203 9807
rect 18459 9764 18466 9802
rect 19231 9774 19285 9868
rect 19313 9863 20116 9868
rect 19313 9807 19322 9863
rect 19378 9861 19402 9863
rect 19458 9861 19482 9863
rect 19538 9861 19562 9863
rect 19618 9861 19642 9863
rect 19698 9861 19722 9863
rect 19778 9861 19802 9863
rect 19858 9861 19882 9863
rect 19938 9861 19962 9863
rect 20018 9861 20116 9863
rect 19394 9809 19402 9861
rect 19458 9809 19470 9861
rect 19714 9809 19722 9861
rect 19778 9809 19790 9861
rect 20034 9815 20116 9861
rect 20034 9809 20057 9815
rect 19378 9807 19402 9809
rect 19458 9807 19482 9809
rect 19538 9807 19562 9809
rect 19618 9807 19642 9809
rect 19698 9807 19722 9809
rect 19778 9807 19802 9809
rect 19858 9807 19882 9809
rect 19938 9807 19962 9809
rect 20018 9807 20057 9809
rect 19313 9802 20057 9807
rect 17434 9716 17436 9746
rect 18200 9718 18205 9764
rect 17380 9704 17436 9716
rect 16550 9687 16616 9690
rect 16550 9684 16557 9687
rect 16609 9684 16616 9687
rect 16550 9628 16555 9684
rect 16611 9628 16616 9684
rect 17380 9662 17382 9704
rect 16644 9652 17382 9662
rect 17434 9662 17436 9704
rect 17464 9708 18205 9718
rect 18261 9708 18405 9764
rect 18461 9718 18466 9764
rect 18494 9768 20022 9774
rect 18494 9746 19232 9768
rect 18461 9708 19202 9718
rect 17464 9699 18207 9708
rect 18259 9699 18407 9708
rect 18459 9699 19202 9708
rect 17464 9690 19202 9699
rect 19230 9716 19232 9746
rect 19284 9746 20022 9768
rect 20050 9764 20057 9802
rect 20109 9764 20116 9815
rect 19284 9716 19286 9746
rect 20050 9718 20055 9764
rect 19230 9704 19286 9716
rect 18200 9687 18466 9690
rect 18200 9684 18207 9687
rect 18259 9684 18407 9687
rect 18459 9684 18466 9687
rect 17434 9652 18172 9662
rect 16644 9640 18172 9652
rect 16644 9634 17382 9640
rect 16550 9623 16616 9628
rect 16550 9604 16557 9623
rect 16609 9606 16616 9623
rect 16609 9604 17352 9606
rect 16550 9548 16555 9604
rect 16611 9578 17352 9604
rect 17380 9588 17382 9634
rect 17434 9634 18172 9640
rect 17434 9588 17436 9634
rect 18200 9628 18205 9684
rect 18261 9628 18405 9684
rect 18461 9628 18466 9684
rect 19230 9662 19232 9704
rect 18494 9652 19232 9662
rect 19284 9662 19286 9704
rect 19314 9708 20055 9718
rect 20111 9708 20116 9764
rect 19314 9699 20057 9708
rect 20109 9699 20116 9708
rect 19314 9690 20116 9699
rect 20050 9687 20116 9690
rect 20050 9684 20057 9687
rect 20109 9684 20116 9687
rect 19284 9652 20022 9662
rect 18494 9640 20022 9652
rect 18494 9634 19232 9640
rect 18200 9623 18466 9628
rect 18200 9606 18207 9623
rect 16611 9548 16616 9578
rect 17380 9576 17436 9588
rect 17464 9604 18207 9606
rect 18259 9604 18407 9623
rect 18459 9606 18466 9623
rect 18459 9604 19202 9606
rect 17464 9578 18205 9604
rect 17380 9550 17382 9576
rect 16550 9524 16557 9548
rect 16609 9524 16616 9548
rect 16550 9468 16555 9524
rect 16611 9494 16616 9524
rect 16644 9524 17382 9550
rect 17434 9550 17436 9576
rect 17434 9524 18172 9550
rect 16644 9522 18172 9524
rect 18200 9548 18205 9578
rect 18261 9548 18405 9604
rect 18461 9578 19202 9604
rect 19230 9588 19232 9634
rect 19284 9634 20022 9640
rect 19284 9588 19286 9634
rect 20050 9628 20055 9684
rect 20111 9628 20116 9684
rect 20050 9623 20116 9628
rect 20050 9606 20057 9623
rect 18461 9548 18466 9578
rect 19230 9576 19286 9588
rect 19314 9604 20057 9606
rect 20109 9604 20116 9623
rect 19314 9578 20055 9604
rect 19230 9550 19232 9576
rect 18200 9524 18207 9548
rect 18259 9524 18407 9548
rect 18459 9524 18466 9548
rect 17380 9512 17436 9522
rect 16611 9468 17352 9494
rect 16550 9444 16557 9468
rect 16609 9466 17352 9468
rect 16609 9444 16616 9466
rect 16550 9388 16555 9444
rect 16611 9388 16616 9444
rect 17380 9460 17382 9512
rect 17434 9460 17436 9512
rect 18200 9494 18205 9524
rect 17464 9468 18205 9494
rect 18261 9468 18405 9524
rect 18461 9494 18466 9524
rect 18494 9524 19232 9550
rect 19284 9550 19286 9576
rect 19284 9524 20022 9550
rect 18494 9522 20022 9524
rect 20050 9548 20055 9578
rect 20111 9548 20116 9604
rect 20050 9524 20057 9548
rect 20109 9524 20116 9548
rect 19230 9512 19286 9522
rect 18461 9468 19202 9494
rect 17464 9466 18207 9468
rect 17380 9448 17436 9460
rect 17380 9438 17382 9448
rect 16644 9410 17382 9438
rect 16550 9379 16557 9388
rect 16609 9382 16616 9388
rect 17380 9396 17382 9410
rect 17434 9438 17436 9448
rect 18200 9444 18207 9466
rect 18259 9444 18407 9468
rect 18459 9466 19202 9468
rect 18459 9444 18466 9466
rect 17434 9410 18172 9438
rect 17434 9396 17436 9410
rect 17380 9384 17436 9396
rect 16609 9379 17352 9382
rect 16550 9367 17352 9379
rect 16550 9364 16557 9367
rect 16609 9364 17352 9367
rect 16550 9308 16555 9364
rect 16611 9354 17352 9364
rect 16611 9308 16616 9354
rect 17380 9332 17382 9384
rect 17434 9332 17436 9384
rect 18200 9388 18205 9444
rect 18261 9388 18405 9444
rect 18461 9388 18466 9444
rect 19230 9460 19232 9512
rect 19284 9460 19286 9512
rect 20050 9494 20055 9524
rect 19314 9468 20055 9494
rect 20111 9468 20116 9524
rect 19314 9466 20057 9468
rect 19230 9448 19286 9460
rect 19230 9438 19232 9448
rect 18494 9410 19232 9438
rect 18200 9382 18207 9388
rect 17464 9379 18207 9382
rect 18259 9379 18407 9388
rect 18459 9382 18466 9388
rect 19230 9396 19232 9410
rect 19284 9438 19286 9448
rect 20050 9444 20057 9466
rect 20109 9444 20116 9468
rect 19284 9410 20022 9438
rect 19284 9396 19286 9410
rect 19230 9384 19286 9396
rect 18459 9379 19202 9382
rect 17464 9367 19202 9379
rect 17464 9364 18207 9367
rect 18259 9364 18407 9367
rect 18459 9364 19202 9367
rect 17464 9354 18205 9364
rect 17380 9326 17436 9332
rect 16550 9303 16616 9308
rect 16550 9284 16557 9303
rect 16609 9284 16616 9303
rect 16644 9320 18172 9326
rect 16644 9298 17382 9320
rect 16550 9228 16555 9284
rect 16611 9270 16616 9284
rect 16611 9242 17352 9270
rect 17380 9268 17382 9298
rect 17434 9298 18172 9320
rect 18200 9308 18205 9354
rect 18261 9308 18405 9364
rect 18461 9354 19202 9364
rect 18461 9308 18466 9354
rect 19230 9332 19232 9384
rect 19284 9332 19286 9384
rect 20050 9388 20055 9444
rect 20111 9388 20116 9444
rect 20050 9382 20057 9388
rect 19314 9379 20057 9382
rect 20109 9379 20116 9388
rect 19314 9367 20116 9379
rect 19314 9364 20057 9367
rect 20109 9364 20116 9367
rect 19314 9354 20055 9364
rect 19230 9326 19286 9332
rect 18200 9303 18466 9308
rect 17434 9268 17436 9298
rect 18200 9284 18207 9303
rect 18259 9284 18407 9303
rect 18459 9284 18466 9303
rect 18494 9320 20022 9326
rect 18494 9298 19232 9320
rect 18200 9270 18205 9284
rect 17380 9256 17436 9268
rect 16611 9228 16616 9242
rect 16550 9204 16557 9228
rect 16609 9204 16616 9228
rect 17380 9214 17382 9256
rect 16550 9148 16555 9204
rect 16611 9148 16616 9204
rect 16550 9139 16616 9148
rect 16644 9204 17382 9214
rect 17434 9214 17436 9256
rect 17464 9242 18205 9270
rect 18200 9228 18205 9242
rect 18261 9228 18405 9284
rect 18461 9270 18466 9284
rect 18461 9242 19202 9270
rect 19230 9268 19232 9298
rect 19284 9298 20022 9320
rect 20050 9308 20055 9354
rect 20111 9308 20116 9364
rect 20050 9303 20116 9308
rect 19284 9268 19286 9298
rect 20050 9284 20057 9303
rect 20109 9284 20116 9303
rect 20050 9270 20055 9284
rect 19230 9256 19286 9268
rect 18461 9228 18466 9242
rect 17434 9204 18172 9214
rect 16644 9192 18172 9204
rect 16644 9140 17382 9192
rect 17434 9140 18172 9192
rect 18200 9204 18207 9228
rect 18259 9204 18407 9228
rect 18459 9204 18466 9228
rect 19230 9214 19232 9256
rect 18200 9148 18205 9204
rect 18261 9148 18405 9204
rect 18461 9148 18466 9204
rect 17380 9112 17436 9140
rect 18200 9139 18466 9148
rect 18494 9204 19232 9214
rect 19284 9214 19286 9256
rect 19314 9242 20055 9270
rect 20050 9228 20055 9242
rect 20111 9228 20116 9284
rect 19284 9204 20022 9214
rect 18494 9192 20022 9204
rect 18494 9140 19232 9192
rect 19284 9140 20022 9192
rect 20050 9204 20057 9228
rect 20109 9204 20116 9228
rect 20050 9148 20055 9204
rect 20111 9148 20116 9204
rect 19230 9112 19286 9140
rect 20050 9139 20116 9148
rect 16624 9111 16740 9112
rect 16550 9110 16740 9111
rect 16796 9110 16820 9112
rect 16876 9110 16900 9112
rect 16956 9110 16980 9112
rect 17036 9110 17060 9112
rect 17116 9110 17140 9112
rect 17196 9110 17220 9112
rect 17276 9110 17300 9112
rect 16550 9058 16655 9110
rect 16707 9058 16719 9110
rect 16899 9058 16900 9110
rect 16963 9058 16975 9110
rect 17036 9058 17039 9110
rect 17219 9058 17220 9110
rect 17283 9058 17295 9110
rect 16550 9057 16740 9058
rect 16624 9056 16740 9057
rect 16796 9056 16820 9058
rect 16876 9056 16900 9058
rect 16956 9056 16980 9058
rect 17036 9056 17060 9058
rect 17116 9056 17140 9058
rect 17196 9056 17220 9058
rect 17276 9056 17300 9058
rect 17356 9056 17380 9112
rect 17436 9056 17460 9112
rect 17516 9110 17540 9112
rect 17596 9110 17620 9112
rect 17676 9110 17700 9112
rect 17756 9110 17780 9112
rect 17836 9110 17860 9112
rect 17916 9110 17940 9112
rect 17996 9110 18020 9112
rect 18076 9111 18192 9112
rect 18474 9111 18590 9112
rect 18076 9110 18590 9111
rect 18646 9110 18670 9112
rect 18726 9110 18750 9112
rect 18806 9110 18830 9112
rect 18886 9110 18910 9112
rect 18966 9110 18990 9112
rect 19046 9110 19070 9112
rect 19126 9110 19150 9112
rect 17521 9058 17533 9110
rect 17596 9058 17597 9110
rect 17777 9058 17780 9110
rect 17841 9058 17853 9110
rect 17916 9058 17917 9110
rect 18097 9058 18109 9110
rect 18161 9058 18505 9110
rect 18557 9058 18569 9110
rect 18749 9058 18750 9110
rect 18813 9058 18825 9110
rect 18886 9058 18889 9110
rect 19069 9058 19070 9110
rect 19133 9058 19145 9110
rect 17516 9056 17540 9058
rect 17596 9056 17620 9058
rect 17676 9056 17700 9058
rect 17756 9056 17780 9058
rect 17836 9056 17860 9058
rect 17916 9056 17940 9058
rect 17996 9056 18020 9058
rect 18076 9057 18590 9058
rect 18076 9056 18192 9057
rect 16550 9020 16616 9029
rect 17380 9028 17436 9056
rect 16550 8964 16555 9020
rect 16611 8964 16616 9020
rect 16550 8940 16557 8964
rect 16609 8940 16616 8964
rect 16644 8976 17382 9028
rect 17434 8976 18172 9028
rect 16644 8964 18172 8976
rect 16644 8954 17382 8964
rect 16550 8884 16555 8940
rect 16611 8926 16616 8940
rect 16611 8898 17352 8926
rect 17380 8912 17382 8954
rect 17434 8954 18172 8964
rect 18200 9020 18266 9029
rect 18200 8964 18205 9020
rect 18261 8964 18266 9020
rect 17434 8912 17436 8954
rect 18200 8940 18207 8964
rect 18259 8940 18266 8964
rect 18200 8926 18205 8940
rect 17380 8900 17436 8912
rect 16611 8884 16616 8898
rect 16550 8865 16557 8884
rect 16609 8865 16616 8884
rect 17380 8870 17382 8900
rect 16550 8860 16616 8865
rect 16550 8804 16555 8860
rect 16611 8814 16616 8860
rect 16644 8848 17382 8870
rect 17434 8870 17436 8900
rect 17464 8898 18205 8926
rect 18200 8884 18205 8898
rect 18261 8884 18266 8940
rect 17434 8848 18172 8870
rect 16644 8842 18172 8848
rect 18200 8865 18207 8884
rect 18259 8865 18266 8884
rect 18200 8860 18266 8865
rect 17380 8836 17436 8842
rect 16611 8804 17352 8814
rect 16550 8801 16557 8804
rect 16609 8801 17352 8804
rect 16550 8789 17352 8801
rect 16550 8780 16557 8789
rect 16609 8786 17352 8789
rect 16609 8780 16616 8786
rect 16550 8724 16555 8780
rect 16611 8724 16616 8780
rect 17380 8784 17382 8836
rect 17434 8784 17436 8836
rect 18200 8814 18205 8860
rect 17464 8804 18205 8814
rect 18261 8804 18266 8860
rect 17464 8801 18207 8804
rect 18259 8801 18266 8804
rect 17464 8789 18266 8801
rect 17464 8786 18207 8789
rect 17380 8772 17436 8784
rect 17380 8758 17382 8772
rect 16644 8730 17382 8758
rect 16550 8700 16557 8724
rect 16609 8702 16616 8724
rect 17380 8720 17382 8730
rect 17434 8758 17436 8772
rect 18200 8780 18207 8786
rect 18259 8780 18266 8789
rect 17434 8730 18172 8758
rect 17434 8720 17436 8730
rect 17380 8708 17436 8720
rect 16609 8700 17352 8702
rect 16550 8644 16555 8700
rect 16611 8674 17352 8700
rect 16611 8644 16616 8674
rect 17380 8656 17382 8708
rect 17434 8656 17436 8708
rect 18200 8724 18205 8780
rect 18261 8724 18266 8780
rect 18200 8702 18207 8724
rect 17464 8700 18207 8702
rect 18259 8700 18266 8724
rect 17464 8674 18205 8700
rect 17380 8646 17436 8656
rect 16550 8620 16557 8644
rect 16609 8620 16616 8644
rect 16550 8564 16555 8620
rect 16611 8590 16616 8620
rect 16644 8644 18172 8646
rect 16644 8618 17382 8644
rect 17380 8592 17382 8618
rect 17434 8618 18172 8644
rect 18200 8644 18205 8674
rect 18261 8644 18266 8700
rect 18200 8620 18207 8644
rect 18259 8620 18266 8644
rect 17434 8592 17436 8618
rect 16611 8564 17352 8590
rect 16550 8545 16557 8564
rect 16609 8562 17352 8564
rect 17380 8580 17436 8592
rect 18200 8590 18205 8620
rect 16609 8545 16616 8562
rect 16550 8540 16616 8545
rect 16550 8484 16555 8540
rect 16611 8484 16616 8540
rect 17380 8534 17382 8580
rect 16644 8528 17382 8534
rect 17434 8534 17436 8580
rect 17464 8564 18205 8590
rect 18261 8564 18266 8620
rect 17464 8562 18207 8564
rect 18200 8545 18207 8562
rect 18259 8545 18266 8564
rect 18200 8540 18266 8545
rect 17434 8528 18172 8534
rect 16644 8516 18172 8528
rect 16644 8506 17382 8516
rect 16550 8481 16557 8484
rect 16609 8481 16616 8484
rect 16550 8478 16616 8481
rect 16550 8469 17352 8478
rect 16550 8460 16557 8469
rect 16609 8460 17352 8469
rect 16550 8404 16555 8460
rect 16611 8450 17352 8460
rect 17380 8464 17382 8506
rect 17434 8506 18172 8516
rect 17434 8464 17436 8506
rect 18200 8484 18205 8540
rect 18261 8484 18266 8540
rect 18200 8481 18207 8484
rect 18259 8481 18266 8484
rect 18200 8478 18266 8481
rect 17380 8452 17436 8464
rect 16611 8404 16616 8450
rect 17380 8422 17382 8452
rect 16550 8353 16557 8404
rect 16609 8366 16616 8404
rect 16644 8400 17382 8422
rect 17434 8422 17436 8452
rect 17464 8469 18266 8478
rect 17464 8460 18207 8469
rect 18259 8460 18266 8469
rect 17464 8450 18205 8460
rect 17434 8400 18172 8422
rect 16644 8394 18172 8400
rect 18200 8404 18205 8450
rect 18261 8404 18266 8460
rect 16609 8361 17353 8366
rect 16609 8359 16648 8361
rect 16704 8359 16728 8361
rect 16784 8359 16808 8361
rect 16864 8359 16888 8361
rect 16944 8359 16968 8361
rect 17024 8359 17048 8361
rect 17104 8359 17128 8361
rect 17184 8359 17208 8361
rect 17264 8359 17288 8361
rect 16609 8353 16638 8359
rect 16550 8307 16638 8353
rect 16882 8307 16888 8359
rect 16946 8307 16958 8359
rect 17202 8307 17208 8359
rect 17266 8307 17278 8359
rect 16550 8305 16648 8307
rect 16704 8305 16728 8307
rect 16784 8305 16808 8307
rect 16864 8305 16888 8307
rect 16944 8305 16968 8307
rect 17024 8305 17048 8307
rect 17104 8305 17128 8307
rect 17184 8305 17208 8307
rect 17264 8305 17288 8307
rect 17344 8305 17353 8361
rect 16550 8300 17353 8305
rect 15800 8250 16500 8300
rect 15800 8220 17290 8250
rect 17381 8220 17435 8394
rect 18200 8366 18207 8404
rect 17463 8361 18207 8366
rect 17463 8305 17472 8361
rect 17528 8359 17552 8361
rect 17608 8359 17632 8361
rect 17688 8359 17712 8361
rect 17768 8359 17792 8361
rect 17848 8359 17872 8361
rect 17928 8359 17952 8361
rect 18008 8359 18032 8361
rect 18088 8359 18112 8361
rect 18168 8359 18207 8361
rect 17544 8307 17552 8359
rect 17608 8307 17620 8359
rect 17864 8307 17872 8359
rect 17928 8307 17940 8359
rect 18184 8353 18207 8359
rect 18259 8353 18266 8404
rect 18184 8307 18266 8353
rect 17528 8305 17552 8307
rect 17608 8305 17632 8307
rect 17688 8305 17712 8307
rect 17768 8305 17792 8307
rect 17848 8305 17872 8307
rect 17928 8305 17952 8307
rect 18008 8305 18032 8307
rect 18088 8305 18112 8307
rect 18168 8305 18266 8307
rect 17463 8300 18266 8305
rect 18300 8220 18370 9057
rect 18474 9056 18590 9057
rect 18646 9056 18670 9058
rect 18726 9056 18750 9058
rect 18806 9056 18830 9058
rect 18886 9056 18910 9058
rect 18966 9056 18990 9058
rect 19046 9056 19070 9058
rect 19126 9056 19150 9058
rect 19206 9056 19230 9112
rect 19286 9056 19310 9112
rect 19366 9110 19390 9112
rect 19446 9110 19470 9112
rect 19526 9110 19550 9112
rect 19606 9110 19630 9112
rect 19686 9110 19710 9112
rect 19766 9110 19790 9112
rect 19846 9110 19870 9112
rect 19926 9111 20042 9112
rect 19926 9110 20230 9111
rect 19371 9058 19383 9110
rect 19446 9058 19447 9110
rect 19627 9058 19630 9110
rect 19691 9058 19703 9110
rect 19766 9058 19767 9110
rect 19947 9058 19959 9110
rect 20011 9058 20230 9110
rect 19366 9056 19390 9058
rect 19446 9056 19470 9058
rect 19526 9056 19550 9058
rect 19606 9056 19630 9058
rect 19686 9056 19710 9058
rect 19766 9056 19790 9058
rect 19846 9056 19870 9058
rect 19926 9057 20230 9058
rect 19926 9056 20042 9057
rect 18400 9020 18466 9029
rect 19230 9028 19286 9056
rect 18400 8964 18405 9020
rect 18461 8964 18466 9020
rect 18400 8940 18407 8964
rect 18459 8940 18466 8964
rect 18494 8976 19232 9028
rect 19284 8976 20022 9028
rect 18494 8964 20022 8976
rect 18494 8954 19232 8964
rect 18400 8884 18405 8940
rect 18461 8926 18466 8940
rect 18461 8898 19202 8926
rect 19230 8912 19232 8954
rect 19284 8954 20022 8964
rect 20050 9020 20116 9029
rect 20050 8964 20055 9020
rect 20111 8964 20116 9020
rect 19284 8912 19286 8954
rect 20050 8940 20057 8964
rect 20109 8940 20116 8964
rect 20050 8926 20055 8940
rect 19230 8900 19286 8912
rect 18461 8884 18466 8898
rect 18400 8865 18407 8884
rect 18459 8865 18466 8884
rect 19230 8870 19232 8900
rect 18400 8860 18466 8865
rect 18400 8804 18405 8860
rect 18461 8814 18466 8860
rect 18494 8848 19232 8870
rect 19284 8870 19286 8900
rect 19314 8898 20055 8926
rect 20050 8884 20055 8898
rect 20111 8884 20116 8940
rect 19284 8848 20022 8870
rect 18494 8842 20022 8848
rect 20050 8865 20057 8884
rect 20109 8865 20116 8884
rect 20050 8860 20116 8865
rect 19230 8836 19286 8842
rect 18461 8804 19202 8814
rect 18400 8801 18407 8804
rect 18459 8801 19202 8804
rect 18400 8789 19202 8801
rect 18400 8780 18407 8789
rect 18459 8786 19202 8789
rect 18459 8780 18466 8786
rect 18400 8724 18405 8780
rect 18461 8724 18466 8780
rect 19230 8784 19232 8836
rect 19284 8784 19286 8836
rect 20050 8814 20055 8860
rect 19314 8804 20055 8814
rect 20111 8804 20116 8860
rect 19314 8801 20057 8804
rect 20109 8801 20116 8804
rect 19314 8789 20116 8801
rect 19314 8786 20057 8789
rect 19230 8772 19286 8784
rect 19230 8758 19232 8772
rect 18494 8730 19232 8758
rect 18400 8700 18407 8724
rect 18459 8702 18466 8724
rect 19230 8720 19232 8730
rect 19284 8758 19286 8772
rect 20050 8780 20057 8786
rect 20109 8780 20116 8789
rect 19284 8730 20022 8758
rect 19284 8720 19286 8730
rect 19230 8708 19286 8720
rect 18459 8700 19202 8702
rect 18400 8644 18405 8700
rect 18461 8674 19202 8700
rect 18461 8644 18466 8674
rect 19230 8656 19232 8708
rect 19284 8656 19286 8708
rect 20050 8724 20055 8780
rect 20111 8724 20116 8780
rect 20050 8702 20057 8724
rect 19314 8700 20057 8702
rect 20109 8700 20116 8724
rect 19314 8674 20055 8700
rect 19230 8646 19286 8656
rect 18400 8620 18407 8644
rect 18459 8620 18466 8644
rect 18400 8564 18405 8620
rect 18461 8590 18466 8620
rect 18494 8644 20022 8646
rect 18494 8618 19232 8644
rect 19230 8592 19232 8618
rect 19284 8618 20022 8644
rect 20050 8644 20055 8674
rect 20111 8644 20116 8700
rect 20050 8620 20057 8644
rect 20109 8620 20116 8644
rect 19284 8592 19286 8618
rect 18461 8564 19202 8590
rect 18400 8545 18407 8564
rect 18459 8562 19202 8564
rect 19230 8580 19286 8592
rect 20050 8590 20055 8620
rect 18459 8545 18466 8562
rect 18400 8540 18466 8545
rect 18400 8484 18405 8540
rect 18461 8484 18466 8540
rect 19230 8534 19232 8580
rect 18494 8528 19232 8534
rect 19284 8534 19286 8580
rect 19314 8564 20055 8590
rect 20111 8564 20116 8620
rect 19314 8562 20057 8564
rect 20050 8545 20057 8562
rect 20109 8545 20116 8564
rect 20050 8540 20116 8545
rect 19284 8528 20022 8534
rect 18494 8516 20022 8528
rect 18494 8506 19232 8516
rect 18400 8481 18407 8484
rect 18459 8481 18466 8484
rect 18400 8478 18466 8481
rect 18400 8469 19202 8478
rect 18400 8460 18407 8469
rect 18459 8460 19202 8469
rect 18400 8404 18405 8460
rect 18461 8450 19202 8460
rect 19230 8464 19232 8506
rect 19284 8506 20022 8516
rect 19284 8464 19286 8506
rect 20050 8484 20055 8540
rect 20111 8484 20116 8540
rect 20050 8481 20057 8484
rect 20109 8481 20116 8484
rect 20050 8478 20116 8481
rect 19230 8452 19286 8464
rect 18461 8404 18466 8450
rect 19230 8422 19232 8452
rect 18400 8353 18407 8404
rect 18459 8366 18466 8404
rect 18494 8400 19232 8422
rect 19284 8422 19286 8452
rect 19314 8469 20116 8478
rect 19314 8460 20057 8469
rect 20109 8460 20116 8469
rect 19314 8450 20055 8460
rect 19284 8400 20022 8422
rect 18494 8394 20022 8400
rect 20050 8404 20055 8450
rect 20111 8404 20116 8460
rect 18459 8361 19203 8366
rect 18459 8359 18498 8361
rect 18554 8359 18578 8361
rect 18634 8359 18658 8361
rect 18714 8359 18738 8361
rect 18794 8359 18818 8361
rect 18874 8359 18898 8361
rect 18954 8359 18978 8361
rect 19034 8359 19058 8361
rect 19114 8359 19138 8361
rect 18459 8353 18488 8359
rect 18400 8307 18488 8353
rect 18732 8307 18738 8359
rect 18796 8307 18808 8359
rect 19052 8307 19058 8359
rect 19116 8307 19128 8359
rect 18400 8305 18498 8307
rect 18554 8305 18578 8307
rect 18634 8305 18658 8307
rect 18714 8305 18738 8307
rect 18794 8305 18818 8307
rect 18874 8305 18898 8307
rect 18954 8305 18978 8307
rect 19034 8305 19058 8307
rect 19114 8305 19138 8307
rect 19194 8305 19203 8361
rect 18400 8300 19203 8305
rect 19231 8220 19285 8394
rect 20050 8366 20057 8404
rect 19313 8361 20057 8366
rect 19313 8305 19322 8361
rect 19378 8359 19402 8361
rect 19458 8359 19482 8361
rect 19538 8359 19562 8361
rect 19618 8359 19642 8361
rect 19698 8359 19722 8361
rect 19778 8359 19802 8361
rect 19858 8359 19882 8361
rect 19938 8359 19962 8361
rect 20018 8359 20057 8361
rect 19394 8307 19402 8359
rect 19458 8307 19470 8359
rect 19714 8307 19722 8359
rect 19778 8307 19790 8359
rect 20034 8353 20057 8359
rect 20109 8353 20116 8404
rect 20034 8307 20116 8353
rect 19378 8305 19402 8307
rect 19458 8305 19482 8307
rect 19538 8305 19562 8307
rect 19618 8305 19642 8307
rect 19698 8305 19722 8307
rect 19778 8305 19802 8307
rect 19858 8305 19882 8307
rect 19938 8305 19962 8307
rect 20018 8305 20116 8307
rect 19313 8300 20116 8305
rect 20160 8220 20230 9057
rect 15800 8120 16510 8220
rect 17260 8120 17290 8220
rect 15800 8110 17290 8120
rect 11860 7050 12654 7070
rect 12480 6990 12654 7050
rect 11860 6970 12654 6990
rect 12980 7050 13240 7070
rect 12980 6990 13000 7050
rect 13220 6990 13240 7050
rect 12980 6970 13240 6990
rect 13540 7050 13800 7070
rect 13540 6990 13560 7050
rect 13780 6990 13800 7050
rect 13540 6970 13800 6990
rect 14100 7050 14380 7070
rect 14100 6990 14140 7050
rect 14320 6990 14380 7050
rect 14100 6970 14380 6990
rect 14660 7050 15500 7070
rect 14660 6970 14680 7050
rect 15480 6970 15500 7050
rect 11860 6958 12088 6970
rect 11774 6844 11830 6858
rect 11774 6792 11776 6844
rect 11828 6792 11830 6844
rect 11774 6780 11830 6792
rect 11774 6728 11776 6780
rect 11828 6728 11830 6780
rect 11774 6716 11830 6728
rect 11774 6664 11776 6716
rect 11828 6664 11830 6716
rect 11774 6652 11830 6664
rect 11774 6600 11776 6652
rect 11828 6600 11830 6652
rect 11774 6588 11830 6600
rect 11774 6536 11776 6588
rect 11828 6536 11830 6588
rect 11774 6524 11830 6536
rect 11774 6472 11776 6524
rect 11828 6472 11830 6524
rect 11774 6460 11830 6472
rect 11774 6408 11776 6460
rect 11828 6408 11830 6460
rect 11774 6396 11830 6408
rect 11774 6344 11776 6396
rect 11828 6344 11830 6396
rect 11774 6332 11830 6344
rect 11774 6280 11776 6332
rect 11828 6280 11830 6332
rect 11774 6268 11830 6280
rect 11774 6216 11776 6268
rect 11828 6216 11830 6268
rect 11774 6204 11830 6216
rect 11774 6152 11776 6204
rect 11828 6152 11830 6204
rect 11774 6140 11830 6152
rect 11774 6088 11776 6140
rect 11828 6088 11830 6140
rect 11774 6076 11830 6088
rect 11774 6024 11776 6076
rect 11828 6024 11830 6076
rect 11774 6012 11830 6024
rect 11774 5960 11776 6012
rect 11828 5960 11830 6012
rect 11774 5948 11830 5960
rect 11774 5896 11776 5948
rect 11828 5896 11830 5948
rect 11774 5750 11830 5896
rect 11860 6810 11916 6958
rect 11860 6758 11862 6810
rect 11914 6758 11916 6810
rect 11860 6746 11916 6758
rect 11860 6694 11862 6746
rect 11914 6694 11916 6746
rect 11860 6682 11916 6694
rect 11860 6630 11862 6682
rect 11914 6630 11916 6682
rect 11860 6618 11916 6630
rect 11860 6566 11862 6618
rect 11914 6566 11916 6618
rect 11860 6554 11916 6566
rect 11860 6502 11862 6554
rect 11914 6502 11916 6554
rect 11860 6490 11916 6502
rect 11860 6438 11862 6490
rect 11914 6438 11916 6490
rect 11860 6426 11916 6438
rect 11860 6374 11862 6426
rect 11914 6374 11916 6426
rect 11860 6362 11916 6374
rect 11860 6310 11862 6362
rect 11914 6310 11916 6362
rect 11860 6298 11916 6310
rect 11860 6246 11862 6298
rect 11914 6246 11916 6298
rect 11860 6234 11916 6246
rect 11860 6182 11862 6234
rect 11914 6182 11916 6234
rect 11860 6170 11916 6182
rect 11860 6118 11862 6170
rect 11914 6118 11916 6170
rect 11860 6106 11916 6118
rect 11860 6054 11862 6106
rect 11914 6054 11916 6106
rect 11860 6042 11916 6054
rect 11860 5990 11862 6042
rect 11914 5990 11916 6042
rect 11860 5978 11916 5990
rect 11860 5926 11862 5978
rect 11914 5926 11916 5978
rect 11860 5914 11916 5926
rect 11860 5862 11862 5914
rect 11914 5862 11916 5914
rect 11860 5848 11916 5862
rect 11946 6844 12002 6858
rect 11946 6792 11948 6844
rect 12000 6792 12002 6844
rect 11946 6780 12002 6792
rect 11946 6728 11948 6780
rect 12000 6728 12002 6780
rect 11946 6716 12002 6728
rect 11946 6664 11948 6716
rect 12000 6664 12002 6716
rect 11946 6652 12002 6664
rect 11946 6600 11948 6652
rect 12000 6600 12002 6652
rect 11946 6588 12002 6600
rect 11946 6536 11948 6588
rect 12000 6536 12002 6588
rect 11946 6524 12002 6536
rect 11946 6472 11948 6524
rect 12000 6472 12002 6524
rect 11946 6460 12002 6472
rect 11946 6408 11948 6460
rect 12000 6408 12002 6460
rect 11946 6396 12002 6408
rect 11946 6344 11948 6396
rect 12000 6344 12002 6396
rect 11946 6332 12002 6344
rect 11946 6280 11948 6332
rect 12000 6280 12002 6332
rect 11946 6268 12002 6280
rect 11946 6216 11948 6268
rect 12000 6216 12002 6268
rect 11946 6204 12002 6216
rect 11946 6152 11948 6204
rect 12000 6152 12002 6204
rect 11946 6140 12002 6152
rect 11946 6088 11948 6140
rect 12000 6088 12002 6140
rect 11946 6076 12002 6088
rect 11946 6024 11948 6076
rect 12000 6024 12002 6076
rect 11946 6012 12002 6024
rect 11946 5960 11948 6012
rect 12000 5960 12002 6012
rect 11946 5948 12002 5960
rect 11946 5896 11948 5948
rect 12000 5896 12002 5948
rect 11946 5750 12002 5896
rect 12032 6810 12088 6958
rect 12426 6958 12654 6970
rect 12032 6758 12034 6810
rect 12086 6758 12088 6810
rect 12032 6746 12088 6758
rect 12032 6694 12034 6746
rect 12086 6694 12088 6746
rect 12032 6682 12088 6694
rect 12032 6630 12034 6682
rect 12086 6630 12088 6682
rect 12032 6618 12088 6630
rect 12032 6566 12034 6618
rect 12086 6566 12088 6618
rect 12032 6554 12088 6566
rect 12032 6502 12034 6554
rect 12086 6502 12088 6554
rect 12032 6490 12088 6502
rect 12032 6438 12034 6490
rect 12086 6438 12088 6490
rect 12032 6426 12088 6438
rect 12032 6374 12034 6426
rect 12086 6374 12088 6426
rect 12032 6362 12088 6374
rect 12032 6310 12034 6362
rect 12086 6310 12088 6362
rect 12032 6298 12088 6310
rect 12032 6246 12034 6298
rect 12086 6246 12088 6298
rect 12032 6234 12088 6246
rect 12032 6182 12034 6234
rect 12086 6182 12088 6234
rect 12032 6170 12088 6182
rect 12032 6118 12034 6170
rect 12086 6118 12088 6170
rect 12032 6106 12088 6118
rect 12032 6054 12034 6106
rect 12086 6054 12088 6106
rect 12032 6042 12088 6054
rect 12032 5990 12034 6042
rect 12086 5990 12088 6042
rect 12032 5978 12088 5990
rect 12032 5926 12034 5978
rect 12086 5926 12088 5978
rect 12032 5914 12088 5926
rect 12032 5862 12034 5914
rect 12086 5862 12088 5914
rect 12032 5848 12088 5862
rect 12118 6844 12174 6858
rect 12118 6792 12120 6844
rect 12172 6792 12174 6844
rect 12118 6780 12174 6792
rect 12118 6728 12120 6780
rect 12172 6728 12174 6780
rect 12118 6716 12174 6728
rect 12118 6664 12120 6716
rect 12172 6664 12174 6716
rect 12118 6652 12174 6664
rect 12118 6600 12120 6652
rect 12172 6600 12174 6652
rect 12118 6588 12174 6600
rect 12118 6536 12120 6588
rect 12172 6536 12174 6588
rect 12118 6524 12174 6536
rect 12118 6472 12120 6524
rect 12172 6472 12174 6524
rect 12118 6460 12174 6472
rect 12118 6408 12120 6460
rect 12172 6408 12174 6460
rect 12118 6396 12174 6408
rect 12118 6344 12120 6396
rect 12172 6344 12174 6396
rect 12118 6332 12174 6344
rect 12118 6280 12120 6332
rect 12172 6280 12174 6332
rect 12118 6268 12174 6280
rect 12118 6216 12120 6268
rect 12172 6216 12174 6268
rect 12118 6204 12174 6216
rect 12118 6152 12120 6204
rect 12172 6152 12174 6204
rect 12118 6140 12174 6152
rect 12118 6088 12120 6140
rect 12172 6088 12174 6140
rect 12118 6076 12174 6088
rect 12118 6024 12120 6076
rect 12172 6024 12174 6076
rect 12118 6012 12174 6024
rect 12118 5960 12120 6012
rect 12172 5960 12174 6012
rect 12118 5948 12174 5960
rect 12118 5896 12120 5948
rect 12172 5896 12174 5948
rect 12118 5750 12174 5896
rect 12340 6844 12396 6858
rect 12340 6792 12342 6844
rect 12394 6792 12396 6844
rect 12340 6780 12396 6792
rect 12340 6728 12342 6780
rect 12394 6728 12396 6780
rect 12340 6716 12396 6728
rect 12340 6664 12342 6716
rect 12394 6664 12396 6716
rect 12340 6652 12396 6664
rect 12340 6600 12342 6652
rect 12394 6600 12396 6652
rect 12340 6588 12396 6600
rect 12340 6536 12342 6588
rect 12394 6536 12396 6588
rect 12340 6524 12396 6536
rect 12340 6472 12342 6524
rect 12394 6472 12396 6524
rect 12340 6460 12396 6472
rect 12340 6408 12342 6460
rect 12394 6408 12396 6460
rect 12340 6396 12396 6408
rect 12340 6344 12342 6396
rect 12394 6344 12396 6396
rect 12340 6332 12396 6344
rect 12340 6280 12342 6332
rect 12394 6280 12396 6332
rect 12340 6268 12396 6280
rect 12340 6216 12342 6268
rect 12394 6216 12396 6268
rect 12340 6204 12396 6216
rect 12340 6152 12342 6204
rect 12394 6152 12396 6204
rect 12340 6140 12396 6152
rect 12340 6088 12342 6140
rect 12394 6088 12396 6140
rect 12340 6076 12396 6088
rect 12340 6024 12342 6076
rect 12394 6024 12396 6076
rect 12340 6012 12396 6024
rect 12340 5960 12342 6012
rect 12394 5960 12396 6012
rect 12340 5948 12396 5960
rect 12340 5896 12342 5948
rect 12394 5896 12396 5948
rect 12340 5750 12396 5896
rect 12426 6810 12482 6958
rect 12426 6758 12428 6810
rect 12480 6758 12482 6810
rect 12426 6746 12482 6758
rect 12426 6694 12428 6746
rect 12480 6694 12482 6746
rect 12426 6682 12482 6694
rect 12426 6630 12428 6682
rect 12480 6630 12482 6682
rect 12426 6618 12482 6630
rect 12426 6566 12428 6618
rect 12480 6566 12482 6618
rect 12426 6554 12482 6566
rect 12426 6502 12428 6554
rect 12480 6502 12482 6554
rect 12426 6490 12482 6502
rect 12426 6438 12428 6490
rect 12480 6438 12482 6490
rect 12426 6426 12482 6438
rect 12426 6374 12428 6426
rect 12480 6374 12482 6426
rect 12426 6362 12482 6374
rect 12426 6310 12428 6362
rect 12480 6310 12482 6362
rect 12426 6298 12482 6310
rect 12426 6246 12428 6298
rect 12480 6246 12482 6298
rect 12426 6234 12482 6246
rect 12426 6182 12428 6234
rect 12480 6182 12482 6234
rect 12426 6170 12482 6182
rect 12426 6118 12428 6170
rect 12480 6118 12482 6170
rect 12426 6106 12482 6118
rect 12426 6054 12428 6106
rect 12480 6054 12482 6106
rect 12426 6042 12482 6054
rect 12426 5990 12428 6042
rect 12480 5990 12482 6042
rect 12426 5978 12482 5990
rect 12426 5926 12428 5978
rect 12480 5926 12482 5978
rect 12426 5914 12482 5926
rect 12426 5862 12428 5914
rect 12480 5862 12482 5914
rect 12426 5848 12482 5862
rect 12512 6844 12568 6858
rect 12512 6792 12514 6844
rect 12566 6792 12568 6844
rect 12512 6780 12568 6792
rect 12512 6728 12514 6780
rect 12566 6728 12568 6780
rect 12512 6716 12568 6728
rect 12512 6664 12514 6716
rect 12566 6664 12568 6716
rect 12512 6652 12568 6664
rect 12512 6600 12514 6652
rect 12566 6600 12568 6652
rect 12512 6588 12568 6600
rect 12512 6536 12514 6588
rect 12566 6536 12568 6588
rect 12512 6524 12568 6536
rect 12512 6472 12514 6524
rect 12566 6472 12568 6524
rect 12512 6460 12568 6472
rect 12512 6408 12514 6460
rect 12566 6408 12568 6460
rect 12512 6396 12568 6408
rect 12512 6344 12514 6396
rect 12566 6344 12568 6396
rect 12512 6332 12568 6344
rect 12512 6280 12514 6332
rect 12566 6280 12568 6332
rect 12512 6268 12568 6280
rect 12512 6216 12514 6268
rect 12566 6216 12568 6268
rect 12512 6204 12568 6216
rect 12512 6152 12514 6204
rect 12566 6152 12568 6204
rect 12512 6140 12568 6152
rect 12512 6088 12514 6140
rect 12566 6088 12568 6140
rect 12512 6076 12568 6088
rect 12512 6024 12514 6076
rect 12566 6024 12568 6076
rect 12512 6012 12568 6024
rect 12512 5960 12514 6012
rect 12566 5960 12568 6012
rect 12512 5948 12568 5960
rect 12512 5896 12514 5948
rect 12566 5896 12568 5948
rect 12512 5750 12568 5896
rect 12598 6810 12654 6958
rect 12992 6958 13220 6970
rect 12598 6758 12600 6810
rect 12652 6758 12654 6810
rect 12598 6746 12654 6758
rect 12598 6694 12600 6746
rect 12652 6694 12654 6746
rect 12598 6682 12654 6694
rect 12598 6630 12600 6682
rect 12652 6630 12654 6682
rect 12598 6618 12654 6630
rect 12598 6566 12600 6618
rect 12652 6566 12654 6618
rect 12598 6554 12654 6566
rect 12598 6502 12600 6554
rect 12652 6502 12654 6554
rect 12598 6490 12654 6502
rect 12598 6438 12600 6490
rect 12652 6438 12654 6490
rect 12598 6426 12654 6438
rect 12598 6374 12600 6426
rect 12652 6374 12654 6426
rect 12598 6362 12654 6374
rect 12598 6310 12600 6362
rect 12652 6310 12654 6362
rect 12598 6298 12654 6310
rect 12598 6246 12600 6298
rect 12652 6246 12654 6298
rect 12598 6234 12654 6246
rect 12598 6182 12600 6234
rect 12652 6182 12654 6234
rect 12598 6170 12654 6182
rect 12598 6118 12600 6170
rect 12652 6118 12654 6170
rect 12598 6106 12654 6118
rect 12598 6054 12600 6106
rect 12652 6054 12654 6106
rect 12598 6042 12654 6054
rect 12598 5990 12600 6042
rect 12652 5990 12654 6042
rect 12598 5978 12654 5990
rect 12598 5926 12600 5978
rect 12652 5926 12654 5978
rect 12598 5914 12654 5926
rect 12598 5862 12600 5914
rect 12652 5862 12654 5914
rect 12598 5848 12654 5862
rect 12684 6844 12740 6858
rect 12684 6792 12686 6844
rect 12738 6792 12740 6844
rect 12684 6780 12740 6792
rect 12684 6728 12686 6780
rect 12738 6728 12740 6780
rect 12684 6716 12740 6728
rect 12684 6664 12686 6716
rect 12738 6664 12740 6716
rect 12684 6652 12740 6664
rect 12684 6600 12686 6652
rect 12738 6600 12740 6652
rect 12684 6588 12740 6600
rect 12684 6536 12686 6588
rect 12738 6536 12740 6588
rect 12684 6524 12740 6536
rect 12684 6472 12686 6524
rect 12738 6472 12740 6524
rect 12684 6460 12740 6472
rect 12684 6408 12686 6460
rect 12738 6408 12740 6460
rect 12684 6396 12740 6408
rect 12684 6344 12686 6396
rect 12738 6344 12740 6396
rect 12684 6332 12740 6344
rect 12684 6280 12686 6332
rect 12738 6280 12740 6332
rect 12684 6268 12740 6280
rect 12684 6216 12686 6268
rect 12738 6216 12740 6268
rect 12684 6204 12740 6216
rect 12684 6152 12686 6204
rect 12738 6152 12740 6204
rect 12684 6140 12740 6152
rect 12684 6088 12686 6140
rect 12738 6088 12740 6140
rect 12684 6076 12740 6088
rect 12684 6024 12686 6076
rect 12738 6024 12740 6076
rect 12684 6012 12740 6024
rect 12684 5960 12686 6012
rect 12738 5960 12740 6012
rect 12684 5948 12740 5960
rect 12684 5896 12686 5948
rect 12738 5896 12740 5948
rect 12684 5750 12740 5896
rect 12906 6844 12962 6858
rect 12906 6792 12908 6844
rect 12960 6792 12962 6844
rect 12906 6780 12962 6792
rect 12906 6728 12908 6780
rect 12960 6728 12962 6780
rect 12906 6716 12962 6728
rect 12906 6664 12908 6716
rect 12960 6664 12962 6716
rect 12906 6652 12962 6664
rect 12906 6600 12908 6652
rect 12960 6600 12962 6652
rect 12906 6588 12962 6600
rect 12906 6536 12908 6588
rect 12960 6536 12962 6588
rect 12906 6524 12962 6536
rect 12906 6472 12908 6524
rect 12960 6472 12962 6524
rect 12906 6460 12962 6472
rect 12906 6408 12908 6460
rect 12960 6408 12962 6460
rect 12906 6396 12962 6408
rect 12906 6344 12908 6396
rect 12960 6344 12962 6396
rect 12906 6332 12962 6344
rect 12906 6280 12908 6332
rect 12960 6280 12962 6332
rect 12906 6268 12962 6280
rect 12906 6216 12908 6268
rect 12960 6216 12962 6268
rect 12906 6204 12962 6216
rect 12906 6152 12908 6204
rect 12960 6152 12962 6204
rect 12906 6140 12962 6152
rect 12906 6088 12908 6140
rect 12960 6088 12962 6140
rect 12906 6076 12962 6088
rect 12906 6024 12908 6076
rect 12960 6024 12962 6076
rect 12906 6012 12962 6024
rect 12906 5960 12908 6012
rect 12960 5960 12962 6012
rect 12906 5948 12962 5960
rect 12906 5896 12908 5948
rect 12960 5896 12962 5948
rect 12906 5750 12962 5896
rect 12992 6810 13048 6958
rect 12992 6758 12994 6810
rect 13046 6758 13048 6810
rect 12992 6746 13048 6758
rect 12992 6694 12994 6746
rect 13046 6694 13048 6746
rect 12992 6682 13048 6694
rect 12992 6630 12994 6682
rect 13046 6630 13048 6682
rect 12992 6618 13048 6630
rect 12992 6566 12994 6618
rect 13046 6566 13048 6618
rect 12992 6554 13048 6566
rect 12992 6502 12994 6554
rect 13046 6502 13048 6554
rect 12992 6490 13048 6502
rect 12992 6438 12994 6490
rect 13046 6438 13048 6490
rect 12992 6426 13048 6438
rect 12992 6374 12994 6426
rect 13046 6374 13048 6426
rect 12992 6362 13048 6374
rect 12992 6310 12994 6362
rect 13046 6310 13048 6362
rect 12992 6298 13048 6310
rect 12992 6246 12994 6298
rect 13046 6246 13048 6298
rect 12992 6234 13048 6246
rect 12992 6182 12994 6234
rect 13046 6182 13048 6234
rect 12992 6170 13048 6182
rect 12992 6118 12994 6170
rect 13046 6118 13048 6170
rect 12992 6106 13048 6118
rect 12992 6054 12994 6106
rect 13046 6054 13048 6106
rect 12992 6042 13048 6054
rect 12992 5990 12994 6042
rect 13046 5990 13048 6042
rect 12992 5978 13048 5990
rect 12992 5926 12994 5978
rect 13046 5926 13048 5978
rect 12992 5914 13048 5926
rect 12992 5862 12994 5914
rect 13046 5862 13048 5914
rect 12992 5848 13048 5862
rect 13078 6844 13134 6858
rect 13078 6792 13080 6844
rect 13132 6792 13134 6844
rect 13078 6780 13134 6792
rect 13078 6728 13080 6780
rect 13132 6728 13134 6780
rect 13078 6716 13134 6728
rect 13078 6664 13080 6716
rect 13132 6664 13134 6716
rect 13078 6652 13134 6664
rect 13078 6600 13080 6652
rect 13132 6600 13134 6652
rect 13078 6588 13134 6600
rect 13078 6536 13080 6588
rect 13132 6536 13134 6588
rect 13078 6524 13134 6536
rect 13078 6472 13080 6524
rect 13132 6472 13134 6524
rect 13078 6460 13134 6472
rect 13078 6408 13080 6460
rect 13132 6408 13134 6460
rect 13078 6396 13134 6408
rect 13078 6344 13080 6396
rect 13132 6344 13134 6396
rect 13078 6332 13134 6344
rect 13078 6280 13080 6332
rect 13132 6280 13134 6332
rect 13078 6268 13134 6280
rect 13078 6216 13080 6268
rect 13132 6216 13134 6268
rect 13078 6204 13134 6216
rect 13078 6152 13080 6204
rect 13132 6152 13134 6204
rect 13078 6140 13134 6152
rect 13078 6088 13080 6140
rect 13132 6088 13134 6140
rect 13078 6076 13134 6088
rect 13078 6024 13080 6076
rect 13132 6024 13134 6076
rect 13078 6012 13134 6024
rect 13078 5960 13080 6012
rect 13132 5960 13134 6012
rect 13078 5948 13134 5960
rect 13078 5896 13080 5948
rect 13132 5896 13134 5948
rect 13078 5750 13134 5896
rect 13164 6810 13220 6958
rect 13558 6958 13786 6970
rect 13164 6758 13166 6810
rect 13218 6758 13220 6810
rect 13164 6746 13220 6758
rect 13164 6694 13166 6746
rect 13218 6694 13220 6746
rect 13164 6682 13220 6694
rect 13164 6630 13166 6682
rect 13218 6630 13220 6682
rect 13164 6618 13220 6630
rect 13164 6566 13166 6618
rect 13218 6566 13220 6618
rect 13164 6554 13220 6566
rect 13164 6502 13166 6554
rect 13218 6502 13220 6554
rect 13164 6490 13220 6502
rect 13164 6438 13166 6490
rect 13218 6438 13220 6490
rect 13164 6426 13220 6438
rect 13164 6374 13166 6426
rect 13218 6374 13220 6426
rect 13164 6362 13220 6374
rect 13164 6310 13166 6362
rect 13218 6310 13220 6362
rect 13164 6298 13220 6310
rect 13164 6246 13166 6298
rect 13218 6246 13220 6298
rect 13164 6234 13220 6246
rect 13164 6182 13166 6234
rect 13218 6182 13220 6234
rect 13164 6170 13220 6182
rect 13164 6118 13166 6170
rect 13218 6118 13220 6170
rect 13164 6106 13220 6118
rect 13164 6054 13166 6106
rect 13218 6054 13220 6106
rect 13164 6042 13220 6054
rect 13164 5990 13166 6042
rect 13218 5990 13220 6042
rect 13164 5978 13220 5990
rect 13164 5926 13166 5978
rect 13218 5926 13220 5978
rect 13164 5914 13220 5926
rect 13164 5862 13166 5914
rect 13218 5862 13220 5914
rect 13164 5848 13220 5862
rect 13250 6844 13306 6858
rect 13250 6792 13252 6844
rect 13304 6792 13306 6844
rect 13250 6780 13306 6792
rect 13250 6728 13252 6780
rect 13304 6728 13306 6780
rect 13250 6716 13306 6728
rect 13250 6664 13252 6716
rect 13304 6664 13306 6716
rect 13250 6652 13306 6664
rect 13250 6600 13252 6652
rect 13304 6600 13306 6652
rect 13250 6588 13306 6600
rect 13250 6536 13252 6588
rect 13304 6536 13306 6588
rect 13250 6524 13306 6536
rect 13250 6472 13252 6524
rect 13304 6472 13306 6524
rect 13250 6460 13306 6472
rect 13250 6408 13252 6460
rect 13304 6408 13306 6460
rect 13250 6396 13306 6408
rect 13250 6344 13252 6396
rect 13304 6344 13306 6396
rect 13250 6332 13306 6344
rect 13250 6280 13252 6332
rect 13304 6280 13306 6332
rect 13250 6268 13306 6280
rect 13250 6216 13252 6268
rect 13304 6216 13306 6268
rect 13250 6204 13306 6216
rect 13250 6152 13252 6204
rect 13304 6152 13306 6204
rect 13250 6140 13306 6152
rect 13250 6088 13252 6140
rect 13304 6088 13306 6140
rect 13250 6076 13306 6088
rect 13250 6024 13252 6076
rect 13304 6024 13306 6076
rect 13250 6012 13306 6024
rect 13250 5960 13252 6012
rect 13304 5960 13306 6012
rect 13250 5948 13306 5960
rect 13250 5896 13252 5948
rect 13304 5896 13306 5948
rect 13250 5750 13306 5896
rect 13472 6844 13528 6858
rect 13472 6792 13474 6844
rect 13526 6792 13528 6844
rect 13472 6780 13528 6792
rect 13472 6728 13474 6780
rect 13526 6728 13528 6780
rect 13472 6716 13528 6728
rect 13472 6664 13474 6716
rect 13526 6664 13528 6716
rect 13472 6652 13528 6664
rect 13472 6600 13474 6652
rect 13526 6600 13528 6652
rect 13472 6588 13528 6600
rect 13472 6536 13474 6588
rect 13526 6536 13528 6588
rect 13472 6524 13528 6536
rect 13472 6472 13474 6524
rect 13526 6472 13528 6524
rect 13472 6460 13528 6472
rect 13472 6408 13474 6460
rect 13526 6408 13528 6460
rect 13472 6396 13528 6408
rect 13472 6344 13474 6396
rect 13526 6344 13528 6396
rect 13472 6332 13528 6344
rect 13472 6280 13474 6332
rect 13526 6280 13528 6332
rect 13472 6268 13528 6280
rect 13472 6216 13474 6268
rect 13526 6216 13528 6268
rect 13472 6204 13528 6216
rect 13472 6152 13474 6204
rect 13526 6152 13528 6204
rect 13472 6140 13528 6152
rect 13472 6088 13474 6140
rect 13526 6088 13528 6140
rect 13472 6076 13528 6088
rect 13472 6024 13474 6076
rect 13526 6024 13528 6076
rect 13472 6012 13528 6024
rect 13472 5960 13474 6012
rect 13526 5960 13528 6012
rect 13472 5948 13528 5960
rect 13472 5896 13474 5948
rect 13526 5896 13528 5948
rect 13472 5750 13528 5896
rect 13558 6810 13614 6958
rect 13558 6758 13560 6810
rect 13612 6758 13614 6810
rect 13558 6746 13614 6758
rect 13558 6694 13560 6746
rect 13612 6694 13614 6746
rect 13558 6682 13614 6694
rect 13558 6630 13560 6682
rect 13612 6630 13614 6682
rect 13558 6618 13614 6630
rect 13558 6566 13560 6618
rect 13612 6566 13614 6618
rect 13558 6554 13614 6566
rect 13558 6502 13560 6554
rect 13612 6502 13614 6554
rect 13558 6490 13614 6502
rect 13558 6438 13560 6490
rect 13612 6438 13614 6490
rect 13558 6426 13614 6438
rect 13558 6374 13560 6426
rect 13612 6374 13614 6426
rect 13558 6362 13614 6374
rect 13558 6310 13560 6362
rect 13612 6310 13614 6362
rect 13558 6298 13614 6310
rect 13558 6246 13560 6298
rect 13612 6246 13614 6298
rect 13558 6234 13614 6246
rect 13558 6182 13560 6234
rect 13612 6182 13614 6234
rect 13558 6170 13614 6182
rect 13558 6118 13560 6170
rect 13612 6118 13614 6170
rect 13558 6106 13614 6118
rect 13558 6054 13560 6106
rect 13612 6054 13614 6106
rect 13558 6042 13614 6054
rect 13558 5990 13560 6042
rect 13612 5990 13614 6042
rect 13558 5978 13614 5990
rect 13558 5926 13560 5978
rect 13612 5926 13614 5978
rect 13558 5914 13614 5926
rect 13558 5862 13560 5914
rect 13612 5862 13614 5914
rect 13558 5848 13614 5862
rect 13644 6844 13700 6858
rect 13644 6792 13646 6844
rect 13698 6792 13700 6844
rect 13644 6780 13700 6792
rect 13644 6728 13646 6780
rect 13698 6728 13700 6780
rect 13644 6716 13700 6728
rect 13644 6664 13646 6716
rect 13698 6664 13700 6716
rect 13644 6652 13700 6664
rect 13644 6600 13646 6652
rect 13698 6600 13700 6652
rect 13644 6588 13700 6600
rect 13644 6536 13646 6588
rect 13698 6536 13700 6588
rect 13644 6524 13700 6536
rect 13644 6472 13646 6524
rect 13698 6472 13700 6524
rect 13644 6460 13700 6472
rect 13644 6408 13646 6460
rect 13698 6408 13700 6460
rect 13644 6396 13700 6408
rect 13644 6344 13646 6396
rect 13698 6344 13700 6396
rect 13644 6332 13700 6344
rect 13644 6280 13646 6332
rect 13698 6280 13700 6332
rect 13644 6268 13700 6280
rect 13644 6216 13646 6268
rect 13698 6216 13700 6268
rect 13644 6204 13700 6216
rect 13644 6152 13646 6204
rect 13698 6152 13700 6204
rect 13644 6140 13700 6152
rect 13644 6088 13646 6140
rect 13698 6088 13700 6140
rect 13644 6076 13700 6088
rect 13644 6024 13646 6076
rect 13698 6024 13700 6076
rect 13644 6012 13700 6024
rect 13644 5960 13646 6012
rect 13698 5960 13700 6012
rect 13644 5948 13700 5960
rect 13644 5896 13646 5948
rect 13698 5896 13700 5948
rect 13644 5750 13700 5896
rect 13730 6810 13786 6958
rect 14124 6958 14352 6970
rect 13730 6758 13732 6810
rect 13784 6758 13786 6810
rect 13730 6746 13786 6758
rect 13730 6694 13732 6746
rect 13784 6694 13786 6746
rect 13730 6682 13786 6694
rect 13730 6630 13732 6682
rect 13784 6630 13786 6682
rect 13730 6618 13786 6630
rect 13730 6566 13732 6618
rect 13784 6566 13786 6618
rect 13730 6554 13786 6566
rect 13730 6502 13732 6554
rect 13784 6502 13786 6554
rect 13730 6490 13786 6502
rect 13730 6438 13732 6490
rect 13784 6438 13786 6490
rect 13730 6426 13786 6438
rect 13730 6374 13732 6426
rect 13784 6374 13786 6426
rect 13730 6362 13786 6374
rect 13730 6310 13732 6362
rect 13784 6310 13786 6362
rect 13730 6298 13786 6310
rect 13730 6246 13732 6298
rect 13784 6246 13786 6298
rect 13730 6234 13786 6246
rect 13730 6182 13732 6234
rect 13784 6182 13786 6234
rect 13730 6170 13786 6182
rect 13730 6118 13732 6170
rect 13784 6118 13786 6170
rect 13730 6106 13786 6118
rect 13730 6054 13732 6106
rect 13784 6054 13786 6106
rect 13730 6042 13786 6054
rect 13730 5990 13732 6042
rect 13784 5990 13786 6042
rect 13730 5978 13786 5990
rect 13730 5926 13732 5978
rect 13784 5926 13786 5978
rect 13730 5914 13786 5926
rect 13730 5862 13732 5914
rect 13784 5862 13786 5914
rect 13730 5848 13786 5862
rect 13816 6844 13872 6858
rect 13816 6792 13818 6844
rect 13870 6792 13872 6844
rect 13816 6780 13872 6792
rect 13816 6728 13818 6780
rect 13870 6728 13872 6780
rect 13816 6716 13872 6728
rect 13816 6664 13818 6716
rect 13870 6664 13872 6716
rect 13816 6652 13872 6664
rect 13816 6600 13818 6652
rect 13870 6600 13872 6652
rect 13816 6588 13872 6600
rect 13816 6536 13818 6588
rect 13870 6536 13872 6588
rect 13816 6524 13872 6536
rect 13816 6472 13818 6524
rect 13870 6472 13872 6524
rect 13816 6460 13872 6472
rect 13816 6408 13818 6460
rect 13870 6408 13872 6460
rect 13816 6396 13872 6408
rect 13816 6344 13818 6396
rect 13870 6344 13872 6396
rect 13816 6332 13872 6344
rect 13816 6280 13818 6332
rect 13870 6280 13872 6332
rect 13816 6268 13872 6280
rect 13816 6216 13818 6268
rect 13870 6216 13872 6268
rect 13816 6204 13872 6216
rect 13816 6152 13818 6204
rect 13870 6152 13872 6204
rect 13816 6140 13872 6152
rect 13816 6088 13818 6140
rect 13870 6088 13872 6140
rect 13816 6076 13872 6088
rect 13816 6024 13818 6076
rect 13870 6024 13872 6076
rect 13816 6012 13872 6024
rect 13816 5960 13818 6012
rect 13870 5960 13872 6012
rect 13816 5948 13872 5960
rect 13816 5896 13818 5948
rect 13870 5896 13872 5948
rect 13816 5750 13872 5896
rect 14038 6844 14094 6858
rect 14038 6792 14040 6844
rect 14092 6792 14094 6844
rect 14038 6780 14094 6792
rect 14038 6728 14040 6780
rect 14092 6728 14094 6780
rect 14038 6716 14094 6728
rect 14038 6664 14040 6716
rect 14092 6664 14094 6716
rect 14038 6652 14094 6664
rect 14038 6600 14040 6652
rect 14092 6600 14094 6652
rect 14038 6588 14094 6600
rect 14038 6536 14040 6588
rect 14092 6536 14094 6588
rect 14038 6524 14094 6536
rect 14038 6472 14040 6524
rect 14092 6472 14094 6524
rect 14038 6460 14094 6472
rect 14038 6408 14040 6460
rect 14092 6408 14094 6460
rect 14038 6396 14094 6408
rect 14038 6344 14040 6396
rect 14092 6344 14094 6396
rect 14038 6332 14094 6344
rect 14038 6280 14040 6332
rect 14092 6280 14094 6332
rect 14038 6268 14094 6280
rect 14038 6216 14040 6268
rect 14092 6216 14094 6268
rect 14038 6204 14094 6216
rect 14038 6152 14040 6204
rect 14092 6152 14094 6204
rect 14038 6140 14094 6152
rect 14038 6088 14040 6140
rect 14092 6088 14094 6140
rect 14038 6076 14094 6088
rect 14038 6024 14040 6076
rect 14092 6024 14094 6076
rect 14038 6012 14094 6024
rect 14038 5960 14040 6012
rect 14092 5960 14094 6012
rect 14038 5948 14094 5960
rect 14038 5896 14040 5948
rect 14092 5896 14094 5948
rect 14038 5750 14094 5896
rect 14124 6810 14180 6958
rect 14124 6758 14126 6810
rect 14178 6758 14180 6810
rect 14124 6746 14180 6758
rect 14124 6694 14126 6746
rect 14178 6694 14180 6746
rect 14124 6682 14180 6694
rect 14124 6630 14126 6682
rect 14178 6630 14180 6682
rect 14124 6618 14180 6630
rect 14124 6566 14126 6618
rect 14178 6566 14180 6618
rect 14124 6554 14180 6566
rect 14124 6502 14126 6554
rect 14178 6502 14180 6554
rect 14124 6490 14180 6502
rect 14124 6438 14126 6490
rect 14178 6438 14180 6490
rect 14124 6426 14180 6438
rect 14124 6374 14126 6426
rect 14178 6374 14180 6426
rect 14124 6362 14180 6374
rect 14124 6310 14126 6362
rect 14178 6310 14180 6362
rect 14124 6298 14180 6310
rect 14124 6246 14126 6298
rect 14178 6246 14180 6298
rect 14124 6234 14180 6246
rect 14124 6182 14126 6234
rect 14178 6182 14180 6234
rect 14124 6170 14180 6182
rect 14124 6118 14126 6170
rect 14178 6118 14180 6170
rect 14124 6106 14180 6118
rect 14124 6054 14126 6106
rect 14178 6054 14180 6106
rect 14124 6042 14180 6054
rect 14124 5990 14126 6042
rect 14178 5990 14180 6042
rect 14124 5978 14180 5990
rect 14124 5926 14126 5978
rect 14178 5926 14180 5978
rect 14124 5914 14180 5926
rect 14124 5862 14126 5914
rect 14178 5862 14180 5914
rect 14124 5848 14180 5862
rect 14210 6844 14266 6858
rect 14210 6792 14212 6844
rect 14264 6792 14266 6844
rect 14210 6780 14266 6792
rect 14210 6728 14212 6780
rect 14264 6728 14266 6780
rect 14210 6716 14266 6728
rect 14210 6664 14212 6716
rect 14264 6664 14266 6716
rect 14210 6652 14266 6664
rect 14210 6600 14212 6652
rect 14264 6600 14266 6652
rect 14210 6588 14266 6600
rect 14210 6536 14212 6588
rect 14264 6536 14266 6588
rect 14210 6524 14266 6536
rect 14210 6472 14212 6524
rect 14264 6472 14266 6524
rect 14210 6460 14266 6472
rect 14210 6408 14212 6460
rect 14264 6408 14266 6460
rect 14210 6396 14266 6408
rect 14210 6344 14212 6396
rect 14264 6344 14266 6396
rect 14210 6332 14266 6344
rect 14210 6280 14212 6332
rect 14264 6280 14266 6332
rect 14210 6268 14266 6280
rect 14210 6216 14212 6268
rect 14264 6216 14266 6268
rect 14210 6204 14266 6216
rect 14210 6152 14212 6204
rect 14264 6152 14266 6204
rect 14210 6140 14266 6152
rect 14210 6088 14212 6140
rect 14264 6088 14266 6140
rect 14210 6076 14266 6088
rect 14210 6024 14212 6076
rect 14264 6024 14266 6076
rect 14210 6012 14266 6024
rect 14210 5960 14212 6012
rect 14264 5960 14266 6012
rect 14210 5948 14266 5960
rect 14210 5896 14212 5948
rect 14264 5896 14266 5948
rect 14210 5750 14266 5896
rect 14296 6810 14352 6958
rect 14660 6950 15500 6970
rect 15800 7000 15960 8110
rect 16060 8100 17290 8110
rect 17380 8180 20230 8220
rect 16060 7000 16070 8100
rect 17380 8080 17420 8180
rect 20140 8080 20230 8180
rect 17380 8040 20230 8080
rect 15800 6980 16070 7000
rect 16195 7901 16247 7971
rect 16195 7821 16247 7849
rect 16195 7741 16247 7769
rect 16195 7661 16247 7689
rect 16195 7581 16247 7609
rect 16195 7501 16247 7529
rect 16195 7421 16247 7449
rect 16195 7341 16247 7369
rect 16195 7261 16247 7289
rect 16195 7181 16247 7209
rect 16195 7101 16247 7129
rect 14296 6758 14298 6810
rect 14350 6758 14352 6810
rect 14296 6746 14352 6758
rect 14296 6694 14298 6746
rect 14350 6694 14352 6746
rect 14296 6682 14352 6694
rect 14296 6630 14298 6682
rect 14350 6630 14352 6682
rect 14296 6618 14352 6630
rect 14296 6566 14298 6618
rect 14350 6566 14352 6618
rect 14296 6554 14352 6566
rect 14296 6502 14298 6554
rect 14350 6502 14352 6554
rect 14296 6490 14352 6502
rect 14296 6438 14298 6490
rect 14350 6438 14352 6490
rect 14296 6426 14352 6438
rect 14296 6374 14298 6426
rect 14350 6374 14352 6426
rect 14296 6362 14352 6374
rect 14296 6310 14298 6362
rect 14350 6310 14352 6362
rect 14296 6298 14352 6310
rect 14296 6246 14298 6298
rect 14350 6246 14352 6298
rect 14296 6234 14352 6246
rect 14296 6182 14298 6234
rect 14350 6182 14352 6234
rect 14296 6170 14352 6182
rect 14296 6118 14298 6170
rect 14350 6118 14352 6170
rect 14296 6106 14352 6118
rect 14296 6054 14298 6106
rect 14350 6054 14352 6106
rect 14296 6042 14352 6054
rect 14296 5990 14298 6042
rect 14350 5990 14352 6042
rect 14296 5978 14352 5990
rect 14296 5926 14298 5978
rect 14350 5926 14352 5978
rect 14296 5914 14352 5926
rect 14296 5862 14298 5914
rect 14350 5862 14352 5914
rect 14296 5848 14352 5862
rect 14382 6844 14438 6858
rect 14382 6792 14384 6844
rect 14436 6792 14438 6844
rect 14382 6780 14438 6792
rect 14382 6728 14384 6780
rect 14436 6728 14438 6780
rect 14382 6716 14438 6728
rect 14382 6664 14384 6716
rect 14436 6664 14438 6716
rect 14382 6652 14438 6664
rect 14382 6600 14384 6652
rect 14436 6600 14438 6652
rect 14382 6588 14438 6600
rect 14382 6536 14384 6588
rect 14436 6536 14438 6588
rect 14382 6524 14438 6536
rect 14382 6472 14384 6524
rect 14436 6472 14438 6524
rect 14382 6460 14438 6472
rect 14382 6408 14384 6460
rect 14436 6408 14438 6460
rect 14382 6396 14438 6408
rect 14382 6344 14384 6396
rect 14436 6344 14438 6396
rect 14382 6332 14438 6344
rect 14382 6280 14384 6332
rect 14436 6280 14438 6332
rect 14382 6268 14438 6280
rect 14382 6216 14384 6268
rect 14436 6216 14438 6268
rect 14382 6204 14438 6216
rect 14382 6152 14384 6204
rect 14436 6152 14438 6204
rect 14382 6140 14438 6152
rect 14382 6088 14384 6140
rect 14436 6088 14438 6140
rect 14382 6076 14438 6088
rect 14382 6024 14384 6076
rect 14436 6024 14438 6076
rect 14382 6012 14438 6024
rect 14382 5960 14384 6012
rect 14436 5960 14438 6012
rect 14382 5948 14438 5960
rect 14382 5896 14384 5948
rect 14436 5896 14438 5948
rect 14382 5750 14438 5896
rect 14604 6844 14660 6858
rect 14604 6792 14606 6844
rect 14658 6792 14660 6844
rect 14604 6780 14660 6792
rect 14604 6728 14606 6780
rect 14658 6728 14660 6780
rect 14604 6716 14660 6728
rect 14604 6664 14606 6716
rect 14658 6664 14660 6716
rect 14604 6652 14660 6664
rect 14604 6600 14606 6652
rect 14658 6600 14660 6652
rect 14604 6588 14660 6600
rect 14604 6536 14606 6588
rect 14658 6536 14660 6588
rect 14604 6524 14660 6536
rect 14604 6472 14606 6524
rect 14658 6472 14660 6524
rect 14604 6460 14660 6472
rect 14604 6408 14606 6460
rect 14658 6408 14660 6460
rect 14604 6396 14660 6408
rect 14604 6344 14606 6396
rect 14658 6344 14660 6396
rect 14604 6332 14660 6344
rect 14604 6280 14606 6332
rect 14658 6280 14660 6332
rect 14604 6268 14660 6280
rect 14604 6216 14606 6268
rect 14658 6216 14660 6268
rect 14604 6204 14660 6216
rect 14604 6152 14606 6204
rect 14658 6152 14660 6204
rect 14604 6140 14660 6152
rect 14604 6088 14606 6140
rect 14658 6088 14660 6140
rect 14604 6076 14660 6088
rect 14604 6024 14606 6076
rect 14658 6024 14660 6076
rect 14604 6012 14660 6024
rect 14604 5960 14606 6012
rect 14658 5960 14660 6012
rect 14604 5948 14660 5960
rect 14604 5896 14606 5948
rect 14658 5896 14660 5948
rect 14604 5750 14660 5896
rect 14690 6810 14746 6950
rect 14690 6758 14692 6810
rect 14744 6758 14746 6810
rect 14690 6746 14746 6758
rect 14690 6694 14692 6746
rect 14744 6694 14746 6746
rect 14690 6682 14746 6694
rect 14690 6630 14692 6682
rect 14744 6630 14746 6682
rect 14690 6618 14746 6630
rect 14690 6566 14692 6618
rect 14744 6566 14746 6618
rect 14690 6554 14746 6566
rect 14690 6502 14692 6554
rect 14744 6502 14746 6554
rect 14690 6490 14746 6502
rect 14690 6438 14692 6490
rect 14744 6438 14746 6490
rect 14690 6426 14746 6438
rect 14690 6374 14692 6426
rect 14744 6374 14746 6426
rect 14690 6362 14746 6374
rect 14690 6310 14692 6362
rect 14744 6310 14746 6362
rect 14690 6298 14746 6310
rect 14690 6246 14692 6298
rect 14744 6246 14746 6298
rect 14690 6234 14746 6246
rect 14690 6182 14692 6234
rect 14744 6182 14746 6234
rect 14690 6170 14746 6182
rect 14690 6118 14692 6170
rect 14744 6118 14746 6170
rect 14690 6106 14746 6118
rect 14690 6054 14692 6106
rect 14744 6054 14746 6106
rect 14690 6042 14746 6054
rect 14690 5990 14692 6042
rect 14744 5990 14746 6042
rect 14690 5978 14746 5990
rect 14690 5926 14692 5978
rect 14744 5926 14746 5978
rect 14690 5914 14746 5926
rect 14690 5862 14692 5914
rect 14744 5862 14746 5914
rect 14690 5848 14746 5862
rect 14776 6844 14832 6858
rect 14776 6792 14778 6844
rect 14830 6792 14832 6844
rect 14776 6780 14832 6792
rect 14776 6728 14778 6780
rect 14830 6728 14832 6780
rect 14776 6716 14832 6728
rect 14776 6664 14778 6716
rect 14830 6664 14832 6716
rect 14776 6652 14832 6664
rect 14776 6600 14778 6652
rect 14830 6600 14832 6652
rect 14776 6588 14832 6600
rect 14776 6536 14778 6588
rect 14830 6536 14832 6588
rect 14776 6524 14832 6536
rect 14776 6472 14778 6524
rect 14830 6472 14832 6524
rect 14776 6460 14832 6472
rect 14776 6408 14778 6460
rect 14830 6408 14832 6460
rect 14776 6396 14832 6408
rect 14776 6344 14778 6396
rect 14830 6344 14832 6396
rect 14776 6332 14832 6344
rect 14776 6280 14778 6332
rect 14830 6280 14832 6332
rect 14776 6268 14832 6280
rect 14776 6216 14778 6268
rect 14830 6216 14832 6268
rect 14776 6204 14832 6216
rect 14776 6152 14778 6204
rect 14830 6152 14832 6204
rect 14776 6140 14832 6152
rect 14776 6088 14778 6140
rect 14830 6088 14832 6140
rect 14776 6076 14832 6088
rect 14776 6024 14778 6076
rect 14830 6024 14832 6076
rect 14776 6012 14832 6024
rect 14776 5960 14778 6012
rect 14830 5960 14832 6012
rect 14776 5948 14832 5960
rect 14776 5896 14778 5948
rect 14830 5896 14832 5948
rect 14776 5750 14832 5896
rect 14862 6810 14918 6950
rect 14862 6758 14864 6810
rect 14916 6758 14918 6810
rect 14862 6746 14918 6758
rect 14862 6694 14864 6746
rect 14916 6694 14918 6746
rect 14862 6682 14918 6694
rect 14862 6630 14864 6682
rect 14916 6630 14918 6682
rect 14862 6618 14918 6630
rect 14862 6566 14864 6618
rect 14916 6566 14918 6618
rect 14862 6554 14918 6566
rect 14862 6502 14864 6554
rect 14916 6502 14918 6554
rect 14862 6490 14918 6502
rect 14862 6438 14864 6490
rect 14916 6438 14918 6490
rect 14862 6426 14918 6438
rect 14862 6374 14864 6426
rect 14916 6374 14918 6426
rect 14862 6362 14918 6374
rect 14862 6310 14864 6362
rect 14916 6310 14918 6362
rect 14862 6298 14918 6310
rect 14862 6246 14864 6298
rect 14916 6246 14918 6298
rect 14862 6234 14918 6246
rect 14862 6182 14864 6234
rect 14916 6182 14918 6234
rect 14862 6170 14918 6182
rect 14862 6118 14864 6170
rect 14916 6118 14918 6170
rect 14862 6106 14918 6118
rect 14862 6054 14864 6106
rect 14916 6054 14918 6106
rect 14862 6042 14918 6054
rect 14862 5990 14864 6042
rect 14916 5990 14918 6042
rect 14862 5978 14918 5990
rect 14862 5926 14864 5978
rect 14916 5926 14918 5978
rect 14862 5914 14918 5926
rect 14862 5862 14864 5914
rect 14916 5862 14918 5914
rect 14862 5848 14918 5862
rect 14948 6844 15004 6858
rect 14948 6792 14950 6844
rect 15002 6792 15004 6844
rect 14948 6780 15004 6792
rect 14948 6728 14950 6780
rect 15002 6728 15004 6780
rect 14948 6716 15004 6728
rect 14948 6664 14950 6716
rect 15002 6664 15004 6716
rect 14948 6652 15004 6664
rect 14948 6600 14950 6652
rect 15002 6600 15004 6652
rect 14948 6588 15004 6600
rect 14948 6536 14950 6588
rect 15002 6536 15004 6588
rect 14948 6524 15004 6536
rect 14948 6472 14950 6524
rect 15002 6472 15004 6524
rect 14948 6460 15004 6472
rect 14948 6408 14950 6460
rect 15002 6408 15004 6460
rect 14948 6396 15004 6408
rect 14948 6344 14950 6396
rect 15002 6344 15004 6396
rect 14948 6332 15004 6344
rect 14948 6280 14950 6332
rect 15002 6280 15004 6332
rect 14948 6268 15004 6280
rect 14948 6216 14950 6268
rect 15002 6216 15004 6268
rect 14948 6204 15004 6216
rect 14948 6152 14950 6204
rect 15002 6152 15004 6204
rect 14948 6140 15004 6152
rect 14948 6088 14950 6140
rect 15002 6088 15004 6140
rect 14948 6076 15004 6088
rect 14948 6024 14950 6076
rect 15002 6024 15004 6076
rect 14948 6012 15004 6024
rect 14948 5960 14950 6012
rect 15002 5960 15004 6012
rect 14948 5948 15004 5960
rect 14948 5896 14950 5948
rect 15002 5896 15004 5948
rect 14948 5750 15004 5896
rect 15170 6844 15226 6858
rect 15170 6792 15172 6844
rect 15224 6792 15226 6844
rect 15170 6780 15226 6792
rect 15170 6728 15172 6780
rect 15224 6728 15226 6780
rect 15170 6716 15226 6728
rect 15170 6664 15172 6716
rect 15224 6664 15226 6716
rect 15170 6652 15226 6664
rect 15170 6600 15172 6652
rect 15224 6600 15226 6652
rect 15170 6588 15226 6600
rect 15170 6536 15172 6588
rect 15224 6536 15226 6588
rect 15170 6524 15226 6536
rect 15170 6472 15172 6524
rect 15224 6472 15226 6524
rect 15170 6460 15226 6472
rect 15170 6408 15172 6460
rect 15224 6408 15226 6460
rect 15170 6396 15226 6408
rect 15170 6344 15172 6396
rect 15224 6344 15226 6396
rect 15170 6332 15226 6344
rect 15170 6280 15172 6332
rect 15224 6280 15226 6332
rect 15170 6268 15226 6280
rect 15170 6216 15172 6268
rect 15224 6216 15226 6268
rect 15170 6204 15226 6216
rect 15170 6152 15172 6204
rect 15224 6152 15226 6204
rect 15170 6140 15226 6152
rect 15170 6088 15172 6140
rect 15224 6088 15226 6140
rect 15170 6076 15226 6088
rect 15170 6024 15172 6076
rect 15224 6024 15226 6076
rect 15170 6012 15226 6024
rect 15170 5960 15172 6012
rect 15224 5960 15226 6012
rect 15170 5948 15226 5960
rect 15170 5896 15172 5948
rect 15224 5896 15226 5948
rect 15170 5750 15226 5896
rect 15256 6810 15312 6950
rect 15256 6758 15258 6810
rect 15310 6758 15312 6810
rect 15256 6746 15312 6758
rect 15256 6694 15258 6746
rect 15310 6694 15312 6746
rect 15256 6682 15312 6694
rect 15256 6630 15258 6682
rect 15310 6630 15312 6682
rect 15256 6618 15312 6630
rect 15256 6566 15258 6618
rect 15310 6566 15312 6618
rect 15256 6554 15312 6566
rect 15256 6502 15258 6554
rect 15310 6502 15312 6554
rect 15256 6490 15312 6502
rect 15256 6438 15258 6490
rect 15310 6438 15312 6490
rect 15256 6426 15312 6438
rect 15256 6374 15258 6426
rect 15310 6374 15312 6426
rect 15256 6362 15312 6374
rect 15256 6310 15258 6362
rect 15310 6310 15312 6362
rect 15256 6298 15312 6310
rect 15256 6246 15258 6298
rect 15310 6246 15312 6298
rect 15256 6234 15312 6246
rect 15256 6182 15258 6234
rect 15310 6182 15312 6234
rect 15256 6170 15312 6182
rect 15256 6118 15258 6170
rect 15310 6118 15312 6170
rect 15256 6106 15312 6118
rect 15256 6054 15258 6106
rect 15310 6054 15312 6106
rect 15256 6042 15312 6054
rect 15256 5990 15258 6042
rect 15310 5990 15312 6042
rect 15256 5978 15312 5990
rect 15256 5926 15258 5978
rect 15310 5926 15312 5978
rect 15256 5914 15312 5926
rect 15256 5862 15258 5914
rect 15310 5862 15312 5914
rect 15256 5848 15312 5862
rect 15342 6844 15398 6858
rect 15342 6792 15344 6844
rect 15396 6792 15398 6844
rect 15342 6780 15398 6792
rect 15342 6728 15344 6780
rect 15396 6728 15398 6780
rect 15342 6716 15398 6728
rect 15342 6664 15344 6716
rect 15396 6664 15398 6716
rect 15342 6652 15398 6664
rect 15342 6600 15344 6652
rect 15396 6600 15398 6652
rect 15342 6588 15398 6600
rect 15342 6536 15344 6588
rect 15396 6536 15398 6588
rect 15342 6524 15398 6536
rect 15342 6472 15344 6524
rect 15396 6472 15398 6524
rect 15342 6460 15398 6472
rect 15342 6408 15344 6460
rect 15396 6408 15398 6460
rect 15342 6396 15398 6408
rect 15342 6344 15344 6396
rect 15396 6344 15398 6396
rect 15342 6332 15398 6344
rect 15342 6280 15344 6332
rect 15396 6280 15398 6332
rect 15342 6268 15398 6280
rect 15342 6216 15344 6268
rect 15396 6216 15398 6268
rect 15342 6204 15398 6216
rect 15342 6152 15344 6204
rect 15396 6152 15398 6204
rect 15342 6140 15398 6152
rect 15342 6088 15344 6140
rect 15396 6088 15398 6140
rect 15342 6076 15398 6088
rect 15342 6024 15344 6076
rect 15396 6024 15398 6076
rect 15342 6012 15398 6024
rect 15342 5960 15344 6012
rect 15396 5960 15398 6012
rect 15342 5948 15398 5960
rect 15342 5896 15344 5948
rect 15396 5896 15398 5948
rect 15342 5750 15398 5896
rect 15428 6810 15484 6950
rect 15428 6758 15430 6810
rect 15482 6758 15484 6810
rect 15428 6746 15484 6758
rect 15428 6694 15430 6746
rect 15482 6694 15484 6746
rect 15428 6682 15484 6694
rect 15428 6630 15430 6682
rect 15482 6630 15484 6682
rect 15428 6618 15484 6630
rect 15428 6566 15430 6618
rect 15482 6566 15484 6618
rect 15428 6554 15484 6566
rect 15428 6502 15430 6554
rect 15482 6502 15484 6554
rect 15428 6490 15484 6502
rect 15428 6438 15430 6490
rect 15482 6438 15484 6490
rect 15428 6426 15484 6438
rect 15428 6374 15430 6426
rect 15482 6374 15484 6426
rect 15428 6362 15484 6374
rect 15428 6310 15430 6362
rect 15482 6310 15484 6362
rect 15428 6298 15484 6310
rect 15428 6246 15430 6298
rect 15482 6246 15484 6298
rect 15428 6234 15484 6246
rect 15428 6182 15430 6234
rect 15482 6182 15484 6234
rect 15428 6170 15484 6182
rect 15428 6118 15430 6170
rect 15482 6118 15484 6170
rect 15428 6106 15484 6118
rect 15428 6054 15430 6106
rect 15482 6054 15484 6106
rect 15428 6042 15484 6054
rect 15428 5990 15430 6042
rect 15482 5990 15484 6042
rect 15428 5978 15484 5990
rect 15428 5926 15430 5978
rect 15482 5926 15484 5978
rect 15428 5914 15484 5926
rect 15428 5862 15430 5914
rect 15482 5862 15484 5914
rect 15428 5848 15484 5862
rect 15514 6844 15570 6858
rect 15514 6792 15516 6844
rect 15568 6792 15570 6844
rect 15514 6780 15570 6792
rect 15514 6728 15516 6780
rect 15568 6728 15570 6780
rect 15514 6716 15570 6728
rect 15514 6664 15516 6716
rect 15568 6664 15570 6716
rect 15514 6652 15570 6664
rect 15514 6600 15516 6652
rect 15568 6600 15570 6652
rect 15514 6588 15570 6600
rect 15514 6536 15516 6588
rect 15568 6536 15570 6588
rect 15514 6524 15570 6536
rect 15514 6472 15516 6524
rect 15568 6472 15570 6524
rect 15514 6460 15570 6472
rect 15514 6408 15516 6460
rect 15568 6408 15570 6460
rect 15514 6396 15570 6408
rect 15800 6400 16050 6980
rect 16195 6941 16247 7049
rect 16367 7901 16419 7971
rect 16367 7821 16419 7849
rect 16367 7741 16419 7769
rect 16367 7661 16419 7689
rect 16367 7581 16419 7609
rect 16367 7501 16419 7529
rect 16367 7421 16419 7449
rect 16367 7341 16419 7369
rect 16367 7261 16419 7289
rect 16367 7181 16419 7209
rect 16367 7101 16419 7129
rect 16367 6941 16419 7049
rect 16539 7901 16591 7971
rect 16539 7821 16591 7849
rect 16539 7741 16591 7769
rect 16539 7661 16591 7689
rect 16539 7581 16591 7609
rect 16539 7501 16591 7529
rect 16539 7421 16591 7449
rect 16539 7341 16591 7369
rect 16539 7261 16591 7289
rect 16539 7181 16591 7209
rect 16539 7101 16591 7129
rect 16539 6941 16591 7049
rect 16711 7901 16763 7971
rect 16711 7821 16763 7849
rect 16711 7741 16763 7769
rect 16711 7661 16763 7689
rect 16711 7581 16763 7609
rect 16711 7501 16763 7529
rect 16711 7421 16763 7449
rect 16711 7341 16763 7369
rect 16711 7261 16763 7289
rect 16711 7181 16763 7209
rect 16711 7101 16763 7129
rect 16711 6941 16763 7049
rect 16883 7901 16935 7971
rect 16883 7821 16935 7849
rect 16883 7741 16935 7769
rect 16883 7661 16935 7689
rect 16883 7581 16935 7609
rect 16883 7501 16935 7529
rect 16883 7421 16935 7449
rect 16883 7341 16935 7369
rect 16883 7261 16935 7289
rect 16883 7181 16935 7209
rect 16883 7101 16935 7129
rect 16883 6941 16935 7049
rect 17055 7901 17107 7971
rect 20160 7940 20230 8040
rect 17055 7821 17107 7849
rect 17055 7741 17107 7769
rect 17055 7661 17107 7689
rect 17055 7581 17107 7609
rect 17055 7501 17107 7529
rect 17055 7421 17107 7449
rect 17055 7341 17107 7369
rect 17055 7261 17107 7289
rect 17055 7181 17107 7209
rect 17055 7101 17107 7129
rect 20050 7930 20230 7940
rect 17055 6941 17107 7049
rect 17692 7109 17758 7118
rect 17692 7053 17697 7109
rect 17753 7053 17758 7109
rect 17692 7047 17699 7053
rect 17751 7047 17758 7053
rect 17692 7035 17758 7047
rect 17692 7029 17699 7035
rect 17751 7029 17758 7035
rect 17170 6990 17340 7010
rect 17170 6941 17180 6990
rect 16129 6870 17180 6941
rect 17330 6870 17340 6990
rect 17692 6973 17697 7029
rect 17753 6973 17758 7029
rect 17692 6964 17758 6973
rect 17864 7109 17930 7118
rect 17864 7053 17869 7109
rect 17925 7053 17930 7109
rect 17864 7047 17871 7053
rect 17923 7047 17930 7053
rect 17864 7035 17930 7047
rect 17864 7029 17871 7035
rect 17923 7029 17930 7035
rect 17864 6973 17869 7029
rect 17925 6973 17930 7029
rect 17864 6964 17930 6973
rect 18036 7109 18102 7118
rect 18036 7053 18041 7109
rect 18097 7053 18102 7109
rect 18036 7047 18043 7053
rect 18095 7047 18102 7053
rect 18036 7035 18102 7047
rect 18036 7029 18043 7035
rect 18095 7029 18102 7035
rect 18036 6973 18041 7029
rect 18097 6973 18102 7029
rect 18036 6964 18102 6973
rect 18208 7109 18274 7118
rect 18208 7053 18213 7109
rect 18269 7053 18274 7109
rect 18208 7047 18215 7053
rect 18267 7047 18274 7053
rect 18208 7035 18274 7047
rect 18208 7029 18215 7035
rect 18267 7029 18274 7035
rect 18208 6973 18213 7029
rect 18269 6973 18274 7029
rect 18208 6964 18274 6973
rect 18380 7109 18446 7118
rect 18380 7053 18385 7109
rect 18441 7053 18446 7109
rect 18380 7047 18387 7053
rect 18439 7047 18446 7053
rect 18380 7035 18446 7047
rect 18380 7029 18387 7035
rect 18439 7029 18446 7035
rect 18380 6973 18385 7029
rect 18441 6973 18446 7029
rect 18380 6964 18446 6973
rect 18552 7109 18618 7118
rect 18552 7053 18557 7109
rect 18613 7053 18618 7109
rect 18552 7047 18559 7053
rect 18611 7047 18618 7053
rect 18552 7035 18618 7047
rect 18552 7029 18559 7035
rect 18611 7029 18618 7035
rect 18552 6973 18557 7029
rect 18613 6973 18618 7029
rect 18552 6964 18618 6973
rect 18724 7109 18790 7118
rect 18724 7053 18729 7109
rect 18785 7053 18790 7109
rect 18724 7047 18731 7053
rect 18783 7047 18790 7053
rect 18724 7035 18790 7047
rect 18724 7029 18731 7035
rect 18783 7029 18790 7035
rect 18724 6973 18729 7029
rect 18785 6973 18790 7029
rect 18724 6964 18790 6973
rect 18896 7109 18962 7118
rect 18896 7053 18901 7109
rect 18957 7053 18962 7109
rect 18896 7047 18903 7053
rect 18955 7047 18962 7053
rect 18896 7035 18962 7047
rect 18896 7029 18903 7035
rect 18955 7029 18962 7035
rect 18896 6973 18901 7029
rect 18957 6973 18962 7029
rect 18896 6964 18962 6973
rect 19068 7109 19134 7118
rect 19068 7053 19073 7109
rect 19129 7053 19134 7109
rect 19068 7047 19075 7053
rect 19127 7047 19134 7053
rect 19068 7035 19134 7047
rect 19068 7029 19075 7035
rect 19127 7029 19134 7035
rect 19068 6973 19073 7029
rect 19129 6973 19134 7029
rect 19068 6964 19134 6973
rect 19240 7109 19306 7118
rect 19240 7053 19245 7109
rect 19301 7053 19306 7109
rect 19240 7047 19247 7053
rect 19299 7047 19306 7053
rect 19240 7035 19306 7047
rect 19240 7029 19247 7035
rect 19299 7029 19306 7035
rect 19240 6973 19245 7029
rect 19301 6973 19306 7029
rect 19240 6964 19306 6973
rect 19412 7109 19478 7118
rect 19412 7053 19417 7109
rect 19473 7053 19478 7109
rect 19412 7047 19419 7053
rect 19471 7047 19478 7053
rect 19412 7035 19478 7047
rect 19412 7029 19419 7035
rect 19471 7029 19478 7035
rect 19412 6973 19417 7029
rect 19473 6973 19478 7029
rect 19412 6964 19478 6973
rect 19584 7109 19650 7118
rect 19584 7053 19589 7109
rect 19645 7053 19650 7109
rect 19584 7047 19591 7053
rect 19643 7047 19650 7053
rect 19584 7035 19650 7047
rect 19584 7029 19591 7035
rect 19643 7029 19650 7035
rect 19584 6973 19589 7029
rect 19645 6973 19650 7029
rect 19584 6964 19650 6973
rect 19756 7109 19822 7118
rect 19756 7053 19761 7109
rect 19817 7053 19822 7109
rect 19756 7047 19763 7053
rect 19815 7047 19822 7053
rect 19756 7035 19822 7047
rect 19756 7029 19763 7035
rect 19815 7029 19822 7035
rect 19756 6973 19761 7029
rect 19817 6973 19822 7029
rect 19756 6964 19822 6973
rect 19928 7109 19994 7118
rect 19928 7053 19933 7109
rect 19989 7053 19994 7109
rect 19928 7047 19935 7053
rect 19987 7047 19994 7053
rect 19928 7035 19994 7047
rect 19928 7029 19935 7035
rect 19987 7029 19994 7035
rect 19928 6973 19933 7029
rect 19989 6973 19994 7029
rect 19928 6964 19994 6973
rect 20050 7000 20060 7930
rect 20180 7900 20230 7930
rect 20180 7000 20300 7900
rect 16129 6861 17340 6870
rect 16130 6860 17340 6861
rect 16130 6820 20010 6830
rect 16130 6810 17440 6820
rect 16130 6750 16140 6810
rect 17130 6750 17440 6810
rect 16130 6720 17440 6750
rect 17590 6720 17680 6820
rect 16130 6710 17680 6720
rect 20000 6710 20010 6820
rect 16130 6690 20010 6710
rect 17650 6500 20000 6510
rect 17650 6490 17660 6500
rect 17330 6480 17660 6490
rect 15514 6344 15516 6396
rect 15568 6344 15570 6396
rect 15514 6332 15570 6344
rect 15514 6280 15516 6332
rect 15568 6280 15570 6332
rect 15514 6268 15570 6280
rect 15514 6216 15516 6268
rect 15568 6216 15570 6268
rect 15514 6204 15570 6216
rect 15514 6152 15516 6204
rect 15568 6152 15570 6204
rect 15514 6140 15570 6152
rect 15514 6088 15516 6140
rect 15568 6088 15570 6140
rect 15514 6076 15570 6088
rect 15514 6024 15516 6076
rect 15568 6024 15570 6076
rect 15514 6012 15570 6024
rect 15514 5960 15516 6012
rect 15568 5960 15570 6012
rect 15514 5948 15570 5960
rect 15514 5896 15516 5948
rect 15568 5896 15570 5948
rect 15514 5750 15570 5896
rect 15900 6180 16050 6400
rect 16130 6470 17660 6480
rect 16130 6410 17180 6470
rect 16130 6350 16140 6410
rect 17170 6370 17180 6410
rect 17330 6390 17660 6470
rect 19980 6390 20000 6500
rect 17330 6380 20000 6390
rect 17330 6370 17340 6380
rect 17170 6360 17340 6370
rect 17170 6350 17210 6360
rect 16130 6340 17210 6350
rect 17400 6330 17600 6340
rect 17400 6310 17440 6330
rect 17190 6300 17440 6310
rect 16130 6299 17440 6300
rect 16129 6230 17440 6299
rect 17590 6230 17600 6330
rect 16129 6220 17600 6230
rect 16129 6219 17197 6220
rect 15900 6160 16110 6180
rect 11600 5730 15700 5750
rect 11600 5670 11620 5730
rect 15680 5670 15700 5730
rect 11600 5650 15700 5670
rect 11840 5580 12680 5590
rect 11840 5570 12410 5580
rect 11840 5510 11860 5570
rect 12100 5520 12410 5570
rect 12670 5520 12680 5580
rect 12100 5510 12420 5520
rect 12660 5510 12680 5520
rect 12960 5580 13240 5590
rect 12960 5520 12970 5580
rect 13230 5520 13240 5580
rect 12960 5510 12980 5520
rect 13220 5510 13240 5520
rect 13540 5580 13820 5590
rect 13540 5520 13550 5580
rect 13810 5520 13820 5580
rect 13540 5510 13560 5520
rect 13800 5510 13820 5520
rect 14100 5580 14380 5590
rect 14100 5520 14110 5580
rect 14370 5520 14380 5580
rect 14100 5510 14120 5520
rect 14360 5510 14380 5520
rect 14680 5580 15520 5590
rect 14680 5520 14690 5580
rect 14950 5570 15520 5580
rect 14950 5520 15260 5570
rect 14680 5510 14700 5520
rect 14940 5510 15260 5520
rect 15500 5510 15520 5570
rect 15900 5470 15960 6160
rect 11640 5460 15960 5470
rect 11640 5380 11650 5460
rect 15690 5440 15960 5460
rect 11640 5300 11920 5380
rect 12280 5300 13220 5380
rect 13580 5300 14320 5380
rect 14680 5300 15540 5380
rect 15880 5300 15960 5440
rect 11640 5280 15960 5300
rect 15900 5050 15960 5280
rect 16100 5076 16110 6160
rect 16195 6111 16247 6219
rect 16195 6031 16247 6059
rect 16195 5951 16247 5979
rect 16195 5871 16247 5899
rect 16195 5791 16247 5819
rect 16195 5711 16247 5739
rect 16195 5631 16247 5659
rect 16195 5551 16247 5579
rect 16195 5471 16247 5499
rect 16195 5391 16247 5419
rect 16195 5311 16247 5339
rect 16195 5189 16247 5259
rect 16367 6111 16419 6219
rect 16367 6031 16419 6059
rect 16367 5951 16419 5979
rect 16367 5871 16419 5899
rect 16367 5791 16419 5819
rect 16367 5711 16419 5739
rect 16367 5631 16419 5659
rect 16367 5551 16419 5579
rect 16367 5471 16419 5499
rect 16367 5391 16419 5419
rect 16367 5311 16419 5339
rect 16367 5189 16419 5259
rect 16539 6111 16591 6219
rect 16539 6031 16591 6059
rect 16539 5951 16591 5979
rect 16539 5871 16591 5899
rect 16539 5791 16591 5819
rect 16539 5711 16591 5739
rect 16539 5631 16591 5659
rect 16539 5551 16591 5579
rect 16539 5471 16591 5499
rect 16539 5391 16591 5419
rect 16539 5311 16591 5339
rect 16539 5189 16591 5259
rect 16711 6111 16763 6219
rect 16711 6031 16763 6059
rect 16711 5951 16763 5979
rect 16711 5871 16763 5899
rect 16711 5791 16763 5819
rect 16711 5711 16763 5739
rect 16711 5631 16763 5659
rect 16711 5551 16763 5579
rect 16711 5471 16763 5499
rect 16711 5391 16763 5419
rect 16711 5311 16763 5339
rect 16711 5189 16763 5259
rect 16883 6111 16935 6219
rect 16883 6031 16935 6059
rect 16883 5951 16935 5979
rect 16883 5871 16935 5899
rect 16883 5791 16935 5819
rect 16883 5711 16935 5739
rect 16883 5631 16935 5659
rect 16883 5551 16935 5579
rect 16883 5471 16935 5499
rect 16883 5391 16935 5419
rect 16883 5311 16935 5339
rect 16883 5189 16935 5259
rect 17055 6111 17107 6219
rect 17674 6217 17740 6226
rect 17674 6161 17679 6217
rect 17735 6161 17740 6217
rect 17674 6155 17681 6161
rect 17733 6155 17740 6161
rect 17674 6143 17740 6155
rect 17674 6137 17681 6143
rect 17733 6137 17740 6143
rect 17674 6081 17679 6137
rect 17735 6081 17740 6137
rect 17674 6072 17740 6081
rect 17846 6217 17912 6226
rect 17846 6161 17851 6217
rect 17907 6161 17912 6217
rect 17846 6155 17853 6161
rect 17905 6155 17912 6161
rect 17846 6143 17912 6155
rect 17846 6137 17853 6143
rect 17905 6137 17912 6143
rect 17846 6081 17851 6137
rect 17907 6081 17912 6137
rect 17846 6072 17912 6081
rect 18018 6217 18084 6226
rect 18018 6161 18023 6217
rect 18079 6161 18084 6217
rect 18018 6155 18025 6161
rect 18077 6155 18084 6161
rect 18018 6143 18084 6155
rect 18018 6137 18025 6143
rect 18077 6137 18084 6143
rect 18018 6081 18023 6137
rect 18079 6081 18084 6137
rect 18018 6072 18084 6081
rect 18190 6217 18256 6226
rect 18190 6161 18195 6217
rect 18251 6161 18256 6217
rect 18190 6155 18197 6161
rect 18249 6155 18256 6161
rect 18190 6143 18256 6155
rect 18190 6137 18197 6143
rect 18249 6137 18256 6143
rect 18190 6081 18195 6137
rect 18251 6081 18256 6137
rect 18190 6072 18256 6081
rect 18362 6217 18428 6226
rect 18362 6161 18367 6217
rect 18423 6161 18428 6217
rect 18362 6155 18369 6161
rect 18421 6155 18428 6161
rect 18362 6143 18428 6155
rect 18362 6137 18369 6143
rect 18421 6137 18428 6143
rect 18362 6081 18367 6137
rect 18423 6081 18428 6137
rect 18362 6072 18428 6081
rect 18534 6217 18600 6226
rect 18534 6161 18539 6217
rect 18595 6161 18600 6217
rect 18534 6155 18541 6161
rect 18593 6155 18600 6161
rect 18534 6143 18600 6155
rect 18534 6137 18541 6143
rect 18593 6137 18600 6143
rect 18534 6081 18539 6137
rect 18595 6081 18600 6137
rect 18534 6072 18600 6081
rect 18706 6217 18772 6226
rect 18706 6161 18711 6217
rect 18767 6161 18772 6217
rect 18706 6155 18713 6161
rect 18765 6155 18772 6161
rect 18706 6143 18772 6155
rect 18706 6137 18713 6143
rect 18765 6137 18772 6143
rect 18706 6081 18711 6137
rect 18767 6081 18772 6137
rect 18706 6072 18772 6081
rect 18878 6217 18944 6226
rect 18878 6161 18883 6217
rect 18939 6161 18944 6217
rect 18878 6155 18885 6161
rect 18937 6155 18944 6161
rect 18878 6143 18944 6155
rect 18878 6137 18885 6143
rect 18937 6137 18944 6143
rect 18878 6081 18883 6137
rect 18939 6081 18944 6137
rect 18878 6072 18944 6081
rect 19050 6217 19116 6226
rect 19050 6161 19055 6217
rect 19111 6161 19116 6217
rect 19050 6155 19057 6161
rect 19109 6155 19116 6161
rect 19050 6143 19116 6155
rect 19050 6137 19057 6143
rect 19109 6137 19116 6143
rect 19050 6081 19055 6137
rect 19111 6081 19116 6137
rect 19050 6072 19116 6081
rect 19222 6217 19288 6226
rect 19222 6161 19227 6217
rect 19283 6161 19288 6217
rect 19222 6155 19229 6161
rect 19281 6155 19288 6161
rect 19222 6143 19288 6155
rect 19222 6137 19229 6143
rect 19281 6137 19288 6143
rect 19222 6081 19227 6137
rect 19283 6081 19288 6137
rect 19222 6072 19288 6081
rect 19394 6217 19460 6226
rect 19394 6161 19399 6217
rect 19455 6161 19460 6217
rect 19394 6155 19401 6161
rect 19453 6155 19460 6161
rect 19394 6143 19460 6155
rect 19394 6137 19401 6143
rect 19453 6137 19460 6143
rect 19394 6081 19399 6137
rect 19455 6081 19460 6137
rect 19394 6072 19460 6081
rect 19566 6217 19632 6226
rect 19566 6161 19571 6217
rect 19627 6161 19632 6217
rect 19566 6155 19573 6161
rect 19625 6155 19632 6161
rect 19566 6143 19632 6155
rect 19566 6137 19573 6143
rect 19625 6137 19632 6143
rect 19566 6081 19571 6137
rect 19627 6081 19632 6137
rect 19566 6072 19632 6081
rect 19738 6217 19804 6226
rect 19738 6161 19743 6217
rect 19799 6161 19804 6217
rect 19738 6155 19745 6161
rect 19797 6155 19804 6161
rect 19738 6143 19804 6155
rect 19738 6137 19745 6143
rect 19797 6137 19804 6143
rect 19738 6081 19743 6137
rect 19799 6081 19804 6137
rect 19738 6072 19804 6081
rect 19910 6217 19976 6226
rect 19910 6161 19915 6217
rect 19971 6161 19976 6217
rect 19910 6155 19917 6161
rect 19969 6155 19976 6161
rect 19910 6143 19976 6155
rect 19910 6137 19917 6143
rect 19969 6137 19976 6143
rect 19910 6081 19915 6137
rect 19971 6081 19976 6137
rect 19910 6072 19976 6081
rect 20050 6190 20300 7000
rect 17055 6031 17107 6059
rect 17055 5951 17107 5979
rect 17055 5871 17107 5899
rect 17055 5791 17107 5819
rect 17055 5711 17107 5739
rect 17055 5631 17107 5659
rect 17055 5551 17107 5579
rect 17055 5471 17107 5499
rect 17055 5391 17107 5419
rect 17055 5311 17107 5339
rect 17055 5189 17107 5259
rect 20050 5260 20060 6190
rect 20180 5260 20300 6190
rect 20050 5250 20300 5260
rect 20060 5140 20300 5250
rect 17380 5100 20300 5140
rect 16100 5050 16111 5076
rect 15900 5039 16111 5050
rect 15900 4818 16577 5039
rect 17380 5000 17420 5100
rect 20140 5000 20300 5100
rect 17380 4960 20300 5000
rect 15900 4813 17353 4818
rect 15900 4811 16648 4813
rect 16704 4811 16728 4813
rect 16784 4811 16808 4813
rect 16864 4811 16888 4813
rect 16944 4811 16968 4813
rect 17024 4811 17048 4813
rect 17104 4811 17128 4813
rect 17184 4811 17208 4813
rect 17264 4811 17288 4813
rect 15900 4781 16638 4811
rect 15909 4765 16638 4781
rect 15909 4714 16557 4765
rect 16609 4759 16638 4765
rect 16882 4759 16888 4811
rect 16946 4759 16958 4811
rect 17202 4759 17208 4811
rect 17266 4759 17278 4811
rect 16609 4757 16648 4759
rect 16704 4757 16728 4759
rect 16784 4757 16808 4759
rect 16864 4757 16888 4759
rect 16944 4757 16968 4759
rect 17024 4757 17048 4759
rect 17104 4757 17128 4759
rect 17184 4757 17208 4759
rect 17264 4757 17288 4759
rect 17344 4757 17353 4813
rect 16609 4752 17353 4757
rect 16609 4714 16616 4752
rect 17381 4724 17435 4960
rect 17463 4813 18266 4818
rect 17463 4757 17472 4813
rect 17528 4811 17552 4813
rect 17608 4811 17632 4813
rect 17688 4811 17712 4813
rect 17768 4811 17792 4813
rect 17848 4811 17872 4813
rect 17928 4811 17952 4813
rect 18008 4811 18032 4813
rect 18088 4811 18112 4813
rect 18168 4811 18266 4813
rect 17544 4759 17552 4811
rect 17608 4759 17620 4811
rect 17864 4759 17872 4811
rect 17928 4759 17940 4811
rect 18184 4765 18266 4811
rect 18184 4759 18207 4765
rect 17528 4757 17552 4759
rect 17608 4757 17632 4759
rect 17688 4757 17712 4759
rect 17768 4757 17792 4759
rect 17848 4757 17872 4759
rect 17928 4757 17952 4759
rect 18008 4757 18032 4759
rect 18088 4757 18112 4759
rect 18168 4757 18207 4759
rect 17463 4752 18207 4757
rect 15909 4658 16555 4714
rect 16611 4668 16616 4714
rect 16644 4718 18172 4724
rect 16644 4696 17382 4718
rect 16611 4658 17352 4668
rect 15909 4649 16557 4658
rect 16609 4649 17352 4658
rect 15909 4640 17352 4649
rect 17380 4666 17382 4696
rect 17434 4696 18172 4718
rect 18200 4714 18207 4752
rect 18259 4714 18266 4765
rect 17434 4666 17436 4696
rect 18200 4668 18205 4714
rect 17380 4654 17436 4666
rect 15909 4637 16616 4640
rect 15909 4634 16557 4637
rect 16609 4634 16616 4637
rect 15909 4626 16555 4634
rect 16550 4578 16555 4626
rect 16611 4578 16616 4634
rect 17380 4612 17382 4654
rect 16644 4602 17382 4612
rect 17434 4612 17436 4654
rect 17464 4658 18205 4668
rect 18261 4658 18266 4714
rect 17464 4649 18207 4658
rect 18259 4649 18266 4658
rect 17464 4640 18266 4649
rect 18200 4637 18266 4640
rect 18200 4634 18207 4637
rect 18259 4634 18266 4637
rect 17434 4602 18172 4612
rect 16644 4590 18172 4602
rect 16644 4584 17382 4590
rect 16550 4573 16616 4578
rect 16550 4554 16557 4573
rect 16609 4556 16616 4573
rect 16609 4554 17352 4556
rect 16550 4498 16555 4554
rect 16611 4528 17352 4554
rect 17380 4538 17382 4584
rect 17434 4584 18172 4590
rect 17434 4538 17436 4584
rect 18200 4578 18205 4634
rect 18261 4578 18266 4634
rect 18200 4573 18266 4578
rect 18200 4556 18207 4573
rect 16611 4498 16616 4528
rect 17380 4526 17436 4538
rect 17464 4554 18207 4556
rect 18259 4554 18266 4573
rect 17464 4528 18205 4554
rect 17380 4500 17382 4526
rect 16550 4474 16557 4498
rect 16609 4474 16616 4498
rect 16550 4418 16555 4474
rect 16611 4444 16616 4474
rect 16644 4474 17382 4500
rect 17434 4500 17436 4526
rect 17434 4474 18172 4500
rect 16644 4472 18172 4474
rect 18200 4498 18205 4528
rect 18261 4498 18266 4554
rect 18200 4474 18207 4498
rect 18259 4474 18266 4498
rect 17380 4462 17436 4472
rect 16611 4418 17352 4444
rect 16550 4394 16557 4418
rect 16609 4416 17352 4418
rect 16609 4394 16616 4416
rect 16550 4338 16555 4394
rect 16611 4338 16616 4394
rect 17380 4410 17382 4462
rect 17434 4410 17436 4462
rect 18200 4444 18205 4474
rect 17464 4418 18205 4444
rect 18261 4418 18266 4474
rect 17464 4416 18207 4418
rect 17380 4398 17436 4410
rect 17380 4388 17382 4398
rect 16644 4360 17382 4388
rect 16550 4329 16557 4338
rect 16609 4332 16616 4338
rect 17380 4346 17382 4360
rect 17434 4388 17436 4398
rect 18200 4394 18207 4416
rect 18259 4394 18266 4418
rect 17434 4360 18172 4388
rect 17434 4346 17436 4360
rect 17380 4334 17436 4346
rect 16609 4329 17352 4332
rect 16550 4317 17352 4329
rect 16550 4314 16557 4317
rect 16609 4314 17352 4317
rect 16550 4258 16555 4314
rect 16611 4304 17352 4314
rect 16611 4258 16616 4304
rect 17380 4282 17382 4334
rect 17434 4282 17436 4334
rect 18200 4338 18205 4394
rect 18261 4338 18266 4394
rect 18200 4332 18207 4338
rect 17464 4329 18207 4332
rect 18259 4329 18266 4338
rect 17464 4317 18266 4329
rect 17464 4314 18207 4317
rect 18259 4314 18266 4317
rect 17464 4304 18205 4314
rect 17380 4276 17436 4282
rect 16550 4253 16616 4258
rect 16550 4234 16557 4253
rect 16609 4234 16616 4253
rect 16644 4270 18172 4276
rect 16644 4248 17382 4270
rect 16550 4178 16555 4234
rect 16611 4220 16616 4234
rect 16611 4192 17352 4220
rect 17380 4218 17382 4248
rect 17434 4248 18172 4270
rect 18200 4258 18205 4304
rect 18261 4258 18266 4314
rect 18200 4253 18266 4258
rect 17434 4218 17436 4248
rect 18200 4234 18207 4253
rect 18259 4234 18266 4253
rect 18200 4220 18205 4234
rect 17380 4206 17436 4218
rect 16611 4178 16616 4192
rect 16550 4154 16557 4178
rect 16609 4154 16616 4178
rect 17380 4164 17382 4206
rect 16550 4098 16555 4154
rect 16611 4098 16616 4154
rect 16550 4089 16616 4098
rect 16644 4154 17382 4164
rect 17434 4164 17436 4206
rect 17464 4192 18205 4220
rect 18200 4178 18205 4192
rect 18261 4178 18266 4234
rect 17434 4154 18172 4164
rect 16644 4142 18172 4154
rect 16644 4090 17382 4142
rect 17434 4090 18172 4142
rect 18200 4154 18207 4178
rect 18259 4154 18266 4178
rect 18200 4098 18205 4154
rect 18261 4098 18266 4154
rect 17380 4062 17436 4090
rect 18200 4089 18266 4098
rect 16624 4061 16740 4062
rect 16550 4060 16740 4061
rect 16796 4060 16820 4062
rect 16876 4060 16900 4062
rect 16956 4060 16980 4062
rect 17036 4060 17060 4062
rect 17116 4060 17140 4062
rect 17196 4060 17220 4062
rect 17276 4060 17300 4062
rect 16550 4008 16655 4060
rect 16707 4008 16719 4060
rect 16899 4008 16900 4060
rect 16963 4008 16975 4060
rect 17036 4008 17039 4060
rect 17219 4008 17220 4060
rect 17283 4008 17295 4060
rect 16550 4007 16740 4008
rect 16624 4006 16740 4007
rect 16796 4006 16820 4008
rect 16876 4006 16900 4008
rect 16956 4006 16980 4008
rect 17036 4006 17060 4008
rect 17116 4006 17140 4008
rect 17196 4006 17220 4008
rect 17276 4006 17300 4008
rect 17356 4006 17380 4062
rect 17436 4006 17460 4062
rect 17516 4060 17540 4062
rect 17596 4060 17620 4062
rect 17676 4060 17700 4062
rect 17756 4060 17780 4062
rect 17836 4060 17860 4062
rect 17916 4060 17940 4062
rect 17996 4060 18020 4062
rect 18076 4061 18192 4062
rect 18298 4061 18368 4960
rect 18400 4813 19203 4818
rect 18400 4811 18498 4813
rect 18554 4811 18578 4813
rect 18634 4811 18658 4813
rect 18714 4811 18738 4813
rect 18794 4811 18818 4813
rect 18874 4811 18898 4813
rect 18954 4811 18978 4813
rect 19034 4811 19058 4813
rect 19114 4811 19138 4813
rect 18400 4765 18488 4811
rect 18400 4714 18407 4765
rect 18459 4759 18488 4765
rect 18732 4759 18738 4811
rect 18796 4759 18808 4811
rect 19052 4759 19058 4811
rect 19116 4759 19128 4811
rect 18459 4757 18498 4759
rect 18554 4757 18578 4759
rect 18634 4757 18658 4759
rect 18714 4757 18738 4759
rect 18794 4757 18818 4759
rect 18874 4757 18898 4759
rect 18954 4757 18978 4759
rect 19034 4757 19058 4759
rect 19114 4757 19138 4759
rect 19194 4757 19203 4813
rect 18459 4752 19203 4757
rect 18459 4714 18466 4752
rect 19231 4724 19285 4960
rect 19313 4813 20116 4818
rect 19313 4757 19322 4813
rect 19378 4811 19402 4813
rect 19458 4811 19482 4813
rect 19538 4811 19562 4813
rect 19618 4811 19642 4813
rect 19698 4811 19722 4813
rect 19778 4811 19802 4813
rect 19858 4811 19882 4813
rect 19938 4811 19962 4813
rect 20018 4811 20116 4813
rect 19394 4759 19402 4811
rect 19458 4759 19470 4811
rect 19714 4759 19722 4811
rect 19778 4759 19790 4811
rect 20034 4765 20116 4811
rect 20034 4759 20057 4765
rect 19378 4757 19402 4759
rect 19458 4757 19482 4759
rect 19538 4757 19562 4759
rect 19618 4757 19642 4759
rect 19698 4757 19722 4759
rect 19778 4757 19802 4759
rect 19858 4757 19882 4759
rect 19938 4757 19962 4759
rect 20018 4757 20057 4759
rect 19313 4752 20057 4757
rect 18400 4658 18405 4714
rect 18461 4668 18466 4714
rect 18494 4718 20022 4724
rect 18494 4696 19232 4718
rect 18461 4658 19202 4668
rect 18400 4649 18407 4658
rect 18459 4649 19202 4658
rect 18400 4640 19202 4649
rect 19230 4666 19232 4696
rect 19284 4696 20022 4718
rect 20050 4714 20057 4752
rect 20109 4714 20116 4765
rect 19284 4666 19286 4696
rect 20050 4668 20055 4714
rect 19230 4654 19286 4666
rect 18400 4637 18466 4640
rect 18400 4634 18407 4637
rect 18459 4634 18466 4637
rect 18400 4578 18405 4634
rect 18461 4578 18466 4634
rect 19230 4612 19232 4654
rect 18494 4602 19232 4612
rect 19284 4612 19286 4654
rect 19314 4658 20055 4668
rect 20111 4658 20116 4714
rect 19314 4649 20057 4658
rect 20109 4649 20116 4658
rect 19314 4640 20116 4649
rect 20050 4637 20116 4640
rect 20050 4634 20057 4637
rect 20109 4634 20116 4637
rect 19284 4602 20022 4612
rect 18494 4590 20022 4602
rect 18494 4584 19232 4590
rect 18400 4573 18466 4578
rect 18400 4554 18407 4573
rect 18459 4556 18466 4573
rect 18459 4554 19202 4556
rect 18400 4498 18405 4554
rect 18461 4528 19202 4554
rect 19230 4538 19232 4584
rect 19284 4584 20022 4590
rect 19284 4538 19286 4584
rect 20050 4578 20055 4634
rect 20111 4578 20116 4634
rect 20050 4573 20116 4578
rect 20050 4556 20057 4573
rect 18461 4498 18466 4528
rect 19230 4526 19286 4538
rect 19314 4554 20057 4556
rect 20109 4554 20116 4573
rect 19314 4528 20055 4554
rect 19230 4500 19232 4526
rect 18400 4474 18407 4498
rect 18459 4474 18466 4498
rect 18400 4418 18405 4474
rect 18461 4444 18466 4474
rect 18494 4474 19232 4500
rect 19284 4500 19286 4526
rect 19284 4474 20022 4500
rect 18494 4472 20022 4474
rect 20050 4498 20055 4528
rect 20111 4498 20116 4554
rect 20050 4474 20057 4498
rect 20109 4474 20116 4498
rect 19230 4462 19286 4472
rect 18461 4418 19202 4444
rect 18400 4394 18407 4418
rect 18459 4416 19202 4418
rect 18459 4394 18466 4416
rect 18400 4338 18405 4394
rect 18461 4338 18466 4394
rect 19230 4410 19232 4462
rect 19284 4410 19286 4462
rect 20050 4444 20055 4474
rect 19314 4418 20055 4444
rect 20111 4418 20116 4474
rect 19314 4416 20057 4418
rect 19230 4398 19286 4410
rect 19230 4388 19232 4398
rect 18494 4360 19232 4388
rect 18400 4329 18407 4338
rect 18459 4332 18466 4338
rect 19230 4346 19232 4360
rect 19284 4388 19286 4398
rect 20050 4394 20057 4416
rect 20109 4394 20116 4418
rect 19284 4360 20022 4388
rect 19284 4346 19286 4360
rect 19230 4334 19286 4346
rect 18459 4329 19202 4332
rect 18400 4317 19202 4329
rect 18400 4314 18407 4317
rect 18459 4314 19202 4317
rect 18400 4258 18405 4314
rect 18461 4304 19202 4314
rect 18461 4258 18466 4304
rect 19230 4282 19232 4334
rect 19284 4282 19286 4334
rect 20050 4338 20055 4394
rect 20111 4338 20116 4394
rect 20050 4332 20057 4338
rect 19314 4329 20057 4332
rect 20109 4329 20116 4338
rect 19314 4317 20116 4329
rect 19314 4314 20057 4317
rect 20109 4314 20116 4317
rect 19314 4304 20055 4314
rect 19230 4276 19286 4282
rect 18400 4253 18466 4258
rect 18400 4234 18407 4253
rect 18459 4234 18466 4253
rect 18494 4270 20022 4276
rect 18494 4248 19232 4270
rect 18400 4178 18405 4234
rect 18461 4220 18466 4234
rect 18461 4192 19202 4220
rect 19230 4218 19232 4248
rect 19284 4248 20022 4270
rect 20050 4258 20055 4304
rect 20111 4258 20116 4314
rect 20050 4253 20116 4258
rect 19284 4218 19286 4248
rect 20050 4234 20057 4253
rect 20109 4234 20116 4253
rect 20050 4220 20055 4234
rect 19230 4206 19286 4218
rect 18461 4178 18466 4192
rect 18400 4154 18407 4178
rect 18459 4154 18466 4178
rect 19230 4164 19232 4206
rect 18400 4098 18405 4154
rect 18461 4098 18466 4154
rect 18400 4089 18466 4098
rect 18494 4154 19232 4164
rect 19284 4164 19286 4206
rect 19314 4192 20055 4220
rect 20050 4178 20055 4192
rect 20111 4178 20116 4234
rect 19284 4154 20022 4164
rect 18494 4142 20022 4154
rect 18494 4090 19232 4142
rect 19284 4090 20022 4142
rect 20050 4154 20057 4178
rect 20109 4154 20116 4178
rect 20050 4098 20055 4154
rect 20111 4098 20116 4154
rect 19230 4062 19286 4090
rect 20050 4089 20116 4098
rect 18474 4061 18590 4062
rect 18076 4060 18590 4061
rect 18646 4060 18670 4062
rect 18726 4060 18750 4062
rect 18806 4060 18830 4062
rect 18886 4060 18910 4062
rect 18966 4060 18990 4062
rect 19046 4060 19070 4062
rect 19126 4060 19150 4062
rect 17521 4008 17533 4060
rect 17596 4008 17597 4060
rect 17777 4008 17780 4060
rect 17841 4008 17853 4060
rect 17916 4008 17917 4060
rect 18097 4008 18109 4060
rect 18161 4008 18505 4060
rect 18557 4008 18569 4060
rect 18749 4008 18750 4060
rect 18813 4008 18825 4060
rect 18886 4008 18889 4060
rect 19069 4008 19070 4060
rect 19133 4008 19145 4060
rect 17516 4006 17540 4008
rect 17596 4006 17620 4008
rect 17676 4006 17700 4008
rect 17756 4006 17780 4008
rect 17836 4006 17860 4008
rect 17916 4006 17940 4008
rect 17996 4006 18020 4008
rect 18076 4007 18590 4008
rect 18076 4006 18192 4007
rect 18474 4006 18590 4007
rect 18646 4006 18670 4008
rect 18726 4006 18750 4008
rect 18806 4006 18830 4008
rect 18886 4006 18910 4008
rect 18966 4006 18990 4008
rect 19046 4006 19070 4008
rect 19126 4006 19150 4008
rect 19206 4006 19230 4062
rect 19286 4006 19310 4062
rect 19366 4060 19390 4062
rect 19446 4060 19470 4062
rect 19526 4060 19550 4062
rect 19606 4060 19630 4062
rect 19686 4060 19710 4062
rect 19766 4060 19790 4062
rect 19846 4060 19870 4062
rect 19926 4061 20042 4062
rect 20150 4061 20300 4960
rect 19926 4060 20300 4061
rect 19371 4008 19383 4060
rect 19446 4008 19447 4060
rect 19627 4008 19630 4060
rect 19691 4008 19703 4060
rect 19766 4008 19767 4060
rect 19947 4008 19959 4060
rect 20011 4008 20300 4060
rect 19366 4006 19390 4008
rect 19446 4006 19470 4008
rect 19526 4006 19550 4008
rect 19606 4006 19630 4008
rect 19686 4006 19710 4008
rect 19766 4006 19790 4008
rect 19846 4006 19870 4008
rect 19926 4007 20300 4008
rect 19926 4006 20042 4007
rect 16550 3970 16616 3979
rect 17380 3978 17436 4006
rect 16550 3914 16555 3970
rect 16611 3914 16616 3970
rect 16550 3890 16557 3914
rect 16609 3890 16616 3914
rect 16644 3926 17382 3978
rect 17434 3926 18172 3978
rect 16644 3914 18172 3926
rect 16644 3904 17382 3914
rect 16550 3834 16555 3890
rect 16611 3876 16616 3890
rect 16611 3848 17352 3876
rect 17380 3862 17382 3904
rect 17434 3904 18172 3914
rect 18200 3970 18466 3979
rect 19230 3978 19286 4006
rect 20150 4005 20300 4007
rect 18200 3914 18205 3970
rect 18261 3914 18405 3970
rect 18461 3914 18466 3970
rect 17434 3862 17436 3904
rect 18200 3890 18207 3914
rect 18259 3890 18407 3914
rect 18459 3890 18466 3914
rect 18494 3926 19232 3978
rect 19284 3926 20022 3978
rect 18494 3914 20022 3926
rect 18494 3904 19232 3914
rect 18200 3876 18205 3890
rect 17380 3850 17436 3862
rect 16611 3834 16616 3848
rect 16550 3815 16557 3834
rect 16609 3815 16616 3834
rect 17380 3820 17382 3850
rect 16550 3810 16616 3815
rect 16550 3754 16555 3810
rect 16611 3764 16616 3810
rect 16644 3798 17382 3820
rect 17434 3820 17436 3850
rect 17464 3848 18205 3876
rect 18200 3834 18205 3848
rect 18261 3834 18405 3890
rect 18461 3876 18466 3890
rect 18461 3848 19202 3876
rect 19230 3862 19232 3904
rect 19284 3904 20022 3914
rect 20050 3970 20116 3979
rect 20050 3914 20055 3970
rect 20111 3914 20116 3970
rect 19284 3862 19286 3904
rect 20050 3890 20057 3914
rect 20109 3890 20116 3914
rect 20050 3876 20055 3890
rect 19230 3850 19286 3862
rect 18461 3834 18466 3848
rect 17434 3798 18172 3820
rect 16644 3792 18172 3798
rect 18200 3815 18207 3834
rect 18259 3815 18407 3834
rect 18459 3815 18466 3834
rect 19230 3820 19232 3850
rect 18200 3810 18466 3815
rect 17380 3786 17436 3792
rect 16611 3754 17352 3764
rect 16550 3751 16557 3754
rect 16609 3751 17352 3754
rect 16550 3739 17352 3751
rect 16550 3730 16557 3739
rect 16609 3736 17352 3739
rect 16609 3730 16616 3736
rect 16550 3674 16555 3730
rect 16611 3674 16616 3730
rect 17380 3734 17382 3786
rect 17434 3734 17436 3786
rect 18200 3764 18205 3810
rect 17464 3754 18205 3764
rect 18261 3754 18405 3810
rect 18461 3764 18466 3810
rect 18494 3798 19232 3820
rect 19284 3820 19286 3850
rect 19314 3848 20055 3876
rect 20050 3834 20055 3848
rect 20111 3834 20116 3890
rect 19284 3798 20022 3820
rect 18494 3792 20022 3798
rect 20050 3815 20057 3834
rect 20109 3815 20116 3834
rect 20050 3810 20116 3815
rect 19230 3786 19286 3792
rect 18461 3754 19202 3764
rect 17464 3751 18207 3754
rect 18259 3751 18407 3754
rect 18459 3751 19202 3754
rect 17464 3739 19202 3751
rect 17464 3736 18207 3739
rect 17380 3722 17436 3734
rect 17380 3708 17382 3722
rect 16644 3680 17382 3708
rect 16550 3650 16557 3674
rect 16609 3652 16616 3674
rect 17380 3670 17382 3680
rect 17434 3708 17436 3722
rect 18200 3730 18207 3736
rect 18259 3730 18407 3739
rect 18459 3736 19202 3739
rect 18459 3730 18466 3736
rect 17434 3680 18172 3708
rect 17434 3670 17436 3680
rect 17380 3658 17436 3670
rect 16609 3650 17352 3652
rect 16550 3594 16555 3650
rect 16611 3624 17352 3650
rect 16611 3594 16616 3624
rect 17380 3606 17382 3658
rect 17434 3606 17436 3658
rect 18200 3674 18205 3730
rect 18261 3674 18405 3730
rect 18461 3674 18466 3730
rect 19230 3734 19232 3786
rect 19284 3734 19286 3786
rect 20050 3764 20055 3810
rect 19314 3754 20055 3764
rect 20111 3754 20116 3810
rect 19314 3751 20057 3754
rect 20109 3751 20116 3754
rect 19314 3739 20116 3751
rect 19314 3736 20057 3739
rect 19230 3722 19286 3734
rect 19230 3708 19232 3722
rect 18494 3680 19232 3708
rect 18200 3652 18207 3674
rect 17464 3650 18207 3652
rect 18259 3650 18407 3674
rect 18459 3652 18466 3674
rect 19230 3670 19232 3680
rect 19284 3708 19286 3722
rect 20050 3730 20057 3736
rect 20109 3730 20116 3739
rect 19284 3680 20022 3708
rect 19284 3670 19286 3680
rect 19230 3658 19286 3670
rect 18459 3650 19202 3652
rect 17464 3624 18205 3650
rect 17380 3596 17436 3606
rect 16550 3570 16557 3594
rect 16609 3570 16616 3594
rect 16550 3514 16555 3570
rect 16611 3540 16616 3570
rect 16644 3594 18172 3596
rect 16644 3568 17382 3594
rect 17380 3542 17382 3568
rect 17434 3568 18172 3594
rect 18200 3594 18205 3624
rect 18261 3594 18405 3650
rect 18461 3624 19202 3650
rect 18461 3594 18466 3624
rect 19230 3606 19232 3658
rect 19284 3606 19286 3658
rect 20050 3674 20055 3730
rect 20111 3674 20116 3730
rect 20050 3652 20057 3674
rect 19314 3650 20057 3652
rect 20109 3650 20116 3674
rect 19314 3624 20055 3650
rect 19230 3596 19286 3606
rect 18200 3570 18207 3594
rect 18259 3570 18407 3594
rect 18459 3570 18466 3594
rect 17434 3542 17436 3568
rect 16611 3514 17352 3540
rect 16550 3495 16557 3514
rect 16609 3512 17352 3514
rect 17380 3530 17436 3542
rect 18200 3540 18205 3570
rect 16609 3495 16616 3512
rect 16550 3490 16616 3495
rect 16550 3434 16555 3490
rect 16611 3434 16616 3490
rect 17380 3484 17382 3530
rect 16644 3478 17382 3484
rect 17434 3484 17436 3530
rect 17464 3514 18205 3540
rect 18261 3514 18405 3570
rect 18461 3540 18466 3570
rect 18494 3594 20022 3596
rect 18494 3568 19232 3594
rect 19230 3542 19232 3568
rect 19284 3568 20022 3594
rect 20050 3594 20055 3624
rect 20111 3594 20116 3650
rect 20050 3570 20057 3594
rect 20109 3570 20116 3594
rect 19284 3542 19286 3568
rect 18461 3514 19202 3540
rect 17464 3512 18207 3514
rect 18200 3495 18207 3512
rect 18259 3495 18407 3514
rect 18459 3512 19202 3514
rect 19230 3530 19286 3542
rect 20050 3540 20055 3570
rect 18459 3495 18466 3512
rect 18200 3490 18466 3495
rect 17434 3478 18172 3484
rect 16644 3466 18172 3478
rect 16644 3456 17382 3466
rect 16550 3431 16557 3434
rect 16609 3431 16616 3434
rect 16550 3428 16616 3431
rect 16550 3419 17352 3428
rect 16550 3410 16557 3419
rect 16609 3410 17352 3419
rect 16550 3354 16555 3410
rect 16611 3400 17352 3410
rect 17380 3414 17382 3456
rect 17434 3456 18172 3466
rect 17434 3414 17436 3456
rect 18200 3434 18205 3490
rect 18261 3434 18405 3490
rect 18461 3434 18466 3490
rect 19230 3484 19232 3530
rect 18494 3478 19232 3484
rect 19284 3484 19286 3530
rect 19314 3514 20055 3540
rect 20111 3514 20116 3570
rect 19314 3512 20057 3514
rect 20050 3495 20057 3512
rect 20109 3495 20116 3514
rect 20050 3490 20116 3495
rect 19284 3478 20022 3484
rect 18494 3466 20022 3478
rect 18494 3456 19232 3466
rect 18200 3431 18207 3434
rect 18259 3431 18407 3434
rect 18459 3431 18466 3434
rect 18200 3428 18466 3431
rect 17380 3402 17436 3414
rect 16611 3354 16616 3400
rect 17380 3372 17382 3402
rect 16550 3303 16557 3354
rect 16609 3316 16616 3354
rect 16644 3350 17382 3372
rect 17434 3372 17436 3402
rect 17464 3419 19202 3428
rect 17464 3410 18207 3419
rect 18259 3410 18407 3419
rect 18459 3410 19202 3419
rect 17464 3400 18205 3410
rect 17434 3350 18172 3372
rect 16644 3344 18172 3350
rect 18200 3354 18205 3400
rect 18261 3354 18405 3410
rect 18461 3400 19202 3410
rect 19230 3414 19232 3456
rect 19284 3456 20022 3466
rect 19284 3414 19286 3456
rect 20050 3434 20055 3490
rect 20111 3434 20116 3490
rect 20050 3431 20057 3434
rect 20109 3431 20116 3434
rect 20050 3428 20116 3431
rect 19230 3402 19286 3414
rect 18461 3354 18466 3400
rect 19230 3372 19232 3402
rect 16609 3311 17353 3316
rect 16609 3309 16648 3311
rect 16704 3309 16728 3311
rect 16784 3309 16808 3311
rect 16864 3309 16888 3311
rect 16944 3309 16968 3311
rect 17024 3309 17048 3311
rect 17104 3309 17128 3311
rect 17184 3309 17208 3311
rect 17264 3309 17288 3311
rect 16609 3303 16638 3309
rect 16550 3257 16638 3303
rect 16882 3257 16888 3309
rect 16946 3257 16958 3309
rect 17202 3257 17208 3309
rect 17266 3257 17278 3309
rect 16550 3255 16648 3257
rect 16704 3255 16728 3257
rect 16784 3255 16808 3257
rect 16864 3255 16888 3257
rect 16944 3255 16968 3257
rect 17024 3255 17048 3257
rect 17104 3255 17128 3257
rect 17184 3255 17208 3257
rect 17264 3255 17288 3257
rect 17344 3255 17353 3311
rect 16550 3250 17353 3255
rect 17381 3250 17435 3344
rect 18200 3316 18207 3354
rect 17463 3311 18207 3316
rect 17463 3255 17472 3311
rect 17528 3309 17552 3311
rect 17608 3309 17632 3311
rect 17688 3309 17712 3311
rect 17768 3309 17792 3311
rect 17848 3309 17872 3311
rect 17928 3309 17952 3311
rect 18008 3309 18032 3311
rect 18088 3309 18112 3311
rect 18168 3309 18207 3311
rect 17544 3257 17552 3309
rect 17608 3257 17620 3309
rect 17864 3257 17872 3309
rect 17928 3257 17940 3309
rect 18184 3303 18207 3309
rect 18259 3303 18407 3354
rect 18459 3316 18466 3354
rect 18494 3350 19232 3372
rect 19284 3372 19286 3402
rect 19314 3419 20116 3428
rect 19314 3410 20057 3419
rect 20109 3410 20116 3419
rect 19314 3400 20055 3410
rect 19284 3350 20022 3372
rect 18494 3344 20022 3350
rect 20050 3354 20055 3400
rect 20111 3354 20116 3410
rect 18459 3311 19203 3316
rect 18459 3309 18498 3311
rect 18554 3309 18578 3311
rect 18634 3309 18658 3311
rect 18714 3309 18738 3311
rect 18794 3309 18818 3311
rect 18874 3309 18898 3311
rect 18954 3309 18978 3311
rect 19034 3309 19058 3311
rect 19114 3309 19138 3311
rect 18459 3303 18488 3309
rect 18184 3257 18488 3303
rect 18732 3257 18738 3309
rect 18796 3257 18808 3309
rect 19052 3257 19058 3309
rect 19116 3257 19128 3309
rect 17528 3255 17552 3257
rect 17608 3255 17632 3257
rect 17688 3255 17712 3257
rect 17768 3255 17792 3257
rect 17848 3255 17872 3257
rect 17928 3255 17952 3257
rect 18008 3255 18032 3257
rect 18088 3255 18112 3257
rect 18168 3255 18498 3257
rect 18554 3255 18578 3257
rect 18634 3255 18658 3257
rect 18714 3255 18738 3257
rect 18794 3255 18818 3257
rect 18874 3255 18898 3257
rect 18954 3255 18978 3257
rect 19034 3255 19058 3257
rect 19114 3255 19138 3257
rect 19194 3255 19203 3311
rect 17463 3250 19203 3255
rect 19231 3250 19285 3344
rect 20050 3316 20057 3354
rect 19313 3311 20057 3316
rect 19313 3255 19322 3311
rect 19378 3309 19402 3311
rect 19458 3309 19482 3311
rect 19538 3309 19562 3311
rect 19618 3309 19642 3311
rect 19698 3309 19722 3311
rect 19778 3309 19802 3311
rect 19858 3309 19882 3311
rect 19938 3309 19962 3311
rect 20018 3309 20057 3311
rect 19394 3257 19402 3309
rect 19458 3257 19470 3309
rect 19714 3257 19722 3309
rect 19778 3257 19790 3309
rect 20034 3303 20057 3309
rect 20109 3303 20116 3354
rect 20034 3257 20116 3303
rect 19378 3255 19402 3257
rect 19458 3255 19482 3257
rect 19538 3255 19562 3257
rect 19618 3255 19642 3257
rect 19698 3255 19722 3257
rect 19778 3255 19802 3257
rect 19858 3255 19882 3257
rect 19938 3255 19962 3257
rect 20018 3255 20116 3257
rect 19313 3250 20116 3255
<< via2 >>
rect 16648 9861 16704 9863
rect 16728 9861 16784 9863
rect 16808 9861 16864 9863
rect 16888 9861 16944 9863
rect 16968 9861 17024 9863
rect 17048 9861 17104 9863
rect 17128 9861 17184 9863
rect 17208 9861 17264 9863
rect 17288 9861 17344 9863
rect 16648 9809 16690 9861
rect 16690 9809 16702 9861
rect 16702 9809 16704 9861
rect 16728 9809 16754 9861
rect 16754 9809 16766 9861
rect 16766 9809 16784 9861
rect 16808 9809 16818 9861
rect 16818 9809 16830 9861
rect 16830 9809 16864 9861
rect 16888 9809 16894 9861
rect 16894 9809 16944 9861
rect 16968 9809 17010 9861
rect 17010 9809 17022 9861
rect 17022 9809 17024 9861
rect 17048 9809 17074 9861
rect 17074 9809 17086 9861
rect 17086 9809 17104 9861
rect 17128 9809 17138 9861
rect 17138 9809 17150 9861
rect 17150 9809 17184 9861
rect 17208 9809 17214 9861
rect 17214 9809 17264 9861
rect 17288 9809 17330 9861
rect 17330 9809 17344 9861
rect 16648 9807 16704 9809
rect 16728 9807 16784 9809
rect 16808 9807 16864 9809
rect 16888 9807 16944 9809
rect 16968 9807 17024 9809
rect 17048 9807 17104 9809
rect 17128 9807 17184 9809
rect 17208 9807 17264 9809
rect 17288 9807 17344 9809
rect 17472 9861 17528 9863
rect 17552 9861 17608 9863
rect 17632 9861 17688 9863
rect 17712 9861 17768 9863
rect 17792 9861 17848 9863
rect 17872 9861 17928 9863
rect 17952 9861 18008 9863
rect 18032 9861 18088 9863
rect 18112 9861 18168 9863
rect 17472 9809 17492 9861
rect 17492 9809 17528 9861
rect 17552 9809 17556 9861
rect 17556 9809 17608 9861
rect 17632 9809 17672 9861
rect 17672 9809 17684 9861
rect 17684 9809 17688 9861
rect 17712 9809 17736 9861
rect 17736 9809 17748 9861
rect 17748 9809 17768 9861
rect 17792 9809 17800 9861
rect 17800 9809 17812 9861
rect 17812 9809 17848 9861
rect 17872 9809 17876 9861
rect 17876 9809 17928 9861
rect 17952 9809 17992 9861
rect 17992 9809 18004 9861
rect 18004 9809 18008 9861
rect 18032 9809 18056 9861
rect 18056 9809 18068 9861
rect 18068 9809 18088 9861
rect 18112 9809 18120 9861
rect 18120 9809 18132 9861
rect 18132 9809 18168 9861
rect 18498 9861 18554 9863
rect 18578 9861 18634 9863
rect 18658 9861 18714 9863
rect 18738 9861 18794 9863
rect 18818 9861 18874 9863
rect 18898 9861 18954 9863
rect 18978 9861 19034 9863
rect 19058 9861 19114 9863
rect 19138 9861 19194 9863
rect 17472 9807 17528 9809
rect 17552 9807 17608 9809
rect 17632 9807 17688 9809
rect 17712 9807 17768 9809
rect 17792 9807 17848 9809
rect 17872 9807 17928 9809
rect 17952 9807 18008 9809
rect 18032 9807 18088 9809
rect 18112 9807 18168 9809
rect 16555 9763 16557 9764
rect 16557 9763 16609 9764
rect 16609 9763 16611 9764
rect 16555 9751 16611 9763
rect 16555 9708 16557 9751
rect 16557 9708 16609 9751
rect 16609 9708 16611 9751
rect 18498 9809 18540 9861
rect 18540 9809 18552 9861
rect 18552 9809 18554 9861
rect 18578 9809 18604 9861
rect 18604 9809 18616 9861
rect 18616 9809 18634 9861
rect 18658 9809 18668 9861
rect 18668 9809 18680 9861
rect 18680 9809 18714 9861
rect 18738 9809 18744 9861
rect 18744 9809 18794 9861
rect 18818 9809 18860 9861
rect 18860 9809 18872 9861
rect 18872 9809 18874 9861
rect 18898 9809 18924 9861
rect 18924 9809 18936 9861
rect 18936 9809 18954 9861
rect 18978 9809 18988 9861
rect 18988 9809 19000 9861
rect 19000 9809 19034 9861
rect 19058 9809 19064 9861
rect 19064 9809 19114 9861
rect 19138 9809 19180 9861
rect 19180 9809 19194 9861
rect 18498 9807 18554 9809
rect 18578 9807 18634 9809
rect 18658 9807 18714 9809
rect 18738 9807 18794 9809
rect 18818 9807 18874 9809
rect 18898 9807 18954 9809
rect 18978 9807 19034 9809
rect 19058 9807 19114 9809
rect 19138 9807 19194 9809
rect 19322 9861 19378 9863
rect 19402 9861 19458 9863
rect 19482 9861 19538 9863
rect 19562 9861 19618 9863
rect 19642 9861 19698 9863
rect 19722 9861 19778 9863
rect 19802 9861 19858 9863
rect 19882 9861 19938 9863
rect 19962 9861 20018 9863
rect 19322 9809 19342 9861
rect 19342 9809 19378 9861
rect 19402 9809 19406 9861
rect 19406 9809 19458 9861
rect 19482 9809 19522 9861
rect 19522 9809 19534 9861
rect 19534 9809 19538 9861
rect 19562 9809 19586 9861
rect 19586 9809 19598 9861
rect 19598 9809 19618 9861
rect 19642 9809 19650 9861
rect 19650 9809 19662 9861
rect 19662 9809 19698 9861
rect 19722 9809 19726 9861
rect 19726 9809 19778 9861
rect 19802 9809 19842 9861
rect 19842 9809 19854 9861
rect 19854 9809 19858 9861
rect 19882 9809 19906 9861
rect 19906 9809 19918 9861
rect 19918 9809 19938 9861
rect 19962 9809 19970 9861
rect 19970 9809 19982 9861
rect 19982 9809 20018 9861
rect 19322 9807 19378 9809
rect 19402 9807 19458 9809
rect 19482 9807 19538 9809
rect 19562 9807 19618 9809
rect 19642 9807 19698 9809
rect 19722 9807 19778 9809
rect 19802 9807 19858 9809
rect 19882 9807 19938 9809
rect 19962 9807 20018 9809
rect 18205 9763 18207 9764
rect 18207 9763 18259 9764
rect 18259 9763 18261 9764
rect 18205 9751 18261 9763
rect 16555 9635 16557 9684
rect 16557 9635 16609 9684
rect 16609 9635 16611 9684
rect 16555 9628 16611 9635
rect 18205 9708 18207 9751
rect 18207 9708 18259 9751
rect 18259 9708 18261 9751
rect 18405 9763 18407 9764
rect 18407 9763 18459 9764
rect 18459 9763 18461 9764
rect 18405 9751 18461 9763
rect 18405 9708 18407 9751
rect 18407 9708 18459 9751
rect 18459 9708 18461 9751
rect 20055 9763 20057 9764
rect 20057 9763 20109 9764
rect 20109 9763 20111 9764
rect 20055 9751 20111 9763
rect 16555 9571 16557 9604
rect 16557 9571 16609 9604
rect 16609 9571 16611 9604
rect 18205 9635 18207 9684
rect 18207 9635 18259 9684
rect 18259 9635 18261 9684
rect 18205 9628 18261 9635
rect 18405 9635 18407 9684
rect 18407 9635 18459 9684
rect 18459 9635 18461 9684
rect 18405 9628 18461 9635
rect 20055 9708 20057 9751
rect 20057 9708 20109 9751
rect 20109 9708 20111 9751
rect 16555 9559 16611 9571
rect 16555 9548 16557 9559
rect 16557 9548 16609 9559
rect 16609 9548 16611 9559
rect 16555 9507 16557 9524
rect 16557 9507 16609 9524
rect 16609 9507 16611 9524
rect 16555 9495 16611 9507
rect 16555 9468 16557 9495
rect 16557 9468 16609 9495
rect 16609 9468 16611 9495
rect 18205 9571 18207 9604
rect 18207 9571 18259 9604
rect 18259 9571 18261 9604
rect 18205 9559 18261 9571
rect 18205 9548 18207 9559
rect 18207 9548 18259 9559
rect 18259 9548 18261 9559
rect 18405 9571 18407 9604
rect 18407 9571 18459 9604
rect 18459 9571 18461 9604
rect 20055 9635 20057 9684
rect 20057 9635 20109 9684
rect 20109 9635 20111 9684
rect 20055 9628 20111 9635
rect 18405 9559 18461 9571
rect 18405 9548 18407 9559
rect 18407 9548 18459 9559
rect 18459 9548 18461 9559
rect 16555 9443 16557 9444
rect 16557 9443 16609 9444
rect 16609 9443 16611 9444
rect 16555 9431 16611 9443
rect 16555 9388 16557 9431
rect 16557 9388 16609 9431
rect 16609 9388 16611 9431
rect 18205 9507 18207 9524
rect 18207 9507 18259 9524
rect 18259 9507 18261 9524
rect 18205 9495 18261 9507
rect 18205 9468 18207 9495
rect 18207 9468 18259 9495
rect 18259 9468 18261 9495
rect 18405 9507 18407 9524
rect 18407 9507 18459 9524
rect 18459 9507 18461 9524
rect 18405 9495 18461 9507
rect 18405 9468 18407 9495
rect 18407 9468 18459 9495
rect 18459 9468 18461 9495
rect 20055 9571 20057 9604
rect 20057 9571 20109 9604
rect 20109 9571 20111 9604
rect 20055 9559 20111 9571
rect 20055 9548 20057 9559
rect 20057 9548 20109 9559
rect 20109 9548 20111 9559
rect 16555 9315 16557 9364
rect 16557 9315 16609 9364
rect 16609 9315 16611 9364
rect 16555 9308 16611 9315
rect 18205 9443 18207 9444
rect 18207 9443 18259 9444
rect 18259 9443 18261 9444
rect 18205 9431 18261 9443
rect 18205 9388 18207 9431
rect 18207 9388 18259 9431
rect 18259 9388 18261 9431
rect 18405 9443 18407 9444
rect 18407 9443 18459 9444
rect 18459 9443 18461 9444
rect 18405 9431 18461 9443
rect 18405 9388 18407 9431
rect 18407 9388 18459 9431
rect 18459 9388 18461 9431
rect 20055 9507 20057 9524
rect 20057 9507 20109 9524
rect 20109 9507 20111 9524
rect 20055 9495 20111 9507
rect 20055 9468 20057 9495
rect 20057 9468 20109 9495
rect 20109 9468 20111 9495
rect 16555 9251 16557 9284
rect 16557 9251 16609 9284
rect 16609 9251 16611 9284
rect 16555 9239 16611 9251
rect 18205 9315 18207 9364
rect 18207 9315 18259 9364
rect 18259 9315 18261 9364
rect 18205 9308 18261 9315
rect 18405 9315 18407 9364
rect 18407 9315 18459 9364
rect 18459 9315 18461 9364
rect 18405 9308 18461 9315
rect 20055 9443 20057 9444
rect 20057 9443 20109 9444
rect 20109 9443 20111 9444
rect 20055 9431 20111 9443
rect 20055 9388 20057 9431
rect 20057 9388 20109 9431
rect 20109 9388 20111 9431
rect 16555 9228 16557 9239
rect 16557 9228 16609 9239
rect 16609 9228 16611 9239
rect 16555 9187 16557 9204
rect 16557 9187 16609 9204
rect 16609 9187 16611 9204
rect 16555 9148 16611 9187
rect 18205 9251 18207 9284
rect 18207 9251 18259 9284
rect 18259 9251 18261 9284
rect 18205 9239 18261 9251
rect 18205 9228 18207 9239
rect 18207 9228 18259 9239
rect 18259 9228 18261 9239
rect 18405 9251 18407 9284
rect 18407 9251 18459 9284
rect 18459 9251 18461 9284
rect 18405 9239 18461 9251
rect 20055 9315 20057 9364
rect 20057 9315 20109 9364
rect 20109 9315 20111 9364
rect 20055 9308 20111 9315
rect 18405 9228 18407 9239
rect 18407 9228 18459 9239
rect 18459 9228 18461 9239
rect 18205 9187 18207 9204
rect 18207 9187 18259 9204
rect 18259 9187 18261 9204
rect 18205 9148 18261 9187
rect 18405 9187 18407 9204
rect 18407 9187 18459 9204
rect 18459 9187 18461 9204
rect 18405 9148 18461 9187
rect 20055 9251 20057 9284
rect 20057 9251 20109 9284
rect 20109 9251 20111 9284
rect 20055 9239 20111 9251
rect 20055 9228 20057 9239
rect 20057 9228 20109 9239
rect 20109 9228 20111 9239
rect 20055 9187 20057 9204
rect 20057 9187 20109 9204
rect 20109 9187 20111 9204
rect 20055 9148 20111 9187
rect 16740 9110 16796 9112
rect 16820 9110 16876 9112
rect 16900 9110 16956 9112
rect 16980 9110 17036 9112
rect 17060 9110 17116 9112
rect 17140 9110 17196 9112
rect 17220 9110 17276 9112
rect 17300 9110 17356 9112
rect 16740 9058 16771 9110
rect 16771 9058 16783 9110
rect 16783 9058 16796 9110
rect 16820 9058 16835 9110
rect 16835 9058 16847 9110
rect 16847 9058 16876 9110
rect 16900 9058 16911 9110
rect 16911 9058 16956 9110
rect 16980 9058 17027 9110
rect 17027 9058 17036 9110
rect 17060 9058 17091 9110
rect 17091 9058 17103 9110
rect 17103 9058 17116 9110
rect 17140 9058 17155 9110
rect 17155 9058 17167 9110
rect 17167 9058 17196 9110
rect 17220 9058 17231 9110
rect 17231 9058 17276 9110
rect 17300 9058 17347 9110
rect 17347 9058 17356 9110
rect 16740 9056 16796 9058
rect 16820 9056 16876 9058
rect 16900 9056 16956 9058
rect 16980 9056 17036 9058
rect 17060 9056 17116 9058
rect 17140 9056 17196 9058
rect 17220 9056 17276 9058
rect 17300 9056 17356 9058
rect 17380 9056 17436 9112
rect 17460 9110 17516 9112
rect 17540 9110 17596 9112
rect 17620 9110 17676 9112
rect 17700 9110 17756 9112
rect 17780 9110 17836 9112
rect 17860 9110 17916 9112
rect 17940 9110 17996 9112
rect 18020 9110 18076 9112
rect 18590 9110 18646 9112
rect 18670 9110 18726 9112
rect 18750 9110 18806 9112
rect 18830 9110 18886 9112
rect 18910 9110 18966 9112
rect 18990 9110 19046 9112
rect 19070 9110 19126 9112
rect 19150 9110 19206 9112
rect 17460 9058 17469 9110
rect 17469 9058 17516 9110
rect 17540 9058 17585 9110
rect 17585 9058 17596 9110
rect 17620 9058 17649 9110
rect 17649 9058 17661 9110
rect 17661 9058 17676 9110
rect 17700 9058 17713 9110
rect 17713 9058 17725 9110
rect 17725 9058 17756 9110
rect 17780 9058 17789 9110
rect 17789 9058 17836 9110
rect 17860 9058 17905 9110
rect 17905 9058 17916 9110
rect 17940 9058 17969 9110
rect 17969 9058 17981 9110
rect 17981 9058 17996 9110
rect 18020 9058 18033 9110
rect 18033 9058 18045 9110
rect 18045 9058 18076 9110
rect 18590 9058 18621 9110
rect 18621 9058 18633 9110
rect 18633 9058 18646 9110
rect 18670 9058 18685 9110
rect 18685 9058 18697 9110
rect 18697 9058 18726 9110
rect 18750 9058 18761 9110
rect 18761 9058 18806 9110
rect 18830 9058 18877 9110
rect 18877 9058 18886 9110
rect 18910 9058 18941 9110
rect 18941 9058 18953 9110
rect 18953 9058 18966 9110
rect 18990 9058 19005 9110
rect 19005 9058 19017 9110
rect 19017 9058 19046 9110
rect 19070 9058 19081 9110
rect 19081 9058 19126 9110
rect 19150 9058 19197 9110
rect 19197 9058 19206 9110
rect 17460 9056 17516 9058
rect 17540 9056 17596 9058
rect 17620 9056 17676 9058
rect 17700 9056 17756 9058
rect 17780 9056 17836 9058
rect 17860 9056 17916 9058
rect 17940 9056 17996 9058
rect 18020 9056 18076 9058
rect 16555 8981 16611 9020
rect 16555 8964 16557 8981
rect 16557 8964 16609 8981
rect 16609 8964 16611 8981
rect 16555 8929 16557 8940
rect 16557 8929 16609 8940
rect 16609 8929 16611 8940
rect 16555 8917 16611 8929
rect 16555 8884 16557 8917
rect 16557 8884 16609 8917
rect 16609 8884 16611 8917
rect 18205 8981 18261 9020
rect 18205 8964 18207 8981
rect 18207 8964 18259 8981
rect 18259 8964 18261 8981
rect 18205 8929 18207 8940
rect 18207 8929 18259 8940
rect 18259 8929 18261 8940
rect 16555 8853 16611 8860
rect 16555 8804 16557 8853
rect 16557 8804 16609 8853
rect 16609 8804 16611 8853
rect 18205 8917 18261 8929
rect 18205 8884 18207 8917
rect 18207 8884 18259 8917
rect 18259 8884 18261 8917
rect 16555 8737 16557 8780
rect 16557 8737 16609 8780
rect 16609 8737 16611 8780
rect 16555 8725 16611 8737
rect 16555 8724 16557 8725
rect 16557 8724 16609 8725
rect 16609 8724 16611 8725
rect 18205 8853 18261 8860
rect 18205 8804 18207 8853
rect 18207 8804 18259 8853
rect 18259 8804 18261 8853
rect 16555 8673 16557 8700
rect 16557 8673 16609 8700
rect 16609 8673 16611 8700
rect 16555 8661 16611 8673
rect 16555 8644 16557 8661
rect 16557 8644 16609 8661
rect 16609 8644 16611 8661
rect 18205 8737 18207 8780
rect 18207 8737 18259 8780
rect 18259 8737 18261 8780
rect 18205 8725 18261 8737
rect 18205 8724 18207 8725
rect 18207 8724 18259 8725
rect 18259 8724 18261 8725
rect 16555 8609 16557 8620
rect 16557 8609 16609 8620
rect 16609 8609 16611 8620
rect 16555 8597 16611 8609
rect 16555 8564 16557 8597
rect 16557 8564 16609 8597
rect 16609 8564 16611 8597
rect 18205 8673 18207 8700
rect 18207 8673 18259 8700
rect 18259 8673 18261 8700
rect 18205 8661 18261 8673
rect 18205 8644 18207 8661
rect 18207 8644 18259 8661
rect 18259 8644 18261 8661
rect 18205 8609 18207 8620
rect 18207 8609 18259 8620
rect 18259 8609 18261 8620
rect 18205 8597 18261 8609
rect 16555 8533 16611 8540
rect 16555 8484 16557 8533
rect 16557 8484 16609 8533
rect 16609 8484 16611 8533
rect 18205 8564 18207 8597
rect 18207 8564 18259 8597
rect 18259 8564 18261 8597
rect 16555 8417 16557 8460
rect 16557 8417 16609 8460
rect 16609 8417 16611 8460
rect 18205 8533 18261 8540
rect 18205 8484 18207 8533
rect 18207 8484 18259 8533
rect 18259 8484 18261 8533
rect 16555 8405 16611 8417
rect 16555 8404 16557 8405
rect 16557 8404 16609 8405
rect 16609 8404 16611 8405
rect 18205 8417 18207 8460
rect 18207 8417 18259 8460
rect 18259 8417 18261 8460
rect 18205 8405 18261 8417
rect 18205 8404 18207 8405
rect 18207 8404 18259 8405
rect 18259 8404 18261 8405
rect 16648 8359 16704 8361
rect 16728 8359 16784 8361
rect 16808 8359 16864 8361
rect 16888 8359 16944 8361
rect 16968 8359 17024 8361
rect 17048 8359 17104 8361
rect 17128 8359 17184 8361
rect 17208 8359 17264 8361
rect 17288 8359 17344 8361
rect 16648 8307 16690 8359
rect 16690 8307 16702 8359
rect 16702 8307 16704 8359
rect 16728 8307 16754 8359
rect 16754 8307 16766 8359
rect 16766 8307 16784 8359
rect 16808 8307 16818 8359
rect 16818 8307 16830 8359
rect 16830 8307 16864 8359
rect 16888 8307 16894 8359
rect 16894 8307 16944 8359
rect 16968 8307 17010 8359
rect 17010 8307 17022 8359
rect 17022 8307 17024 8359
rect 17048 8307 17074 8359
rect 17074 8307 17086 8359
rect 17086 8307 17104 8359
rect 17128 8307 17138 8359
rect 17138 8307 17150 8359
rect 17150 8307 17184 8359
rect 17208 8307 17214 8359
rect 17214 8307 17264 8359
rect 17288 8307 17330 8359
rect 17330 8307 17344 8359
rect 16648 8305 16704 8307
rect 16728 8305 16784 8307
rect 16808 8305 16864 8307
rect 16888 8305 16944 8307
rect 16968 8305 17024 8307
rect 17048 8305 17104 8307
rect 17128 8305 17184 8307
rect 17208 8305 17264 8307
rect 17288 8305 17344 8307
rect 17472 8359 17528 8361
rect 17552 8359 17608 8361
rect 17632 8359 17688 8361
rect 17712 8359 17768 8361
rect 17792 8359 17848 8361
rect 17872 8359 17928 8361
rect 17952 8359 18008 8361
rect 18032 8359 18088 8361
rect 18112 8359 18168 8361
rect 17472 8307 17492 8359
rect 17492 8307 17528 8359
rect 17552 8307 17556 8359
rect 17556 8307 17608 8359
rect 17632 8307 17672 8359
rect 17672 8307 17684 8359
rect 17684 8307 17688 8359
rect 17712 8307 17736 8359
rect 17736 8307 17748 8359
rect 17748 8307 17768 8359
rect 17792 8307 17800 8359
rect 17800 8307 17812 8359
rect 17812 8307 17848 8359
rect 17872 8307 17876 8359
rect 17876 8307 17928 8359
rect 17952 8307 17992 8359
rect 17992 8307 18004 8359
rect 18004 8307 18008 8359
rect 18032 8307 18056 8359
rect 18056 8307 18068 8359
rect 18068 8307 18088 8359
rect 18112 8307 18120 8359
rect 18120 8307 18132 8359
rect 18132 8307 18168 8359
rect 17472 8305 17528 8307
rect 17552 8305 17608 8307
rect 17632 8305 17688 8307
rect 17712 8305 17768 8307
rect 17792 8305 17848 8307
rect 17872 8305 17928 8307
rect 17952 8305 18008 8307
rect 18032 8305 18088 8307
rect 18112 8305 18168 8307
rect 18590 9056 18646 9058
rect 18670 9056 18726 9058
rect 18750 9056 18806 9058
rect 18830 9056 18886 9058
rect 18910 9056 18966 9058
rect 18990 9056 19046 9058
rect 19070 9056 19126 9058
rect 19150 9056 19206 9058
rect 19230 9056 19286 9112
rect 19310 9110 19366 9112
rect 19390 9110 19446 9112
rect 19470 9110 19526 9112
rect 19550 9110 19606 9112
rect 19630 9110 19686 9112
rect 19710 9110 19766 9112
rect 19790 9110 19846 9112
rect 19870 9110 19926 9112
rect 19310 9058 19319 9110
rect 19319 9058 19366 9110
rect 19390 9058 19435 9110
rect 19435 9058 19446 9110
rect 19470 9058 19499 9110
rect 19499 9058 19511 9110
rect 19511 9058 19526 9110
rect 19550 9058 19563 9110
rect 19563 9058 19575 9110
rect 19575 9058 19606 9110
rect 19630 9058 19639 9110
rect 19639 9058 19686 9110
rect 19710 9058 19755 9110
rect 19755 9058 19766 9110
rect 19790 9058 19819 9110
rect 19819 9058 19831 9110
rect 19831 9058 19846 9110
rect 19870 9058 19883 9110
rect 19883 9058 19895 9110
rect 19895 9058 19926 9110
rect 19310 9056 19366 9058
rect 19390 9056 19446 9058
rect 19470 9056 19526 9058
rect 19550 9056 19606 9058
rect 19630 9056 19686 9058
rect 19710 9056 19766 9058
rect 19790 9056 19846 9058
rect 19870 9056 19926 9058
rect 18405 8981 18461 9020
rect 18405 8964 18407 8981
rect 18407 8964 18459 8981
rect 18459 8964 18461 8981
rect 18405 8929 18407 8940
rect 18407 8929 18459 8940
rect 18459 8929 18461 8940
rect 18405 8917 18461 8929
rect 18405 8884 18407 8917
rect 18407 8884 18459 8917
rect 18459 8884 18461 8917
rect 20055 8981 20111 9020
rect 20055 8964 20057 8981
rect 20057 8964 20109 8981
rect 20109 8964 20111 8981
rect 20055 8929 20057 8940
rect 20057 8929 20109 8940
rect 20109 8929 20111 8940
rect 18405 8853 18461 8860
rect 18405 8804 18407 8853
rect 18407 8804 18459 8853
rect 18459 8804 18461 8853
rect 20055 8917 20111 8929
rect 20055 8884 20057 8917
rect 20057 8884 20109 8917
rect 20109 8884 20111 8917
rect 18405 8737 18407 8780
rect 18407 8737 18459 8780
rect 18459 8737 18461 8780
rect 18405 8725 18461 8737
rect 18405 8724 18407 8725
rect 18407 8724 18459 8725
rect 18459 8724 18461 8725
rect 20055 8853 20111 8860
rect 20055 8804 20057 8853
rect 20057 8804 20109 8853
rect 20109 8804 20111 8853
rect 18405 8673 18407 8700
rect 18407 8673 18459 8700
rect 18459 8673 18461 8700
rect 18405 8661 18461 8673
rect 18405 8644 18407 8661
rect 18407 8644 18459 8661
rect 18459 8644 18461 8661
rect 20055 8737 20057 8780
rect 20057 8737 20109 8780
rect 20109 8737 20111 8780
rect 20055 8725 20111 8737
rect 20055 8724 20057 8725
rect 20057 8724 20109 8725
rect 20109 8724 20111 8725
rect 18405 8609 18407 8620
rect 18407 8609 18459 8620
rect 18459 8609 18461 8620
rect 18405 8597 18461 8609
rect 18405 8564 18407 8597
rect 18407 8564 18459 8597
rect 18459 8564 18461 8597
rect 20055 8673 20057 8700
rect 20057 8673 20109 8700
rect 20109 8673 20111 8700
rect 20055 8661 20111 8673
rect 20055 8644 20057 8661
rect 20057 8644 20109 8661
rect 20109 8644 20111 8661
rect 20055 8609 20057 8620
rect 20057 8609 20109 8620
rect 20109 8609 20111 8620
rect 20055 8597 20111 8609
rect 18405 8533 18461 8540
rect 18405 8484 18407 8533
rect 18407 8484 18459 8533
rect 18459 8484 18461 8533
rect 20055 8564 20057 8597
rect 20057 8564 20109 8597
rect 20109 8564 20111 8597
rect 18405 8417 18407 8460
rect 18407 8417 18459 8460
rect 18459 8417 18461 8460
rect 20055 8533 20111 8540
rect 20055 8484 20057 8533
rect 20057 8484 20109 8533
rect 20109 8484 20111 8533
rect 18405 8405 18461 8417
rect 18405 8404 18407 8405
rect 18407 8404 18459 8405
rect 18459 8404 18461 8405
rect 20055 8417 20057 8460
rect 20057 8417 20109 8460
rect 20109 8417 20111 8460
rect 20055 8405 20111 8417
rect 20055 8404 20057 8405
rect 20057 8404 20109 8405
rect 20109 8404 20111 8405
rect 18498 8359 18554 8361
rect 18578 8359 18634 8361
rect 18658 8359 18714 8361
rect 18738 8359 18794 8361
rect 18818 8359 18874 8361
rect 18898 8359 18954 8361
rect 18978 8359 19034 8361
rect 19058 8359 19114 8361
rect 19138 8359 19194 8361
rect 18498 8307 18540 8359
rect 18540 8307 18552 8359
rect 18552 8307 18554 8359
rect 18578 8307 18604 8359
rect 18604 8307 18616 8359
rect 18616 8307 18634 8359
rect 18658 8307 18668 8359
rect 18668 8307 18680 8359
rect 18680 8307 18714 8359
rect 18738 8307 18744 8359
rect 18744 8307 18794 8359
rect 18818 8307 18860 8359
rect 18860 8307 18872 8359
rect 18872 8307 18874 8359
rect 18898 8307 18924 8359
rect 18924 8307 18936 8359
rect 18936 8307 18954 8359
rect 18978 8307 18988 8359
rect 18988 8307 19000 8359
rect 19000 8307 19034 8359
rect 19058 8307 19064 8359
rect 19064 8307 19114 8359
rect 19138 8307 19180 8359
rect 19180 8307 19194 8359
rect 18498 8305 18554 8307
rect 18578 8305 18634 8307
rect 18658 8305 18714 8307
rect 18738 8305 18794 8307
rect 18818 8305 18874 8307
rect 18898 8305 18954 8307
rect 18978 8305 19034 8307
rect 19058 8305 19114 8307
rect 19138 8305 19194 8307
rect 19322 8359 19378 8361
rect 19402 8359 19458 8361
rect 19482 8359 19538 8361
rect 19562 8359 19618 8361
rect 19642 8359 19698 8361
rect 19722 8359 19778 8361
rect 19802 8359 19858 8361
rect 19882 8359 19938 8361
rect 19962 8359 20018 8361
rect 19322 8307 19342 8359
rect 19342 8307 19378 8359
rect 19402 8307 19406 8359
rect 19406 8307 19458 8359
rect 19482 8307 19522 8359
rect 19522 8307 19534 8359
rect 19534 8307 19538 8359
rect 19562 8307 19586 8359
rect 19586 8307 19598 8359
rect 19598 8307 19618 8359
rect 19642 8307 19650 8359
rect 19650 8307 19662 8359
rect 19662 8307 19698 8359
rect 19722 8307 19726 8359
rect 19726 8307 19778 8359
rect 19802 8307 19842 8359
rect 19842 8307 19854 8359
rect 19854 8307 19858 8359
rect 19882 8307 19906 8359
rect 19906 8307 19918 8359
rect 19918 8307 19938 8359
rect 19962 8307 19970 8359
rect 19970 8307 19982 8359
rect 19982 8307 20018 8359
rect 19322 8305 19378 8307
rect 19402 8305 19458 8307
rect 19482 8305 19538 8307
rect 19562 8305 19618 8307
rect 19642 8305 19698 8307
rect 19722 8305 19778 8307
rect 19802 8305 19858 8307
rect 19882 8305 19938 8307
rect 19962 8305 20018 8307
rect 11860 6990 12480 7050
rect 13000 6990 13220 7050
rect 13560 6990 13780 7050
rect 14140 6990 14320 7050
rect 14680 6970 15480 7050
rect 17697 7099 17753 7109
rect 17697 7053 17699 7099
rect 17699 7053 17751 7099
rect 17751 7053 17753 7099
rect 17180 6870 17330 6990
rect 17697 6983 17699 7029
rect 17699 6983 17751 7029
rect 17751 6983 17753 7029
rect 17697 6973 17753 6983
rect 17869 7099 17925 7109
rect 17869 7053 17871 7099
rect 17871 7053 17923 7099
rect 17923 7053 17925 7099
rect 17869 6983 17871 7029
rect 17871 6983 17923 7029
rect 17923 6983 17925 7029
rect 17869 6973 17925 6983
rect 18041 7099 18097 7109
rect 18041 7053 18043 7099
rect 18043 7053 18095 7099
rect 18095 7053 18097 7099
rect 18041 6983 18043 7029
rect 18043 6983 18095 7029
rect 18095 6983 18097 7029
rect 18041 6973 18097 6983
rect 18213 7099 18269 7109
rect 18213 7053 18215 7099
rect 18215 7053 18267 7099
rect 18267 7053 18269 7099
rect 18213 6983 18215 7029
rect 18215 6983 18267 7029
rect 18267 6983 18269 7029
rect 18213 6973 18269 6983
rect 18385 7099 18441 7109
rect 18385 7053 18387 7099
rect 18387 7053 18439 7099
rect 18439 7053 18441 7099
rect 18385 6983 18387 7029
rect 18387 6983 18439 7029
rect 18439 6983 18441 7029
rect 18385 6973 18441 6983
rect 18557 7099 18613 7109
rect 18557 7053 18559 7099
rect 18559 7053 18611 7099
rect 18611 7053 18613 7099
rect 18557 6983 18559 7029
rect 18559 6983 18611 7029
rect 18611 6983 18613 7029
rect 18557 6973 18613 6983
rect 18729 7099 18785 7109
rect 18729 7053 18731 7099
rect 18731 7053 18783 7099
rect 18783 7053 18785 7099
rect 18729 6983 18731 7029
rect 18731 6983 18783 7029
rect 18783 6983 18785 7029
rect 18729 6973 18785 6983
rect 18901 7099 18957 7109
rect 18901 7053 18903 7099
rect 18903 7053 18955 7099
rect 18955 7053 18957 7099
rect 18901 6983 18903 7029
rect 18903 6983 18955 7029
rect 18955 6983 18957 7029
rect 18901 6973 18957 6983
rect 19073 7099 19129 7109
rect 19073 7053 19075 7099
rect 19075 7053 19127 7099
rect 19127 7053 19129 7099
rect 19073 6983 19075 7029
rect 19075 6983 19127 7029
rect 19127 6983 19129 7029
rect 19073 6973 19129 6983
rect 19245 7099 19301 7109
rect 19245 7053 19247 7099
rect 19247 7053 19299 7099
rect 19299 7053 19301 7099
rect 19245 6983 19247 7029
rect 19247 6983 19299 7029
rect 19299 6983 19301 7029
rect 19245 6973 19301 6983
rect 19417 7099 19473 7109
rect 19417 7053 19419 7099
rect 19419 7053 19471 7099
rect 19471 7053 19473 7099
rect 19417 6983 19419 7029
rect 19419 6983 19471 7029
rect 19471 6983 19473 7029
rect 19417 6973 19473 6983
rect 19589 7099 19645 7109
rect 19589 7053 19591 7099
rect 19591 7053 19643 7099
rect 19643 7053 19645 7099
rect 19589 6983 19591 7029
rect 19591 6983 19643 7029
rect 19643 6983 19645 7029
rect 19589 6973 19645 6983
rect 19761 7099 19817 7109
rect 19761 7053 19763 7099
rect 19763 7053 19815 7099
rect 19815 7053 19817 7099
rect 19761 6983 19763 7029
rect 19763 6983 19815 7029
rect 19815 6983 19817 7029
rect 19761 6973 19817 6983
rect 19933 7099 19989 7109
rect 19933 7053 19935 7099
rect 19935 7053 19987 7099
rect 19987 7053 19989 7099
rect 19933 6983 19935 7029
rect 19935 6983 19987 7029
rect 19987 6983 19989 7029
rect 19933 6973 19989 6983
rect 17440 6720 17590 6820
rect 17180 6370 17330 6470
rect 17440 6230 17590 6330
rect 11620 5670 15680 5730
rect 12410 5570 12670 5580
rect 12410 5520 12420 5570
rect 12420 5520 12660 5570
rect 12660 5520 12670 5570
rect 12970 5570 13230 5580
rect 12970 5520 12980 5570
rect 12980 5520 13220 5570
rect 13220 5520 13230 5570
rect 13550 5570 13810 5580
rect 13550 5520 13560 5570
rect 13560 5520 13800 5570
rect 13800 5520 13810 5570
rect 14110 5570 14370 5580
rect 14110 5520 14120 5570
rect 14120 5520 14360 5570
rect 14360 5520 14370 5570
rect 14690 5570 14950 5580
rect 14690 5520 14700 5570
rect 14700 5520 14940 5570
rect 14940 5520 14950 5570
rect 11920 5380 12280 5420
rect 13220 5380 13580 5420
rect 14320 5380 14680 5420
rect 15540 5380 15690 5440
rect 15690 5380 15880 5440
rect 11920 5300 12280 5380
rect 13220 5300 13580 5380
rect 14320 5300 14680 5380
rect 15540 5300 15880 5380
rect 17679 6207 17735 6217
rect 17679 6161 17681 6207
rect 17681 6161 17733 6207
rect 17733 6161 17735 6207
rect 17679 6091 17681 6137
rect 17681 6091 17733 6137
rect 17733 6091 17735 6137
rect 17679 6081 17735 6091
rect 17851 6207 17907 6217
rect 17851 6161 17853 6207
rect 17853 6161 17905 6207
rect 17905 6161 17907 6207
rect 17851 6091 17853 6137
rect 17853 6091 17905 6137
rect 17905 6091 17907 6137
rect 17851 6081 17907 6091
rect 18023 6207 18079 6217
rect 18023 6161 18025 6207
rect 18025 6161 18077 6207
rect 18077 6161 18079 6207
rect 18023 6091 18025 6137
rect 18025 6091 18077 6137
rect 18077 6091 18079 6137
rect 18023 6081 18079 6091
rect 18195 6207 18251 6217
rect 18195 6161 18197 6207
rect 18197 6161 18249 6207
rect 18249 6161 18251 6207
rect 18195 6091 18197 6137
rect 18197 6091 18249 6137
rect 18249 6091 18251 6137
rect 18195 6081 18251 6091
rect 18367 6207 18423 6217
rect 18367 6161 18369 6207
rect 18369 6161 18421 6207
rect 18421 6161 18423 6207
rect 18367 6091 18369 6137
rect 18369 6091 18421 6137
rect 18421 6091 18423 6137
rect 18367 6081 18423 6091
rect 18539 6207 18595 6217
rect 18539 6161 18541 6207
rect 18541 6161 18593 6207
rect 18593 6161 18595 6207
rect 18539 6091 18541 6137
rect 18541 6091 18593 6137
rect 18593 6091 18595 6137
rect 18539 6081 18595 6091
rect 18711 6207 18767 6217
rect 18711 6161 18713 6207
rect 18713 6161 18765 6207
rect 18765 6161 18767 6207
rect 18711 6091 18713 6137
rect 18713 6091 18765 6137
rect 18765 6091 18767 6137
rect 18711 6081 18767 6091
rect 18883 6207 18939 6217
rect 18883 6161 18885 6207
rect 18885 6161 18937 6207
rect 18937 6161 18939 6207
rect 18883 6091 18885 6137
rect 18885 6091 18937 6137
rect 18937 6091 18939 6137
rect 18883 6081 18939 6091
rect 19055 6207 19111 6217
rect 19055 6161 19057 6207
rect 19057 6161 19109 6207
rect 19109 6161 19111 6207
rect 19055 6091 19057 6137
rect 19057 6091 19109 6137
rect 19109 6091 19111 6137
rect 19055 6081 19111 6091
rect 19227 6207 19283 6217
rect 19227 6161 19229 6207
rect 19229 6161 19281 6207
rect 19281 6161 19283 6207
rect 19227 6091 19229 6137
rect 19229 6091 19281 6137
rect 19281 6091 19283 6137
rect 19227 6081 19283 6091
rect 19399 6207 19455 6217
rect 19399 6161 19401 6207
rect 19401 6161 19453 6207
rect 19453 6161 19455 6207
rect 19399 6091 19401 6137
rect 19401 6091 19453 6137
rect 19453 6091 19455 6137
rect 19399 6081 19455 6091
rect 19571 6207 19627 6217
rect 19571 6161 19573 6207
rect 19573 6161 19625 6207
rect 19625 6161 19627 6207
rect 19571 6091 19573 6137
rect 19573 6091 19625 6137
rect 19625 6091 19627 6137
rect 19571 6081 19627 6091
rect 19743 6207 19799 6217
rect 19743 6161 19745 6207
rect 19745 6161 19797 6207
rect 19797 6161 19799 6207
rect 19743 6091 19745 6137
rect 19745 6091 19797 6137
rect 19797 6091 19799 6137
rect 19743 6081 19799 6091
rect 19915 6207 19971 6217
rect 19915 6161 19917 6207
rect 19917 6161 19969 6207
rect 19969 6161 19971 6207
rect 19915 6091 19917 6137
rect 19917 6091 19969 6137
rect 19969 6091 19971 6137
rect 19915 6081 19971 6091
rect 16648 4811 16704 4813
rect 16728 4811 16784 4813
rect 16808 4811 16864 4813
rect 16888 4811 16944 4813
rect 16968 4811 17024 4813
rect 17048 4811 17104 4813
rect 17128 4811 17184 4813
rect 17208 4811 17264 4813
rect 17288 4811 17344 4813
rect 16648 4759 16690 4811
rect 16690 4759 16702 4811
rect 16702 4759 16704 4811
rect 16728 4759 16754 4811
rect 16754 4759 16766 4811
rect 16766 4759 16784 4811
rect 16808 4759 16818 4811
rect 16818 4759 16830 4811
rect 16830 4759 16864 4811
rect 16888 4759 16894 4811
rect 16894 4759 16944 4811
rect 16968 4759 17010 4811
rect 17010 4759 17022 4811
rect 17022 4759 17024 4811
rect 17048 4759 17074 4811
rect 17074 4759 17086 4811
rect 17086 4759 17104 4811
rect 17128 4759 17138 4811
rect 17138 4759 17150 4811
rect 17150 4759 17184 4811
rect 17208 4759 17214 4811
rect 17214 4759 17264 4811
rect 17288 4759 17330 4811
rect 17330 4759 17344 4811
rect 16648 4757 16704 4759
rect 16728 4757 16784 4759
rect 16808 4757 16864 4759
rect 16888 4757 16944 4759
rect 16968 4757 17024 4759
rect 17048 4757 17104 4759
rect 17128 4757 17184 4759
rect 17208 4757 17264 4759
rect 17288 4757 17344 4759
rect 17472 4811 17528 4813
rect 17552 4811 17608 4813
rect 17632 4811 17688 4813
rect 17712 4811 17768 4813
rect 17792 4811 17848 4813
rect 17872 4811 17928 4813
rect 17952 4811 18008 4813
rect 18032 4811 18088 4813
rect 18112 4811 18168 4813
rect 17472 4759 17492 4811
rect 17492 4759 17528 4811
rect 17552 4759 17556 4811
rect 17556 4759 17608 4811
rect 17632 4759 17672 4811
rect 17672 4759 17684 4811
rect 17684 4759 17688 4811
rect 17712 4759 17736 4811
rect 17736 4759 17748 4811
rect 17748 4759 17768 4811
rect 17792 4759 17800 4811
rect 17800 4759 17812 4811
rect 17812 4759 17848 4811
rect 17872 4759 17876 4811
rect 17876 4759 17928 4811
rect 17952 4759 17992 4811
rect 17992 4759 18004 4811
rect 18004 4759 18008 4811
rect 18032 4759 18056 4811
rect 18056 4759 18068 4811
rect 18068 4759 18088 4811
rect 18112 4759 18120 4811
rect 18120 4759 18132 4811
rect 18132 4759 18168 4811
rect 17472 4757 17528 4759
rect 17552 4757 17608 4759
rect 17632 4757 17688 4759
rect 17712 4757 17768 4759
rect 17792 4757 17848 4759
rect 17872 4757 17928 4759
rect 17952 4757 18008 4759
rect 18032 4757 18088 4759
rect 18112 4757 18168 4759
rect 16555 4713 16557 4714
rect 16557 4713 16609 4714
rect 16609 4713 16611 4714
rect 16555 4701 16611 4713
rect 16555 4658 16557 4701
rect 16557 4658 16609 4701
rect 16609 4658 16611 4701
rect 18205 4713 18207 4714
rect 18207 4713 18259 4714
rect 18259 4713 18261 4714
rect 18205 4701 18261 4713
rect 16555 4585 16557 4634
rect 16557 4585 16609 4634
rect 16609 4585 16611 4634
rect 16555 4578 16611 4585
rect 18205 4658 18207 4701
rect 18207 4658 18259 4701
rect 18259 4658 18261 4701
rect 16555 4521 16557 4554
rect 16557 4521 16609 4554
rect 16609 4521 16611 4554
rect 18205 4585 18207 4634
rect 18207 4585 18259 4634
rect 18259 4585 18261 4634
rect 18205 4578 18261 4585
rect 16555 4509 16611 4521
rect 16555 4498 16557 4509
rect 16557 4498 16609 4509
rect 16609 4498 16611 4509
rect 16555 4457 16557 4474
rect 16557 4457 16609 4474
rect 16609 4457 16611 4474
rect 16555 4445 16611 4457
rect 16555 4418 16557 4445
rect 16557 4418 16609 4445
rect 16609 4418 16611 4445
rect 18205 4521 18207 4554
rect 18207 4521 18259 4554
rect 18259 4521 18261 4554
rect 18205 4509 18261 4521
rect 18205 4498 18207 4509
rect 18207 4498 18259 4509
rect 18259 4498 18261 4509
rect 16555 4393 16557 4394
rect 16557 4393 16609 4394
rect 16609 4393 16611 4394
rect 16555 4381 16611 4393
rect 16555 4338 16557 4381
rect 16557 4338 16609 4381
rect 16609 4338 16611 4381
rect 18205 4457 18207 4474
rect 18207 4457 18259 4474
rect 18259 4457 18261 4474
rect 18205 4445 18261 4457
rect 18205 4418 18207 4445
rect 18207 4418 18259 4445
rect 18259 4418 18261 4445
rect 16555 4265 16557 4314
rect 16557 4265 16609 4314
rect 16609 4265 16611 4314
rect 16555 4258 16611 4265
rect 18205 4393 18207 4394
rect 18207 4393 18259 4394
rect 18259 4393 18261 4394
rect 18205 4381 18261 4393
rect 18205 4338 18207 4381
rect 18207 4338 18259 4381
rect 18259 4338 18261 4381
rect 16555 4201 16557 4234
rect 16557 4201 16609 4234
rect 16609 4201 16611 4234
rect 16555 4189 16611 4201
rect 18205 4265 18207 4314
rect 18207 4265 18259 4314
rect 18259 4265 18261 4314
rect 18205 4258 18261 4265
rect 16555 4178 16557 4189
rect 16557 4178 16609 4189
rect 16609 4178 16611 4189
rect 16555 4137 16557 4154
rect 16557 4137 16609 4154
rect 16609 4137 16611 4154
rect 16555 4098 16611 4137
rect 18205 4201 18207 4234
rect 18207 4201 18259 4234
rect 18259 4201 18261 4234
rect 18205 4189 18261 4201
rect 18205 4178 18207 4189
rect 18207 4178 18259 4189
rect 18259 4178 18261 4189
rect 18205 4137 18207 4154
rect 18207 4137 18259 4154
rect 18259 4137 18261 4154
rect 18205 4098 18261 4137
rect 16740 4060 16796 4062
rect 16820 4060 16876 4062
rect 16900 4060 16956 4062
rect 16980 4060 17036 4062
rect 17060 4060 17116 4062
rect 17140 4060 17196 4062
rect 17220 4060 17276 4062
rect 17300 4060 17356 4062
rect 16740 4008 16771 4060
rect 16771 4008 16783 4060
rect 16783 4008 16796 4060
rect 16820 4008 16835 4060
rect 16835 4008 16847 4060
rect 16847 4008 16876 4060
rect 16900 4008 16911 4060
rect 16911 4008 16956 4060
rect 16980 4008 17027 4060
rect 17027 4008 17036 4060
rect 17060 4008 17091 4060
rect 17091 4008 17103 4060
rect 17103 4008 17116 4060
rect 17140 4008 17155 4060
rect 17155 4008 17167 4060
rect 17167 4008 17196 4060
rect 17220 4008 17231 4060
rect 17231 4008 17276 4060
rect 17300 4008 17347 4060
rect 17347 4008 17356 4060
rect 16740 4006 16796 4008
rect 16820 4006 16876 4008
rect 16900 4006 16956 4008
rect 16980 4006 17036 4008
rect 17060 4006 17116 4008
rect 17140 4006 17196 4008
rect 17220 4006 17276 4008
rect 17300 4006 17356 4008
rect 17380 4006 17436 4062
rect 17460 4060 17516 4062
rect 17540 4060 17596 4062
rect 17620 4060 17676 4062
rect 17700 4060 17756 4062
rect 17780 4060 17836 4062
rect 17860 4060 17916 4062
rect 17940 4060 17996 4062
rect 18020 4060 18076 4062
rect 18498 4811 18554 4813
rect 18578 4811 18634 4813
rect 18658 4811 18714 4813
rect 18738 4811 18794 4813
rect 18818 4811 18874 4813
rect 18898 4811 18954 4813
rect 18978 4811 19034 4813
rect 19058 4811 19114 4813
rect 19138 4811 19194 4813
rect 18498 4759 18540 4811
rect 18540 4759 18552 4811
rect 18552 4759 18554 4811
rect 18578 4759 18604 4811
rect 18604 4759 18616 4811
rect 18616 4759 18634 4811
rect 18658 4759 18668 4811
rect 18668 4759 18680 4811
rect 18680 4759 18714 4811
rect 18738 4759 18744 4811
rect 18744 4759 18794 4811
rect 18818 4759 18860 4811
rect 18860 4759 18872 4811
rect 18872 4759 18874 4811
rect 18898 4759 18924 4811
rect 18924 4759 18936 4811
rect 18936 4759 18954 4811
rect 18978 4759 18988 4811
rect 18988 4759 19000 4811
rect 19000 4759 19034 4811
rect 19058 4759 19064 4811
rect 19064 4759 19114 4811
rect 19138 4759 19180 4811
rect 19180 4759 19194 4811
rect 18498 4757 18554 4759
rect 18578 4757 18634 4759
rect 18658 4757 18714 4759
rect 18738 4757 18794 4759
rect 18818 4757 18874 4759
rect 18898 4757 18954 4759
rect 18978 4757 19034 4759
rect 19058 4757 19114 4759
rect 19138 4757 19194 4759
rect 19322 4811 19378 4813
rect 19402 4811 19458 4813
rect 19482 4811 19538 4813
rect 19562 4811 19618 4813
rect 19642 4811 19698 4813
rect 19722 4811 19778 4813
rect 19802 4811 19858 4813
rect 19882 4811 19938 4813
rect 19962 4811 20018 4813
rect 19322 4759 19342 4811
rect 19342 4759 19378 4811
rect 19402 4759 19406 4811
rect 19406 4759 19458 4811
rect 19482 4759 19522 4811
rect 19522 4759 19534 4811
rect 19534 4759 19538 4811
rect 19562 4759 19586 4811
rect 19586 4759 19598 4811
rect 19598 4759 19618 4811
rect 19642 4759 19650 4811
rect 19650 4759 19662 4811
rect 19662 4759 19698 4811
rect 19722 4759 19726 4811
rect 19726 4759 19778 4811
rect 19802 4759 19842 4811
rect 19842 4759 19854 4811
rect 19854 4759 19858 4811
rect 19882 4759 19906 4811
rect 19906 4759 19918 4811
rect 19918 4759 19938 4811
rect 19962 4759 19970 4811
rect 19970 4759 19982 4811
rect 19982 4759 20018 4811
rect 19322 4757 19378 4759
rect 19402 4757 19458 4759
rect 19482 4757 19538 4759
rect 19562 4757 19618 4759
rect 19642 4757 19698 4759
rect 19722 4757 19778 4759
rect 19802 4757 19858 4759
rect 19882 4757 19938 4759
rect 19962 4757 20018 4759
rect 18405 4713 18407 4714
rect 18407 4713 18459 4714
rect 18459 4713 18461 4714
rect 18405 4701 18461 4713
rect 18405 4658 18407 4701
rect 18407 4658 18459 4701
rect 18459 4658 18461 4701
rect 20055 4713 20057 4714
rect 20057 4713 20109 4714
rect 20109 4713 20111 4714
rect 20055 4701 20111 4713
rect 18405 4585 18407 4634
rect 18407 4585 18459 4634
rect 18459 4585 18461 4634
rect 18405 4578 18461 4585
rect 20055 4658 20057 4701
rect 20057 4658 20109 4701
rect 20109 4658 20111 4701
rect 18405 4521 18407 4554
rect 18407 4521 18459 4554
rect 18459 4521 18461 4554
rect 20055 4585 20057 4634
rect 20057 4585 20109 4634
rect 20109 4585 20111 4634
rect 20055 4578 20111 4585
rect 18405 4509 18461 4521
rect 18405 4498 18407 4509
rect 18407 4498 18459 4509
rect 18459 4498 18461 4509
rect 18405 4457 18407 4474
rect 18407 4457 18459 4474
rect 18459 4457 18461 4474
rect 18405 4445 18461 4457
rect 18405 4418 18407 4445
rect 18407 4418 18459 4445
rect 18459 4418 18461 4445
rect 20055 4521 20057 4554
rect 20057 4521 20109 4554
rect 20109 4521 20111 4554
rect 20055 4509 20111 4521
rect 20055 4498 20057 4509
rect 20057 4498 20109 4509
rect 20109 4498 20111 4509
rect 18405 4393 18407 4394
rect 18407 4393 18459 4394
rect 18459 4393 18461 4394
rect 18405 4381 18461 4393
rect 18405 4338 18407 4381
rect 18407 4338 18459 4381
rect 18459 4338 18461 4381
rect 20055 4457 20057 4474
rect 20057 4457 20109 4474
rect 20109 4457 20111 4474
rect 20055 4445 20111 4457
rect 20055 4418 20057 4445
rect 20057 4418 20109 4445
rect 20109 4418 20111 4445
rect 18405 4265 18407 4314
rect 18407 4265 18459 4314
rect 18459 4265 18461 4314
rect 18405 4258 18461 4265
rect 20055 4393 20057 4394
rect 20057 4393 20109 4394
rect 20109 4393 20111 4394
rect 20055 4381 20111 4393
rect 20055 4338 20057 4381
rect 20057 4338 20109 4381
rect 20109 4338 20111 4381
rect 18405 4201 18407 4234
rect 18407 4201 18459 4234
rect 18459 4201 18461 4234
rect 18405 4189 18461 4201
rect 20055 4265 20057 4314
rect 20057 4265 20109 4314
rect 20109 4265 20111 4314
rect 20055 4258 20111 4265
rect 18405 4178 18407 4189
rect 18407 4178 18459 4189
rect 18459 4178 18461 4189
rect 18405 4137 18407 4154
rect 18407 4137 18459 4154
rect 18459 4137 18461 4154
rect 18405 4098 18461 4137
rect 20055 4201 20057 4234
rect 20057 4201 20109 4234
rect 20109 4201 20111 4234
rect 20055 4189 20111 4201
rect 20055 4178 20057 4189
rect 20057 4178 20109 4189
rect 20109 4178 20111 4189
rect 20055 4137 20057 4154
rect 20057 4137 20109 4154
rect 20109 4137 20111 4154
rect 20055 4098 20111 4137
rect 18590 4060 18646 4062
rect 18670 4060 18726 4062
rect 18750 4060 18806 4062
rect 18830 4060 18886 4062
rect 18910 4060 18966 4062
rect 18990 4060 19046 4062
rect 19070 4060 19126 4062
rect 19150 4060 19206 4062
rect 17460 4008 17469 4060
rect 17469 4008 17516 4060
rect 17540 4008 17585 4060
rect 17585 4008 17596 4060
rect 17620 4008 17649 4060
rect 17649 4008 17661 4060
rect 17661 4008 17676 4060
rect 17700 4008 17713 4060
rect 17713 4008 17725 4060
rect 17725 4008 17756 4060
rect 17780 4008 17789 4060
rect 17789 4008 17836 4060
rect 17860 4008 17905 4060
rect 17905 4008 17916 4060
rect 17940 4008 17969 4060
rect 17969 4008 17981 4060
rect 17981 4008 17996 4060
rect 18020 4008 18033 4060
rect 18033 4008 18045 4060
rect 18045 4008 18076 4060
rect 18590 4008 18621 4060
rect 18621 4008 18633 4060
rect 18633 4008 18646 4060
rect 18670 4008 18685 4060
rect 18685 4008 18697 4060
rect 18697 4008 18726 4060
rect 18750 4008 18761 4060
rect 18761 4008 18806 4060
rect 18830 4008 18877 4060
rect 18877 4008 18886 4060
rect 18910 4008 18941 4060
rect 18941 4008 18953 4060
rect 18953 4008 18966 4060
rect 18990 4008 19005 4060
rect 19005 4008 19017 4060
rect 19017 4008 19046 4060
rect 19070 4008 19081 4060
rect 19081 4008 19126 4060
rect 19150 4008 19197 4060
rect 19197 4008 19206 4060
rect 17460 4006 17516 4008
rect 17540 4006 17596 4008
rect 17620 4006 17676 4008
rect 17700 4006 17756 4008
rect 17780 4006 17836 4008
rect 17860 4006 17916 4008
rect 17940 4006 17996 4008
rect 18020 4006 18076 4008
rect 18590 4006 18646 4008
rect 18670 4006 18726 4008
rect 18750 4006 18806 4008
rect 18830 4006 18886 4008
rect 18910 4006 18966 4008
rect 18990 4006 19046 4008
rect 19070 4006 19126 4008
rect 19150 4006 19206 4008
rect 19230 4006 19286 4062
rect 19310 4060 19366 4062
rect 19390 4060 19446 4062
rect 19470 4060 19526 4062
rect 19550 4060 19606 4062
rect 19630 4060 19686 4062
rect 19710 4060 19766 4062
rect 19790 4060 19846 4062
rect 19870 4060 19926 4062
rect 19310 4008 19319 4060
rect 19319 4008 19366 4060
rect 19390 4008 19435 4060
rect 19435 4008 19446 4060
rect 19470 4008 19499 4060
rect 19499 4008 19511 4060
rect 19511 4008 19526 4060
rect 19550 4008 19563 4060
rect 19563 4008 19575 4060
rect 19575 4008 19606 4060
rect 19630 4008 19639 4060
rect 19639 4008 19686 4060
rect 19710 4008 19755 4060
rect 19755 4008 19766 4060
rect 19790 4008 19819 4060
rect 19819 4008 19831 4060
rect 19831 4008 19846 4060
rect 19870 4008 19883 4060
rect 19883 4008 19895 4060
rect 19895 4008 19926 4060
rect 19310 4006 19366 4008
rect 19390 4006 19446 4008
rect 19470 4006 19526 4008
rect 19550 4006 19606 4008
rect 19630 4006 19686 4008
rect 19710 4006 19766 4008
rect 19790 4006 19846 4008
rect 19870 4006 19926 4008
rect 16555 3931 16611 3970
rect 16555 3914 16557 3931
rect 16557 3914 16609 3931
rect 16609 3914 16611 3931
rect 16555 3879 16557 3890
rect 16557 3879 16609 3890
rect 16609 3879 16611 3890
rect 16555 3867 16611 3879
rect 16555 3834 16557 3867
rect 16557 3834 16609 3867
rect 16609 3834 16611 3867
rect 18205 3931 18261 3970
rect 18205 3914 18207 3931
rect 18207 3914 18259 3931
rect 18259 3914 18261 3931
rect 18405 3931 18461 3970
rect 18405 3914 18407 3931
rect 18407 3914 18459 3931
rect 18459 3914 18461 3931
rect 18205 3879 18207 3890
rect 18207 3879 18259 3890
rect 18259 3879 18261 3890
rect 16555 3803 16611 3810
rect 16555 3754 16557 3803
rect 16557 3754 16609 3803
rect 16609 3754 16611 3803
rect 18205 3867 18261 3879
rect 18205 3834 18207 3867
rect 18207 3834 18259 3867
rect 18259 3834 18261 3867
rect 18405 3879 18407 3890
rect 18407 3879 18459 3890
rect 18459 3879 18461 3890
rect 18405 3867 18461 3879
rect 18405 3834 18407 3867
rect 18407 3834 18459 3867
rect 18459 3834 18461 3867
rect 20055 3931 20111 3970
rect 20055 3914 20057 3931
rect 20057 3914 20109 3931
rect 20109 3914 20111 3931
rect 20055 3879 20057 3890
rect 20057 3879 20109 3890
rect 20109 3879 20111 3890
rect 16555 3687 16557 3730
rect 16557 3687 16609 3730
rect 16609 3687 16611 3730
rect 16555 3675 16611 3687
rect 16555 3674 16557 3675
rect 16557 3674 16609 3675
rect 16609 3674 16611 3675
rect 18205 3803 18261 3810
rect 18205 3754 18207 3803
rect 18207 3754 18259 3803
rect 18259 3754 18261 3803
rect 18405 3803 18461 3810
rect 18405 3754 18407 3803
rect 18407 3754 18459 3803
rect 18459 3754 18461 3803
rect 20055 3867 20111 3879
rect 20055 3834 20057 3867
rect 20057 3834 20109 3867
rect 20109 3834 20111 3867
rect 16555 3623 16557 3650
rect 16557 3623 16609 3650
rect 16609 3623 16611 3650
rect 16555 3611 16611 3623
rect 16555 3594 16557 3611
rect 16557 3594 16609 3611
rect 16609 3594 16611 3611
rect 18205 3687 18207 3730
rect 18207 3687 18259 3730
rect 18259 3687 18261 3730
rect 18205 3675 18261 3687
rect 18205 3674 18207 3675
rect 18207 3674 18259 3675
rect 18259 3674 18261 3675
rect 18405 3687 18407 3730
rect 18407 3687 18459 3730
rect 18459 3687 18461 3730
rect 18405 3675 18461 3687
rect 18405 3674 18407 3675
rect 18407 3674 18459 3675
rect 18459 3674 18461 3675
rect 20055 3803 20111 3810
rect 20055 3754 20057 3803
rect 20057 3754 20109 3803
rect 20109 3754 20111 3803
rect 16555 3559 16557 3570
rect 16557 3559 16609 3570
rect 16609 3559 16611 3570
rect 16555 3547 16611 3559
rect 16555 3514 16557 3547
rect 16557 3514 16609 3547
rect 16609 3514 16611 3547
rect 18205 3623 18207 3650
rect 18207 3623 18259 3650
rect 18259 3623 18261 3650
rect 18205 3611 18261 3623
rect 18205 3594 18207 3611
rect 18207 3594 18259 3611
rect 18259 3594 18261 3611
rect 18405 3623 18407 3650
rect 18407 3623 18459 3650
rect 18459 3623 18461 3650
rect 18405 3611 18461 3623
rect 18405 3594 18407 3611
rect 18407 3594 18459 3611
rect 18459 3594 18461 3611
rect 20055 3687 20057 3730
rect 20057 3687 20109 3730
rect 20109 3687 20111 3730
rect 20055 3675 20111 3687
rect 20055 3674 20057 3675
rect 20057 3674 20109 3675
rect 20109 3674 20111 3675
rect 18205 3559 18207 3570
rect 18207 3559 18259 3570
rect 18259 3559 18261 3570
rect 18205 3547 18261 3559
rect 16555 3483 16611 3490
rect 16555 3434 16557 3483
rect 16557 3434 16609 3483
rect 16609 3434 16611 3483
rect 18205 3514 18207 3547
rect 18207 3514 18259 3547
rect 18259 3514 18261 3547
rect 18405 3559 18407 3570
rect 18407 3559 18459 3570
rect 18459 3559 18461 3570
rect 18405 3547 18461 3559
rect 18405 3514 18407 3547
rect 18407 3514 18459 3547
rect 18459 3514 18461 3547
rect 20055 3623 20057 3650
rect 20057 3623 20109 3650
rect 20109 3623 20111 3650
rect 20055 3611 20111 3623
rect 20055 3594 20057 3611
rect 20057 3594 20109 3611
rect 20109 3594 20111 3611
rect 20055 3559 20057 3570
rect 20057 3559 20109 3570
rect 20109 3559 20111 3570
rect 20055 3547 20111 3559
rect 16555 3367 16557 3410
rect 16557 3367 16609 3410
rect 16609 3367 16611 3410
rect 18205 3483 18261 3490
rect 18205 3434 18207 3483
rect 18207 3434 18259 3483
rect 18259 3434 18261 3483
rect 18405 3483 18461 3490
rect 18405 3434 18407 3483
rect 18407 3434 18459 3483
rect 18459 3434 18461 3483
rect 20055 3514 20057 3547
rect 20057 3514 20109 3547
rect 20109 3514 20111 3547
rect 16555 3355 16611 3367
rect 16555 3354 16557 3355
rect 16557 3354 16609 3355
rect 16609 3354 16611 3355
rect 18205 3367 18207 3410
rect 18207 3367 18259 3410
rect 18259 3367 18261 3410
rect 18205 3355 18261 3367
rect 18205 3354 18207 3355
rect 18207 3354 18259 3355
rect 18259 3354 18261 3355
rect 18405 3367 18407 3410
rect 18407 3367 18459 3410
rect 18459 3367 18461 3410
rect 20055 3483 20111 3490
rect 20055 3434 20057 3483
rect 20057 3434 20109 3483
rect 20109 3434 20111 3483
rect 18405 3355 18461 3367
rect 18405 3354 18407 3355
rect 18407 3354 18459 3355
rect 18459 3354 18461 3355
rect 16648 3309 16704 3311
rect 16728 3309 16784 3311
rect 16808 3309 16864 3311
rect 16888 3309 16944 3311
rect 16968 3309 17024 3311
rect 17048 3309 17104 3311
rect 17128 3309 17184 3311
rect 17208 3309 17264 3311
rect 17288 3309 17344 3311
rect 16648 3257 16690 3309
rect 16690 3257 16702 3309
rect 16702 3257 16704 3309
rect 16728 3257 16754 3309
rect 16754 3257 16766 3309
rect 16766 3257 16784 3309
rect 16808 3257 16818 3309
rect 16818 3257 16830 3309
rect 16830 3257 16864 3309
rect 16888 3257 16894 3309
rect 16894 3257 16944 3309
rect 16968 3257 17010 3309
rect 17010 3257 17022 3309
rect 17022 3257 17024 3309
rect 17048 3257 17074 3309
rect 17074 3257 17086 3309
rect 17086 3257 17104 3309
rect 17128 3257 17138 3309
rect 17138 3257 17150 3309
rect 17150 3257 17184 3309
rect 17208 3257 17214 3309
rect 17214 3257 17264 3309
rect 17288 3257 17330 3309
rect 17330 3257 17344 3309
rect 16648 3255 16704 3257
rect 16728 3255 16784 3257
rect 16808 3255 16864 3257
rect 16888 3255 16944 3257
rect 16968 3255 17024 3257
rect 17048 3255 17104 3257
rect 17128 3255 17184 3257
rect 17208 3255 17264 3257
rect 17288 3255 17344 3257
rect 17472 3309 17528 3311
rect 17552 3309 17608 3311
rect 17632 3309 17688 3311
rect 17712 3309 17768 3311
rect 17792 3309 17848 3311
rect 17872 3309 17928 3311
rect 17952 3309 18008 3311
rect 18032 3309 18088 3311
rect 18112 3309 18168 3311
rect 17472 3257 17492 3309
rect 17492 3257 17528 3309
rect 17552 3257 17556 3309
rect 17556 3257 17608 3309
rect 17632 3257 17672 3309
rect 17672 3257 17684 3309
rect 17684 3257 17688 3309
rect 17712 3257 17736 3309
rect 17736 3257 17748 3309
rect 17748 3257 17768 3309
rect 17792 3257 17800 3309
rect 17800 3257 17812 3309
rect 17812 3257 17848 3309
rect 17872 3257 17876 3309
rect 17876 3257 17928 3309
rect 17952 3257 17992 3309
rect 17992 3257 18004 3309
rect 18004 3257 18008 3309
rect 18032 3257 18056 3309
rect 18056 3257 18068 3309
rect 18068 3257 18088 3309
rect 18112 3257 18120 3309
rect 18120 3257 18132 3309
rect 18132 3257 18168 3309
rect 20055 3367 20057 3410
rect 20057 3367 20109 3410
rect 20109 3367 20111 3410
rect 20055 3355 20111 3367
rect 20055 3354 20057 3355
rect 20057 3354 20109 3355
rect 20109 3354 20111 3355
rect 18498 3309 18554 3311
rect 18578 3309 18634 3311
rect 18658 3309 18714 3311
rect 18738 3309 18794 3311
rect 18818 3309 18874 3311
rect 18898 3309 18954 3311
rect 18978 3309 19034 3311
rect 19058 3309 19114 3311
rect 19138 3309 19194 3311
rect 18498 3257 18540 3309
rect 18540 3257 18552 3309
rect 18552 3257 18554 3309
rect 18578 3257 18604 3309
rect 18604 3257 18616 3309
rect 18616 3257 18634 3309
rect 18658 3257 18668 3309
rect 18668 3257 18680 3309
rect 18680 3257 18714 3309
rect 18738 3257 18744 3309
rect 18744 3257 18794 3309
rect 18818 3257 18860 3309
rect 18860 3257 18872 3309
rect 18872 3257 18874 3309
rect 18898 3257 18924 3309
rect 18924 3257 18936 3309
rect 18936 3257 18954 3309
rect 18978 3257 18988 3309
rect 18988 3257 19000 3309
rect 19000 3257 19034 3309
rect 19058 3257 19064 3309
rect 19064 3257 19114 3309
rect 19138 3257 19180 3309
rect 19180 3257 19194 3309
rect 17472 3255 17528 3257
rect 17552 3255 17608 3257
rect 17632 3255 17688 3257
rect 17712 3255 17768 3257
rect 17792 3255 17848 3257
rect 17872 3255 17928 3257
rect 17952 3255 18008 3257
rect 18032 3255 18088 3257
rect 18112 3255 18168 3257
rect 18498 3255 18554 3257
rect 18578 3255 18634 3257
rect 18658 3255 18714 3257
rect 18738 3255 18794 3257
rect 18818 3255 18874 3257
rect 18898 3255 18954 3257
rect 18978 3255 19034 3257
rect 19058 3255 19114 3257
rect 19138 3255 19194 3257
rect 19322 3309 19378 3311
rect 19402 3309 19458 3311
rect 19482 3309 19538 3311
rect 19562 3309 19618 3311
rect 19642 3309 19698 3311
rect 19722 3309 19778 3311
rect 19802 3309 19858 3311
rect 19882 3309 19938 3311
rect 19962 3309 20018 3311
rect 19322 3257 19342 3309
rect 19342 3257 19378 3309
rect 19402 3257 19406 3309
rect 19406 3257 19458 3309
rect 19482 3257 19522 3309
rect 19522 3257 19534 3309
rect 19534 3257 19538 3309
rect 19562 3257 19586 3309
rect 19586 3257 19598 3309
rect 19598 3257 19618 3309
rect 19642 3257 19650 3309
rect 19650 3257 19662 3309
rect 19662 3257 19698 3309
rect 19722 3257 19726 3309
rect 19726 3257 19778 3309
rect 19802 3257 19842 3309
rect 19842 3257 19854 3309
rect 19854 3257 19858 3309
rect 19882 3257 19906 3309
rect 19906 3257 19918 3309
rect 19918 3257 19938 3309
rect 19962 3257 19970 3309
rect 19970 3257 19982 3309
rect 19982 3257 20018 3309
rect 19322 3255 19378 3257
rect 19402 3255 19458 3257
rect 19482 3255 19538 3257
rect 19562 3255 19618 3257
rect 19642 3255 19698 3257
rect 19722 3255 19778 3257
rect 19802 3255 19858 3257
rect 19882 3255 19938 3257
rect 19962 3255 20018 3257
<< metal3 >>
rect 15300 10700 16400 10800
rect 15300 9900 15400 10700
rect 16300 9900 16400 10700
rect 15300 9400 16400 9900
rect 16550 9863 18266 9868
rect 16550 9807 16648 9863
rect 16704 9807 16728 9863
rect 16784 9807 16808 9863
rect 16864 9807 16888 9863
rect 16944 9807 16968 9863
rect 17024 9807 17048 9863
rect 17104 9807 17128 9863
rect 17184 9807 17208 9863
rect 17264 9807 17288 9863
rect 17344 9807 17472 9863
rect 17528 9807 17552 9863
rect 17608 9807 17632 9863
rect 17688 9807 17712 9863
rect 17768 9807 17792 9863
rect 17848 9807 17872 9863
rect 17928 9807 17952 9863
rect 18008 9807 18032 9863
rect 18088 9807 18112 9863
rect 18168 9807 18266 9863
rect 16550 9802 18266 9807
rect 16550 9764 16616 9802
rect 16550 9708 16555 9764
rect 16611 9708 16616 9764
rect 16550 9684 16616 9708
rect 16550 9628 16555 9684
rect 16611 9628 16616 9684
rect 16550 9604 16616 9628
rect 16550 9548 16555 9604
rect 16611 9548 16616 9604
rect 16550 9524 16616 9548
rect 16550 9468 16555 9524
rect 16611 9468 16616 9524
rect 16550 9444 16616 9468
rect 16550 9388 16555 9444
rect 16611 9388 16616 9444
rect 16550 9364 16616 9388
rect 16550 9308 16555 9364
rect 16611 9308 16616 9364
rect 16550 9284 16616 9308
rect 16550 9228 16555 9284
rect 16611 9228 16616 9284
rect 16550 9204 16616 9228
rect 11600 7100 12500 9200
rect 12750 7100 13250 9200
rect 13500 7100 13800 9200
rect 14050 7100 14350 8200
rect 14600 7100 16300 9200
rect 16550 9148 16555 9204
rect 16611 9148 16616 9204
rect 16550 9020 16616 9148
rect 16550 8964 16555 9020
rect 16611 8964 16616 9020
rect 16550 8940 16616 8964
rect 16550 8884 16555 8940
rect 16611 8884 16616 8940
rect 16550 8860 16616 8884
rect 16550 8804 16555 8860
rect 16611 8804 16616 8860
rect 16550 8780 16616 8804
rect 16550 8724 16555 8780
rect 16611 8724 16616 8780
rect 16550 8700 16616 8724
rect 16550 8644 16555 8700
rect 16611 8644 16616 8700
rect 16550 8620 16616 8644
rect 16550 8564 16555 8620
rect 16611 8564 16616 8620
rect 16550 8540 16616 8564
rect 16550 8484 16555 8540
rect 16611 8484 16616 8540
rect 16550 8460 16616 8484
rect 16550 8404 16555 8460
rect 16611 8404 16616 8460
rect 16676 9117 16754 9742
rect 16814 9177 16892 9802
rect 16952 9642 17030 9742
rect 16952 9117 16953 9642
rect 17090 9177 17168 9802
rect 17228 9643 17306 9742
rect 17305 9117 17306 9643
rect 17369 9177 17447 9802
rect 17510 9643 17588 9742
rect 17587 9117 17588 9643
rect 17648 9177 17726 9802
rect 17786 9643 17864 9742
rect 17863 9117 17864 9643
rect 17924 9177 18002 9802
rect 18200 9764 18266 9802
rect 18062 9643 18140 9742
rect 16676 9112 16811 9117
rect 16676 9056 16740 9112
rect 16796 9056 16811 9112
rect 16676 9051 16811 9056
rect 16676 8426 16754 9051
rect 16550 8366 16616 8404
rect 16814 8366 16892 8991
rect 16952 8426 17030 9051
rect 17090 8366 17168 8991
rect 17228 8426 17306 9051
rect 17369 8366 17447 8991
rect 17510 8426 17588 9051
rect 17648 8366 17726 8991
rect 17786 8426 17864 9051
rect 17924 8366 18002 8991
rect 18062 8426 18140 9051
rect 18200 9708 18205 9764
rect 18261 9708 18266 9764
rect 18200 9684 18266 9708
rect 18200 9628 18205 9684
rect 18261 9628 18266 9684
rect 18200 9604 18266 9628
rect 18200 9548 18205 9604
rect 18261 9548 18266 9604
rect 18200 9524 18266 9548
rect 18200 9468 18205 9524
rect 18261 9468 18266 9524
rect 18200 9444 18266 9468
rect 18200 9388 18205 9444
rect 18261 9388 18266 9444
rect 18200 9364 18266 9388
rect 18200 9308 18205 9364
rect 18261 9308 18266 9364
rect 18200 9284 18266 9308
rect 18200 9228 18205 9284
rect 18261 9228 18266 9284
rect 18200 9204 18266 9228
rect 18200 9148 18205 9204
rect 18261 9148 18266 9204
rect 18200 9020 18266 9148
rect 18200 8964 18205 9020
rect 18261 8964 18266 9020
rect 18200 8940 18266 8964
rect 18200 8884 18205 8940
rect 18261 8884 18266 8940
rect 18200 8860 18266 8884
rect 18200 8804 18205 8860
rect 18261 8804 18266 8860
rect 18200 8780 18266 8804
rect 18200 8724 18205 8780
rect 18261 8724 18266 8780
rect 18200 8700 18266 8724
rect 18200 8644 18205 8700
rect 18261 8644 18266 8700
rect 18200 8620 18266 8644
rect 18200 8564 18205 8620
rect 18261 8564 18266 8620
rect 18200 8540 18266 8564
rect 18200 8484 18205 8540
rect 18261 8484 18266 8540
rect 18200 8460 18266 8484
rect 18200 8404 18205 8460
rect 18261 8404 18266 8460
rect 18200 8366 18266 8404
rect 16550 8361 18266 8366
rect 16550 8305 16648 8361
rect 16704 8305 16728 8361
rect 16784 8305 16808 8361
rect 16864 8305 16888 8361
rect 16944 8305 16968 8361
rect 17024 8305 17048 8361
rect 17104 8305 17128 8361
rect 17184 8305 17208 8361
rect 17264 8305 17288 8361
rect 17344 8305 17472 8361
rect 17528 8305 17552 8361
rect 17608 8305 17632 8361
rect 17688 8305 17712 8361
rect 17768 8305 17792 8361
rect 17848 8305 17872 8361
rect 17928 8305 17952 8361
rect 18008 8305 18032 8361
rect 18088 8305 18112 8361
rect 18168 8305 18266 8361
rect 16550 8300 18266 8305
rect 18400 9863 20116 9868
rect 18400 9807 18498 9863
rect 18554 9807 18578 9863
rect 18634 9807 18658 9863
rect 18714 9807 18738 9863
rect 18794 9807 18818 9863
rect 18874 9807 18898 9863
rect 18954 9807 18978 9863
rect 19034 9807 19058 9863
rect 19114 9807 19138 9863
rect 19194 9807 19322 9863
rect 19378 9807 19402 9863
rect 19458 9807 19482 9863
rect 19538 9807 19562 9863
rect 19618 9807 19642 9863
rect 19698 9807 19722 9863
rect 19778 9807 19802 9863
rect 19858 9807 19882 9863
rect 19938 9807 19962 9863
rect 20018 9807 20116 9863
rect 18400 9802 20116 9807
rect 18400 9764 18466 9802
rect 18400 9708 18405 9764
rect 18461 9708 18466 9764
rect 18400 9684 18466 9708
rect 18400 9628 18405 9684
rect 18461 9628 18466 9684
rect 18400 9604 18466 9628
rect 18400 9548 18405 9604
rect 18461 9548 18466 9604
rect 18400 9524 18466 9548
rect 18400 9468 18405 9524
rect 18461 9468 18466 9524
rect 18400 9444 18466 9468
rect 18400 9388 18405 9444
rect 18461 9388 18466 9444
rect 18400 9364 18466 9388
rect 18400 9308 18405 9364
rect 18461 9308 18466 9364
rect 18400 9284 18466 9308
rect 18400 9228 18405 9284
rect 18461 9228 18466 9284
rect 18400 9204 18466 9228
rect 18400 9148 18405 9204
rect 18461 9148 18466 9204
rect 18400 9020 18466 9148
rect 18400 8964 18405 9020
rect 18461 8964 18466 9020
rect 18400 8940 18466 8964
rect 18400 8884 18405 8940
rect 18461 8884 18466 8940
rect 18400 8860 18466 8884
rect 18400 8804 18405 8860
rect 18461 8804 18466 8860
rect 18400 8780 18466 8804
rect 18400 8724 18405 8780
rect 18461 8724 18466 8780
rect 18400 8700 18466 8724
rect 18400 8644 18405 8700
rect 18461 8644 18466 8700
rect 18400 8620 18466 8644
rect 18400 8564 18405 8620
rect 18461 8564 18466 8620
rect 18400 8540 18466 8564
rect 18400 8484 18405 8540
rect 18461 8484 18466 8540
rect 18400 8460 18466 8484
rect 18400 8404 18405 8460
rect 18461 8404 18466 8460
rect 18526 9642 18604 9742
rect 18664 9177 18742 9802
rect 18802 9642 18880 9742
rect 18940 9177 19018 9802
rect 19078 9642 19156 9742
rect 19219 9177 19297 9802
rect 19360 9642 19438 9742
rect 19498 9177 19576 9802
rect 19636 9642 19714 9742
rect 19774 9177 19852 9802
rect 20050 9764 20116 9802
rect 19912 9117 19990 9742
rect 19714 9112 19990 9117
rect 19766 9056 19790 9112
rect 19846 9056 19870 9112
rect 19926 9056 19990 9112
rect 19714 9051 19990 9056
rect 18526 8426 18604 9051
rect 18400 8366 18466 8404
rect 18664 8366 18742 8991
rect 18802 8426 18880 9051
rect 18940 8366 19018 8991
rect 19078 8426 19156 9051
rect 19219 8366 19297 8991
rect 19360 8426 19438 9051
rect 19498 8366 19576 8991
rect 19636 8426 19714 9051
rect 19774 8366 19852 8991
rect 19912 8426 19990 9051
rect 20050 9708 20055 9764
rect 20111 9708 20116 9764
rect 20050 9684 20116 9708
rect 20050 9628 20055 9684
rect 20111 9628 20116 9684
rect 20050 9604 20116 9628
rect 20050 9548 20055 9604
rect 20111 9548 20116 9604
rect 20050 9524 20116 9548
rect 20050 9468 20055 9524
rect 20111 9468 20116 9524
rect 20050 9444 20116 9468
rect 20050 9388 20055 9444
rect 20111 9388 20116 9444
rect 20050 9364 20116 9388
rect 20050 9308 20055 9364
rect 20111 9308 20116 9364
rect 20050 9284 20116 9308
rect 20050 9228 20055 9284
rect 20111 9228 20116 9284
rect 20050 9204 20116 9228
rect 20050 9148 20055 9204
rect 20111 9148 20116 9204
rect 20050 9020 20116 9148
rect 20050 8964 20055 9020
rect 20111 8964 20116 9020
rect 20050 8940 20116 8964
rect 20050 8884 20055 8940
rect 20111 8884 20116 8940
rect 20050 8860 20116 8884
rect 20050 8804 20055 8860
rect 20111 8804 20116 8860
rect 20050 8780 20116 8804
rect 20050 8724 20055 8780
rect 20111 8724 20116 8780
rect 20050 8700 20116 8724
rect 20050 8644 20055 8700
rect 20111 8644 20116 8700
rect 20050 8620 20116 8644
rect 20050 8564 20055 8620
rect 20111 8564 20116 8620
rect 20050 8540 20116 8564
rect 20050 8484 20055 8540
rect 20111 8484 20116 8540
rect 20050 8460 20116 8484
rect 20050 8404 20055 8460
rect 20111 8404 20116 8460
rect 20050 8366 20116 8404
rect 18400 8361 20116 8366
rect 18400 8305 18498 8361
rect 18554 8305 18578 8361
rect 18634 8305 18658 8361
rect 18714 8305 18738 8361
rect 18794 8305 18818 8361
rect 18874 8305 18898 8361
rect 18954 8305 18978 8361
rect 19034 8305 19058 8361
rect 19114 8305 19138 8361
rect 19194 8305 19322 8361
rect 19378 8305 19402 8361
rect 19458 8305 19482 8361
rect 19538 8305 19562 8361
rect 19618 8305 19642 8361
rect 19698 8305 19722 8361
rect 19778 8305 19802 8361
rect 19858 8305 19882 8361
rect 19938 8305 19962 8361
rect 20018 8305 20116 8361
rect 18400 8300 20116 8305
rect 17692 7109 17758 7118
rect 11820 7050 12500 7100
rect 11820 6990 11860 7050
rect 12480 6990 12500 7050
rect 11820 6970 12500 6990
rect 12980 7050 13240 7100
rect 12980 6990 13000 7050
rect 13220 6990 13240 7050
rect 12980 6970 13240 6990
rect 13540 7050 13800 7100
rect 13540 6990 13560 7050
rect 13780 6990 13800 7050
rect 13540 6970 13800 6990
rect 14100 7050 14350 7100
rect 14100 6990 14140 7050
rect 14320 6990 14350 7050
rect 14100 6950 14350 6990
rect 14650 7050 15500 7100
rect 14650 6970 14680 7050
rect 15480 6970 15500 7050
rect 17692 7053 17697 7109
rect 17753 7053 17758 7109
rect 17692 7030 17758 7053
rect 17864 7109 17930 7118
rect 17864 7053 17869 7109
rect 17925 7053 17930 7109
rect 17864 7030 17930 7053
rect 18036 7109 18102 7118
rect 18036 7053 18041 7109
rect 18097 7053 18102 7109
rect 18036 7030 18102 7053
rect 18208 7109 18274 7118
rect 18208 7053 18213 7109
rect 18269 7053 18274 7109
rect 18208 7030 18274 7053
rect 18380 7109 18446 7118
rect 18380 7053 18385 7109
rect 18441 7053 18446 7109
rect 18380 7030 18446 7053
rect 18552 7109 18618 7118
rect 18552 7053 18557 7109
rect 18613 7053 18618 7109
rect 18552 7030 18618 7053
rect 18724 7109 18790 7118
rect 18724 7053 18729 7109
rect 18785 7053 18790 7109
rect 18724 7030 18790 7053
rect 18896 7109 18962 7118
rect 18896 7053 18901 7109
rect 18957 7053 18962 7109
rect 18896 7030 18962 7053
rect 19068 7109 19134 7118
rect 19068 7053 19073 7109
rect 19129 7053 19134 7109
rect 19068 7030 19134 7053
rect 19240 7109 19306 7118
rect 19240 7053 19245 7109
rect 19301 7053 19306 7109
rect 19240 7030 19306 7053
rect 19412 7109 19478 7118
rect 19412 7053 19417 7109
rect 19473 7053 19478 7109
rect 19412 7030 19478 7053
rect 19584 7109 19650 7118
rect 19584 7053 19589 7109
rect 19645 7053 19650 7109
rect 19584 7030 19650 7053
rect 19756 7109 19822 7118
rect 19756 7053 19761 7109
rect 19817 7053 19822 7109
rect 19756 7030 19822 7053
rect 19928 7109 19994 7118
rect 19928 7053 19933 7109
rect 19989 7053 19994 7109
rect 19928 7030 19994 7053
rect 14650 6950 15500 6970
rect 17170 7029 19994 7030
rect 17170 7000 17697 7029
rect 17170 6990 17200 7000
rect 17300 6990 17697 7000
rect 17170 6870 17180 6990
rect 17330 6973 17697 6990
rect 17753 6973 17869 7029
rect 17925 6973 18041 7029
rect 18097 6973 18213 7029
rect 18269 6973 18385 7029
rect 18441 6973 18557 7029
rect 18613 6973 18729 7029
rect 18785 6973 18901 7029
rect 18957 6973 19073 7029
rect 19129 6973 19245 7029
rect 19301 6973 19417 7029
rect 19473 6973 19589 7029
rect 19645 6973 19761 7029
rect 19817 6973 19933 7029
rect 19989 6973 19994 7029
rect 17330 6970 19994 6973
rect 17330 6910 17450 6970
rect 17692 6964 17930 6970
rect 18036 6964 18274 6970
rect 18380 6964 18618 6970
rect 18724 6964 18962 6970
rect 19068 6964 19306 6970
rect 19412 6964 19650 6970
rect 19756 6964 19994 6970
rect 17330 6870 17340 6910
rect 17170 6470 17200 6870
rect 17300 6470 17340 6870
rect 17170 6370 17180 6470
rect 17330 6370 17340 6470
rect 17170 6360 17340 6370
rect 17430 6820 17600 6830
rect 17430 6720 17440 6820
rect 17590 6720 17600 6820
rect 17430 6330 17460 6720
rect 17560 6330 17600 6720
rect 15650 6250 16000 6300
rect 17430 6250 17440 6330
rect 15650 5950 15700 6250
rect 11450 5730 15700 5950
rect 11450 5670 11620 5730
rect 15680 5700 15700 5730
rect 15950 5700 16000 6250
rect 17410 6230 17440 6250
rect 17590 6230 17600 6330
rect 17410 6220 17460 6230
rect 17340 6200 17460 6220
rect 17560 6220 17600 6230
rect 17674 6220 17912 6226
rect 18018 6220 18256 6226
rect 18362 6220 18600 6226
rect 18706 6220 18944 6226
rect 19050 6220 19288 6226
rect 19394 6220 19632 6226
rect 19738 6220 19976 6226
rect 17560 6217 19976 6220
rect 17560 6200 17679 6217
rect 17340 6161 17679 6200
rect 17735 6161 17851 6217
rect 17907 6161 18023 6217
rect 18079 6161 18195 6217
rect 18251 6161 18367 6217
rect 18423 6161 18539 6217
rect 18595 6161 18711 6217
rect 18767 6161 18883 6217
rect 18939 6161 19055 6217
rect 19111 6161 19227 6217
rect 19283 6161 19399 6217
rect 19455 6161 19571 6217
rect 19627 6161 19743 6217
rect 19799 6161 19915 6217
rect 19971 6161 19976 6217
rect 17340 6160 19976 6161
rect 17674 6137 17740 6160
rect 17674 6081 17679 6137
rect 17735 6081 17740 6137
rect 17674 6072 17740 6081
rect 17846 6137 17912 6160
rect 17846 6081 17851 6137
rect 17907 6081 17912 6137
rect 17846 6072 17912 6081
rect 18018 6137 18084 6160
rect 18018 6081 18023 6137
rect 18079 6081 18084 6137
rect 18018 6072 18084 6081
rect 18190 6137 18256 6160
rect 18190 6081 18195 6137
rect 18251 6081 18256 6137
rect 18190 6072 18256 6081
rect 18362 6137 18428 6160
rect 18362 6081 18367 6137
rect 18423 6081 18428 6137
rect 18362 6072 18428 6081
rect 18534 6137 18600 6160
rect 18534 6081 18539 6137
rect 18595 6081 18600 6137
rect 18534 6072 18600 6081
rect 18706 6137 18772 6160
rect 18706 6081 18711 6137
rect 18767 6081 18772 6137
rect 18706 6072 18772 6081
rect 18878 6137 18944 6160
rect 18878 6081 18883 6137
rect 18939 6081 18944 6137
rect 18878 6072 18944 6081
rect 19050 6137 19116 6160
rect 19050 6081 19055 6137
rect 19111 6081 19116 6137
rect 19050 6072 19116 6081
rect 19222 6137 19288 6160
rect 19222 6081 19227 6137
rect 19283 6081 19288 6137
rect 19222 6072 19288 6081
rect 19394 6137 19460 6160
rect 19394 6081 19399 6137
rect 19455 6081 19460 6137
rect 19394 6072 19460 6081
rect 19566 6137 19632 6160
rect 19566 6081 19571 6137
rect 19627 6081 19632 6137
rect 19566 6072 19632 6081
rect 19738 6137 19804 6160
rect 19738 6081 19743 6137
rect 19799 6081 19804 6137
rect 19738 6072 19804 6081
rect 19910 6137 19976 6160
rect 19910 6081 19915 6137
rect 19971 6081 19976 6137
rect 19910 6072 19976 6081
rect 15680 5670 16000 5700
rect 11450 5650 16000 5670
rect 12400 5580 12680 5590
rect 12960 5580 13240 5590
rect 12400 5520 12410 5580
rect 12670 5520 12680 5580
rect 12400 5480 12680 5520
rect 11900 5420 12300 5460
rect 11900 5300 11920 5420
rect 12280 5300 12300 5420
rect 11900 5200 12300 5300
rect 12500 2860 12680 5480
rect 12860 5520 12970 5580
rect 13230 5520 13240 5580
rect 12860 5510 13240 5520
rect 13540 5580 13820 5590
rect 14100 5580 14380 5590
rect 13540 5520 13550 5580
rect 13810 5520 13880 5580
rect 13540 5510 13880 5520
rect 12860 5480 13140 5510
rect 12860 2860 13040 5480
rect 13200 5420 13600 5440
rect 13200 5300 13220 5420
rect 13580 5300 13600 5420
rect 13200 5200 13600 5300
rect 13700 2860 13880 5510
rect 14060 5520 14110 5580
rect 14370 5520 14380 5580
rect 14060 5510 14380 5520
rect 14680 5580 14960 5590
rect 14680 5520 14690 5580
rect 14950 5520 14980 5580
rect 14680 5510 14980 5520
rect 14060 2860 14240 5510
rect 14300 5420 14700 5440
rect 14300 5300 14320 5420
rect 14680 5300 14700 5420
rect 14300 5200 14700 5300
rect 14800 2860 14980 5510
rect 15500 5440 15960 5460
rect 15500 5300 15540 5440
rect 15880 5300 15960 5440
rect 15500 5200 15960 5300
rect 16550 4813 18266 4818
rect 16550 4757 16648 4813
rect 16704 4757 16728 4813
rect 16784 4757 16808 4813
rect 16864 4757 16888 4813
rect 16944 4757 16968 4813
rect 17024 4757 17048 4813
rect 17104 4757 17128 4813
rect 17184 4757 17208 4813
rect 17264 4757 17288 4813
rect 17344 4757 17472 4813
rect 17528 4757 17552 4813
rect 17608 4757 17632 4813
rect 17688 4757 17712 4813
rect 17768 4757 17792 4813
rect 17848 4757 17872 4813
rect 17928 4757 17952 4813
rect 18008 4757 18032 4813
rect 18088 4757 18112 4813
rect 18168 4757 18266 4813
rect 16550 4752 18266 4757
rect 16550 4714 16616 4752
rect 16550 4658 16555 4714
rect 16611 4658 16616 4714
rect 16550 4634 16616 4658
rect 16550 4578 16555 4634
rect 16611 4578 16616 4634
rect 16550 4554 16616 4578
rect 16550 4498 16555 4554
rect 16611 4498 16616 4554
rect 16550 4474 16616 4498
rect 16550 4418 16555 4474
rect 16611 4418 16616 4474
rect 16550 4394 16616 4418
rect 16550 4338 16555 4394
rect 16611 4338 16616 4394
rect 16550 4314 16616 4338
rect 16550 4258 16555 4314
rect 16611 4258 16616 4314
rect 16550 4234 16616 4258
rect 16550 4178 16555 4234
rect 16611 4178 16616 4234
rect 16550 4154 16616 4178
rect 16550 4098 16555 4154
rect 16611 4098 16616 4154
rect 16550 3970 16616 4098
rect 16550 3914 16555 3970
rect 16611 3914 16616 3970
rect 16550 3890 16616 3914
rect 16550 3834 16555 3890
rect 16611 3834 16616 3890
rect 16550 3810 16616 3834
rect 16550 3754 16555 3810
rect 16611 3754 16616 3810
rect 16550 3730 16616 3754
rect 16550 3674 16555 3730
rect 16611 3674 16616 3730
rect 16550 3650 16616 3674
rect 16550 3594 16555 3650
rect 16611 3594 16616 3650
rect 16550 3570 16616 3594
rect 16550 3514 16555 3570
rect 16611 3514 16616 3570
rect 16550 3490 16616 3514
rect 16550 3434 16555 3490
rect 16611 3434 16616 3490
rect 16550 3410 16616 3434
rect 16550 3354 16555 3410
rect 16611 3354 16616 3410
rect 16676 4067 16754 4692
rect 16814 4127 16892 4752
rect 16952 4067 17030 4692
rect 17090 4127 17168 4752
rect 17228 4067 17306 4692
rect 17369 4127 17447 4752
rect 17510 4067 17588 4692
rect 17648 4127 17726 4752
rect 17786 4067 17864 4692
rect 17924 4127 18002 4752
rect 18200 4714 18266 4752
rect 18062 4067 18140 4692
rect 18130 4005 18140 4067
rect 16676 3376 16754 3476
rect 16550 3316 16616 3354
rect 16814 3316 16892 3941
rect 16952 3376 17030 3476
rect 17090 3316 17168 3941
rect 17228 3376 17306 3476
rect 17369 3316 17447 3941
rect 17510 3376 17588 3476
rect 17648 3316 17726 3941
rect 17786 3376 17864 3476
rect 17924 3316 18002 3941
rect 18062 3376 18140 3475
rect 18200 4658 18205 4714
rect 18261 4658 18266 4714
rect 18200 4634 18266 4658
rect 18200 4578 18205 4634
rect 18261 4578 18266 4634
rect 18200 4554 18266 4578
rect 18200 4498 18205 4554
rect 18261 4498 18266 4554
rect 18200 4474 18266 4498
rect 18200 4418 18205 4474
rect 18261 4418 18266 4474
rect 18200 4394 18266 4418
rect 18200 4338 18205 4394
rect 18261 4338 18266 4394
rect 18200 4314 18266 4338
rect 18200 4258 18205 4314
rect 18261 4258 18266 4314
rect 18200 4234 18266 4258
rect 18200 4178 18205 4234
rect 18261 4178 18266 4234
rect 18200 4154 18266 4178
rect 18200 4098 18205 4154
rect 18261 4098 18266 4154
rect 18200 3970 18266 4098
rect 18200 3914 18205 3970
rect 18261 3914 18266 3970
rect 18200 3890 18266 3914
rect 18200 3834 18205 3890
rect 18261 3834 18266 3890
rect 18200 3810 18266 3834
rect 18200 3754 18205 3810
rect 18261 3754 18266 3810
rect 18200 3730 18266 3754
rect 18200 3674 18205 3730
rect 18261 3674 18266 3730
rect 18200 3650 18266 3674
rect 18200 3594 18205 3650
rect 18261 3594 18266 3650
rect 18200 3570 18266 3594
rect 18200 3514 18205 3570
rect 18261 3514 18266 3570
rect 18200 3490 18266 3514
rect 18200 3434 18205 3490
rect 18261 3434 18266 3490
rect 18200 3410 18266 3434
rect 18200 3354 18205 3410
rect 18261 3354 18266 3410
rect 18200 3316 18266 3354
rect 16550 3311 18266 3316
rect 16550 3255 16648 3311
rect 16704 3255 16728 3311
rect 16784 3255 16808 3311
rect 16864 3255 16888 3311
rect 16944 3255 16968 3311
rect 17024 3255 17048 3311
rect 17104 3255 17128 3311
rect 17184 3255 17208 3311
rect 17264 3255 17288 3311
rect 17344 3255 17472 3311
rect 17528 3255 17552 3311
rect 17608 3255 17632 3311
rect 17688 3255 17712 3311
rect 17768 3255 17792 3311
rect 17848 3255 17872 3311
rect 17928 3255 17952 3311
rect 18008 3255 18032 3311
rect 18088 3255 18112 3311
rect 18168 3255 18266 3311
rect 16550 3250 18266 3255
rect 18400 4813 20116 4818
rect 18400 4757 18498 4813
rect 18554 4757 18578 4813
rect 18634 4757 18658 4813
rect 18714 4757 18738 4813
rect 18794 4757 18818 4813
rect 18874 4757 18898 4813
rect 18954 4757 18978 4813
rect 19034 4757 19058 4813
rect 19114 4757 19138 4813
rect 19194 4757 19322 4813
rect 19378 4757 19402 4813
rect 19458 4757 19482 4813
rect 19538 4757 19562 4813
rect 19618 4757 19642 4813
rect 19698 4757 19722 4813
rect 19778 4757 19802 4813
rect 19858 4757 19882 4813
rect 19938 4757 19962 4813
rect 20018 4757 20116 4813
rect 18400 4752 20116 4757
rect 18400 4714 18466 4752
rect 18400 4658 18405 4714
rect 18461 4658 18466 4714
rect 18400 4634 18466 4658
rect 18400 4578 18405 4634
rect 18461 4578 18466 4634
rect 18400 4554 18466 4578
rect 18400 4498 18405 4554
rect 18461 4498 18466 4554
rect 18400 4474 18466 4498
rect 18400 4418 18405 4474
rect 18461 4418 18466 4474
rect 18400 4394 18466 4418
rect 18400 4338 18405 4394
rect 18461 4338 18466 4394
rect 18400 4314 18466 4338
rect 18400 4258 18405 4314
rect 18461 4258 18466 4314
rect 18400 4234 18466 4258
rect 18400 4178 18405 4234
rect 18461 4178 18466 4234
rect 18400 4154 18466 4178
rect 18400 4098 18405 4154
rect 18461 4098 18466 4154
rect 18400 3970 18466 4098
rect 18400 3914 18405 3970
rect 18461 3914 18466 3970
rect 18400 3890 18466 3914
rect 18400 3834 18405 3890
rect 18461 3834 18466 3890
rect 18400 3810 18466 3834
rect 18400 3754 18405 3810
rect 18461 3754 18466 3810
rect 18400 3730 18466 3754
rect 18400 3674 18405 3730
rect 18461 3674 18466 3730
rect 18400 3650 18466 3674
rect 18400 3594 18405 3650
rect 18461 3594 18466 3650
rect 18400 3570 18466 3594
rect 18400 3514 18405 3570
rect 18461 3514 18466 3570
rect 18400 3490 18466 3514
rect 18400 3434 18405 3490
rect 18461 3434 18466 3490
rect 18400 3410 18466 3434
rect 18400 3354 18405 3410
rect 18461 3354 18466 3410
rect 18526 4067 18604 4692
rect 18664 4127 18742 4752
rect 18802 4067 18880 4692
rect 18940 4127 19018 4752
rect 19078 4067 19156 4692
rect 19219 4127 19297 4752
rect 19360 4067 19438 4692
rect 19498 4127 19576 4752
rect 19636 4067 19714 4692
rect 19774 4127 19852 4752
rect 20050 4714 20116 4752
rect 19912 4067 19990 4692
rect 19713 4062 19990 4067
rect 19766 4006 19790 4062
rect 19846 4006 19870 4062
rect 19926 4006 19990 4062
rect 19713 4005 19990 4006
rect 19714 4001 19990 4005
rect 18526 3376 18604 3475
rect 18400 3316 18466 3354
rect 18664 3316 18742 3941
rect 18802 3376 18880 3475
rect 18940 3316 19018 3941
rect 19078 3376 19156 3475
rect 19219 3316 19297 3941
rect 19360 3376 19438 3475
rect 19498 3316 19576 3941
rect 19636 3376 19714 3475
rect 19774 3316 19852 3941
rect 19912 3376 19990 4001
rect 20050 4658 20055 4714
rect 20111 4658 20116 4714
rect 20050 4634 20116 4658
rect 20050 4578 20055 4634
rect 20111 4578 20116 4634
rect 20050 4554 20116 4578
rect 20050 4498 20055 4554
rect 20111 4498 20116 4554
rect 20050 4474 20116 4498
rect 20050 4418 20055 4474
rect 20111 4418 20116 4474
rect 20050 4394 20116 4418
rect 20050 4338 20055 4394
rect 20111 4338 20116 4394
rect 20050 4314 20116 4338
rect 20050 4258 20055 4314
rect 20111 4258 20116 4314
rect 20050 4234 20116 4258
rect 20050 4178 20055 4234
rect 20111 4178 20116 4234
rect 20050 4154 20116 4178
rect 20050 4098 20055 4154
rect 20111 4098 20116 4154
rect 20050 3970 20116 4098
rect 20050 3914 20055 3970
rect 20111 3914 20116 3970
rect 20050 3890 20116 3914
rect 20050 3834 20055 3890
rect 20111 3834 20116 3890
rect 20050 3810 20116 3834
rect 20050 3754 20055 3810
rect 20111 3754 20116 3810
rect 20050 3730 20116 3754
rect 20050 3674 20055 3730
rect 20111 3674 20116 3730
rect 20050 3650 20116 3674
rect 20050 3594 20055 3650
rect 20111 3594 20116 3650
rect 20050 3570 20116 3594
rect 20050 3514 20055 3570
rect 20111 3514 20116 3570
rect 20050 3490 20116 3514
rect 20050 3434 20055 3490
rect 20111 3434 20116 3490
rect 20050 3410 20116 3434
rect 20050 3354 20055 3410
rect 20111 3354 20116 3410
rect 20050 3316 20116 3354
rect 18400 3311 20116 3316
rect 18400 3255 18498 3311
rect 18554 3255 18578 3311
rect 18634 3255 18658 3311
rect 18714 3255 18738 3311
rect 18794 3255 18818 3311
rect 18874 3255 18898 3311
rect 18954 3255 18978 3311
rect 19034 3255 19058 3311
rect 19114 3255 19138 3311
rect 19194 3255 19322 3311
rect 19378 3255 19402 3311
rect 19458 3255 19482 3311
rect 19538 3255 19562 3311
rect 19618 3255 19642 3311
rect 19698 3255 19722 3311
rect 19778 3255 19802 3311
rect 19858 3255 19882 3311
rect 19938 3255 19962 3311
rect 20018 3255 20116 3311
rect 18400 3250 20116 3255
<< via3 >>
rect 15400 9900 16300 10700
rect 16953 9117 17030 9642
rect 17228 9117 17305 9643
rect 17510 9117 17587 9643
rect 17786 9117 17863 9643
rect 18062 9117 18140 9643
rect 16811 9112 18140 9117
rect 16811 9056 16820 9112
rect 16820 9056 16876 9112
rect 16876 9056 16900 9112
rect 16900 9056 16956 9112
rect 16956 9056 16980 9112
rect 16980 9056 17036 9112
rect 17036 9056 17060 9112
rect 17060 9056 17116 9112
rect 17116 9056 17140 9112
rect 17140 9056 17196 9112
rect 17196 9056 17220 9112
rect 17220 9056 17276 9112
rect 17276 9056 17300 9112
rect 17300 9056 17356 9112
rect 17356 9056 17380 9112
rect 17380 9056 17436 9112
rect 17436 9056 17460 9112
rect 17460 9056 17516 9112
rect 17516 9056 17540 9112
rect 17540 9056 17596 9112
rect 17596 9056 17620 9112
rect 17620 9056 17676 9112
rect 17676 9056 17700 9112
rect 17700 9056 17756 9112
rect 17756 9056 17780 9112
rect 17780 9056 17836 9112
rect 17836 9056 17860 9112
rect 17860 9056 17916 9112
rect 17916 9056 17940 9112
rect 17940 9056 17996 9112
rect 17996 9056 18020 9112
rect 18020 9056 18076 9112
rect 18076 9056 18140 9112
rect 16811 9051 18140 9056
rect 18526 9117 18604 9642
rect 18802 9117 18880 9642
rect 19078 9117 19156 9642
rect 19360 9117 19438 9642
rect 19636 9117 19714 9642
rect 18526 9112 19714 9117
rect 18526 9056 18590 9112
rect 18590 9056 18646 9112
rect 18646 9056 18670 9112
rect 18670 9056 18726 9112
rect 18726 9056 18750 9112
rect 18750 9056 18806 9112
rect 18806 9056 18830 9112
rect 18830 9056 18886 9112
rect 18886 9056 18910 9112
rect 18910 9056 18966 9112
rect 18966 9056 18990 9112
rect 18990 9056 19046 9112
rect 19046 9056 19070 9112
rect 19070 9056 19126 9112
rect 19126 9056 19150 9112
rect 19150 9056 19206 9112
rect 19206 9056 19230 9112
rect 19230 9056 19286 9112
rect 19286 9056 19310 9112
rect 19310 9056 19366 9112
rect 19366 9056 19390 9112
rect 19390 9056 19446 9112
rect 19446 9056 19470 9112
rect 19470 9056 19526 9112
rect 19526 9056 19550 9112
rect 19550 9056 19606 9112
rect 19606 9056 19630 9112
rect 19630 9056 19686 9112
rect 19686 9056 19710 9112
rect 19710 9056 19714 9112
rect 18526 9051 19714 9056
rect 17200 6990 17300 7000
rect 17200 6870 17300 6990
rect 17200 6470 17300 6870
rect 17200 6450 17300 6470
rect 17460 6720 17560 6760
rect 17460 6330 17560 6720
rect 15700 5700 15950 6250
rect 17460 6230 17560 6330
rect 17460 6200 17560 6230
rect 11920 5300 12280 5420
rect 13220 5300 13580 5420
rect 14320 5300 14680 5420
rect 15540 5300 15880 5440
rect 16676 4062 18130 4067
rect 16676 4006 16740 4062
rect 16740 4006 16796 4062
rect 16796 4006 16820 4062
rect 16820 4006 16876 4062
rect 16876 4006 16900 4062
rect 16900 4006 16956 4062
rect 16956 4006 16980 4062
rect 16980 4006 17036 4062
rect 17036 4006 17060 4062
rect 17060 4006 17116 4062
rect 17116 4006 17140 4062
rect 17140 4006 17196 4062
rect 17196 4006 17220 4062
rect 17220 4006 17276 4062
rect 17276 4006 17300 4062
rect 17300 4006 17356 4062
rect 17356 4006 17380 4062
rect 17380 4006 17436 4062
rect 17436 4006 17460 4062
rect 17460 4006 17516 4062
rect 17516 4006 17540 4062
rect 17540 4006 17596 4062
rect 17596 4006 17620 4062
rect 17620 4006 17676 4062
rect 17676 4006 17700 4062
rect 17700 4006 17756 4062
rect 17756 4006 17780 4062
rect 17780 4006 17836 4062
rect 17836 4006 17860 4062
rect 17860 4006 17916 4062
rect 17916 4006 17940 4062
rect 17940 4006 17996 4062
rect 17996 4006 18020 4062
rect 18020 4006 18076 4062
rect 18076 4006 18130 4062
rect 16676 4005 18130 4006
rect 16676 4001 18140 4005
rect 16676 3476 16754 4001
rect 16952 3476 17030 4001
rect 17228 3476 17306 4001
rect 17510 3476 17588 4001
rect 17786 3476 17864 4001
rect 18062 3475 18140 4001
rect 18526 4062 19713 4067
rect 18526 4006 18590 4062
rect 18590 4006 18646 4062
rect 18646 4006 18670 4062
rect 18670 4006 18726 4062
rect 18726 4006 18750 4062
rect 18750 4006 18806 4062
rect 18806 4006 18830 4062
rect 18830 4006 18886 4062
rect 18886 4006 18910 4062
rect 18910 4006 18966 4062
rect 18966 4006 18990 4062
rect 18990 4006 19046 4062
rect 19046 4006 19070 4062
rect 19070 4006 19126 4062
rect 19126 4006 19150 4062
rect 19150 4006 19206 4062
rect 19206 4006 19230 4062
rect 19230 4006 19286 4062
rect 19286 4006 19310 4062
rect 19310 4006 19366 4062
rect 19366 4006 19390 4062
rect 19390 4006 19446 4062
rect 19446 4006 19470 4062
rect 19470 4006 19526 4062
rect 19526 4006 19550 4062
rect 19550 4006 19606 4062
rect 19606 4006 19630 4062
rect 19630 4006 19686 4062
rect 19686 4006 19710 4062
rect 19710 4006 19713 4062
rect 18526 4005 19713 4006
rect 18526 4001 19714 4005
rect 18526 3475 18604 4001
rect 18802 3475 18880 4001
rect 19078 3475 19156 4001
rect 19360 3475 19438 4001
rect 19636 3475 19714 4001
<< mimcap >>
rect 11650 9100 12450 9150
rect 11650 7200 11700 9100
rect 12400 7200 12450 9100
rect 11650 7150 12450 7200
rect 12800 9100 13200 9150
rect 12800 7200 12850 9100
rect 13150 7200 13200 9100
rect 12800 7150 13200 7200
rect 13550 9100 13750 9150
rect 13550 7200 13600 9100
rect 13700 7200 13750 9100
rect 14650 9100 16250 9150
rect 13550 7150 13750 7200
rect 14100 8100 14300 8150
rect 14100 7200 14150 8100
rect 14250 7200 14300 8100
rect 14100 7150 14300 7200
rect 14650 7200 14700 9100
rect 16200 7200 16250 9100
rect 14650 7150 16250 7200
<< mimcapcontact >>
rect 11700 7200 12400 9100
rect 12850 7200 13150 9100
rect 13600 7200 13700 9100
rect 14150 7200 14250 8100
rect 14700 7200 16200 9100
<< metal4 >>
rect 21400 16400 25400 16600
rect 21400 13400 21600 16400
rect 21000 12400 21600 13400
rect 25200 12400 25400 16400
rect 17700 11400 18500 11800
rect 15700 10800 18500 11400
rect 10000 10700 18500 10800
rect 10000 10600 15400 10700
rect 10100 9900 15400 10600
rect 16300 10000 18500 10700
rect 16300 9900 16500 10000
rect 10100 9600 16500 9900
rect 16700 9700 19900 9800
rect 10100 8300 11100 9600
rect 16700 9300 16800 9700
rect 19800 9300 19900 9700
rect 21000 9500 25400 12400
rect 11600 9100 12500 9200
rect 10100 6400 10700 8300
rect 11000 7400 11400 8000
rect 11600 7400 11700 9100
rect 11000 7200 11700 7400
rect 12400 7400 12500 9100
rect 12750 9100 13250 9200
rect 12750 7400 12850 9100
rect 12400 7200 12850 7400
rect 13150 7400 13250 9100
rect 13500 9100 13800 9200
rect 13500 7400 13600 9100
rect 13150 7200 13600 7400
rect 13700 7400 13800 9100
rect 14600 9100 16300 9200
rect 14050 8100 14350 8200
rect 14050 7400 14150 8100
rect 13700 7200 14150 7400
rect 14250 7400 14350 8100
rect 14600 7400 14700 9100
rect 14250 7200 14700 7400
rect 16200 7400 16300 9100
rect 16700 9117 16953 9300
rect 17030 9117 17228 9300
rect 17305 9117 17510 9300
rect 17587 9117 17786 9300
rect 17863 9117 18062 9300
rect 16700 9051 16811 9117
rect 18140 9051 18526 9300
rect 18604 9117 18802 9300
rect 18880 9117 19078 9300
rect 19156 9117 19360 9300
rect 19438 9117 19636 9300
rect 19714 9051 19900 9300
rect 16700 9000 19900 9051
rect 20300 8600 25400 9500
rect 17100 8200 25400 8600
rect 17100 8000 21100 8200
rect 17200 7800 21100 8000
rect 17200 7400 17800 7800
rect 16200 7200 17800 7400
rect 11000 7100 17800 7200
rect 11000 6700 11400 7100
rect 17150 7000 17350 7100
rect 17150 6450 17200 7000
rect 17300 6450 17350 7000
rect 17150 6400 17350 6450
rect 17440 6760 17620 6800
rect 10100 3600 11100 6400
rect 15650 6250 16000 6300
rect 15650 5700 15700 6250
rect 15950 6050 16000 6250
rect 17440 6200 17460 6760
rect 17560 6200 17620 6760
rect 17440 6050 17620 6200
rect 15950 5750 17620 6050
rect 15950 5700 17800 5750
rect 15650 5650 17800 5700
rect 15500 5440 16100 5460
rect 11900 5420 12300 5440
rect 11900 5300 11920 5420
rect 12280 5300 12300 5420
rect 11900 3600 12300 5300
rect 13200 5420 13600 5440
rect 13200 5300 13220 5420
rect 13580 5300 13600 5420
rect 13200 3600 13600 5300
rect 14300 5420 14700 5440
rect 14300 5300 14320 5420
rect 14680 5300 14700 5420
rect 14300 3600 14700 5300
rect 15500 5300 15540 5440
rect 15880 5300 16100 5440
rect 15500 5200 16100 5300
rect 17200 5400 17800 5650
rect 17200 5200 21100 5400
rect 15500 3600 16300 5200
rect 17100 4800 21100 5200
rect 17100 4600 25400 4800
rect 20300 4200 25400 4600
rect 10100 3100 16300 3600
rect 16500 4067 19900 4100
rect 16500 3800 16676 4067
rect 18130 4005 18526 4067
rect 19713 4005 19900 4067
rect 16754 3800 16952 4001
rect 17030 3800 17228 4001
rect 17306 3800 17510 4001
rect 17588 3800 17786 4001
rect 17864 3800 18062 4001
rect 18140 3800 18526 4005
rect 18604 3800 18802 4001
rect 18880 3800 19078 4001
rect 19156 3800 19360 4001
rect 19438 3800 19636 4001
rect 19714 3800 19900 4005
rect 16500 3400 16600 3800
rect 19800 3400 19900 3800
rect 20300 4088 34600 4200
rect 20300 3600 30712 4088
rect 16500 3300 19900 3400
rect 10100 3000 18500 3100
rect 15500 1800 18500 3000
rect 17700 1400 18500 1800
rect 21000 312 30712 3600
rect 34488 312 34600 4088
rect 21000 200 34600 312
<< via4 >>
rect 21600 12400 25200 16400
rect 16800 9643 19800 9700
rect 16800 9642 17228 9643
rect 16800 9300 16953 9642
rect 16953 9300 17030 9642
rect 17030 9300 17228 9642
rect 17228 9300 17305 9643
rect 17305 9300 17510 9643
rect 17510 9300 17587 9643
rect 17587 9300 17786 9643
rect 17786 9300 17863 9643
rect 17863 9300 18062 9643
rect 18062 9300 18140 9643
rect 18140 9642 19800 9643
rect 18140 9300 18526 9642
rect 18526 9300 18604 9642
rect 18604 9300 18802 9642
rect 18802 9300 18880 9642
rect 18880 9300 19078 9642
rect 19078 9300 19156 9642
rect 19156 9300 19360 9642
rect 19360 9300 19438 9642
rect 19438 9300 19636 9642
rect 19636 9300 19714 9642
rect 19714 9300 19800 9642
rect 16600 3476 16676 3800
rect 16676 3476 16754 3800
rect 16754 3476 16952 3800
rect 16952 3476 17030 3800
rect 17030 3476 17228 3800
rect 17228 3476 17306 3800
rect 17306 3476 17510 3800
rect 17510 3476 17588 3800
rect 17588 3476 17786 3800
rect 17786 3476 17864 3800
rect 17864 3476 18062 3800
rect 16600 3475 18062 3476
rect 18062 3475 18140 3800
rect 18140 3475 18526 3800
rect 18526 3475 18604 3800
rect 18604 3475 18802 3800
rect 18802 3475 18880 3800
rect 18880 3475 19078 3800
rect 19078 3475 19156 3800
rect 19156 3475 19360 3800
rect 19360 3475 19438 3800
rect 19438 3475 19636 3800
rect 19636 3475 19714 3800
rect 19714 3475 19800 3800
rect 16600 3400 19800 3475
rect 30712 312 34488 4088
<< metal5 >>
tri 32220 27200 36220 31200 se
rect 36220 27200 57580 31200
tri 57580 27200 61580 31200 sw
tri 30000 24980 32220 27200 se
rect 32220 26600 37277 27200
tri 37277 26600 37877 27200 nw
tri 55923 26600 56523 27200 ne
rect 56523 26600 61580 27200
rect 32220 25751 36428 26600
tri 36428 25751 37277 26600 nw
tri 37277 25751 38126 26600 se
rect 38126 25751 55674 26600
tri 55674 25751 56523 26600 sw
tri 56523 25751 57372 26600 ne
rect 57372 25751 61580 26600
rect 32220 24980 35579 25751
tri 28469 23449 30000 24980 se
rect 30000 24902 35579 24980
tri 35579 24902 36428 25751 nw
tri 36428 24902 37277 25751 se
rect 37277 24902 56523 25751
tri 56523 24902 57372 25751 sw
tri 57372 24902 58221 25751 ne
rect 58221 24902 61580 25751
rect 30000 24298 34975 24902
tri 34975 24298 35579 24902 nw
tri 35824 24298 36428 24902 se
rect 36428 24298 57372 24902
tri 57372 24298 57976 24902 sw
tri 58221 24298 58825 24902 ne
rect 58825 24298 61580 24902
rect 30000 23449 34126 24298
tri 34126 23449 34975 24298 nw
tri 34975 23449 35824 24298 se
rect 35824 23449 57976 24298
tri 57976 23449 58825 24298 sw
tri 58825 23449 59674 24298 ne
rect 59674 23449 61580 24298
tri 25400 20380 28469 23449 se
rect 28469 22600 33277 23449
tri 33277 22600 34126 23449 nw
tri 34126 22600 34975 23449 se
rect 34975 22600 58825 23449
tri 58825 22600 59674 23449 sw
tri 59674 22600 60523 23449 ne
rect 60523 22600 61580 23449
tri 61580 22600 66180 27200 sw
rect 28469 21751 32428 22600
tri 32428 21751 33277 22600 nw
tri 33277 21751 34126 22600 se
rect 28469 20902 31579 21751
tri 31579 20902 32428 21751 nw
tri 32428 20902 33277 21751 se
rect 33277 20902 34126 21751
rect 28469 20380 30849 20902
tri 24343 19323 25400 20380 se
rect 25400 20172 30849 20380
tri 30849 20172 31579 20902 nw
tri 31698 20172 32428 20902 se
rect 32428 20172 34126 20902
rect 25400 19323 30000 20172
tri 30000 19323 30849 20172 nw
tri 30849 19323 31698 20172 se
rect 31698 19323 34126 20172
tri 21420 16400 24343 19323 se
rect 24343 18474 29151 19323
tri 29151 18474 30000 19323 nw
tri 30000 18474 30849 19323 se
rect 30849 18474 34126 19323
rect 24343 17625 28302 18474
tri 28302 17625 29151 18474 nw
tri 29151 17625 30000 18474 se
rect 30000 17625 34126 18474
rect 24343 16943 27620 17625
tri 27620 16943 28302 17625 nw
tri 28469 16943 29151 17625 se
rect 29151 16943 34126 17625
tri 34126 16943 39783 22600 nw
tri 54017 16943 59674 22600 ne
tri 59674 21751 60523 22600 sw
tri 60523 21751 61372 22600 ne
rect 61372 21751 66180 22600
rect 59674 20902 60523 21751
tri 60523 20902 61372 21751 sw
tri 61372 20902 62221 21751 ne
rect 62221 20902 66180 21751
rect 59674 20172 61372 20902
tri 61372 20172 62102 20902 sw
tri 62221 20172 62951 20902 ne
rect 62951 20172 66180 20902
rect 59674 19323 62102 20172
tri 62102 19323 62951 20172 sw
tri 62951 19323 63800 20172 ne
rect 63800 19323 66180 20172
rect 59674 18474 62951 19323
tri 62951 18474 63800 19323 sw
tri 63800 18474 64649 19323 ne
rect 64649 18474 66180 19323
tri 66180 18474 70306 22600 sw
rect 59674 17625 63800 18474
tri 63800 17625 64649 18474 sw
tri 64649 17625 65498 18474 ne
rect 65498 17625 70306 18474
rect 59674 16943 64649 17625
rect 24343 16400 26877 16943
tri 21400 16380 21420 16400 se
rect 21420 16380 21600 16400
rect 21400 12400 21600 16380
rect 25200 16200 26877 16400
tri 26877 16200 27620 16943 nw
tri 27726 16200 28469 16943 se
rect 28469 16200 30000 16943
rect 25200 15351 26028 16200
tri 26028 15351 26877 16200 nw
tri 26877 15351 27726 16200 se
rect 27726 15351 30000 16200
rect 25200 12400 25400 15351
tri 25400 14723 26028 15351 nw
tri 26249 14723 26877 15351 se
rect 26877 14723 30000 15351
rect 21400 12200 25400 12400
tri 26000 14474 26249 14723 se
rect 26249 14474 30000 14723
rect 10000 10000 19900 10600
rect 10100 9700 19900 10000
rect 10100 9600 16800 9700
rect 10100 5200 11100 9600
rect 16600 9300 16800 9600
rect 19800 9300 19900 9700
rect 16600 9200 19900 9300
rect 10100 4800 16300 5200
rect 10100 4400 11100 4800
rect 11900 4400 12300 4800
rect 13100 4400 13500 4800
rect 14300 4400 14700 4800
rect 15500 4400 16300 4800
rect 10100 4000 16300 4400
rect 10100 3600 11100 4000
rect 11900 3600 12300 4000
rect 13100 3600 13500 4000
rect 14300 3600 14700 4000
rect 15500 3900 16300 4000
rect 15500 3800 19900 3900
rect 15500 3600 16600 3800
rect 10100 3400 16600 3600
rect 19800 3400 19900 3800
rect 10100 3200 19900 3400
rect 15500 2600 19900 3200
rect 26000 -270 30000 14474
tri 30000 12817 34126 16943 nw
tri 59674 12817 63800 16943 ne
rect 63800 16776 64649 16943
tri 64649 16776 65498 17625 sw
tri 65498 16776 66347 17625 ne
rect 66347 16776 70306 17625
rect 63800 16172 65498 16776
tri 65498 16172 66102 16776 sw
tri 66347 16172 66951 16776 ne
rect 66951 16380 70306 16776
tri 70306 16380 72400 18474 sw
rect 66951 16172 72400 16380
rect 63800 15323 66102 16172
tri 66102 15323 66951 16172 sw
tri 66951 15323 67800 16172 ne
rect 67800 15323 72400 16172
rect 63800 14474 66951 15323
tri 66951 14474 67800 15323 sw
tri 67800 14723 68400 15323 ne
rect 30600 4088 34600 4200
tri 30000 -270 30600 330 sw
rect 30600 312 30712 4088
rect 34488 312 34600 4088
rect 30600 200 34600 312
tri 30978 -270 31448 200 ne
rect 31448 -270 34600 200
rect 26000 -1118 30600 -270
tri 30600 -1118 31448 -270 sw
tri 31448 -1118 32296 -270 ne
rect 32296 -1118 34600 -270
rect 26000 -1327 31448 -1118
tri 26000 -6200 30873 -1327 ne
rect 30873 -1726 31448 -1327
tri 31448 -1726 32056 -1118 sw
tri 32296 -1726 32904 -1118 ne
rect 32904 -1726 34600 -1118
rect 30873 -2574 32056 -1726
tri 32056 -2574 32904 -1726 sw
tri 32904 -2574 33752 -1726 ne
rect 33752 -2574 34600 -1726
rect 30873 -3422 32904 -2574
tri 32904 -3422 33752 -2574 sw
tri 33752 -3422 34600 -2574 ne
tri 34600 -3422 40257 2235 sw
tri 61022 -543 63800 2235 se
rect 63800 578 67800 14474
rect 63800 -270 66952 578
tri 66952 -270 67800 578 nw
tri 67800 -270 68400 330 se
rect 68400 -270 72400 15323
rect 63800 -543 66679 -270
tri 66679 -543 66952 -270 nw
tri 67527 -543 67800 -270 se
rect 67800 -543 72400 -270
tri 58143 -3422 61022 -543 se
rect 61022 -1391 65831 -543
tri 65831 -1391 66679 -543 nw
tri 66679 -1391 67527 -543 se
rect 67527 -1327 72400 -543
rect 67527 -1391 68400 -1327
rect 61022 -1726 65496 -1391
tri 65496 -1726 65831 -1391 nw
tri 66344 -1726 66679 -1391 se
rect 66679 -1726 68400 -1391
rect 61022 -2574 64648 -1726
tri 64648 -2574 65496 -1726 nw
tri 65496 -2574 66344 -1726 se
rect 66344 -2574 68400 -1726
rect 61022 -3422 63800 -2574
tri 63800 -3422 64648 -2574 nw
tri 64648 -3422 65496 -2574 se
rect 65496 -3422 68400 -2574
rect 30873 -4270 33752 -3422
tri 33752 -4270 34600 -3422 sw
tri 34600 -4270 35448 -3422 ne
rect 35448 -4270 40257 -3422
rect 30873 -5118 34600 -4270
tri 34600 -5118 35448 -4270 sw
tri 35448 -5118 36296 -4270 ne
rect 36296 -5118 40257 -4270
rect 30873 -5352 35448 -5118
tri 35448 -5352 35682 -5118 sw
tri 36296 -5352 36530 -5118 ne
rect 36530 -5352 40257 -5118
rect 30873 -6200 35682 -5352
tri 35682 -6200 36530 -5352 sw
tri 36530 -6200 37378 -5352 ne
rect 37378 -6200 40257 -5352
tri 40257 -6200 43035 -3422 sw
tri 55365 -6200 58143 -3422 se
rect 58143 -4270 62952 -3422
tri 62952 -4270 63800 -3422 nw
tri 63800 -4270 64648 -3422 se
rect 64648 -4270 68400 -3422
rect 58143 -5118 62104 -4270
tri 62104 -5118 62952 -4270 nw
tri 62952 -5118 63800 -4270 se
rect 63800 -5118 68400 -4270
rect 58143 -5352 61870 -5118
tri 61870 -5352 62104 -5118 nw
tri 62718 -5352 62952 -5118 se
rect 62952 -5327 68400 -5118
tri 68400 -5327 72400 -1327 nw
rect 62952 -5352 63800 -5327
rect 58143 -6200 61022 -5352
tri 61022 -6200 61870 -5352 nw
tri 61870 -6200 62718 -5352 se
rect 62718 -6200 63800 -5352
tri 30873 -10800 35473 -6200 ne
rect 35473 -7048 36530 -6200
tri 36530 -7048 37378 -6200 sw
tri 37378 -7048 38226 -6200 ne
rect 38226 -7048 60174 -6200
tri 60174 -7048 61022 -6200 nw
tri 61022 -7048 61870 -6200 se
rect 61870 -7048 63800 -6200
rect 35473 -7896 37378 -7048
tri 37378 -7896 38226 -7048 sw
tri 38226 -7896 39074 -7048 ne
rect 39074 -7896 59326 -7048
tri 59326 -7896 60174 -7048 nw
tri 60174 -7896 61022 -7048 se
rect 61022 -7896 63800 -7048
rect 35473 -8504 38226 -7896
tri 38226 -8504 38834 -7896 sw
tri 39074 -8504 39682 -7896 ne
rect 39682 -8504 58718 -7896
tri 58718 -8504 59326 -7896 nw
tri 59566 -8504 60174 -7896 se
rect 60174 -8504 63800 -7896
rect 35473 -9352 38834 -8504
tri 38834 -9352 39682 -8504 sw
tri 39682 -9352 40530 -8504 ne
rect 40530 -9352 57870 -8504
tri 57870 -9352 58718 -8504 nw
tri 58718 -9352 59566 -8504 se
rect 59566 -9352 63800 -8504
rect 35473 -10200 39682 -9352
tri 39682 -10200 40530 -9352 sw
tri 40530 -10200 41378 -9352 ne
rect 41378 -10200 57022 -9352
tri 57022 -10200 57870 -9352 nw
tri 57870 -10200 58718 -9352 se
rect 58718 -9927 63800 -9352
tri 63800 -9927 68400 -5327 nw
rect 58718 -10200 58927 -9927
rect 35473 -10800 40530 -10200
tri 40530 -10800 41130 -10200 sw
tri 57270 -10800 57870 -10200 se
rect 57870 -10800 58927 -10200
tri 35473 -14800 39473 -10800 ne
rect 39473 -14800 58927 -10800
tri 58927 -14800 63800 -9927 nw
<< end >>
