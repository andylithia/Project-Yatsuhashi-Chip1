magic
tech sky130A
magscale 1 2
timestamp 1658628487
<< error_s >>
rect 487 1224 511 1244
rect 485 1190 511 1224
rect 487 1178 511 1190
rect 515 1178 549 1244
rect 837 1224 861 1244
rect 835 1190 861 1224
rect 837 1178 861 1190
rect 865 1178 899 1244
rect 519 1174 549 1178
rect 869 1174 899 1178
rect 354 1144 355 1156
rect 348 150 364 1144
rect 376 1140 434 1152
rect 376 1098 441 1140
rect 493 1098 533 1140
rect 592 1132 650 1152
rect 671 1144 672 1156
rect 704 1144 705 1156
rect 585 1098 650 1132
rect 376 1072 434 1098
rect 376 1026 441 1072
rect 493 1026 533 1072
rect 592 1060 650 1098
rect 585 1026 650 1060
rect 376 1004 434 1026
rect 376 954 441 1004
rect 493 954 533 1004
rect 592 988 650 1026
rect 585 954 650 988
rect 376 936 434 954
rect 376 882 441 936
rect 493 882 533 936
rect 592 916 650 954
rect 585 882 650 916
rect 376 868 434 882
rect 376 810 441 868
rect 493 810 533 868
rect 592 844 650 882
rect 585 810 650 844
rect 376 800 434 810
rect 376 738 441 800
rect 493 738 533 800
rect 592 772 650 810
rect 585 738 650 772
rect 376 732 434 738
rect 376 666 441 732
rect 493 666 533 732
rect 592 700 650 738
rect 585 666 650 700
rect 376 664 434 666
rect 376 630 441 664
rect 493 630 533 664
rect 376 628 434 630
rect 592 628 650 666
rect 376 562 441 628
rect 493 592 533 628
rect 585 594 650 628
rect 376 556 434 562
rect 376 494 441 556
rect 484 540 542 592
rect 592 556 650 594
rect 493 528 533 540
rect 376 484 434 494
rect 376 426 441 484
rect 484 476 542 528
rect 585 522 650 556
rect 592 484 650 522
rect 493 464 533 476
rect 376 412 434 426
rect 484 412 542 464
rect 585 450 650 484
rect 592 412 650 450
rect 376 358 441 412
rect 493 400 533 412
rect 376 340 434 358
rect 484 348 542 400
rect 585 378 650 412
rect 592 340 650 378
rect 376 290 441 340
rect 493 336 533 340
rect 376 268 434 290
rect 484 284 542 336
rect 585 306 650 340
rect 376 222 441 268
rect 376 196 434 222
rect 484 220 542 272
rect 592 268 650 306
rect 585 234 650 268
rect 376 162 441 196
rect 350 100 366 150
rect 376 142 434 162
rect 484 156 542 208
rect 592 196 650 234
rect 585 162 650 196
rect 493 154 533 156
rect 592 142 650 162
rect 662 150 678 1144
rect 698 150 714 1144
rect 726 1140 784 1152
rect 726 1098 791 1140
rect 843 1098 883 1140
rect 942 1132 1000 1152
rect 1021 1144 1022 1156
rect 935 1098 1000 1132
rect 726 1072 784 1098
rect 726 1026 791 1072
rect 843 1026 883 1072
rect 942 1060 1000 1098
rect 935 1026 1000 1060
rect 726 1004 784 1026
rect 726 954 791 1004
rect 843 954 883 1004
rect 942 988 1000 1026
rect 935 954 1000 988
rect 726 936 784 954
rect 726 882 791 936
rect 843 882 883 936
rect 942 916 1000 954
rect 935 882 1000 916
rect 726 868 784 882
rect 726 810 791 868
rect 843 810 883 868
rect 942 844 1000 882
rect 935 810 1000 844
rect 726 800 784 810
rect 726 738 791 800
rect 843 738 883 800
rect 942 772 1000 810
rect 935 738 1000 772
rect 726 732 784 738
rect 726 666 791 732
rect 843 666 883 732
rect 942 700 1000 738
rect 935 666 1000 700
rect 726 664 784 666
rect 726 630 791 664
rect 843 630 883 664
rect 726 628 784 630
rect 942 628 1000 666
rect 726 562 791 628
rect 843 592 883 628
rect 935 594 1000 628
rect 726 556 784 562
rect 726 494 791 556
rect 834 540 892 592
rect 942 556 1000 594
rect 843 528 883 540
rect 726 484 784 494
rect 726 426 791 484
rect 834 476 892 528
rect 935 522 1000 556
rect 942 484 1000 522
rect 843 464 883 476
rect 726 412 784 426
rect 834 412 892 464
rect 935 450 1000 484
rect 942 412 1000 450
rect 726 358 791 412
rect 843 400 883 412
rect 726 340 784 358
rect 834 348 892 400
rect 935 378 1000 412
rect 942 340 1000 378
rect 726 290 791 340
rect 843 336 883 340
rect 726 268 784 290
rect 834 284 892 336
rect 935 306 1000 340
rect 726 222 791 268
rect 726 196 784 222
rect 834 220 892 272
rect 942 268 1000 306
rect 935 234 1000 268
rect 726 162 791 196
rect 477 120 482 142
rect 544 120 549 142
rect 671 138 672 150
rect 519 116 549 120
rect 487 104 511 116
rect 485 70 511 104
rect 487 50 511 70
rect 515 50 549 116
rect 700 100 716 150
rect 726 142 784 162
rect 834 156 892 208
rect 942 196 1000 234
rect 935 162 1000 196
rect 843 154 883 156
rect 942 142 1000 162
rect 1012 150 1028 1144
rect 827 120 832 142
rect 894 120 899 142
rect 1021 138 1022 150
rect 869 116 899 120
rect 837 104 861 116
rect 835 70 861 104
rect 837 50 861 70
rect 865 50 899 116
rect 1050 100 1066 150
<< metal2 >>
rect 338 361 350 597
rect 688 361 700 597
rect 1038 361 1050 597
rect 338 100 350 336
rect 688 100 700 336
rect 1038 100 1050 336
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_0 ../SKY130A_rf
timestamp 1649977179
transform 1 0 0 0 1 50
box 0 0 676 1194
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_1
timestamp 1649977179
transform 1 0 700 0 1 50
box 0 0 676 1194
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_2
timestamp 1649977179
transform 1 0 350 0 1 50
box 0 0 676 1194
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_3
timestamp 1649977179
transform 1 0 1540 0 1 654
box 0 0 676 1194
<< end >>
