** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA1.sch
**.subckt LNA1
XM1 net7 vgate1 net1 GND sky130_fd_pr__nfet_01v8 L=L W=W nf=NF ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=M m=M
Ldeg1 net1 GND 0.9n m=1
Li1 net8 net7 3n m=1
V1 net2 GND 1.8
XM2 vbias1 vbias1 GND GND sky130_fd_pr__nfet_01v8 L=L W=W nf=NF ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=M m=M
R1 vbias1 vgate1 10k m=1
I0 net2 vbias1 50u
C1 vbias1 GND 10p m=1
V2 net3 GND dc 0 ac 0 portnum 1 z0 50
C2 net5 net3 1p m=1
V3 net4 GND dc 0 ac 0 portnum 2 z0 200
Lg1 vgate1 net5 0.3n m=1
XM3 net6 net2 net8 GND sky130_fd_pr__nfet_01v8 L=L W=W2 nf=NF ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=M m=M
Li2 net2 net6 1n m=1
C4 net4 net6 10p m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.param L=0.3
.param W=40
.param W2=50
.param NF=1
.param M=1
.op
.sp dec 100 1e9 100e9 0
.control
run
display
plot db(S_1_1) db(S_1_2) db(S_2_2) db(S_2_1)
plot S_1_1 smithgrid
print @m.xm1.msky130_fd_pr__nfet_01v8[id]
print @m.xm1.msky130_fd_pr__nfet_01v8[vgs]
print @m.xm1.msky130_fd_pr__nfet_01v8[vds]
print @m.xm3.msky130_fd_pr__nfet_01v8[vgs]
print @m.xm3.msky130_fd_pr__nfet_01v8[vds]
print @m.xm3.msky130_fd_pr__nfet_01v8[id]
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
