magic
tech sky130B
magscale 1 2
timestamp 1661314321
<< metal4 >>
rect -19900 -4112 -6100 -4000
rect -19900 -7888 -19788 -4112
rect -16012 -7888 -9988 -4112
rect -6212 -7888 -6100 -4112
rect -19900 -8000 -6100 -7888
<< via4 >>
rect -19788 -7888 -16012 -4112
rect -9988 -7888 -6212 -4112
<< metal5 >>
tri -10700 17642 -9342 19000 se
rect -9342 17642 4742 19000
tri 4742 17642 6100 19000 sw
tri -13342 15000 -10700 17642 se
rect -10700 15000 6100 17642
tri 6100 15000 8742 17642 sw
tri -15300 13042 -13342 15000 se
rect -13342 14400 -8285 15000
tri -8285 14400 -7685 15000 nw
tri 3085 14400 3685 15000 ne
rect 3685 14400 8742 15000
rect -13342 13551 -9134 14400
tri -9134 13551 -8285 14400 nw
tri -8285 13551 -7436 14400 se
rect -7436 13551 2836 14400
tri 2836 13551 3685 14400 sw
tri 3685 13551 4534 14400 ne
rect 4534 13551 8742 14400
rect -13342 13042 -9851 13551
tri -16357 11985 -15300 13042 se
rect -15300 12834 -9851 13042
tri -9851 12834 -9134 13551 nw
tri -9002 12834 -8285 13551 se
rect -8285 12834 3685 13551
rect -15300 11985 -10700 12834
tri -10700 11985 -9851 12834 nw
tri -9851 11985 -9002 12834 se
rect -9002 12702 3685 12834
tri 3685 12702 4534 13551 sw
tri 4534 12702 5383 13551 ne
rect 5383 12702 8742 13551
rect -9002 12098 4534 12702
tri 4534 12098 5138 12702 sw
tri 5383 12098 5987 12702 ne
rect 5987 12098 8742 12702
rect -9002 11985 5138 12098
tri -19300 9042 -16357 11985 se
rect -16357 11136 -11549 11985
tri -11549 11136 -10700 11985 nw
tri -10700 11136 -9851 11985 se
rect -9851 11249 5138 11985
tri 5138 11249 5987 12098 sw
tri 5987 11249 6836 12098 ne
rect 6836 11249 8742 12098
rect -9851 11136 5987 11249
tri 5987 11136 6100 11249 sw
tri 6836 11136 6949 11249 ne
rect 6949 11136 8742 11249
rect -16357 10400 -12285 11136
tri -12285 10400 -11549 11136 nw
tri -11436 10400 -10700 11136 se
rect -10700 10400 6100 11136
tri 6100 10400 6836 11136 sw
tri 6949 10400 7685 11136 ne
rect 7685 10400 8742 11136
tri 8742 10400 13342 15000 sw
rect -16357 9551 -13134 10400
tri -13134 9551 -12285 10400 nw
tri -12285 9551 -11436 10400 se
rect -11436 9551 -8179 10400
rect -16357 9042 -13836 9551
rect -19300 8849 -13836 9042
tri -13836 8849 -13134 9551 nw
tri -12987 8849 -12285 9551 se
rect -12285 8849 -8179 9551
rect -19300 8000 -14685 8849
tri -14685 8000 -13836 8849 nw
tri -13836 8000 -12987 8849 se
rect -12987 8000 -8179 8849
tri -8179 8000 -5779 10400 nw
tri 1179 8000 3579 10400 ne
rect 3579 9551 6836 10400
tri 6836 9551 7685 10400 sw
tri 7685 9551 8534 10400 ne
rect 8534 9551 13342 10400
rect 3579 8834 7685 9551
tri 7685 8834 8402 9551 sw
tri 8534 8834 9251 9551 ne
rect 9251 9042 13342 9551
tri 13342 9042 14700 10400 sw
rect 9251 8834 14700 9042
rect 3579 8000 8402 8834
rect -23300 7985 -14700 8000
tri -14700 7985 -14685 8000 nw
tri -13851 7985 -13836 8000 se
rect -13836 7985 -10700 8000
rect -23300 4000 -15300 7985
tri -15300 7385 -14700 7985 nw
tri -14451 7385 -13851 7985 se
rect -13851 7385 -10700 7985
tri -14700 7136 -14451 7385 se
rect -14451 7136 -10700 7385
rect -19900 -4112 -15900 -4000
rect -19900 -7888 -19788 -4112
rect -16012 -7888 -15900 -4112
rect -19900 -8000 -15900 -7888
rect -14700 -9332 -10700 7136
tri -10700 5479 -8179 8000 nw
tri 3579 5479 6100 8000 ne
rect 6100 7985 8402 8000
tri 8402 7985 9251 8834 sw
tri 9251 7985 10100 8834 ne
rect 10100 7985 14700 8834
rect 6100 7385 9251 7985
tri 9251 7385 9851 7985 sw
tri 10100 7385 10700 7985 ne
rect 6100 7136 9851 7385
tri 9851 7136 10100 7385 sw
rect -10100 -4112 -6100 -4000
rect -10100 -7888 -9988 -4112
rect -6212 -7888 -6100 -4112
rect -10100 -8484 -6100 -7888
tri -10100 -8732 -9852 -8484 ne
rect -9852 -8732 -6100 -8484
tri -10700 -9332 -10100 -8732 sw
tri -9852 -9332 -9252 -8732 ne
rect -9252 -9332 -6100 -8732
rect -14700 -9552 -10100 -9332
tri -10100 -9552 -9880 -9332 sw
tri -9252 -9552 -9032 -9332 ne
rect -9032 -9552 -6100 -9332
rect -14700 -10389 -9880 -9552
tri -14700 -10400 -14689 -10389 ne
rect -14689 -10400 -9880 -10389
tri -9880 -10400 -9032 -9552 sw
tri -9032 -10400 -8184 -9552 ne
rect -8184 -10400 -6100 -9552
tri -6100 -10400 -2527 -6827 sw
tri 2527 -10400 6100 -6827 se
rect 6100 -8484 10100 7136
rect 6100 -8732 9852 -8484
tri 9852 -8732 10100 -8484 nw
rect 6100 -9332 9252 -8732
tri 9252 -9332 9852 -8732 nw
tri 10100 -9332 10700 -8732 se
rect 10700 -9332 14700 7985
rect 6100 -9552 9032 -9332
tri 9032 -9552 9252 -9332 nw
tri 9880 -9552 10100 -9332 se
rect 10100 -9552 14700 -9332
rect 6100 -10400 8184 -9552
tri 8184 -10400 9032 -9552 nw
tri 9032 -10400 9880 -9552 se
rect 9880 -10389 14700 -9552
rect 9880 -10400 11757 -10389
tri -14689 -15000 -10089 -10400 ne
rect -10089 -11248 -9032 -10400
tri -9032 -11248 -8184 -10400 sw
tri -8184 -11248 -7336 -10400 ne
rect -7336 -11248 7336 -10400
tri 7336 -11248 8184 -10400 nw
tri 8184 -11248 9032 -10400 se
rect 9032 -11248 11757 -10400
rect -10089 -12096 -8184 -11248
tri -8184 -12096 -7336 -11248 sw
tri -7336 -12096 -6488 -11248 ne
rect -6488 -11636 6948 -11248
tri 6948 -11636 7336 -11248 nw
tri 7796 -11636 8184 -11248 se
rect 8184 -11636 11757 -11248
rect -6488 -12096 6100 -11636
rect -10089 -12704 -7336 -12096
tri -7336 -12704 -6728 -12096 sw
tri -6488 -12704 -5880 -12096 ne
rect -5880 -12484 6100 -12096
tri 6100 -12484 6948 -11636 nw
tri 6948 -12484 7796 -11636 se
rect 7796 -12484 11757 -11636
rect -5880 -12704 5252 -12484
rect -10089 -13552 -6728 -12704
tri -6728 -13552 -5880 -12704 sw
tri -5880 -13552 -5032 -12704 ne
rect -5032 -13332 5252 -12704
tri 5252 -13332 6100 -12484 nw
tri 6100 -13332 6948 -12484 se
rect 6948 -13332 11757 -12484
tri 11757 -13332 14700 -10389 nw
rect -5032 -13552 5032 -13332
tri 5032 -13552 5252 -13332 nw
tri 5880 -13552 6100 -13332 se
rect 6100 -13552 10700 -13332
rect -10089 -14400 -5880 -13552
tri -5880 -14400 -5032 -13552 sw
tri -5032 -14400 -4184 -13552 ne
rect -4184 -14400 4184 -13552
tri 4184 -14400 5032 -13552 nw
tri 5032 -14400 5880 -13552 se
rect 5880 -14389 10700 -13552
tri 10700 -14389 11757 -13332 nw
rect 5880 -14400 10089 -14389
rect -10089 -15000 -5032 -14400
tri -5032 -15000 -4432 -14400 sw
tri 4432 -15000 5032 -14400 se
rect 5032 -15000 10089 -14400
tri 10089 -15000 10700 -14389 nw
tri -10089 -18989 -6100 -15000 ne
rect -6100 -18989 6100 -15000
tri 6100 -18989 10089 -15000 nw
tri -6100 -19000 -6089 -18989 ne
rect -6089 -19000 6089 -18989
tri 6089 -19000 6100 -18989 nw
<< end >>
