magic
tech sky130B
magscale 1 2
timestamp 1662239336
<< nwell >>
rect 9400 400 9422 1269
rect -200 -620 9422 400
rect -200 -700 -80 -620
rect -60 -700 9422 -620
<< locali >>
rect -80 1660 9320 1680
rect -80 1540 -60 1660
rect 9300 1540 9320 1660
rect -80 1520 9320 1540
rect -400 1440 -160 1480
rect -400 300 -380 1440
rect -220 300 -160 1440
rect -400 280 -160 300
rect 9360 1440 9600 1480
rect 9360 300 9420 1440
rect 9580 300 9600 1440
rect 9360 280 9600 300
rect -400 -640 -160 -600
rect -400 -1780 -380 -640
rect -220 -1780 -160 -640
rect -400 -1800 -160 -1780
rect 9360 -660 9600 -620
rect 9360 -1800 9420 -660
rect 9580 -1800 9600 -660
rect 9360 -1820 9600 -1800
rect -100 -1860 9300 -1840
rect -100 -1980 -80 -1860
rect 9280 -1980 9300 -1860
rect -100 -2000 9300 -1980
<< viali >>
rect -60 1540 9300 1660
rect -380 300 -220 1440
rect 9420 300 9580 1440
rect -380 -1780 -220 -640
rect 9420 -1800 9580 -660
rect -80 -1980 9280 -1860
<< metal1 >>
rect -80 1660 9320 1680
rect -80 1540 -60 1660
rect 9300 1540 9320 1660
rect -80 1520 9320 1540
rect -400 1440 -200 1480
rect -400 300 -380 1440
rect -220 300 -200 1440
rect -80 1420 0 1520
rect -80 420 0 440
rect 180 1420 260 1520
rect 180 420 260 440
rect 440 1420 520 1440
rect 440 420 520 440
rect 700 1420 780 1520
rect 700 420 780 440
rect 960 1420 1040 1440
rect 960 420 1040 440
rect 1220 1420 1300 1520
rect 1220 420 1300 440
rect 1480 1420 1560 1440
rect 1480 420 1560 440
rect 1740 1420 1820 1520
rect 1740 420 1820 440
rect 2000 1420 2080 1440
rect 2000 420 2080 440
rect 2240 1420 2320 1520
rect 2240 420 2320 440
rect 2500 1420 2580 1440
rect 2500 420 2580 440
rect 2760 1420 2840 1520
rect 2760 420 2840 440
rect 3020 1420 3100 1440
rect 3020 420 3100 440
rect 3280 1420 3360 1520
rect 3280 420 3360 440
rect 3540 1420 3620 1440
rect 3540 420 3620 440
rect 3800 1420 3880 1520
rect 3800 420 3880 440
rect 4060 1420 4140 1440
rect 4060 420 4140 440
rect 4320 1420 4400 1520
rect 4320 420 4400 440
rect 4580 1420 4660 1440
rect 4580 420 4660 440
rect 4820 1420 4900 1520
rect 4820 420 4900 440
rect 5080 1420 5160 1440
rect 5080 420 5160 440
rect 5340 1420 5420 1520
rect 5340 420 5420 440
rect 5600 1420 5680 1440
rect 5600 420 5680 440
rect 5860 1420 5940 1520
rect 5860 420 5940 440
rect 6120 1420 6200 1440
rect 6120 420 6200 440
rect 6380 1420 6460 1520
rect 6380 420 6460 440
rect 6640 1420 6720 1440
rect 6640 420 6720 440
rect 6900 1420 6980 1520
rect 6900 420 6980 440
rect 7160 1420 7240 1440
rect 7160 420 7240 440
rect 7400 1420 7480 1520
rect 7400 420 7480 440
rect 7660 1420 7740 1440
rect 7660 420 7740 440
rect 7920 1420 8000 1520
rect 7920 420 8000 440
rect 8180 1420 8260 1440
rect 8180 420 8260 440
rect 8440 1420 8520 1520
rect 8440 420 8520 440
rect 8700 1420 8780 1440
rect 8700 420 8780 440
rect 8960 1420 9040 1520
rect 8960 420 9040 440
rect 9220 1420 9300 1520
rect 9220 420 9300 440
rect 9400 1440 9600 1460
rect -20 300 0 380
rect 180 300 200 380
rect 240 300 260 380
rect 440 300 460 380
rect 500 300 520 380
rect 700 300 720 380
rect 760 300 780 380
rect 960 300 980 380
rect 1020 300 1040 380
rect 1220 300 1240 380
rect 1280 300 1300 380
rect 1480 300 1500 380
rect 1540 300 1560 380
rect 1740 300 1760 380
rect 1800 300 1820 380
rect 2000 300 2020 380
rect 2060 300 2080 380
rect 2260 300 2272 380
rect 2308 300 2320 380
rect 2500 300 2520 380
rect 2560 300 2580 380
rect 2760 300 2780 380
rect 2820 300 2840 380
rect 3020 300 3040 380
rect 3080 300 3100 380
rect 3280 300 3300 380
rect 3340 300 3360 380
rect 3540 300 3560 380
rect 3600 300 3620 380
rect 3800 300 3820 380
rect 3860 300 3880 380
rect 4060 300 4080 380
rect 4120 300 4140 380
rect 4320 300 4340 380
rect 4380 300 4400 380
rect 4580 300 4660 380
rect 4840 300 4860 380
rect 4888 300 4900 380
rect 5080 300 5100 380
rect 5140 300 5160 380
rect 5340 300 5360 380
rect 5400 300 5420 380
rect 5600 300 5620 380
rect 5660 300 5680 380
rect 5860 300 5880 380
rect 5920 300 5940 380
rect 6120 300 6140 380
rect 6180 300 6200 380
rect 6380 300 6400 380
rect 6440 300 6460 380
rect 6640 300 6660 380
rect 6700 300 6720 380
rect 6900 300 6920 380
rect 6960 300 6980 380
rect 7160 300 7180 380
rect 7220 300 7240 380
rect 7420 300 7432 380
rect 7468 300 7480 380
rect 7660 300 7680 380
rect 7720 300 7740 380
rect 7920 300 7940 380
rect 7980 300 8000 380
rect 8180 300 8200 380
rect 8240 300 8260 380
rect 8440 300 8460 380
rect 8500 300 8520 380
rect 8700 300 8720 380
rect 8760 300 8780 380
rect 8960 300 8980 380
rect 9020 300 9040 380
rect 9220 300 9240 380
rect 9400 300 9420 1440
rect 9580 300 9600 1440
rect -400 -640 -200 300
rect -400 -1780 -380 -640
rect -220 -1780 -200 -640
rect -20 -700 0 -620
rect 180 -700 200 -620
rect 240 -700 260 -620
rect 440 -700 460 -620
rect 500 -700 520 -620
rect 700 -700 720 -620
rect 760 -700 780 -620
rect 960 -700 980 -620
rect 1020 -700 1040 -620
rect 1220 -700 1240 -620
rect 1280 -700 1300 -620
rect 1480 -700 1500 -620
rect 1540 -700 1560 -620
rect 1740 -700 1760 -620
rect 1800 -700 1820 -620
rect 2000 -700 2020 -620
rect 2060 -700 2080 -620
rect 2260 -700 2280 -620
rect 2320 -700 2340 -620
rect 2520 -700 2540 -620
rect 2580 -700 2600 -620
rect 2780 -700 2792 -620
rect 2828 -700 2840 -620
rect 3020 -700 3040 -620
rect 3080 -700 3100 -620
rect 3280 -700 3300 -620
rect 3340 -700 3360 -620
rect 3540 -700 3560 -620
rect 3600 -700 3620 -620
rect 3800 -700 3820 -620
rect 3860 -700 3880 -620
rect 4060 -700 4080 -620
rect 4120 -700 4140 -620
rect 4320 -700 4340 -620
rect 4380 -700 4400 -620
rect 4580 -700 4660 -620
rect 4840 -700 4852 -620
rect 4888 -700 4900 -620
rect 5080 -700 5100 -620
rect 5140 -700 5160 -620
rect 5340 -700 5360 -620
rect 5400 -700 5420 -620
rect 5600 -700 5620 -620
rect 5660 -700 5680 -620
rect 5860 -700 5880 -620
rect 5920 -700 5940 -620
rect 6120 -700 6140 -620
rect 6180 -700 6200 -620
rect 6380 -700 6400 -620
rect 6440 -700 6460 -620
rect 6640 -700 6660 -620
rect 6700 -700 6720 -620
rect 6900 -700 6912 -620
rect 6948 -700 6960 -620
rect 7140 -700 7160 -620
rect 7200 -700 7220 -620
rect 7400 -700 7420 -620
rect 7460 -700 7480 -620
rect 7660 -700 7680 -620
rect 7720 -700 7740 -620
rect 7920 -700 7940 -620
rect 7980 -700 8000 -620
rect 8180 -700 8200 -620
rect 8240 -700 8260 -620
rect 8440 -700 8460 -620
rect 8500 -700 8520 -620
rect 8700 -700 8720 -620
rect 8760 -700 8780 -620
rect 8960 -700 8980 -620
rect 9020 -700 9040 -620
rect 9220 -700 9240 -620
rect 9400 -660 9600 300
rect -400 -1800 -200 -1780
rect -80 -760 0 -740
rect -80 -1840 0 -1740
rect 180 -760 260 -740
rect 180 -1840 260 -1740
rect 440 -760 520 -740
rect 440 -1760 520 -1740
rect 700 -760 780 -740
rect 700 -1840 780 -1740
rect 960 -760 1040 -740
rect 960 -1760 1040 -1740
rect 1220 -760 1300 -740
rect 1220 -1840 1300 -1740
rect 1480 -760 1560 -740
rect 1480 -1760 1560 -1740
rect 1740 -760 1820 -740
rect 1740 -1840 1820 -1740
rect 2000 -760 2080 -740
rect 2000 -1760 2080 -1740
rect 2260 -760 2340 -740
rect 2260 -1840 2340 -1740
rect 2520 -760 2600 -740
rect 2520 -1760 2600 -1740
rect 2760 -760 2840 -740
rect 2760 -1840 2840 -1740
rect 3020 -760 3100 -740
rect 3020 -1760 3100 -1740
rect 3280 -760 3360 -740
rect 3280 -1840 3360 -1740
rect 3540 -760 3620 -740
rect 3540 -1760 3620 -1740
rect 3800 -760 3880 -740
rect 3800 -1840 3880 -1740
rect 4060 -760 4140 -740
rect 4060 -1760 4140 -1740
rect 4320 -760 4400 -740
rect 4320 -1840 4400 -1740
rect 4580 -760 4660 -740
rect 4580 -1760 4660 -1740
rect 4820 -760 4900 -740
rect 4820 -1840 4900 -1740
rect 5080 -760 5160 -740
rect 5080 -1760 5160 -1740
rect 5340 -760 5420 -740
rect 5340 -1840 5420 -1740
rect 5600 -760 5680 -740
rect 5600 -1760 5680 -1740
rect 5860 -760 5940 -740
rect 5860 -1840 5940 -1740
rect 6120 -760 6200 -740
rect 6120 -1760 6200 -1740
rect 6380 -760 6460 -740
rect 6380 -1840 6460 -1740
rect 6640 -760 6720 -740
rect 6640 -1760 6720 -1740
rect 6880 -760 6960 -740
rect 6880 -1840 6960 -1740
rect 7140 -760 7220 -740
rect 7140 -1760 7220 -1740
rect 7400 -760 7480 -740
rect 7400 -1840 7480 -1740
rect 7660 -760 7740 -740
rect 7660 -1760 7740 -1740
rect 7920 -760 8000 -740
rect 7920 -1840 8000 -1740
rect 8180 -760 8260 -740
rect 8180 -1760 8260 -1740
rect 8440 -760 8520 -740
rect 8440 -1840 8520 -1740
rect 8700 -760 8780 -740
rect 8700 -1760 8780 -1740
rect 8960 -760 9040 -740
rect 8960 -1840 9040 -1740
rect 9220 -760 9300 -740
rect 9220 -1840 9300 -1740
rect 9400 -1800 9420 -660
rect 9580 -1800 9600 -660
rect 9400 -1820 9600 -1800
rect -100 -1860 9300 -1840
rect -100 -1980 -80 -1860
rect 9280 -1980 9300 -1860
rect -100 -2000 9300 -1980
<< via1 >>
rect -60 1540 9300 1660
rect -380 300 -220 1440
rect -80 440 0 1420
rect 180 440 260 1420
rect 440 440 520 1420
rect 700 440 780 1420
rect 960 440 1040 1420
rect 1220 440 1300 1420
rect 1480 440 1560 1420
rect 1740 440 1820 1420
rect 2000 440 2080 1420
rect 2240 440 2320 1420
rect 2500 440 2580 1420
rect 2760 440 2840 1420
rect 3020 440 3100 1420
rect 3280 440 3360 1420
rect 3540 440 3620 1420
rect 3800 440 3880 1420
rect 4060 440 4140 1420
rect 4320 440 4400 1420
rect 4580 440 4660 1420
rect 4820 440 4900 1420
rect 5080 440 5160 1420
rect 5340 440 5420 1420
rect 5600 440 5680 1420
rect 5860 440 5940 1420
rect 6120 440 6200 1420
rect 6380 440 6460 1420
rect 6640 440 6720 1420
rect 6900 440 6980 1420
rect 7160 440 7240 1420
rect 7400 440 7480 1420
rect 7660 440 7740 1420
rect 7920 440 8000 1420
rect 8180 440 8260 1420
rect 8440 440 8520 1420
rect 8700 440 8780 1420
rect 8960 440 9040 1420
rect 9220 440 9300 1420
rect 0 300 180 380
rect 260 300 440 380
rect 520 300 700 380
rect 780 300 960 380
rect 1040 300 1220 380
rect 1300 300 1480 380
rect 1560 300 1740 380
rect 1820 300 2000 380
rect 2080 300 2260 380
rect 2320 300 2500 380
rect 2580 300 2760 380
rect 2840 300 3020 380
rect 3100 300 3280 380
rect 3360 300 3540 380
rect 3620 300 3800 380
rect 3880 300 4060 380
rect 4140 300 4320 380
rect 4400 300 4580 380
rect 4660 300 4840 380
rect 4900 300 5080 380
rect 5160 300 5340 380
rect 5420 300 5600 380
rect 5680 300 5860 380
rect 5940 300 6120 380
rect 6200 300 6380 380
rect 6460 300 6640 380
rect 6720 300 6900 380
rect 6980 300 7160 380
rect 7240 300 7420 380
rect 7480 300 7660 380
rect 7740 300 7920 380
rect 8000 300 8180 380
rect 8260 300 8440 380
rect 8520 300 8700 380
rect 8780 300 8960 380
rect 9040 300 9220 380
rect 9420 300 9580 1440
rect -380 -1780 -220 -640
rect 0 -700 180 -620
rect 260 -700 440 -620
rect 520 -700 700 -620
rect 780 -700 960 -620
rect 1040 -700 1220 -620
rect 1300 -700 1480 -620
rect 1560 -700 1740 -620
rect 1820 -700 2000 -620
rect 2080 -700 2260 -620
rect 2340 -700 2520 -620
rect 2600 -700 2780 -620
rect 2840 -700 3020 -620
rect 3100 -700 3280 -620
rect 3360 -700 3540 -620
rect 3620 -700 3800 -620
rect 3880 -700 4060 -620
rect 4140 -700 4320 -620
rect 4400 -700 4580 -620
rect 4660 -700 4840 -620
rect 4900 -700 5080 -620
rect 5160 -700 5340 -620
rect 5420 -700 5600 -620
rect 5680 -700 5860 -620
rect 5940 -700 6120 -620
rect 6200 -700 6380 -620
rect 6460 -700 6640 -620
rect 6720 -700 6900 -620
rect 6960 -700 7140 -620
rect 7220 -700 7400 -620
rect 7480 -700 7660 -620
rect 7740 -700 7920 -620
rect 8000 -700 8180 -620
rect 8260 -700 8440 -620
rect 8520 -700 8700 -620
rect 8780 -700 8960 -620
rect 9040 -700 9220 -620
rect -80 -1740 0 -760
rect 180 -1740 260 -760
rect 440 -1740 520 -760
rect 700 -1740 780 -760
rect 960 -1740 1040 -760
rect 1220 -1740 1300 -760
rect 1480 -1740 1560 -760
rect 1740 -1740 1820 -760
rect 2000 -1740 2080 -760
rect 2260 -1740 2340 -760
rect 2520 -1740 2600 -760
rect 2760 -1740 2840 -760
rect 3020 -1740 3100 -760
rect 3280 -1740 3360 -760
rect 3540 -1740 3620 -760
rect 3800 -1740 3880 -760
rect 4060 -1740 4140 -760
rect 4320 -1740 4400 -760
rect 4580 -1740 4660 -760
rect 4820 -1740 4900 -760
rect 5080 -1740 5160 -760
rect 5340 -1740 5420 -760
rect 5600 -1740 5680 -760
rect 5860 -1740 5940 -760
rect 6120 -1740 6200 -760
rect 6380 -1740 6460 -760
rect 6640 -1740 6720 -760
rect 6880 -1740 6960 -760
rect 7140 -1740 7220 -760
rect 7400 -1740 7480 -760
rect 7660 -1740 7740 -760
rect 7920 -1740 8000 -760
rect 8180 -1740 8260 -760
rect 8440 -1740 8520 -760
rect 8700 -1740 8780 -760
rect 8960 -1740 9040 -760
rect 9220 -1740 9300 -760
rect 9420 -1800 9580 -660
rect -80 -1980 9280 -1860
<< metal2 >>
rect -400 1660 9600 1680
rect -400 1540 -60 1660
rect 9300 1540 9600 1660
rect -400 1520 9600 1540
rect -400 1440 -200 1520
rect 9400 1440 9600 1520
rect -400 300 -380 1440
rect -220 300 -200 1440
rect -80 1420 0 1440
rect 180 1420 260 1440
rect -80 300 0 440
rect 160 440 180 460
rect 440 1420 520 1440
rect 160 420 260 440
rect 420 530 440 540
rect 700 1420 780 1440
rect 520 530 540 540
rect 420 430 430 530
rect 530 430 540 530
rect 420 420 540 430
rect 960 1420 1040 1440
rect 700 420 780 440
rect 940 530 960 540
rect 1220 1420 1300 1440
rect 1040 530 1060 540
rect 940 430 950 530
rect 1050 430 1060 530
rect 940 420 1060 430
rect 1480 1420 1560 1440
rect 1220 420 1300 440
rect 1460 530 1480 540
rect 1740 1420 1820 1440
rect 1560 530 1580 540
rect 1460 430 1470 530
rect 1570 430 1580 530
rect 1460 420 1580 430
rect 2000 1420 2080 1440
rect 1740 420 1820 440
rect 1980 530 2000 540
rect 2240 1420 2320 1440
rect 2080 530 2100 540
rect 1980 430 1990 530
rect 2090 430 2100 530
rect 1980 420 2100 430
rect 2500 1420 2580 1440
rect 2240 420 2320 440
rect 2480 530 2500 540
rect 2760 1420 2840 1440
rect 2580 530 2600 540
rect 2480 430 2490 530
rect 2590 430 2600 530
rect 2480 420 2600 430
rect 3020 1420 3100 1440
rect 2760 420 2840 440
rect 3000 530 3020 540
rect 3280 1420 3360 1440
rect 3100 530 3120 540
rect 3000 430 3010 530
rect 3110 430 3120 530
rect 3000 420 3120 430
rect 3540 1420 3620 1440
rect 3280 420 3360 440
rect 3520 530 3540 540
rect 3800 1420 3880 1440
rect 3620 530 3640 540
rect 3520 430 3530 530
rect 3630 430 3640 530
rect 3520 420 3640 430
rect 4060 1420 4140 1440
rect 3800 420 3880 440
rect 4040 530 4060 540
rect 4320 1420 4400 1440
rect 4140 530 4160 540
rect 4040 430 4050 530
rect 4150 430 4160 530
rect 4040 420 4160 430
rect 4580 1420 4660 1440
rect 4320 420 4400 440
rect 4560 530 4580 540
rect 4820 1420 4900 1440
rect 4660 530 4680 540
rect 4560 430 4570 530
rect 4670 430 4680 530
rect 160 380 200 420
rect 4560 380 4680 430
rect 5080 1420 5160 1440
rect 4820 420 4900 440
rect 5060 530 5080 540
rect 5340 1420 5420 1440
rect 5160 530 5180 540
rect 5060 430 5070 530
rect 5170 430 5180 530
rect 5060 420 5180 430
rect 5600 1420 5680 1440
rect 5340 420 5420 440
rect 5580 530 5600 540
rect 5860 1420 5940 1440
rect 5680 530 5700 540
rect 5580 430 5590 530
rect 5690 430 5700 530
rect 5580 420 5700 430
rect 6120 1420 6200 1440
rect 5860 420 5940 440
rect 6100 530 6120 540
rect 6380 1420 6460 1440
rect 6200 530 6220 540
rect 6100 430 6110 530
rect 6210 430 6220 530
rect 6100 420 6220 430
rect 6640 1420 6720 1440
rect 6380 420 6460 440
rect 6620 530 6640 540
rect 6900 1420 6980 1440
rect 6720 530 6740 540
rect 6620 430 6630 530
rect 6730 430 6740 530
rect 6620 420 6740 430
rect 7160 1420 7240 1440
rect 6900 420 6980 440
rect 7140 530 7160 540
rect 7400 1420 7480 1440
rect 7240 530 7260 540
rect 7140 430 7150 530
rect 7250 430 7260 530
rect 7140 420 7260 430
rect 7660 1420 7740 1440
rect 7400 420 7480 440
rect 7640 530 7660 540
rect 7920 1420 8000 1440
rect 7740 530 7760 540
rect 7640 430 7650 530
rect 7750 430 7760 530
rect 7640 420 7760 430
rect 8180 1420 8260 1440
rect 7920 420 8000 440
rect 8160 530 8180 540
rect 8440 1420 8520 1440
rect 8260 530 8280 540
rect 8160 430 8170 530
rect 8270 430 8280 530
rect 8160 420 8280 430
rect 8700 1420 8780 1440
rect 8440 420 8520 440
rect 8680 530 8700 540
rect 8960 1420 9040 1440
rect 8780 530 8800 540
rect 8680 430 8690 530
rect 8790 430 8800 530
rect 8680 420 8800 430
rect 9220 1420 9300 1440
rect 9040 440 9060 480
rect 8960 420 9060 440
rect 9020 380 9060 420
rect 180 300 200 380
rect 240 300 260 380
rect 440 300 520 380
rect 700 300 780 380
rect 960 300 1040 380
rect 1220 300 1300 380
rect 1480 300 1560 380
rect 1740 300 1820 380
rect 2000 300 2080 380
rect 2260 300 2320 380
rect 2500 300 2580 380
rect 2760 300 2840 380
rect 3020 300 3100 380
rect 3280 300 3360 380
rect 3540 300 3620 380
rect 3800 300 3880 380
rect 4060 300 4140 380
rect 4320 300 4400 380
rect 4580 300 4660 380
rect 4840 300 4900 380
rect 5080 300 5160 380
rect 5340 300 5420 380
rect 5600 300 5680 380
rect 5860 300 5940 380
rect 6120 300 6200 380
rect 6380 300 6460 380
rect 6640 300 6720 380
rect 6900 300 6980 380
rect 7160 300 7240 380
rect 7420 300 7480 380
rect 7660 300 7740 380
rect 7920 300 8000 380
rect 8180 300 8260 380
rect 8440 300 8520 380
rect 8700 300 8780 380
rect 8960 300 8980 380
rect 9020 300 9040 380
rect 9220 300 9300 440
rect 9400 300 9420 1440
rect 9580 300 9600 1440
rect -400 280 -200 300
rect 9400 280 9600 300
rect -420 190 9400 200
rect -420 120 3530 190
rect 3630 180 5070 190
rect 3630 120 4050 180
rect -420 110 4050 120
rect 4150 120 5070 180
rect 5170 180 6110 190
rect 5170 120 5330 180
rect 4150 110 5330 120
rect 5430 120 6110 180
rect 6210 120 9400 190
rect 5430 110 9400 120
rect -420 100 9400 110
rect -420 50 9400 60
rect -420 -20 1990 50
rect 2090 40 6630 50
rect 2090 -20 2510 40
rect -420 -30 2510 -20
rect 2610 -30 6110 40
rect 6210 -20 6630 40
rect 6730 40 9400 50
rect 6730 -20 6870 40
rect 6210 -30 6870 -20
rect 6970 -30 9400 40
rect -420 -40 9400 -30
rect -420 -90 9400 -80
rect -420 -100 950 -90
rect -420 -170 430 -100
rect 530 -170 950 -100
rect 1050 -170 1470 -90
rect 1570 -170 7650 -90
rect 7750 -170 8170 -90
rect 8270 -160 8690 -90
rect 8790 -160 9400 -90
rect 8270 -170 9400 -160
rect -420 -180 9400 -170
rect -420 -230 9400 -220
rect -420 -240 2230 -230
rect -420 -310 1990 -240
rect 2090 -300 2230 -240
rect 2330 -240 7150 -230
rect 2330 -300 3010 -240
rect 2090 -310 3010 -300
rect 3110 -310 6630 -240
rect 6730 -300 7150 -240
rect 7250 -300 9400 -230
rect 6730 -310 9400 -300
rect -420 -320 9400 -310
rect -420 -370 9400 -360
rect -420 -440 2750 -370
rect 2850 -380 3790 -370
rect 2850 -440 3530 -380
rect -420 -450 3530 -440
rect 3630 -440 3790 -380
rect 3890 -380 5590 -370
rect 3890 -440 5070 -380
rect 3630 -450 5070 -440
rect 5170 -440 5590 -380
rect 5690 -440 9400 -370
rect 5170 -450 9400 -440
rect -420 -460 9400 -450
rect -400 -640 -200 -600
rect -400 -1780 -380 -640
rect -220 -1780 -200 -640
rect -80 -760 0 -620
rect 180 -700 200 -620
rect 240 -700 260 -620
rect 440 -700 520 -620
rect 700 -700 780 -620
rect 960 -700 1040 -620
rect 1220 -700 1300 -620
rect 1480 -700 1560 -620
rect 1740 -700 1820 -620
rect 2000 -700 2080 -620
rect 2260 -700 2340 -620
rect 2520 -700 2600 -620
rect 2780 -700 2840 -620
rect 3020 -700 3100 -620
rect 3280 -700 3360 -620
rect 3540 -700 3620 -620
rect 3800 -700 3880 -620
rect 4060 -700 4140 -620
rect 4320 -700 4400 -620
rect 4580 -700 4660 -620
rect 4840 -700 4900 -620
rect 5080 -700 5160 -620
rect 5340 -700 5420 -620
rect 5600 -700 5680 -620
rect 5860 -700 5940 -620
rect 6120 -700 6200 -620
rect 6380 -700 6460 -620
rect 6640 -700 6720 -620
rect 6900 -700 6960 -620
rect 7140 -700 7220 -620
rect 7400 -700 7480 -620
rect 7660 -700 7740 -620
rect 7920 -700 8000 -620
rect 8180 -700 8260 -620
rect 8440 -700 8520 -620
rect 8700 -700 8780 -620
rect 8960 -700 8980 -620
rect 9020 -700 9040 -620
rect 160 -740 200 -700
rect 160 -760 260 -740
rect 160 -780 180 -760
rect -80 -1760 0 -1740
rect 420 -750 540 -740
rect 420 -850 430 -750
rect 530 -850 540 -750
rect 420 -860 440 -850
rect 180 -1760 260 -1740
rect 520 -860 540 -850
rect 700 -760 780 -740
rect 440 -1760 520 -1740
rect 940 -750 1060 -740
rect 940 -850 950 -750
rect 1050 -850 1060 -750
rect 940 -860 960 -850
rect 700 -1760 780 -1740
rect 1040 -860 1060 -850
rect 1220 -760 1300 -740
rect 960 -1760 1040 -1740
rect 1460 -750 1580 -740
rect 1460 -850 1470 -750
rect 1570 -850 1580 -750
rect 1460 -860 1480 -850
rect 1220 -1760 1300 -1740
rect 1560 -860 1580 -850
rect 1740 -760 1820 -740
rect 1480 -1760 1560 -1740
rect 1980 -750 2100 -740
rect 1980 -850 1990 -750
rect 2090 -850 2100 -750
rect 1980 -860 2000 -850
rect 1740 -1760 1820 -1740
rect 2080 -860 2100 -850
rect 2260 -760 2340 -740
rect 2000 -1760 2080 -1740
rect 2500 -750 2620 -740
rect 2500 -850 2510 -750
rect 2610 -850 2620 -750
rect 2500 -860 2520 -850
rect 2260 -1760 2340 -1740
rect 2600 -860 2620 -850
rect 2760 -760 2840 -740
rect 2520 -1760 2600 -1740
rect 3000 -750 3120 -740
rect 3000 -850 3010 -750
rect 3110 -850 3120 -750
rect 3000 -860 3020 -850
rect 2760 -1760 2840 -1740
rect 3100 -860 3120 -850
rect 3280 -760 3360 -740
rect 3020 -1760 3100 -1740
rect 3520 -750 3640 -740
rect 3520 -850 3530 -750
rect 3630 -850 3640 -750
rect 3520 -860 3540 -850
rect 3280 -1760 3360 -1740
rect 3620 -860 3640 -850
rect 3800 -760 3880 -740
rect 3540 -1760 3620 -1740
rect 4040 -750 4160 -740
rect 4040 -850 4050 -750
rect 4150 -850 4160 -750
rect 4040 -860 4060 -850
rect 3800 -1760 3880 -1740
rect 4140 -860 4160 -850
rect 4320 -760 4400 -740
rect 4060 -1760 4140 -1740
rect 4560 -750 4680 -700
rect 9020 -740 9060 -700
rect 4560 -850 4570 -750
rect 4670 -850 4680 -750
rect 4560 -860 4580 -850
rect 4320 -1760 4400 -1740
rect 4660 -860 4680 -850
rect 4820 -760 4900 -740
rect 4580 -1760 4660 -1740
rect 5060 -750 5180 -740
rect 5060 -850 5070 -750
rect 5170 -850 5180 -750
rect 5060 -860 5080 -850
rect 4820 -1760 4900 -1740
rect 5160 -860 5180 -850
rect 5340 -760 5420 -740
rect 5080 -1760 5160 -1740
rect 5580 -750 5700 -740
rect 5580 -850 5590 -750
rect 5690 -850 5700 -750
rect 5580 -860 5600 -850
rect 5340 -1760 5420 -1740
rect 5680 -860 5700 -850
rect 5860 -760 5940 -740
rect 5600 -1760 5680 -1740
rect 6100 -750 6220 -740
rect 6100 -850 6110 -750
rect 6210 -850 6220 -750
rect 6100 -860 6120 -850
rect 5860 -1760 5940 -1740
rect 6200 -860 6220 -850
rect 6380 -760 6460 -740
rect 6120 -1760 6200 -1740
rect 6620 -750 6740 -740
rect 6620 -850 6630 -750
rect 6730 -850 6740 -750
rect 6620 -860 6640 -850
rect 6380 -1760 6460 -1740
rect 6720 -860 6740 -850
rect 6880 -760 6960 -740
rect 6640 -1760 6720 -1740
rect 7120 -750 7240 -740
rect 7120 -850 7130 -750
rect 7230 -850 7240 -750
rect 7120 -860 7140 -850
rect 6880 -1760 6960 -1740
rect 7220 -860 7240 -850
rect 7400 -760 7480 -740
rect 7140 -1760 7220 -1740
rect 7640 -750 7760 -740
rect 7640 -850 7650 -750
rect 7750 -850 7760 -750
rect 7640 -860 7660 -850
rect 7400 -1760 7480 -1740
rect 7740 -860 7760 -850
rect 7920 -760 8000 -740
rect 7660 -1760 7740 -1740
rect 8160 -750 8280 -740
rect 8160 -850 8170 -750
rect 8270 -850 8280 -750
rect 8160 -860 8180 -850
rect 7920 -1760 8000 -1740
rect 8260 -860 8280 -850
rect 8440 -760 8520 -740
rect 8180 -1760 8260 -1740
rect 8680 -750 8800 -740
rect 8680 -850 8690 -750
rect 8790 -850 8800 -750
rect 8680 -860 8700 -850
rect 8440 -1760 8520 -1740
rect 8780 -860 8800 -850
rect 8960 -760 9060 -740
rect 8700 -1760 8780 -1740
rect 9040 -780 9060 -760
rect 9220 -760 9300 -620
rect 8960 -1760 9040 -1740
rect 9220 -1760 9300 -1740
rect 9400 -660 9600 -600
rect -400 -1840 -200 -1780
rect 9400 -1800 9420 -660
rect 9580 -1800 9600 -660
rect 9400 -1840 9600 -1800
rect -400 -1860 9600 -1840
rect -400 -1980 -80 -1860
rect 9280 -1980 9600 -1860
rect -400 -2000 9600 -1980
<< via2 >>
rect 430 440 440 530
rect 440 440 520 530
rect 520 440 530 530
rect 430 430 530 440
rect 950 440 960 530
rect 960 440 1040 530
rect 1040 440 1050 530
rect 950 430 1050 440
rect 1470 440 1480 530
rect 1480 440 1560 530
rect 1560 440 1570 530
rect 1470 430 1570 440
rect 1990 440 2000 530
rect 2000 440 2080 530
rect 2080 440 2090 530
rect 1990 430 2090 440
rect 2490 440 2500 530
rect 2500 440 2580 530
rect 2580 440 2590 530
rect 2490 430 2590 440
rect 3010 440 3020 530
rect 3020 440 3100 530
rect 3100 440 3110 530
rect 3010 430 3110 440
rect 3530 440 3540 530
rect 3540 440 3620 530
rect 3620 440 3630 530
rect 3530 430 3630 440
rect 4050 440 4060 530
rect 4060 440 4140 530
rect 4140 440 4150 530
rect 4050 430 4150 440
rect 4570 440 4580 530
rect 4580 440 4660 530
rect 4660 440 4670 530
rect 4570 430 4670 440
rect 5070 440 5080 530
rect 5080 440 5160 530
rect 5160 440 5170 530
rect 5070 430 5170 440
rect 5590 440 5600 530
rect 5600 440 5680 530
rect 5680 440 5690 530
rect 5590 430 5690 440
rect 6110 440 6120 530
rect 6120 440 6200 530
rect 6200 440 6210 530
rect 6110 430 6210 440
rect 6630 440 6640 530
rect 6640 440 6720 530
rect 6720 440 6730 530
rect 6630 430 6730 440
rect 7150 440 7160 530
rect 7160 440 7240 530
rect 7240 440 7250 530
rect 7150 430 7250 440
rect 7650 440 7660 530
rect 7660 440 7740 530
rect 7740 440 7750 530
rect 7650 430 7750 440
rect 8170 440 8180 530
rect 8180 440 8260 530
rect 8260 440 8270 530
rect 8170 430 8270 440
rect 8690 440 8700 530
rect 8700 440 8780 530
rect 8780 440 8790 530
rect 8690 430 8790 440
rect 3530 120 3630 190
rect 4050 110 4150 180
rect 5070 120 5170 190
rect 5330 110 5430 180
rect 6110 120 6210 190
rect 1990 -20 2090 50
rect 2510 -30 2610 40
rect 6110 -30 6210 40
rect 6630 -20 6730 50
rect 6870 -30 6970 40
rect 430 -170 530 -100
rect 950 -170 1050 -90
rect 1470 -170 1570 -90
rect 7650 -170 7750 -90
rect 8170 -170 8270 -90
rect 8690 -160 8790 -90
rect 1990 -310 2090 -240
rect 2230 -300 2330 -230
rect 3010 -310 3110 -240
rect 6630 -310 6730 -240
rect 7150 -300 7250 -230
rect 2750 -440 2850 -370
rect 3530 -450 3630 -380
rect 3790 -440 3890 -370
rect 5070 -450 5170 -380
rect 5590 -440 5690 -370
rect 430 -760 530 -750
rect 430 -850 440 -760
rect 440 -850 520 -760
rect 520 -850 530 -760
rect 950 -760 1050 -750
rect 950 -850 960 -760
rect 960 -850 1040 -760
rect 1040 -850 1050 -760
rect 1470 -760 1570 -750
rect 1470 -850 1480 -760
rect 1480 -850 1560 -760
rect 1560 -850 1570 -760
rect 1990 -760 2090 -750
rect 1990 -850 2000 -760
rect 2000 -850 2080 -760
rect 2080 -850 2090 -760
rect 2510 -760 2610 -750
rect 2510 -850 2520 -760
rect 2520 -850 2600 -760
rect 2600 -850 2610 -760
rect 3010 -760 3110 -750
rect 3010 -850 3020 -760
rect 3020 -850 3100 -760
rect 3100 -850 3110 -760
rect 3530 -760 3630 -750
rect 3530 -850 3540 -760
rect 3540 -850 3620 -760
rect 3620 -850 3630 -760
rect 4050 -760 4150 -750
rect 4050 -850 4060 -760
rect 4060 -850 4140 -760
rect 4140 -850 4150 -760
rect 4570 -760 4670 -750
rect 4570 -850 4580 -760
rect 4580 -850 4660 -760
rect 4660 -850 4670 -760
rect 5070 -760 5170 -750
rect 5070 -850 5080 -760
rect 5080 -850 5160 -760
rect 5160 -850 5170 -760
rect 5590 -760 5690 -750
rect 5590 -850 5600 -760
rect 5600 -850 5680 -760
rect 5680 -850 5690 -760
rect 6110 -760 6210 -750
rect 6110 -850 6120 -760
rect 6120 -850 6200 -760
rect 6200 -850 6210 -760
rect 6630 -760 6730 -750
rect 6630 -850 6640 -760
rect 6640 -850 6720 -760
rect 6720 -850 6730 -760
rect 7130 -760 7230 -750
rect 7130 -850 7140 -760
rect 7140 -850 7220 -760
rect 7220 -850 7230 -760
rect 7650 -760 7750 -750
rect 7650 -850 7660 -760
rect 7660 -850 7740 -760
rect 7740 -850 7750 -760
rect 8170 -760 8270 -750
rect 8170 -850 8180 -760
rect 8180 -850 8260 -760
rect 8260 -850 8270 -760
rect 8690 -760 8790 -750
rect 8690 -850 8700 -760
rect 8700 -850 8780 -760
rect 8780 -850 8790 -760
<< metal3 >>
rect 420 530 540 540
rect 420 430 430 530
rect 530 430 540 530
rect 420 420 540 430
rect 940 530 1060 540
rect 940 430 950 530
rect 1050 430 1060 530
rect 940 -90 1060 430
rect 420 -100 540 -90
rect 420 -170 430 -100
rect 530 -170 540 -100
rect 420 -750 540 -170
rect 420 -850 430 -750
rect 530 -850 540 -750
rect 420 -860 540 -850
rect 940 -170 950 -90
rect 1050 -170 1060 -90
rect 940 -750 1060 -170
rect 940 -850 950 -750
rect 1050 -850 1060 -750
rect 940 -860 1060 -850
rect 1460 530 1580 540
rect 1460 430 1470 530
rect 1570 430 1580 530
rect 1460 -90 1580 430
rect 1980 530 2100 540
rect 1980 430 1990 530
rect 2090 430 2100 530
rect 1980 50 2100 430
rect 2480 530 2600 540
rect 2480 430 2490 530
rect 2590 430 2600 530
rect 2480 300 2600 430
rect 3000 530 3120 540
rect 3000 430 3010 530
rect 3110 430 3120 530
rect 3000 300 3120 430
rect 1980 -20 1990 50
rect 2090 -20 2100 50
rect 1980 -30 2100 -20
rect 2220 220 2600 300
rect 2740 220 3120 300
rect 3520 530 3640 540
rect 3520 430 3530 530
rect 3630 430 3640 530
rect 1460 -170 1470 -90
rect 1570 -170 1580 -90
rect 1460 -750 1580 -170
rect 2220 -230 2340 220
rect 1460 -850 1470 -750
rect 1570 -850 1580 -750
rect 1460 -860 1580 -850
rect 1980 -240 2100 -230
rect 1980 -310 1990 -240
rect 2090 -310 2100 -240
rect 2220 -300 2230 -230
rect 2330 -300 2340 -230
rect 2220 -310 2340 -300
rect 2500 40 2620 50
rect 2500 -30 2510 40
rect 2610 -30 2620 40
rect 1980 -750 2100 -310
rect 1980 -850 1990 -750
rect 2090 -850 2100 -750
rect 1980 -860 2100 -850
rect 2500 -750 2620 -30
rect 2740 -370 2860 220
rect 3520 190 3640 430
rect 4040 530 4160 540
rect 4040 430 4050 530
rect 4150 430 4160 530
rect 4040 330 4160 430
rect 3520 120 3530 190
rect 3630 120 3640 190
rect 3520 110 3640 120
rect 3780 250 4160 330
rect 4560 530 4680 540
rect 4560 430 4570 530
rect 4670 430 4680 530
rect 2740 -440 2750 -370
rect 2850 -440 2860 -370
rect 2740 -450 2860 -440
rect 3000 -240 3120 -230
rect 3000 -310 3010 -240
rect 3110 -310 3120 -240
rect 2500 -850 2510 -750
rect 2610 -850 2620 -750
rect 2500 -860 2620 -850
rect 3000 -750 3120 -310
rect 3780 -370 3900 250
rect 3000 -850 3010 -750
rect 3110 -850 3120 -750
rect 3000 -860 3120 -850
rect 3520 -380 3640 -370
rect 3520 -450 3530 -380
rect 3630 -450 3640 -380
rect 3780 -440 3790 -370
rect 3890 -440 3900 -370
rect 3780 -450 3900 -440
rect 4040 180 4160 190
rect 4040 110 4050 180
rect 4150 110 4160 180
rect 3520 -750 3640 -450
rect 3520 -850 3530 -750
rect 3630 -850 3640 -750
rect 3520 -860 3640 -850
rect 4040 -750 4160 110
rect 4040 -850 4050 -750
rect 4150 -850 4160 -750
rect 4040 -860 4160 -850
rect 4560 -750 4680 430
rect 5060 530 5180 540
rect 5060 430 5070 530
rect 5170 430 5180 530
rect 5060 190 5180 430
rect 5580 530 5700 540
rect 5580 430 5590 530
rect 5690 430 5700 530
rect 5060 120 5070 190
rect 5170 120 5180 190
rect 5060 110 5180 120
rect 5320 180 5440 190
rect 5320 110 5330 180
rect 5430 110 5440 180
rect 4560 -850 4570 -750
rect 4670 -850 4680 -750
rect 4560 -2040 4680 -850
rect 5060 -380 5180 -370
rect 5060 -450 5070 -380
rect 5170 -450 5180 -380
rect 5060 -750 5180 -450
rect 5320 -540 5440 110
rect 5580 -370 5700 430
rect 6100 530 6220 540
rect 6100 430 6110 530
rect 6210 430 6220 530
rect 6100 190 6220 430
rect 6100 120 6110 190
rect 6210 120 6220 190
rect 6100 110 6220 120
rect 6620 530 6740 540
rect 6620 430 6630 530
rect 6730 430 6740 530
rect 6620 50 6740 430
rect 7140 530 7260 540
rect 7140 430 7150 530
rect 7250 430 7260 530
rect 5580 -440 5590 -370
rect 5690 -440 5700 -370
rect 5580 -450 5700 -440
rect 6100 40 6220 50
rect 6100 -30 6110 40
rect 6210 -30 6220 40
rect 6620 -20 6630 50
rect 6730 -20 6740 50
rect 6620 -30 6740 -20
rect 6860 40 6980 50
rect 6860 -30 6870 40
rect 6970 -30 6980 40
rect 5320 -620 5700 -540
rect 5060 -850 5070 -750
rect 5170 -850 5180 -750
rect 5060 -860 5180 -850
rect 5580 -750 5700 -620
rect 5580 -850 5590 -750
rect 5690 -850 5700 -750
rect 5580 -860 5700 -850
rect 6100 -750 6220 -30
rect 6100 -850 6110 -750
rect 6210 -850 6220 -750
rect 6100 -860 6220 -850
rect 6620 -240 6740 -230
rect 6620 -310 6630 -240
rect 6730 -310 6740 -240
rect 6620 -750 6740 -310
rect 6860 -540 6980 -30
rect 7140 -230 7260 430
rect 7140 -300 7150 -230
rect 7250 -300 7260 -230
rect 7140 -310 7260 -300
rect 7640 530 7760 540
rect 7640 430 7650 530
rect 7750 430 7760 530
rect 7640 -90 7760 430
rect 7640 -170 7650 -90
rect 7750 -170 7760 -90
rect 6860 -620 7240 -540
rect 6620 -850 6630 -750
rect 6730 -850 6740 -750
rect 6620 -860 6740 -850
rect 7120 -750 7240 -620
rect 7120 -850 7130 -750
rect 7230 -850 7240 -750
rect 7120 -860 7240 -850
rect 7640 -750 7760 -170
rect 7640 -850 7650 -750
rect 7750 -850 7760 -750
rect 7640 -860 7760 -850
rect 8160 530 8280 540
rect 8160 430 8170 530
rect 8270 430 8280 530
rect 8160 -90 8280 430
rect 8160 -170 8170 -90
rect 8270 -170 8280 -90
rect 8680 530 8800 540
rect 8680 430 8690 530
rect 8790 430 8800 530
rect 8680 -90 8800 430
rect 8680 -160 8690 -90
rect 8790 -160 8800 -90
rect 8680 -170 8800 -160
rect 8160 -750 8280 -170
rect 8160 -850 8170 -750
rect 8270 -850 8280 -750
rect 8160 -860 8280 -850
rect 8680 -750 8800 -740
rect 8680 -850 8690 -750
rect 8790 -850 8800 -750
rect 8680 -860 8800 -850
use sky130_fd_pr__pfet_01v8_VM83GD  sky130_fd_pr__pfet_01v8_VM83GD_0
timestamp 1662234432
transform 1 0 4611 0 1 884
box -4811 -684 4811 684
use sky130_fd_pr__pfet_01v8_VM83GD  sky130_fd_pr__pfet_01v8_VM83GD_1
timestamp 1662234432
transform 1 0 4611 0 -1 -1216
box -4811 -684 4811 684
<< labels >>
rlabel metal3 4560 -2040 4680 -2020 1 IREF
rlabel metal2 -420 100 -400 200 1 A
rlabel metal2 -420 -40 -400 60 1 B
rlabel metal2 -420 -180 -400 -80 1 R
rlabel metal2 -420 -320 -400 -220 1 C
rlabel metal2 -420 -460 -400 -360 1 D
rlabel metal2 -400 1540 -200 1680 1 VHI
<< end >>
