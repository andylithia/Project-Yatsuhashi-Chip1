magic
tech sky130B
timestamp 1660526289
use octa_1p2n_2_0  octa_1p2n_2_0_0
timestamp 1660526289
transform 1 0 -10000 0 1 -10000
box -15900 -11500 11600 11500
<< end >>
