magic
tech sky130A
timestamp 1658635850
use 2  2_0
timestamp 1649977179
transform 1 0 -7 0 1 0
box 7 0 394 694
<< end >>
