magic
tech sky130B
magscale 1 2
timestamp 1663719933
<< pwell >>
rect -2569 -3258 2569 3258
<< mvnmos >>
rect -2341 -3000 -2241 3000
rect -2183 -3000 -2083 3000
rect -2025 -3000 -1925 3000
rect -1867 -3000 -1767 3000
rect -1709 -3000 -1609 3000
rect -1551 -3000 -1451 3000
rect -1393 -3000 -1293 3000
rect -1235 -3000 -1135 3000
rect -1077 -3000 -977 3000
rect -919 -3000 -819 3000
rect -761 -3000 -661 3000
rect -603 -3000 -503 3000
rect -445 -3000 -345 3000
rect -287 -3000 -187 3000
rect -129 -3000 -29 3000
rect 29 -3000 129 3000
rect 187 -3000 287 3000
rect 345 -3000 445 3000
rect 503 -3000 603 3000
rect 661 -3000 761 3000
rect 819 -3000 919 3000
rect 977 -3000 1077 3000
rect 1135 -3000 1235 3000
rect 1293 -3000 1393 3000
rect 1451 -3000 1551 3000
rect 1609 -3000 1709 3000
rect 1767 -3000 1867 3000
rect 1925 -3000 2025 3000
rect 2083 -3000 2183 3000
rect 2241 -3000 2341 3000
<< mvndiff >>
rect -2399 2988 -2341 3000
rect -2399 -2988 -2387 2988
rect -2353 -2988 -2341 2988
rect -2399 -3000 -2341 -2988
rect -2241 2988 -2183 3000
rect -2241 -2988 -2229 2988
rect -2195 -2988 -2183 2988
rect -2241 -3000 -2183 -2988
rect -2083 2988 -2025 3000
rect -2083 -2988 -2071 2988
rect -2037 -2988 -2025 2988
rect -2083 -3000 -2025 -2988
rect -1925 2988 -1867 3000
rect -1925 -2988 -1913 2988
rect -1879 -2988 -1867 2988
rect -1925 -3000 -1867 -2988
rect -1767 2988 -1709 3000
rect -1767 -2988 -1755 2988
rect -1721 -2988 -1709 2988
rect -1767 -3000 -1709 -2988
rect -1609 2988 -1551 3000
rect -1609 -2988 -1597 2988
rect -1563 -2988 -1551 2988
rect -1609 -3000 -1551 -2988
rect -1451 2988 -1393 3000
rect -1451 -2988 -1439 2988
rect -1405 -2988 -1393 2988
rect -1451 -3000 -1393 -2988
rect -1293 2988 -1235 3000
rect -1293 -2988 -1281 2988
rect -1247 -2988 -1235 2988
rect -1293 -3000 -1235 -2988
rect -1135 2988 -1077 3000
rect -1135 -2988 -1123 2988
rect -1089 -2988 -1077 2988
rect -1135 -3000 -1077 -2988
rect -977 2988 -919 3000
rect -977 -2988 -965 2988
rect -931 -2988 -919 2988
rect -977 -3000 -919 -2988
rect -819 2988 -761 3000
rect -819 -2988 -807 2988
rect -773 -2988 -761 2988
rect -819 -3000 -761 -2988
rect -661 2988 -603 3000
rect -661 -2988 -649 2988
rect -615 -2988 -603 2988
rect -661 -3000 -603 -2988
rect -503 2988 -445 3000
rect -503 -2988 -491 2988
rect -457 -2988 -445 2988
rect -503 -3000 -445 -2988
rect -345 2988 -287 3000
rect -345 -2988 -333 2988
rect -299 -2988 -287 2988
rect -345 -3000 -287 -2988
rect -187 2988 -129 3000
rect -187 -2988 -175 2988
rect -141 -2988 -129 2988
rect -187 -3000 -129 -2988
rect -29 2988 29 3000
rect -29 -2988 -17 2988
rect 17 -2988 29 2988
rect -29 -3000 29 -2988
rect 129 2988 187 3000
rect 129 -2988 141 2988
rect 175 -2988 187 2988
rect 129 -3000 187 -2988
rect 287 2988 345 3000
rect 287 -2988 299 2988
rect 333 -2988 345 2988
rect 287 -3000 345 -2988
rect 445 2988 503 3000
rect 445 -2988 457 2988
rect 491 -2988 503 2988
rect 445 -3000 503 -2988
rect 603 2988 661 3000
rect 603 -2988 615 2988
rect 649 -2988 661 2988
rect 603 -3000 661 -2988
rect 761 2988 819 3000
rect 761 -2988 773 2988
rect 807 -2988 819 2988
rect 761 -3000 819 -2988
rect 919 2988 977 3000
rect 919 -2988 931 2988
rect 965 -2988 977 2988
rect 919 -3000 977 -2988
rect 1077 2988 1135 3000
rect 1077 -2988 1089 2988
rect 1123 -2988 1135 2988
rect 1077 -3000 1135 -2988
rect 1235 2988 1293 3000
rect 1235 -2988 1247 2988
rect 1281 -2988 1293 2988
rect 1235 -3000 1293 -2988
rect 1393 2988 1451 3000
rect 1393 -2988 1405 2988
rect 1439 -2988 1451 2988
rect 1393 -3000 1451 -2988
rect 1551 2988 1609 3000
rect 1551 -2988 1563 2988
rect 1597 -2988 1609 2988
rect 1551 -3000 1609 -2988
rect 1709 2988 1767 3000
rect 1709 -2988 1721 2988
rect 1755 -2988 1767 2988
rect 1709 -3000 1767 -2988
rect 1867 2988 1925 3000
rect 1867 -2988 1879 2988
rect 1913 -2988 1925 2988
rect 1867 -3000 1925 -2988
rect 2025 2988 2083 3000
rect 2025 -2988 2037 2988
rect 2071 -2988 2083 2988
rect 2025 -3000 2083 -2988
rect 2183 2988 2241 3000
rect 2183 -2988 2195 2988
rect 2229 -2988 2241 2988
rect 2183 -3000 2241 -2988
rect 2341 2988 2399 3000
rect 2341 -2988 2353 2988
rect 2387 -2988 2399 2988
rect 2341 -3000 2399 -2988
<< mvndiffc >>
rect -2387 -2988 -2353 2988
rect -2229 -2988 -2195 2988
rect -2071 -2988 -2037 2988
rect -1913 -2988 -1879 2988
rect -1755 -2988 -1721 2988
rect -1597 -2988 -1563 2988
rect -1439 -2988 -1405 2988
rect -1281 -2988 -1247 2988
rect -1123 -2988 -1089 2988
rect -965 -2988 -931 2988
rect -807 -2988 -773 2988
rect -649 -2988 -615 2988
rect -491 -2988 -457 2988
rect -333 -2988 -299 2988
rect -175 -2988 -141 2988
rect -17 -2988 17 2988
rect 141 -2988 175 2988
rect 299 -2988 333 2988
rect 457 -2988 491 2988
rect 615 -2988 649 2988
rect 773 -2988 807 2988
rect 931 -2988 965 2988
rect 1089 -2988 1123 2988
rect 1247 -2988 1281 2988
rect 1405 -2988 1439 2988
rect 1563 -2988 1597 2988
rect 1721 -2988 1755 2988
rect 1879 -2988 1913 2988
rect 2037 -2988 2071 2988
rect 2195 -2988 2229 2988
rect 2353 -2988 2387 2988
<< mvpsubdiff >>
rect -2533 3210 2533 3222
rect -2533 3176 -2425 3210
rect 2425 3176 2533 3210
rect -2533 3164 2533 3176
rect -2533 3114 -2475 3164
rect -2533 -3114 -2521 3114
rect -2487 -3114 -2475 3114
rect 2475 3114 2533 3164
rect -2533 -3164 -2475 -3114
rect 2475 -3114 2487 3114
rect 2521 -3114 2533 3114
rect 2475 -3164 2533 -3114
rect -2533 -3176 2533 -3164
rect -2533 -3210 -2425 -3176
rect 2425 -3210 2533 -3176
rect -2533 -3222 2533 -3210
<< mvpsubdiffcont >>
rect -2425 3176 2425 3210
rect -2521 -3114 -2487 3114
rect 2487 -3114 2521 3114
rect -2425 -3210 2425 -3176
<< poly >>
rect -2341 3072 -2241 3088
rect -2341 3038 -2325 3072
rect -2257 3038 -2241 3072
rect -2341 3000 -2241 3038
rect -2183 3072 -2083 3088
rect -2183 3038 -2167 3072
rect -2099 3038 -2083 3072
rect -2183 3000 -2083 3038
rect -2025 3072 -1925 3088
rect -2025 3038 -2009 3072
rect -1941 3038 -1925 3072
rect -2025 3000 -1925 3038
rect -1867 3072 -1767 3088
rect -1867 3038 -1851 3072
rect -1783 3038 -1767 3072
rect -1867 3000 -1767 3038
rect -1709 3072 -1609 3088
rect -1709 3038 -1693 3072
rect -1625 3038 -1609 3072
rect -1709 3000 -1609 3038
rect -1551 3072 -1451 3088
rect -1551 3038 -1535 3072
rect -1467 3038 -1451 3072
rect -1551 3000 -1451 3038
rect -1393 3072 -1293 3088
rect -1393 3038 -1377 3072
rect -1309 3038 -1293 3072
rect -1393 3000 -1293 3038
rect -1235 3072 -1135 3088
rect -1235 3038 -1219 3072
rect -1151 3038 -1135 3072
rect -1235 3000 -1135 3038
rect -1077 3072 -977 3088
rect -1077 3038 -1061 3072
rect -993 3038 -977 3072
rect -1077 3000 -977 3038
rect -919 3072 -819 3088
rect -919 3038 -903 3072
rect -835 3038 -819 3072
rect -919 3000 -819 3038
rect -761 3072 -661 3088
rect -761 3038 -745 3072
rect -677 3038 -661 3072
rect -761 3000 -661 3038
rect -603 3072 -503 3088
rect -603 3038 -587 3072
rect -519 3038 -503 3072
rect -603 3000 -503 3038
rect -445 3072 -345 3088
rect -445 3038 -429 3072
rect -361 3038 -345 3072
rect -445 3000 -345 3038
rect -287 3072 -187 3088
rect -287 3038 -271 3072
rect -203 3038 -187 3072
rect -287 3000 -187 3038
rect -129 3072 -29 3088
rect -129 3038 -113 3072
rect -45 3038 -29 3072
rect -129 3000 -29 3038
rect 29 3072 129 3088
rect 29 3038 45 3072
rect 113 3038 129 3072
rect 29 3000 129 3038
rect 187 3072 287 3088
rect 187 3038 203 3072
rect 271 3038 287 3072
rect 187 3000 287 3038
rect 345 3072 445 3088
rect 345 3038 361 3072
rect 429 3038 445 3072
rect 345 3000 445 3038
rect 503 3072 603 3088
rect 503 3038 519 3072
rect 587 3038 603 3072
rect 503 3000 603 3038
rect 661 3072 761 3088
rect 661 3038 677 3072
rect 745 3038 761 3072
rect 661 3000 761 3038
rect 819 3072 919 3088
rect 819 3038 835 3072
rect 903 3038 919 3072
rect 819 3000 919 3038
rect 977 3072 1077 3088
rect 977 3038 993 3072
rect 1061 3038 1077 3072
rect 977 3000 1077 3038
rect 1135 3072 1235 3088
rect 1135 3038 1151 3072
rect 1219 3038 1235 3072
rect 1135 3000 1235 3038
rect 1293 3072 1393 3088
rect 1293 3038 1309 3072
rect 1377 3038 1393 3072
rect 1293 3000 1393 3038
rect 1451 3072 1551 3088
rect 1451 3038 1467 3072
rect 1535 3038 1551 3072
rect 1451 3000 1551 3038
rect 1609 3072 1709 3088
rect 1609 3038 1625 3072
rect 1693 3038 1709 3072
rect 1609 3000 1709 3038
rect 1767 3072 1867 3088
rect 1767 3038 1783 3072
rect 1851 3038 1867 3072
rect 1767 3000 1867 3038
rect 1925 3072 2025 3088
rect 1925 3038 1941 3072
rect 2009 3038 2025 3072
rect 1925 3000 2025 3038
rect 2083 3072 2183 3088
rect 2083 3038 2099 3072
rect 2167 3038 2183 3072
rect 2083 3000 2183 3038
rect 2241 3072 2341 3088
rect 2241 3038 2257 3072
rect 2325 3038 2341 3072
rect 2241 3000 2341 3038
rect -2341 -3038 -2241 -3000
rect -2341 -3072 -2325 -3038
rect -2257 -3072 -2241 -3038
rect -2341 -3088 -2241 -3072
rect -2183 -3038 -2083 -3000
rect -2183 -3072 -2167 -3038
rect -2099 -3072 -2083 -3038
rect -2183 -3088 -2083 -3072
rect -2025 -3038 -1925 -3000
rect -2025 -3072 -2009 -3038
rect -1941 -3072 -1925 -3038
rect -2025 -3088 -1925 -3072
rect -1867 -3038 -1767 -3000
rect -1867 -3072 -1851 -3038
rect -1783 -3072 -1767 -3038
rect -1867 -3088 -1767 -3072
rect -1709 -3038 -1609 -3000
rect -1709 -3072 -1693 -3038
rect -1625 -3072 -1609 -3038
rect -1709 -3088 -1609 -3072
rect -1551 -3038 -1451 -3000
rect -1551 -3072 -1535 -3038
rect -1467 -3072 -1451 -3038
rect -1551 -3088 -1451 -3072
rect -1393 -3038 -1293 -3000
rect -1393 -3072 -1377 -3038
rect -1309 -3072 -1293 -3038
rect -1393 -3088 -1293 -3072
rect -1235 -3038 -1135 -3000
rect -1235 -3072 -1219 -3038
rect -1151 -3072 -1135 -3038
rect -1235 -3088 -1135 -3072
rect -1077 -3038 -977 -3000
rect -1077 -3072 -1061 -3038
rect -993 -3072 -977 -3038
rect -1077 -3088 -977 -3072
rect -919 -3038 -819 -3000
rect -919 -3072 -903 -3038
rect -835 -3072 -819 -3038
rect -919 -3088 -819 -3072
rect -761 -3038 -661 -3000
rect -761 -3072 -745 -3038
rect -677 -3072 -661 -3038
rect -761 -3088 -661 -3072
rect -603 -3038 -503 -3000
rect -603 -3072 -587 -3038
rect -519 -3072 -503 -3038
rect -603 -3088 -503 -3072
rect -445 -3038 -345 -3000
rect -445 -3072 -429 -3038
rect -361 -3072 -345 -3038
rect -445 -3088 -345 -3072
rect -287 -3038 -187 -3000
rect -287 -3072 -271 -3038
rect -203 -3072 -187 -3038
rect -287 -3088 -187 -3072
rect -129 -3038 -29 -3000
rect -129 -3072 -113 -3038
rect -45 -3072 -29 -3038
rect -129 -3088 -29 -3072
rect 29 -3038 129 -3000
rect 29 -3072 45 -3038
rect 113 -3072 129 -3038
rect 29 -3088 129 -3072
rect 187 -3038 287 -3000
rect 187 -3072 203 -3038
rect 271 -3072 287 -3038
rect 187 -3088 287 -3072
rect 345 -3038 445 -3000
rect 345 -3072 361 -3038
rect 429 -3072 445 -3038
rect 345 -3088 445 -3072
rect 503 -3038 603 -3000
rect 503 -3072 519 -3038
rect 587 -3072 603 -3038
rect 503 -3088 603 -3072
rect 661 -3038 761 -3000
rect 661 -3072 677 -3038
rect 745 -3072 761 -3038
rect 661 -3088 761 -3072
rect 819 -3038 919 -3000
rect 819 -3072 835 -3038
rect 903 -3072 919 -3038
rect 819 -3088 919 -3072
rect 977 -3038 1077 -3000
rect 977 -3072 993 -3038
rect 1061 -3072 1077 -3038
rect 977 -3088 1077 -3072
rect 1135 -3038 1235 -3000
rect 1135 -3072 1151 -3038
rect 1219 -3072 1235 -3038
rect 1135 -3088 1235 -3072
rect 1293 -3038 1393 -3000
rect 1293 -3072 1309 -3038
rect 1377 -3072 1393 -3038
rect 1293 -3088 1393 -3072
rect 1451 -3038 1551 -3000
rect 1451 -3072 1467 -3038
rect 1535 -3072 1551 -3038
rect 1451 -3088 1551 -3072
rect 1609 -3038 1709 -3000
rect 1609 -3072 1625 -3038
rect 1693 -3072 1709 -3038
rect 1609 -3088 1709 -3072
rect 1767 -3038 1867 -3000
rect 1767 -3072 1783 -3038
rect 1851 -3072 1867 -3038
rect 1767 -3088 1867 -3072
rect 1925 -3038 2025 -3000
rect 1925 -3072 1941 -3038
rect 2009 -3072 2025 -3038
rect 1925 -3088 2025 -3072
rect 2083 -3038 2183 -3000
rect 2083 -3072 2099 -3038
rect 2167 -3072 2183 -3038
rect 2083 -3088 2183 -3072
rect 2241 -3038 2341 -3000
rect 2241 -3072 2257 -3038
rect 2325 -3072 2341 -3038
rect 2241 -3088 2341 -3072
<< polycont >>
rect -2325 3038 -2257 3072
rect -2167 3038 -2099 3072
rect -2009 3038 -1941 3072
rect -1851 3038 -1783 3072
rect -1693 3038 -1625 3072
rect -1535 3038 -1467 3072
rect -1377 3038 -1309 3072
rect -1219 3038 -1151 3072
rect -1061 3038 -993 3072
rect -903 3038 -835 3072
rect -745 3038 -677 3072
rect -587 3038 -519 3072
rect -429 3038 -361 3072
rect -271 3038 -203 3072
rect -113 3038 -45 3072
rect 45 3038 113 3072
rect 203 3038 271 3072
rect 361 3038 429 3072
rect 519 3038 587 3072
rect 677 3038 745 3072
rect 835 3038 903 3072
rect 993 3038 1061 3072
rect 1151 3038 1219 3072
rect 1309 3038 1377 3072
rect 1467 3038 1535 3072
rect 1625 3038 1693 3072
rect 1783 3038 1851 3072
rect 1941 3038 2009 3072
rect 2099 3038 2167 3072
rect 2257 3038 2325 3072
rect -2325 -3072 -2257 -3038
rect -2167 -3072 -2099 -3038
rect -2009 -3072 -1941 -3038
rect -1851 -3072 -1783 -3038
rect -1693 -3072 -1625 -3038
rect -1535 -3072 -1467 -3038
rect -1377 -3072 -1309 -3038
rect -1219 -3072 -1151 -3038
rect -1061 -3072 -993 -3038
rect -903 -3072 -835 -3038
rect -745 -3072 -677 -3038
rect -587 -3072 -519 -3038
rect -429 -3072 -361 -3038
rect -271 -3072 -203 -3038
rect -113 -3072 -45 -3038
rect 45 -3072 113 -3038
rect 203 -3072 271 -3038
rect 361 -3072 429 -3038
rect 519 -3072 587 -3038
rect 677 -3072 745 -3038
rect 835 -3072 903 -3038
rect 993 -3072 1061 -3038
rect 1151 -3072 1219 -3038
rect 1309 -3072 1377 -3038
rect 1467 -3072 1535 -3038
rect 1625 -3072 1693 -3038
rect 1783 -3072 1851 -3038
rect 1941 -3072 2009 -3038
rect 2099 -3072 2167 -3038
rect 2257 -3072 2325 -3038
<< locali >>
rect -2521 3176 -2425 3210
rect 2425 3176 2521 3210
rect -2521 3114 -2487 3176
rect 2487 3114 2521 3176
rect -2341 3038 -2325 3072
rect -2257 3038 -2241 3072
rect -2183 3038 -2167 3072
rect -2099 3038 -2083 3072
rect -2025 3038 -2009 3072
rect -1941 3038 -1925 3072
rect -1867 3038 -1851 3072
rect -1783 3038 -1767 3072
rect -1709 3038 -1693 3072
rect -1625 3038 -1609 3072
rect -1551 3038 -1535 3072
rect -1467 3038 -1451 3072
rect -1393 3038 -1377 3072
rect -1309 3038 -1293 3072
rect -1235 3038 -1219 3072
rect -1151 3038 -1135 3072
rect -1077 3038 -1061 3072
rect -993 3038 -977 3072
rect -919 3038 -903 3072
rect -835 3038 -819 3072
rect -761 3038 -745 3072
rect -677 3038 -661 3072
rect -603 3038 -587 3072
rect -519 3038 -503 3072
rect -445 3038 -429 3072
rect -361 3038 -345 3072
rect -287 3038 -271 3072
rect -203 3038 -187 3072
rect -129 3038 -113 3072
rect -45 3038 -29 3072
rect 29 3038 45 3072
rect 113 3038 129 3072
rect 187 3038 203 3072
rect 271 3038 287 3072
rect 345 3038 361 3072
rect 429 3038 445 3072
rect 503 3038 519 3072
rect 587 3038 603 3072
rect 661 3038 677 3072
rect 745 3038 761 3072
rect 819 3038 835 3072
rect 903 3038 919 3072
rect 977 3038 993 3072
rect 1061 3038 1077 3072
rect 1135 3038 1151 3072
rect 1219 3038 1235 3072
rect 1293 3038 1309 3072
rect 1377 3038 1393 3072
rect 1451 3038 1467 3072
rect 1535 3038 1551 3072
rect 1609 3038 1625 3072
rect 1693 3038 1709 3072
rect 1767 3038 1783 3072
rect 1851 3038 1867 3072
rect 1925 3038 1941 3072
rect 2009 3038 2025 3072
rect 2083 3038 2099 3072
rect 2167 3038 2183 3072
rect 2241 3038 2257 3072
rect 2325 3038 2341 3072
rect -2387 2988 -2353 3004
rect -2387 -3004 -2353 -2988
rect -2229 2988 -2195 3004
rect -2229 -3004 -2195 -2988
rect -2071 2988 -2037 3004
rect -2071 -3004 -2037 -2988
rect -1913 2988 -1879 3004
rect -1913 -3004 -1879 -2988
rect -1755 2988 -1721 3004
rect -1755 -3004 -1721 -2988
rect -1597 2988 -1563 3004
rect -1597 -3004 -1563 -2988
rect -1439 2988 -1405 3004
rect -1439 -3004 -1405 -2988
rect -1281 2988 -1247 3004
rect -1281 -3004 -1247 -2988
rect -1123 2988 -1089 3004
rect -1123 -3004 -1089 -2988
rect -965 2988 -931 3004
rect -965 -3004 -931 -2988
rect -807 2988 -773 3004
rect -807 -3004 -773 -2988
rect -649 2988 -615 3004
rect -649 -3004 -615 -2988
rect -491 2988 -457 3004
rect -491 -3004 -457 -2988
rect -333 2988 -299 3004
rect -333 -3004 -299 -2988
rect -175 2988 -141 3004
rect -175 -3004 -141 -2988
rect -17 2988 17 3004
rect -17 -3004 17 -2988
rect 141 2988 175 3004
rect 141 -3004 175 -2988
rect 299 2988 333 3004
rect 299 -3004 333 -2988
rect 457 2988 491 3004
rect 457 -3004 491 -2988
rect 615 2988 649 3004
rect 615 -3004 649 -2988
rect 773 2988 807 3004
rect 773 -3004 807 -2988
rect 931 2988 965 3004
rect 931 -3004 965 -2988
rect 1089 2988 1123 3004
rect 1089 -3004 1123 -2988
rect 1247 2988 1281 3004
rect 1247 -3004 1281 -2988
rect 1405 2988 1439 3004
rect 1405 -3004 1439 -2988
rect 1563 2988 1597 3004
rect 1563 -3004 1597 -2988
rect 1721 2988 1755 3004
rect 1721 -3004 1755 -2988
rect 1879 2988 1913 3004
rect 1879 -3004 1913 -2988
rect 2037 2988 2071 3004
rect 2037 -3004 2071 -2988
rect 2195 2988 2229 3004
rect 2195 -3004 2229 -2988
rect 2353 2988 2387 3004
rect 2353 -3004 2387 -2988
rect -2341 -3072 -2325 -3038
rect -2257 -3072 -2241 -3038
rect -2183 -3072 -2167 -3038
rect -2099 -3072 -2083 -3038
rect -2025 -3072 -2009 -3038
rect -1941 -3072 -1925 -3038
rect -1867 -3072 -1851 -3038
rect -1783 -3072 -1767 -3038
rect -1709 -3072 -1693 -3038
rect -1625 -3072 -1609 -3038
rect -1551 -3072 -1535 -3038
rect -1467 -3072 -1451 -3038
rect -1393 -3072 -1377 -3038
rect -1309 -3072 -1293 -3038
rect -1235 -3072 -1219 -3038
rect -1151 -3072 -1135 -3038
rect -1077 -3072 -1061 -3038
rect -993 -3072 -977 -3038
rect -919 -3072 -903 -3038
rect -835 -3072 -819 -3038
rect -761 -3072 -745 -3038
rect -677 -3072 -661 -3038
rect -603 -3072 -587 -3038
rect -519 -3072 -503 -3038
rect -445 -3072 -429 -3038
rect -361 -3072 -345 -3038
rect -287 -3072 -271 -3038
rect -203 -3072 -187 -3038
rect -129 -3072 -113 -3038
rect -45 -3072 -29 -3038
rect 29 -3072 45 -3038
rect 113 -3072 129 -3038
rect 187 -3072 203 -3038
rect 271 -3072 287 -3038
rect 345 -3072 361 -3038
rect 429 -3072 445 -3038
rect 503 -3072 519 -3038
rect 587 -3072 603 -3038
rect 661 -3072 677 -3038
rect 745 -3072 761 -3038
rect 819 -3072 835 -3038
rect 903 -3072 919 -3038
rect 977 -3072 993 -3038
rect 1061 -3072 1077 -3038
rect 1135 -3072 1151 -3038
rect 1219 -3072 1235 -3038
rect 1293 -3072 1309 -3038
rect 1377 -3072 1393 -3038
rect 1451 -3072 1467 -3038
rect 1535 -3072 1551 -3038
rect 1609 -3072 1625 -3038
rect 1693 -3072 1709 -3038
rect 1767 -3072 1783 -3038
rect 1851 -3072 1867 -3038
rect 1925 -3072 1941 -3038
rect 2009 -3072 2025 -3038
rect 2083 -3072 2099 -3038
rect 2167 -3072 2183 -3038
rect 2241 -3072 2257 -3038
rect 2325 -3072 2341 -3038
rect -2521 -3176 -2487 -3114
rect 2487 -3176 2521 -3114
rect -2521 -3210 -2425 -3176
rect 2425 -3210 2521 -3176
<< viali >>
rect -2325 3038 -2257 3072
rect -2167 3038 -2099 3072
rect -2009 3038 -1941 3072
rect -1851 3038 -1783 3072
rect -1693 3038 -1625 3072
rect -1535 3038 -1467 3072
rect -1377 3038 -1309 3072
rect -1219 3038 -1151 3072
rect -1061 3038 -993 3072
rect -903 3038 -835 3072
rect -745 3038 -677 3072
rect -587 3038 -519 3072
rect -429 3038 -361 3072
rect -271 3038 -203 3072
rect -113 3038 -45 3072
rect 45 3038 113 3072
rect 203 3038 271 3072
rect 361 3038 429 3072
rect 519 3038 587 3072
rect 677 3038 745 3072
rect 835 3038 903 3072
rect 993 3038 1061 3072
rect 1151 3038 1219 3072
rect 1309 3038 1377 3072
rect 1467 3038 1535 3072
rect 1625 3038 1693 3072
rect 1783 3038 1851 3072
rect 1941 3038 2009 3072
rect 2099 3038 2167 3072
rect 2257 3038 2325 3072
rect -2387 -2988 -2353 2988
rect -2229 -2988 -2195 2988
rect -2071 -2988 -2037 2988
rect -1913 -2988 -1879 2988
rect -1755 -2988 -1721 2988
rect -1597 -2988 -1563 2988
rect -1439 -2988 -1405 2988
rect -1281 -2988 -1247 2988
rect -1123 -2988 -1089 2988
rect -965 -2988 -931 2988
rect -807 -2988 -773 2988
rect -649 -2988 -615 2988
rect -491 -2988 -457 2988
rect -333 -2988 -299 2988
rect -175 -2988 -141 2988
rect -17 -2988 17 2988
rect 141 -2988 175 2988
rect 299 -2988 333 2988
rect 457 -2988 491 2988
rect 615 -2988 649 2988
rect 773 -2988 807 2988
rect 931 -2988 965 2988
rect 1089 -2988 1123 2988
rect 1247 -2988 1281 2988
rect 1405 -2988 1439 2988
rect 1563 -2988 1597 2988
rect 1721 -2988 1755 2988
rect 1879 -2988 1913 2988
rect 2037 -2988 2071 2988
rect 2195 -2988 2229 2988
rect 2353 -2988 2387 2988
rect -2325 -3072 -2257 -3038
rect -2167 -3072 -2099 -3038
rect -2009 -3072 -1941 -3038
rect -1851 -3072 -1783 -3038
rect -1693 -3072 -1625 -3038
rect -1535 -3072 -1467 -3038
rect -1377 -3072 -1309 -3038
rect -1219 -3072 -1151 -3038
rect -1061 -3072 -993 -3038
rect -903 -3072 -835 -3038
rect -745 -3072 -677 -3038
rect -587 -3072 -519 -3038
rect -429 -3072 -361 -3038
rect -271 -3072 -203 -3038
rect -113 -3072 -45 -3038
rect 45 -3072 113 -3038
rect 203 -3072 271 -3038
rect 361 -3072 429 -3038
rect 519 -3072 587 -3038
rect 677 -3072 745 -3038
rect 835 -3072 903 -3038
rect 993 -3072 1061 -3038
rect 1151 -3072 1219 -3038
rect 1309 -3072 1377 -3038
rect 1467 -3072 1535 -3038
rect 1625 -3072 1693 -3038
rect 1783 -3072 1851 -3038
rect 1941 -3072 2009 -3038
rect 2099 -3072 2167 -3038
rect 2257 -3072 2325 -3038
<< metal1 >>
rect -2337 3072 -2245 3078
rect -2337 3038 -2325 3072
rect -2257 3038 -2245 3072
rect -2337 3032 -2245 3038
rect -2179 3072 -2087 3078
rect -2179 3038 -2167 3072
rect -2099 3038 -2087 3072
rect -2179 3032 -2087 3038
rect -2021 3072 -1929 3078
rect -2021 3038 -2009 3072
rect -1941 3038 -1929 3072
rect -2021 3032 -1929 3038
rect -1863 3072 -1771 3078
rect -1863 3038 -1851 3072
rect -1783 3038 -1771 3072
rect -1863 3032 -1771 3038
rect -1705 3072 -1613 3078
rect -1705 3038 -1693 3072
rect -1625 3038 -1613 3072
rect -1705 3032 -1613 3038
rect -1547 3072 -1455 3078
rect -1547 3038 -1535 3072
rect -1467 3038 -1455 3072
rect -1547 3032 -1455 3038
rect -1389 3072 -1297 3078
rect -1389 3038 -1377 3072
rect -1309 3038 -1297 3072
rect -1389 3032 -1297 3038
rect -1231 3072 -1139 3078
rect -1231 3038 -1219 3072
rect -1151 3038 -1139 3072
rect -1231 3032 -1139 3038
rect -1073 3072 -981 3078
rect -1073 3038 -1061 3072
rect -993 3038 -981 3072
rect -1073 3032 -981 3038
rect -915 3072 -823 3078
rect -915 3038 -903 3072
rect -835 3038 -823 3072
rect -915 3032 -823 3038
rect -757 3072 -665 3078
rect -757 3038 -745 3072
rect -677 3038 -665 3072
rect -757 3032 -665 3038
rect -599 3072 -507 3078
rect -599 3038 -587 3072
rect -519 3038 -507 3072
rect -599 3032 -507 3038
rect -441 3072 -349 3078
rect -441 3038 -429 3072
rect -361 3038 -349 3072
rect -441 3032 -349 3038
rect -283 3072 -191 3078
rect -283 3038 -271 3072
rect -203 3038 -191 3072
rect -283 3032 -191 3038
rect -125 3072 -33 3078
rect -125 3038 -113 3072
rect -45 3038 -33 3072
rect -125 3032 -33 3038
rect 33 3072 125 3078
rect 33 3038 45 3072
rect 113 3038 125 3072
rect 33 3032 125 3038
rect 191 3072 283 3078
rect 191 3038 203 3072
rect 271 3038 283 3072
rect 191 3032 283 3038
rect 349 3072 441 3078
rect 349 3038 361 3072
rect 429 3038 441 3072
rect 349 3032 441 3038
rect 507 3072 599 3078
rect 507 3038 519 3072
rect 587 3038 599 3072
rect 507 3032 599 3038
rect 665 3072 757 3078
rect 665 3038 677 3072
rect 745 3038 757 3072
rect 665 3032 757 3038
rect 823 3072 915 3078
rect 823 3038 835 3072
rect 903 3038 915 3072
rect 823 3032 915 3038
rect 981 3072 1073 3078
rect 981 3038 993 3072
rect 1061 3038 1073 3072
rect 981 3032 1073 3038
rect 1139 3072 1231 3078
rect 1139 3038 1151 3072
rect 1219 3038 1231 3072
rect 1139 3032 1231 3038
rect 1297 3072 1389 3078
rect 1297 3038 1309 3072
rect 1377 3038 1389 3072
rect 1297 3032 1389 3038
rect 1455 3072 1547 3078
rect 1455 3038 1467 3072
rect 1535 3038 1547 3072
rect 1455 3032 1547 3038
rect 1613 3072 1705 3078
rect 1613 3038 1625 3072
rect 1693 3038 1705 3072
rect 1613 3032 1705 3038
rect 1771 3072 1863 3078
rect 1771 3038 1783 3072
rect 1851 3038 1863 3072
rect 1771 3032 1863 3038
rect 1929 3072 2021 3078
rect 1929 3038 1941 3072
rect 2009 3038 2021 3072
rect 1929 3032 2021 3038
rect 2087 3072 2179 3078
rect 2087 3038 2099 3072
rect 2167 3038 2179 3072
rect 2087 3032 2179 3038
rect 2245 3072 2337 3078
rect 2245 3038 2257 3072
rect 2325 3038 2337 3072
rect 2245 3032 2337 3038
rect -2393 2988 -2347 3000
rect -2393 -2988 -2387 2988
rect -2353 -2988 -2347 2988
rect -2393 -3000 -2347 -2988
rect -2235 2988 -2189 3000
rect -2235 -2988 -2229 2988
rect -2195 -2988 -2189 2988
rect -2235 -3000 -2189 -2988
rect -2077 2988 -2031 3000
rect -2077 -2988 -2071 2988
rect -2037 -2988 -2031 2988
rect -2077 -3000 -2031 -2988
rect -1919 2988 -1873 3000
rect -1919 -2988 -1913 2988
rect -1879 -2988 -1873 2988
rect -1919 -3000 -1873 -2988
rect -1761 2988 -1715 3000
rect -1761 -2988 -1755 2988
rect -1721 -2988 -1715 2988
rect -1761 -3000 -1715 -2988
rect -1603 2988 -1557 3000
rect -1603 -2988 -1597 2988
rect -1563 -2988 -1557 2988
rect -1603 -3000 -1557 -2988
rect -1445 2988 -1399 3000
rect -1445 -2988 -1439 2988
rect -1405 -2988 -1399 2988
rect -1445 -3000 -1399 -2988
rect -1287 2988 -1241 3000
rect -1287 -2988 -1281 2988
rect -1247 -2988 -1241 2988
rect -1287 -3000 -1241 -2988
rect -1129 2988 -1083 3000
rect -1129 -2988 -1123 2988
rect -1089 -2988 -1083 2988
rect -1129 -3000 -1083 -2988
rect -971 2988 -925 3000
rect -971 -2988 -965 2988
rect -931 -2988 -925 2988
rect -971 -3000 -925 -2988
rect -813 2988 -767 3000
rect -813 -2988 -807 2988
rect -773 -2988 -767 2988
rect -813 -3000 -767 -2988
rect -655 2988 -609 3000
rect -655 -2988 -649 2988
rect -615 -2988 -609 2988
rect -655 -3000 -609 -2988
rect -497 2988 -451 3000
rect -497 -2988 -491 2988
rect -457 -2988 -451 2988
rect -497 -3000 -451 -2988
rect -339 2988 -293 3000
rect -339 -2988 -333 2988
rect -299 -2988 -293 2988
rect -339 -3000 -293 -2988
rect -181 2988 -135 3000
rect -181 -2988 -175 2988
rect -141 -2988 -135 2988
rect -181 -3000 -135 -2988
rect -23 2988 23 3000
rect -23 -2988 -17 2988
rect 17 -2988 23 2988
rect -23 -3000 23 -2988
rect 135 2988 181 3000
rect 135 -2988 141 2988
rect 175 -2988 181 2988
rect 135 -3000 181 -2988
rect 293 2988 339 3000
rect 293 -2988 299 2988
rect 333 -2988 339 2988
rect 293 -3000 339 -2988
rect 451 2988 497 3000
rect 451 -2988 457 2988
rect 491 -2988 497 2988
rect 451 -3000 497 -2988
rect 609 2988 655 3000
rect 609 -2988 615 2988
rect 649 -2988 655 2988
rect 609 -3000 655 -2988
rect 767 2988 813 3000
rect 767 -2988 773 2988
rect 807 -2988 813 2988
rect 767 -3000 813 -2988
rect 925 2988 971 3000
rect 925 -2988 931 2988
rect 965 -2988 971 2988
rect 925 -3000 971 -2988
rect 1083 2988 1129 3000
rect 1083 -2988 1089 2988
rect 1123 -2988 1129 2988
rect 1083 -3000 1129 -2988
rect 1241 2988 1287 3000
rect 1241 -2988 1247 2988
rect 1281 -2988 1287 2988
rect 1241 -3000 1287 -2988
rect 1399 2988 1445 3000
rect 1399 -2988 1405 2988
rect 1439 -2988 1445 2988
rect 1399 -3000 1445 -2988
rect 1557 2988 1603 3000
rect 1557 -2988 1563 2988
rect 1597 -2988 1603 2988
rect 1557 -3000 1603 -2988
rect 1715 2988 1761 3000
rect 1715 -2988 1721 2988
rect 1755 -2988 1761 2988
rect 1715 -3000 1761 -2988
rect 1873 2988 1919 3000
rect 1873 -2988 1879 2988
rect 1913 -2988 1919 2988
rect 1873 -3000 1919 -2988
rect 2031 2988 2077 3000
rect 2031 -2988 2037 2988
rect 2071 -2988 2077 2988
rect 2031 -3000 2077 -2988
rect 2189 2988 2235 3000
rect 2189 -2988 2195 2988
rect 2229 -2988 2235 2988
rect 2189 -3000 2235 -2988
rect 2347 2988 2393 3000
rect 2347 -2988 2353 2988
rect 2387 -2988 2393 2988
rect 2347 -3000 2393 -2988
rect -2337 -3038 -2245 -3032
rect -2337 -3072 -2325 -3038
rect -2257 -3072 -2245 -3038
rect -2337 -3078 -2245 -3072
rect -2179 -3038 -2087 -3032
rect -2179 -3072 -2167 -3038
rect -2099 -3072 -2087 -3038
rect -2179 -3078 -2087 -3072
rect -2021 -3038 -1929 -3032
rect -2021 -3072 -2009 -3038
rect -1941 -3072 -1929 -3038
rect -2021 -3078 -1929 -3072
rect -1863 -3038 -1771 -3032
rect -1863 -3072 -1851 -3038
rect -1783 -3072 -1771 -3038
rect -1863 -3078 -1771 -3072
rect -1705 -3038 -1613 -3032
rect -1705 -3072 -1693 -3038
rect -1625 -3072 -1613 -3038
rect -1705 -3078 -1613 -3072
rect -1547 -3038 -1455 -3032
rect -1547 -3072 -1535 -3038
rect -1467 -3072 -1455 -3038
rect -1547 -3078 -1455 -3072
rect -1389 -3038 -1297 -3032
rect -1389 -3072 -1377 -3038
rect -1309 -3072 -1297 -3038
rect -1389 -3078 -1297 -3072
rect -1231 -3038 -1139 -3032
rect -1231 -3072 -1219 -3038
rect -1151 -3072 -1139 -3038
rect -1231 -3078 -1139 -3072
rect -1073 -3038 -981 -3032
rect -1073 -3072 -1061 -3038
rect -993 -3072 -981 -3038
rect -1073 -3078 -981 -3072
rect -915 -3038 -823 -3032
rect -915 -3072 -903 -3038
rect -835 -3072 -823 -3038
rect -915 -3078 -823 -3072
rect -757 -3038 -665 -3032
rect -757 -3072 -745 -3038
rect -677 -3072 -665 -3038
rect -757 -3078 -665 -3072
rect -599 -3038 -507 -3032
rect -599 -3072 -587 -3038
rect -519 -3072 -507 -3038
rect -599 -3078 -507 -3072
rect -441 -3038 -349 -3032
rect -441 -3072 -429 -3038
rect -361 -3072 -349 -3038
rect -441 -3078 -349 -3072
rect -283 -3038 -191 -3032
rect -283 -3072 -271 -3038
rect -203 -3072 -191 -3038
rect -283 -3078 -191 -3072
rect -125 -3038 -33 -3032
rect -125 -3072 -113 -3038
rect -45 -3072 -33 -3038
rect -125 -3078 -33 -3072
rect 33 -3038 125 -3032
rect 33 -3072 45 -3038
rect 113 -3072 125 -3038
rect 33 -3078 125 -3072
rect 191 -3038 283 -3032
rect 191 -3072 203 -3038
rect 271 -3072 283 -3038
rect 191 -3078 283 -3072
rect 349 -3038 441 -3032
rect 349 -3072 361 -3038
rect 429 -3072 441 -3038
rect 349 -3078 441 -3072
rect 507 -3038 599 -3032
rect 507 -3072 519 -3038
rect 587 -3072 599 -3038
rect 507 -3078 599 -3072
rect 665 -3038 757 -3032
rect 665 -3072 677 -3038
rect 745 -3072 757 -3038
rect 665 -3078 757 -3072
rect 823 -3038 915 -3032
rect 823 -3072 835 -3038
rect 903 -3072 915 -3038
rect 823 -3078 915 -3072
rect 981 -3038 1073 -3032
rect 981 -3072 993 -3038
rect 1061 -3072 1073 -3038
rect 981 -3078 1073 -3072
rect 1139 -3038 1231 -3032
rect 1139 -3072 1151 -3038
rect 1219 -3072 1231 -3038
rect 1139 -3078 1231 -3072
rect 1297 -3038 1389 -3032
rect 1297 -3072 1309 -3038
rect 1377 -3072 1389 -3038
rect 1297 -3078 1389 -3072
rect 1455 -3038 1547 -3032
rect 1455 -3072 1467 -3038
rect 1535 -3072 1547 -3038
rect 1455 -3078 1547 -3072
rect 1613 -3038 1705 -3032
rect 1613 -3072 1625 -3038
rect 1693 -3072 1705 -3038
rect 1613 -3078 1705 -3072
rect 1771 -3038 1863 -3032
rect 1771 -3072 1783 -3038
rect 1851 -3072 1863 -3038
rect 1771 -3078 1863 -3072
rect 1929 -3038 2021 -3032
rect 1929 -3072 1941 -3038
rect 2009 -3072 2021 -3038
rect 1929 -3078 2021 -3072
rect 2087 -3038 2179 -3032
rect 2087 -3072 2099 -3038
rect 2167 -3072 2179 -3038
rect 2087 -3078 2179 -3072
rect 2245 -3038 2337 -3032
rect 2245 -3072 2257 -3038
rect 2325 -3072 2337 -3038
rect 2245 -3078 2337 -3072
<< properties >>
string FIXED_BBOX -2504 -3193 2504 3193
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 30 l 0.50 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
