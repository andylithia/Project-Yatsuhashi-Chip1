magic
tech sky130B
magscale 1 2
timestamp 1659297343
<< psubdiff >>
rect 592 156 744 1166
rect 1252 156 1404 1166
<< metal1 >>
rect 570 1270 770 1280
rect 570 1258 580 1270
rect 165 1210 580 1258
rect 760 1258 770 1270
rect 1230 1270 1430 1280
rect 1230 1258 1240 1270
rect 760 1210 1240 1258
rect 1420 1258 1430 1270
rect 1420 1210 1831 1258
rect 165 1192 1831 1210
rect 0 1140 80 1150
rect 0 180 10 1140
rect 70 180 80 1140
rect 0 170 80 180
rect 592 952 744 1158
rect 592 370 598 952
rect 738 370 744 952
rect 592 164 744 370
rect 1252 952 1404 1158
rect 1252 370 1258 952
rect 1398 370 1404 952
rect 1252 164 1404 370
rect 1920 1140 2000 1150
rect 1920 180 1930 1140
rect 1990 180 2000 1140
rect 1920 170 2000 180
rect 506 120 1495 130
rect 506 64 580 120
rect 570 60 580 64
rect 760 64 1240 120
rect 760 60 770 64
rect 570 50 770 60
rect 1230 60 1240 64
rect 1420 64 1495 120
rect 1420 60 1430 64
rect 1230 50 1430 60
<< via1 >>
rect 580 1210 760 1270
rect 1240 1210 1420 1270
rect 10 180 70 1140
rect 598 370 738 952
rect 1258 370 1398 952
rect 1930 180 1990 1140
rect 580 60 760 120
rect 1240 60 1420 120
<< metal2 >>
rect 220 1370 460 1380
rect 220 1280 230 1370
rect 450 1280 460 1370
rect 880 1370 1120 1380
rect 220 1270 460 1280
rect 570 1300 770 1310
rect 570 1210 580 1300
rect 760 1210 770 1300
rect 880 1280 890 1370
rect 1110 1280 1120 1370
rect 1540 1370 1780 1380
rect 880 1270 1120 1280
rect 1230 1300 1430 1310
rect 570 1200 770 1210
rect 1230 1210 1240 1300
rect 1420 1210 1430 1300
rect 1540 1280 1550 1370
rect 1770 1280 1780 1370
rect 1540 1270 1780 1280
rect 1230 1200 1430 1210
rect 0 1140 80 1150
rect 0 750 10 1140
rect 0 180 10 610
rect 70 180 80 1140
rect 1920 1140 2000 1150
rect 592 952 744 980
rect 592 370 598 952
rect 738 370 744 952
rect 592 340 744 370
rect 1252 952 1404 980
rect 1252 370 1258 952
rect 1398 370 1404 952
rect 1252 340 1404 370
rect 0 170 80 180
rect 1920 180 1930 1140
rect 1990 750 2000 1140
rect 1990 180 2000 610
rect 1920 170 2000 180
rect 570 120 770 130
rect 220 40 460 50
rect 220 -50 230 40
rect 450 -50 460 40
rect 570 30 580 120
rect 760 30 770 120
rect 1230 120 1430 130
rect 570 20 770 30
rect 880 40 1120 50
rect 220 -60 460 -50
rect 880 -50 890 40
rect 1110 -50 1120 40
rect 1230 30 1240 120
rect 1420 30 1430 120
rect 1230 20 1430 30
rect 1540 40 1780 50
rect 880 -60 1120 -50
rect 1540 -50 1550 40
rect 1770 -50 1780 40
rect 1540 -60 1780 -50
<< via2 >>
rect 230 1280 450 1370
rect 580 1270 760 1300
rect 580 1210 760 1270
rect 890 1280 1110 1370
rect 1240 1270 1420 1300
rect 1240 1210 1420 1270
rect 1550 1280 1770 1370
rect 0 610 10 750
rect 10 610 70 750
rect 600 620 730 740
rect 1260 620 1390 740
rect 1930 610 1990 750
rect 1990 610 2000 750
rect 230 -50 450 40
rect 580 60 760 120
rect 580 30 760 60
rect 890 -50 1110 40
rect 1240 60 1420 120
rect 1240 30 1420 60
rect 1550 -50 1770 40
<< metal3 >>
rect 220 1490 1780 1500
rect 220 1390 240 1490
rect 1760 1390 1780 1490
rect 220 1380 1780 1390
rect 220 1370 460 1380
rect 220 1280 230 1370
rect 450 1280 460 1370
rect 880 1370 1120 1380
rect 220 1270 460 1280
rect 570 1300 770 1310
rect 570 1210 580 1300
rect 760 1210 770 1300
rect 880 1280 890 1370
rect 1110 1280 1120 1370
rect 1540 1370 1780 1380
rect 880 1270 1120 1280
rect 1230 1300 1430 1310
rect 570 1130 770 1210
rect 1230 1210 1240 1300
rect 1420 1210 1430 1300
rect 1540 1280 1550 1370
rect 1770 1280 1780 1370
rect 1540 1270 1780 1280
rect 1230 1130 1430 1210
rect 570 970 1430 1130
rect -10 750 80 760
rect -10 610 0 750
rect 70 610 80 750
rect -10 600 80 610
rect 592 740 744 760
rect 592 620 600 740
rect 730 620 744 740
rect 592 600 744 620
rect 1252 740 1404 760
rect 1252 620 1260 740
rect 1390 620 1404 740
rect 1252 600 1404 620
rect 1920 750 2010 760
rect 1920 610 1930 750
rect 2000 610 2010 750
rect 1920 600 2010 610
rect 570 200 1430 360
rect 570 120 770 200
rect 220 40 460 50
rect 220 -50 230 40
rect 450 -50 460 40
rect 570 30 580 120
rect 760 30 770 120
rect 1230 120 1430 200
rect 570 20 770 30
rect 880 40 1120 50
rect 220 -60 460 -50
rect 880 -50 890 40
rect 1110 -50 1120 40
rect 1230 30 1240 120
rect 1420 30 1430 120
rect 1230 20 1430 30
rect 1540 40 1780 50
rect 880 -60 1120 -50
rect 1540 -50 1550 40
rect 1770 -50 1780 40
rect 1540 -60 1780 -50
rect 220 -70 1780 -60
rect 220 -170 240 -70
rect 1760 -170 1780 -70
rect 220 -180 1780 -170
<< via3 >>
rect 240 1390 1760 1490
rect 0 610 70 750
rect 600 620 730 740
rect 1260 620 1390 740
rect 1930 610 2000 750
rect 240 -170 1760 -70
<< metal4 >>
rect 220 1490 1780 1500
rect 220 1390 240 1490
rect 1760 1390 1780 1490
rect 220 1380 1780 1390
rect -10 750 80 760
rect 1920 750 2010 760
rect -10 610 0 750
rect 70 740 1930 750
rect 70 620 600 740
rect 730 620 1260 740
rect 1390 620 1930 740
rect 70 610 1930 620
rect 2000 610 2010 750
rect -10 600 80 610
rect 1920 600 2010 610
rect 220 -70 1780 -60
rect 220 -170 240 -70
rect 1760 -170 1780 -70
rect 220 -180 1780 -170
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_0
timestamp 1659146707
transform 1 0 0 0 1 64
box 0 -64 676 1258
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_1
timestamp 1659146707
transform 1 0 660 0 1 64
box 0 -64 676 1258
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2
timestamp 1659146707
transform 1 0 1320 0 1 64
box 0 -64 676 1258
<< labels >>
rlabel metal3 570 970 1430 1130 1 G1
rlabel metal3 570 200 1430 360 1 G2
rlabel metal4 -10 600 90 760 1 SUB
rlabel metal4 220 1380 1780 1500 1 SD1
rlabel metal4 220 -180 1780 -60 1 SD2
<< end >>
