magic
tech sky130B
timestamp 1659241375
<< metal4 >>
rect 6100 3950 6800 4000
rect -200 3750 4550 3800
rect -200 3050 -150 3750
rect 450 3050 4550 3750
rect -200 3000 4550 3050
rect 3850 -100 4550 3000
rect 6100 3250 6150 3950
rect 6750 3250 6800 3950
rect 6100 -100 6800 3250
<< via4 >>
rect -150 3050 450 3750
rect 6150 3250 6750 3950
<< metal5 >>
rect 0 9500 10000 10000
rect 0 3950 500 9500
rect -50 3900 500 3950
rect -100 3850 500 3900
rect -150 3800 500 3850
rect -200 3750 500 3800
rect -200 3050 -150 3750
rect 450 3050 500 3750
rect -200 3000 500 3050
rect 800 8700 9200 9200
rect 800 500 1300 8700
rect 1600 7900 8400 8400
rect 1600 1300 2100 7900
rect 2400 7100 7600 7600
rect 2400 2100 2900 7100
rect 3200 6300 6800 6800
rect 3200 2900 3700 6300
rect 6300 4150 6800 6300
rect 6250 4100 6800 4150
rect 6200 4050 6800 4100
rect 6150 4000 6800 4050
rect 6100 3950 6800 4000
rect 6100 3250 6150 3950
rect 6750 3250 6800 3950
rect 6100 3200 6800 3250
rect 7100 2900 7600 7100
rect 3200 2400 7600 2900
rect 7900 2100 8400 7900
rect 2400 1600 8400 2100
rect 8700 1300 9200 8700
rect 1600 800 9200 1300
rect 9500 500 10000 9500
rect 800 0 10000 500
<< labels >>
rlabel metal4 3850 -100 4550 0 1 A
rlabel metal4 6100 -100 6800 0 1 B
<< end >>
