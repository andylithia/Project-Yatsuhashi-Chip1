magic
tech sky130B
magscale 1 2
timestamp 1660705385
<< locali >>
rect 1430 9590 1530 9620
rect 678 9488 1320 9522
rect 1430 7830 1440 9590
rect 1500 7830 1530 9590
rect 582 7778 1224 7812
rect 1430 7710 1530 7830
rect 430 7700 1530 7710
rect 430 7650 470 7700
rect 1430 7650 1530 7700
rect 430 7640 1530 7650
<< viali >>
rect 1440 7830 1500 9590
rect 470 7650 1430 7700
<< metal1 >>
rect 1430 9590 1530 9620
rect 660 9550 1320 9560
rect 660 9490 670 9550
rect 1310 9490 1320 9550
rect 660 9480 1320 9490
rect 540 9410 600 9450
rect 540 7850 600 7890
rect 630 9410 690 9450
rect 630 7850 690 7890
rect 730 9410 790 9450
rect 730 7850 790 7890
rect 830 9410 890 9450
rect 830 7850 890 7890
rect 920 9410 980 9450
rect 920 7850 980 7890
rect 1020 9410 1080 9450
rect 1020 7850 1080 7890
rect 1110 9410 1170 9450
rect 1110 7850 1170 7890
rect 1210 9410 1270 9450
rect 1210 7850 1270 7890
rect 1310 9410 1370 9450
rect 1310 7850 1370 7890
rect 1430 7830 1440 9590
rect 1500 7830 1530 9590
rect 570 7810 1230 7820
rect 570 7750 580 7810
rect 1220 7750 1230 7810
rect 570 7740 1230 7750
rect 1430 7710 1530 7830
rect 430 7700 1530 7710
rect 430 7650 470 7700
rect 1430 7650 1530 7700
rect 430 7640 1530 7650
<< via1 >>
rect 670 9490 1310 9550
rect 540 7890 600 9410
rect 630 7890 690 9410
rect 730 7890 790 9410
rect 830 7890 890 9410
rect 920 7890 980 9410
rect 1020 7890 1080 9410
rect 1110 7890 1170 9410
rect 1210 7890 1270 9410
rect 1310 7890 1370 9410
rect 580 7750 1220 7810
<< metal2 >>
rect 630 9550 1320 9560
rect 630 9490 670 9550
rect 1310 9490 1320 9550
rect 630 9480 1320 9490
rect 540 9410 600 9450
rect 540 7850 600 7890
rect 630 9410 690 9480
rect 630 7820 690 7890
rect 730 9410 790 9450
rect 730 7850 790 7890
rect 830 9410 890 9480
rect 830 7820 890 7890
rect 920 9410 980 9450
rect 920 7850 980 7890
rect 1020 9410 1080 9480
rect 1020 7820 1080 7890
rect 1110 9410 1170 9450
rect 1110 7850 1170 7890
rect 1210 9410 1270 9480
rect 1210 7820 1270 7890
rect 1310 9410 1370 9450
rect 1310 7850 1370 7890
rect 570 7810 1270 7820
rect 570 7750 580 7810
rect 1220 7750 1270 7810
rect 570 7740 1270 7750
<< via2 >>
rect 670 9490 1310 9550
rect 540 8270 600 9030
rect 730 8270 790 9030
rect 920 8270 980 9030
rect 1110 8270 1170 9030
rect 1310 8270 1370 9030
rect 580 7750 1220 7810
<< metal3 >>
rect 340 9550 1320 9560
rect 340 9490 670 9550
rect 1310 9490 1320 9550
rect 340 9480 1320 9490
rect 340 7820 420 9480
rect 1500 9060 1560 9100
rect 1440 9050 1560 9060
rect 520 9030 1560 9050
rect 520 8270 540 9030
rect 600 8980 730 9030
rect 600 8700 620 8980
rect 710 8700 730 8980
rect 600 8620 730 8700
rect 600 8320 620 8620
rect 710 8320 730 8620
rect 600 8270 730 8320
rect 790 8980 920 9030
rect 790 8700 810 8980
rect 900 8700 920 8980
rect 790 8620 920 8700
rect 790 8320 810 8620
rect 900 8320 920 8620
rect 790 8270 920 8320
rect 980 8980 1110 9030
rect 980 8700 1000 8980
rect 1090 8700 1110 8980
rect 980 8620 1110 8700
rect 980 8320 1000 8620
rect 1090 8320 1110 8620
rect 980 8270 1110 8320
rect 1170 8980 1310 9030
rect 1170 8700 1190 8980
rect 1290 8700 1310 8980
rect 1170 8620 1310 8700
rect 1170 8320 1190 8620
rect 1290 8320 1310 8620
rect 1170 8270 1310 8320
rect 1370 8980 1560 9030
rect 1370 8700 1390 8980
rect 1460 8700 1560 8980
rect 1370 8620 1560 8700
rect 1370 8320 1390 8620
rect 1460 8320 1560 8620
rect 1370 8270 1560 8320
rect 520 8250 1560 8270
rect 1440 8240 1560 8250
rect 340 7810 1230 7820
rect 340 7750 580 7810
rect 1220 7750 1230 7810
rect 340 7740 1230 7750
rect 1460 7640 1560 8240
rect 1500 7600 1560 7640
use sky130_fd_pr__nfet_01v8_6H2JGK  sky130_fd_pr__nfet_01v8_6H2JGK_0
timestamp 1660448881
transform 1 0 951 0 1 8650
box -551 -1010 551 1010
<< labels >>
rlabel metal3 420 9480 1320 9560 1 IREF_L
rlabel metal3 1500 7600 1560 9100 1 GND
<< end >>
