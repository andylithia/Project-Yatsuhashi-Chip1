magic
tech sky130A
magscale 1 2
timestamp 1665269856
<< metal4 >>
rect -64700 -7112 -33500 -7000
rect -64700 -13888 -64588 -7112
rect -57812 -13888 -40388 -7112
rect -33612 -13888 -33500 -7112
rect -64700 -14000 -33500 -13888
<< via4 >>
rect -64588 -13888 -57812 -7112
rect -40388 -13888 -33612 -7112
<< metal5 >>
tri -31400 51962 -30862 52500 se
rect -30862 51962 23062 52500
tri 23062 51962 23600 52500 sw
tri -37862 45500 -31400 51962 se
rect -31400 45500 23600 51962
tri 23600 45500 30062 51962 sw
tri -41300 42062 -37862 45500 se
rect -37862 44700 -28762 45500
tri -28762 44700 -27962 45500 nw
tri 20162 44700 20962 45500 ne
rect 20962 44700 30062 45500
rect -37862 43569 -29893 44700
tri -29893 43569 -28762 44700 nw
tri -28762 43569 -27631 44700 se
rect -27631 43569 19831 44700
tri 19831 43569 20962 44700 sw
tri 20962 43569 22093 44700 ne
rect 22093 43569 30062 44700
rect -37862 43193 -30269 43569
tri -30269 43193 -29893 43569 nw
tri -29138 43193 -28762 43569 se
rect -28762 43193 20962 43569
rect -37862 42062 -31400 43193
tri -31400 42062 -30269 43193 nw
tri -30269 42062 -29138 43193 se
rect -29138 42438 20962 43193
tri 20962 42438 22093 43569 sw
tri 22093 42438 23224 43569 ne
rect 23224 42438 30062 43569
rect -29138 42062 22093 42438
tri -49100 34262 -41300 42062 se
rect -41300 40931 -32531 42062
tri -32531 40931 -31400 42062 nw
tri -31400 40931 -30269 42062 se
rect -30269 41307 22093 42062
tri 22093 41307 23224 42438 sw
tri 23224 41307 24355 42438 ne
rect 24355 41307 30062 42438
rect -30269 41093 23224 41307
tri 23224 41093 23438 41307 sw
tri 24355 41093 24569 41307 ne
rect 24569 41093 30062 41307
rect -30269 40931 23438 41093
tri 23438 40931 23600 41093 sw
tri 24569 40931 24731 41093 ne
rect 24731 40931 30062 41093
rect -41300 39800 -33662 40931
tri -33662 39800 -32531 40931 nw
tri -32531 39800 -31400 40931 se
rect -31400 39962 23600 40931
tri 23600 39962 24569 40931 sw
tri 24731 39962 25700 40931 ne
rect 25700 39962 30062 40931
rect -31400 39800 24569 39962
rect -41300 38831 -34631 39800
tri -34631 38831 -33662 39800 nw
tri -33500 38831 -32531 39800 se
rect -32531 38831 24569 39800
tri 24569 38831 25700 39962 sw
tri 25700 38831 26831 39962 ne
rect 26831 38831 30062 39962
rect -41300 37700 -35762 38831
tri -35762 37700 -34631 38831 nw
tri -34631 37700 -33500 38831 se
rect -33500 37700 25700 38831
tri 25700 37700 26831 38831 sw
tri 26831 37700 27962 38831 ne
rect 27962 37700 30062 38831
tri 30062 37700 37862 45500 sw
rect -41300 36569 -36893 37700
tri -36893 36569 -35762 37700 nw
tri -35762 36569 -34631 37700 se
rect -34631 36900 -25531 37700
tri -25531 36900 -24731 37700 nw
tri 16931 36900 17731 37700 ne
rect 17731 36900 26831 37700
rect -34631 36569 -26662 36900
rect -41300 35438 -38024 36569
tri -38024 35438 -36893 36569 nw
tri -36893 35438 -35762 36569 se
rect -35762 35769 -26662 36569
tri -26662 35769 -25531 36900 nw
tri -25531 35769 -24400 36900 se
rect -24400 35769 16600 36900
tri 16600 35769 17731 36900 sw
tri 17731 35769 18862 36900 ne
rect 18862 36569 26831 36900
tri 26831 36569 27962 37700 sw
tri 27962 36569 29093 37700 ne
rect 29093 36569 37862 37700
rect 18862 35769 27962 36569
rect -35762 35438 -27793 35769
rect -41300 34424 -39038 35438
tri -39038 34424 -38024 35438 nw
tri -37907 34424 -36893 35438 se
rect -36893 34638 -27793 35438
tri -27793 34638 -26662 35769 nw
tri -26662 34638 -25531 35769 se
rect -25531 34638 17731 35769
tri 17731 34638 18862 35769 sw
tri 18862 34638 19993 35769 ne
rect 19993 35438 27962 35769
tri 27962 35438 29093 36569 sw
tri 29093 35438 30224 36569 ne
rect 30224 35438 37862 36569
rect 19993 34638 29093 35438
rect -36893 34424 -28924 34638
rect -41300 34262 -40169 34424
tri -51200 32162 -49100 34262 se
rect -49100 33293 -40169 34262
tri -40169 33293 -39038 34424 nw
tri -39038 33293 -37907 34424 se
rect -37907 33507 -28924 34424
tri -28924 33507 -27793 34638 nw
tri -27793 33507 -26662 34638 se
rect -26662 33507 18862 34638
tri 18862 33507 19993 34638 sw
tri 19993 33507 21124 34638 ne
rect 21124 34307 29093 34638
tri 29093 34307 30224 35438 sw
tri 30224 34307 31355 35438 ne
rect 31355 34307 37862 35438
rect 21124 33507 30224 34307
rect -37907 33293 -29138 33507
tri -29138 33293 -28924 33507 nw
tri -28007 33293 -27793 33507 se
rect -27793 33293 19993 33507
tri 19993 33293 20207 33507 sw
tri 21124 33293 21338 33507 ne
rect 21338 33293 30224 33507
tri 30224 33293 31238 34307 sw
tri 31355 33293 32369 34307 ne
rect 32369 33293 37862 34307
rect -49100 32162 -41300 33293
tri -41300 32162 -40169 33293 nw
tri -40169 32162 -39038 33293 se
rect -39038 32162 -30269 33293
tri -30269 32162 -29138 33293 nw
tri -29138 32162 -28007 33293 se
rect -28007 32162 20207 33293
tri 20207 32162 21338 33293 sw
tri 21338 32162 22469 33293 ne
rect 22469 32162 31238 33293
tri 31238 32162 32369 33293 sw
tri 32369 32162 33500 33293 ne
rect 33500 32162 37862 33293
tri -56900 26462 -51200 32162 se
rect -51200 31031 -42431 32162
tri -42431 31031 -41300 32162 nw
tri -41300 31031 -40169 32162 se
rect -40169 31031 -31400 32162
tri -31400 31031 -30269 32162 nw
tri -30269 31031 -29138 32162 se
rect -29138 31031 21338 32162
tri 21338 31031 22469 32162 sw
tri 22469 31031 23600 32162 ne
rect 23600 31031 32369 32162
tri 32369 31031 33500 32162 sw
tri 33500 31031 34631 32162 ne
rect 34631 31031 37862 32162
rect -51200 29900 -43562 31031
tri -43562 29900 -42431 31031 nw
tri -42431 29900 -41300 31031 se
rect -41300 29900 -32531 31031
tri -32531 29900 -31400 31031 nw
tri -31400 29900 -30269 31031 se
rect -30269 29900 22469 31031
tri 22469 29900 23600 31031 sw
tri 23600 29900 24731 31031 ne
rect 24731 29900 33500 31031
tri 33500 29900 34631 31031 sw
tri 34631 29900 35762 31031 ne
rect 35762 29900 37862 31031
tri 37862 29900 45662 37700 sw
rect -51200 28769 -44693 29900
tri -44693 28769 -43562 29900 nw
tri -43562 28769 -42431 29900 se
rect -42431 28769 -33662 29900
tri -33662 28769 -32531 29900 nw
tri -32531 28769 -31400 29900 se
rect -51200 27638 -45824 28769
tri -45824 27638 -44693 28769 nw
tri -44693 27638 -43562 28769 se
rect -43562 27638 -34793 28769
tri -34793 27638 -33662 28769 nw
tri -33662 27638 -32531 28769 se
rect -32531 27638 -31400 28769
rect -51200 26624 -46838 27638
tri -46838 26624 -45824 27638 nw
tri -45707 26624 -44693 27638 se
rect -44693 26624 -35924 27638
rect -51200 26462 -47969 26624
tri -59000 24362 -56900 26462 se
rect -56900 25493 -47969 26462
tri -47969 25493 -46838 26624 nw
tri -46838 25493 -45707 26624 se
rect -45707 26507 -35924 26624
tri -35924 26507 -34793 27638 nw
tri -34793 26507 -33662 27638 se
rect -33662 26507 -31400 27638
rect -45707 25493 -37055 26507
rect -56900 24362 -49100 25493
tri -49100 24362 -47969 25493 nw
tri -47969 24362 -46838 25493 se
rect -46838 25376 -37055 25493
tri -37055 25376 -35924 26507 nw
tri -35924 25376 -34793 26507 se
rect -34793 25376 -31400 26507
rect -46838 24524 -37907 25376
tri -37907 24524 -37055 25376 nw
tri -36776 24524 -35924 25376 se
rect -35924 24524 -31400 25376
rect -46838 24362 -39038 24524
tri -63900 19462 -59000 24362 se
rect -59000 23231 -50231 24362
tri -50231 23231 -49100 24362 nw
tri -49100 23231 -47969 24362 se
rect -47969 23393 -39038 24362
tri -39038 23393 -37907 24524 nw
tri -37907 23393 -36776 24524 se
rect -36776 23393 -31400 24524
rect -47969 23231 -40169 23393
rect -59000 22100 -51362 23231
tri -51362 22100 -50231 23231 nw
tri -50231 22100 -49100 23231 se
rect -49100 22262 -40169 23231
tri -40169 22262 -39038 23393 nw
tri -39038 22262 -37907 23393 se
rect -37907 22262 -31400 23393
rect -49100 22100 -41300 22262
rect -59000 21131 -52331 22100
tri -52331 21131 -51362 22100 nw
tri -51200 21131 -50231 22100 se
rect -50231 21131 -41300 22100
tri -41300 21131 -40169 22262 nw
tri -40169 21131 -39038 22262 se
rect -39038 21131 -31400 22262
rect -59000 20000 -53462 21131
tri -53462 20000 -52331 21131 nw
tri -52331 20000 -51200 21131 se
rect -51200 20000 -42431 21131
tri -42431 20000 -41300 21131 nw
tri -41300 20000 -40169 21131 se
rect -40169 20000 -31400 21131
tri -31400 20000 -21500 29900 nw
tri 13700 20000 23600 29900 ne
tri 23600 28769 24731 29900 sw
tri 24731 28769 25862 29900 ne
rect 25862 28769 34631 29900
tri 34631 28769 35762 29900 sw
tri 35762 28769 36893 29900 ne
rect 36893 28769 45662 29900
rect 23600 27638 24731 28769
tri 24731 27638 25862 28769 sw
tri 25862 27638 26993 28769 ne
rect 26993 27638 35762 28769
tri 35762 27638 36893 28769 sw
tri 36893 27638 38024 28769 ne
rect 38024 27638 45662 28769
rect 23600 26507 25862 27638
tri 25862 26507 26993 27638 sw
tri 26993 26507 28124 27638 ne
rect 28124 26507 36893 27638
tri 36893 26507 38024 27638 sw
tri 38024 26507 39155 27638 ne
rect 39155 26507 45662 27638
rect 23600 25376 26993 26507
tri 26993 25376 28124 26507 sw
tri 28124 25376 29255 26507 ne
rect 29255 25376 38024 26507
tri 38024 25376 39155 26507 sw
tri 39155 25376 40286 26507 ne
rect 40286 25376 45662 26507
rect 23600 24524 28124 25376
tri 28124 24524 28976 25376 sw
tri 29255 24524 30107 25376 ne
rect 30107 24524 39155 25376
tri 39155 24524 40007 25376 sw
tri 40286 24524 41138 25376 ne
rect 41138 24524 45662 25376
rect 23600 23393 28976 24524
tri 28976 23393 30107 24524 sw
tri 30107 23393 31238 24524 ne
rect 31238 23393 40007 24524
tri 40007 23393 41138 24524 sw
tri 41138 23393 42269 24524 ne
rect 42269 23393 45662 24524
rect 23600 22262 30107 23393
tri 30107 22262 31238 23393 sw
tri 31238 22262 32369 23393 ne
rect 32369 22262 41138 23393
tri 41138 22262 42269 23393 sw
tri 42269 22262 43400 23393 ne
rect 43400 22262 45662 23393
rect 23600 21131 31238 22262
tri 31238 21131 32369 22262 sw
tri 32369 21131 33500 22262 ne
rect 33500 21131 42269 22262
tri 42269 21131 43400 22262 sw
tri 43400 21131 44531 22262 ne
rect 44531 21131 45662 22262
rect 23600 20000 32369 21131
tri 32369 20000 33500 21131 sw
tri 33500 20000 34631 21131 ne
rect 34631 20000 43400 21131
tri 43400 20000 44531 21131 sw
tri 44531 20000 45662 21131 ne
tri 45662 20000 55562 29900 sw
rect -59000 19462 -54593 20000
rect -63900 18869 -54593 19462
tri -54593 18869 -53462 20000 nw
tri -53462 18869 -52331 20000 se
rect -52331 18869 -43562 20000
tri -43562 18869 -42431 20000 nw
tri -42431 18869 -41300 20000 se
rect -41300 18869 -37400 20000
rect -63900 18493 -54969 18869
tri -54969 18493 -54593 18869 nw
tri -53838 18493 -53462 18869 se
rect -53462 18493 -44693 18869
rect -63900 17362 -56100 18493
tri -56100 17362 -54969 18493 nw
tri -54969 17362 -53838 18493 se
rect -53838 17738 -44693 18493
tri -44693 17738 -43562 18869 nw
tri -43562 17738 -42431 18869 se
rect -42431 17738 -37400 18869
rect -53838 17362 -45824 17738
rect -63900 14000 -56900 17362
tri -56900 16562 -56100 17362 nw
tri -55769 16562 -54969 17362 se
rect -54969 16607 -45824 17362
tri -45824 16607 -44693 17738 nw
tri -44693 16607 -43562 17738 se
rect -43562 16607 -37400 17738
rect -54969 16562 -46038 16607
rect -70900 7000 -56900 14000
tri -56100 16231 -55769 16562 se
rect -55769 16393 -46038 16562
tri -46038 16393 -45824 16607 nw
tri -44907 16393 -44693 16607 se
rect -44693 16393 -37400 16607
rect -55769 16231 -47169 16393
rect -56100 15262 -47169 16231
tri -47169 15262 -46038 16393 nw
tri -46038 15262 -44907 16393 se
rect -44907 15262 -37400 16393
rect -56100 14131 -48300 15262
tri -48300 14131 -47169 15262 nw
tri -47169 14131 -46038 15262 se
rect -46038 14131 -37400 15262
rect -56100 14000 -48431 14131
tri -48431 14000 -48300 14131 nw
tri -47300 14000 -47169 14131 se
rect -47169 14000 -37400 14131
tri -37400 14000 -31400 20000 nw
tri 23600 14000 29600 20000 ne
rect 29600 18869 33500 20000
tri 33500 18869 34631 20000 sw
tri 34631 18869 35762 20000 ne
rect 35762 18869 44531 20000
tri 44531 18869 45662 20000 sw
tri 45662 18869 46793 20000 ne
rect 46793 19462 55562 20000
tri 55562 19462 56100 20000 sw
rect 46793 18869 56100 19462
rect 29600 17738 34631 18869
tri 34631 17738 35762 18869 sw
tri 35762 17738 36893 18869 ne
rect 36893 18493 45662 18869
tri 45662 18493 46038 18869 sw
tri 46793 18493 47169 18869 ne
rect 47169 18493 56100 18869
rect 36893 17738 46038 18493
rect 29600 16607 35762 17738
tri 35762 16607 36893 17738 sw
tri 36893 16607 38024 17738 ne
rect 38024 17362 46038 17738
tri 46038 17362 47169 18493 sw
tri 47169 17362 48300 18493 ne
rect 48300 17362 56100 18493
rect 38024 16607 47169 17362
rect 29600 16393 36893 16607
tri 36893 16393 37107 16607 sw
tri 38024 16393 38238 16607 ne
rect 38238 16562 47169 16607
tri 47169 16562 47969 17362 sw
tri 48300 16562 49100 17362 ne
rect 38238 16393 47969 16562
rect 29600 15262 37107 16393
tri 37107 15262 38238 16393 sw
tri 38238 15262 39369 16393 ne
rect 39369 16231 47969 16393
tri 47969 16231 48300 16562 sw
rect 39369 15262 48300 16231
rect 29600 14131 38238 15262
tri 38238 14131 39369 15262 sw
tri 39369 14131 40500 15262 ne
rect 40500 14131 48300 15262
rect 29600 14000 39369 14131
rect -64700 -7112 -57700 -7000
rect -64700 -13888 -64588 -7112
rect -57812 -13888 -57700 -7112
rect -64700 -14000 -57700 -13888
rect -56100 -19647 -49100 14000
tri -49100 13331 -48431 14000 nw
tri -47969 13331 -47300 14000 se
rect -47300 13331 -41300 14000
tri -48300 13000 -47969 13331 se
rect -47969 13000 -41300 13331
rect -48300 -16416 -41300 13000
tri -41300 10100 -37400 14000 nw
tri 29600 10100 33500 14000 ne
rect 33500 13331 39369 14000
tri 39369 13331 40169 14131 sw
tri 40500 13331 41300 14131 ne
rect 33500 13000 40169 13331
tri 40169 13000 40500 13331 sw
rect -40500 -7112 -33500 -7000
rect -40500 -13888 -40388 -7112
rect -33612 -13888 -33500 -7112
rect -40500 -15284 -33500 -13888
tri -40500 -15616 -40168 -15284 ne
rect -40168 -15616 -33500 -15284
tri -41300 -16416 -40500 -15616 sw
tri -40168 -16416 -39368 -15616 ne
rect -39368 -16416 -33500 -15616
rect -48300 -17548 -40500 -16416
tri -40500 -17548 -39368 -16416 sw
tri -39368 -17548 -38236 -16416 ne
rect -38236 -17548 -33500 -16416
rect -48300 -18515 -39368 -17548
tri -48300 -18847 -47968 -18515 ne
rect -47968 -18680 -39368 -18515
tri -39368 -18680 -38236 -17548 sw
tri -38236 -18680 -37104 -17548 ne
rect -37104 -18680 -33500 -17548
rect -47968 -18847 -38236 -18680
tri -49100 -19647 -48300 -18847 sw
tri -47968 -19647 -47168 -18847 ne
rect -47168 -18888 -38236 -18847
tri -38236 -18888 -38028 -18680 sw
tri -37104 -18888 -36896 -18680 ne
rect -36896 -18888 -33500 -18680
rect -47168 -19647 -38028 -18888
rect -56100 -20779 -48300 -19647
tri -48300 -20779 -47168 -19647 sw
tri -47168 -20779 -46036 -19647 ne
rect -46036 -20020 -38028 -19647
tri -38028 -20020 -36896 -18888 sw
tri -36896 -20020 -35764 -18888 ne
rect -35764 -20020 -33500 -18888
rect -46036 -20779 -36896 -20020
rect -56100 -21152 -47168 -20779
tri -47168 -21152 -46795 -20779 sw
tri -46036 -21152 -45663 -20779 ne
rect -45663 -21152 -36896 -20779
tri -36896 -21152 -35764 -20020 sw
tri -35764 -21152 -34632 -20020 ne
rect -34632 -21152 -33500 -20020
rect -56100 -21746 -46795 -21152
tri -56100 -22284 -55562 -21746 ne
rect -55562 -22284 -46795 -21746
tri -46795 -22284 -45663 -21152 sw
tri -45663 -22284 -44531 -21152 ne
rect -44531 -22284 -35764 -21152
tri -35764 -22284 -34632 -21152 sw
tri -34632 -22284 -33500 -21152 ne
tri -33500 -22284 -23601 -12385 sw
tri 25884 -20001 33500 -12385 se
rect 33500 -15284 40500 13000
rect 33500 -15616 40168 -15284
tri 40168 -15616 40500 -15284 nw
rect 33500 -16416 39368 -15616
tri 39368 -16416 40168 -15616 nw
tri 40500 -16416 41300 -15616 se
rect 41300 -16416 48300 14131
rect 33500 -17548 38236 -16416
tri 38236 -17548 39368 -16416 nw
tri 39368 -17548 40500 -16416 se
rect 40500 -17548 48300 -16416
rect 33500 -17737 38047 -17548
tri 38047 -17737 38236 -17548 nw
tri 39179 -17737 39368 -17548 se
rect 39368 -17737 48300 -17548
rect 33500 -18869 36915 -17737
tri 36915 -18869 38047 -17737 nw
tri 38047 -18869 39179 -17737 se
rect 39179 -18515 48300 -17737
rect 39179 -18847 47968 -18515
tri 47968 -18847 48300 -18515 nw
rect 39179 -18869 47168 -18847
rect 33500 -20001 35783 -18869
tri 35783 -20001 36915 -18869 nw
tri 36915 -20001 38047 -18869 se
rect 38047 -19647 47168 -18869
tri 47168 -19647 47968 -18847 nw
tri 48300 -19647 49100 -18847 se
rect 49100 -19647 56100 17362
rect 38047 -20001 46036 -19647
tri 23601 -22284 25884 -20001 se
rect 25884 -21133 34651 -20001
tri 34651 -21133 35783 -20001 nw
tri 35783 -21133 36915 -20001 se
rect 36915 -20779 46036 -20001
tri 46036 -20779 47168 -19647 nw
tri 47168 -20779 48300 -19647 se
rect 48300 -20779 56100 -19647
rect 36915 -21133 45663 -20779
rect 25884 -21152 34632 -21133
tri 34632 -21152 34651 -21133 nw
tri 35764 -21152 35783 -21133 se
rect 35783 -21152 45663 -21133
tri 45663 -21152 46036 -20779 nw
tri 46795 -21152 47168 -20779 se
rect 47168 -21152 56100 -20779
rect 25884 -22284 33500 -21152
tri 33500 -22284 34632 -21152 nw
tri 34632 -22284 35764 -21152 se
rect 35764 -22284 44531 -21152
tri 44531 -22284 45663 -21152 nw
tri 45663 -22284 46795 -21152 se
rect 46795 -21746 56100 -21152
rect 46795 -22284 51199 -21746
tri -55562 -29900 -47946 -22284 ne
rect -47946 -23416 -45663 -22284
tri -45663 -23416 -44531 -22284 sw
tri -44531 -23416 -43399 -22284 ne
rect -43399 -23416 -34632 -22284
tri -34632 -23416 -33500 -22284 sw
tri -33500 -23416 -32368 -22284 ne
rect -32368 -23416 -23601 -22284
rect -47946 -24548 -44531 -23416
tri -44531 -24548 -43399 -23416 sw
tri -43399 -24548 -42267 -23416 ne
rect -42267 -24548 -33500 -23416
tri -33500 -24548 -32368 -23416 sw
tri -32368 -24548 -31236 -23416 ne
rect -31236 -24548 -23601 -23416
rect -47946 -25680 -43399 -24548
tri -43399 -25680 -42267 -24548 sw
tri -42267 -25680 -41135 -24548 ne
rect -41135 -25680 -32368 -24548
tri -32368 -25680 -31236 -24548 sw
tri -31236 -25680 -30104 -24548 ne
rect -30104 -25680 -23601 -24548
rect -47946 -26504 -42267 -25680
tri -42267 -26504 -41443 -25680 sw
tri -41135 -26504 -40311 -25680 ne
rect -40311 -26504 -31236 -25680
tri -31236 -26504 -30412 -25680 sw
tri -30104 -26504 -29280 -25680 ne
rect -29280 -26504 -23601 -25680
rect -47946 -27636 -41443 -26504
tri -41443 -27636 -40311 -26504 sw
tri -40311 -27636 -39179 -26504 ne
rect -39179 -27636 -30412 -26504
tri -30412 -27636 -29280 -26504 sw
tri -29280 -27636 -28148 -26504 ne
rect -28148 -27636 -23601 -26504
rect -47946 -28768 -40311 -27636
tri -40311 -28768 -39179 -27636 sw
tri -39179 -28768 -38047 -27636 ne
rect -38047 -28768 -29280 -27636
tri -29280 -28768 -28148 -27636 sw
tri -28148 -28768 -27016 -27636 ne
rect -27016 -28768 -23601 -27636
rect -47946 -29900 -39179 -28768
tri -39179 -29900 -38047 -28768 sw
tri -38047 -29900 -36915 -28768 ne
rect -36915 -29900 -28148 -28768
tri -28148 -29900 -27016 -28768 sw
tri -27016 -29900 -25884 -28768 ne
rect -25884 -29900 -23601 -28768
tri -23601 -29900 -15985 -22284 sw
tri 15985 -29900 23601 -22284 se
rect 23601 -23416 32368 -22284
tri 32368 -23416 33500 -22284 nw
tri 33500 -23416 34632 -22284 se
rect 34632 -23416 43399 -22284
tri 43399 -23416 44531 -22284 nw
tri 44531 -23416 45663 -22284 se
rect 45663 -23416 51199 -22284
rect 23601 -24548 31236 -23416
tri 31236 -24548 32368 -23416 nw
tri 32368 -24548 33500 -23416 se
rect 33500 -24383 42432 -23416
tri 42432 -24383 43399 -23416 nw
tri 43564 -24383 44531 -23416 se
rect 44531 -24383 51199 -23416
rect 33500 -24548 41300 -24383
rect 23601 -25680 30104 -24548
tri 30104 -25680 31236 -24548 nw
tri 31236 -25680 32368 -24548 se
rect 32368 -25515 41300 -24548
tri 41300 -25515 42432 -24383 nw
tri 42432 -25515 43564 -24383 se
rect 43564 -25515 51199 -24383
rect 32368 -25680 40168 -25515
rect 23601 -26504 29280 -25680
tri 29280 -26504 30104 -25680 nw
tri 30412 -26504 31236 -25680 se
rect 31236 -26504 40168 -25680
rect 23601 -27636 28148 -26504
tri 28148 -27636 29280 -26504 nw
tri 29280 -27636 30412 -26504 se
rect 30412 -26647 40168 -26504
tri 40168 -26647 41300 -25515 nw
tri 41300 -26647 42432 -25515 se
rect 42432 -26647 51199 -25515
tri 51199 -26647 56100 -21746 nw
rect 30412 -27636 39036 -26647
rect 23601 -28768 27016 -27636
tri 27016 -28768 28148 -27636 nw
tri 28148 -28768 29280 -27636 se
rect 29280 -27779 39036 -27636
tri 39036 -27779 40168 -26647 nw
tri 40168 -27779 41300 -26647 se
rect 41300 -27779 49100 -26647
rect 29280 -28768 38047 -27779
tri 38047 -28768 39036 -27779 nw
tri 39179 -28768 40168 -27779 se
rect 40168 -28746 49100 -27779
tri 49100 -28746 51199 -26647 nw
rect 40168 -28768 43399 -28746
rect 23601 -29900 25884 -28768
tri 25884 -29900 27016 -28768 nw
tri 27016 -29900 28148 -28768 se
rect 28148 -29900 36915 -28768
tri 36915 -29900 38047 -28768 nw
tri 38047 -29900 39179 -28768 se
rect 39179 -29900 43399 -28768
tri -47946 -37700 -40146 -29900 ne
rect -40146 -31032 -38047 -29900
tri -38047 -31032 -36915 -29900 sw
tri -36915 -31032 -35783 -29900 ne
rect -35783 -31032 -27016 -29900
tri -27016 -31032 -25884 -29900 sw
tri -25884 -31032 -24752 -29900 ne
rect -24752 -31032 24752 -29900
tri 24752 -31032 25884 -29900 nw
tri 25884 -31032 27016 -29900 se
rect 27016 -31032 35783 -29900
tri 35783 -31032 36915 -29900 nw
tri 36915 -31032 38047 -29900 se
rect 38047 -31032 43399 -29900
rect -40146 -32164 -36915 -31032
tri -36915 -32164 -35783 -31032 sw
tri -35783 -32164 -34651 -31032 ne
rect -34651 -32164 -25884 -31032
tri -25884 -32164 -24752 -31032 sw
tri -24752 -32164 -23620 -31032 ne
rect -23620 -32164 23620 -31032
tri 23620 -32164 24752 -31032 nw
tri 24752 -32164 25884 -31032 se
rect 25884 -32164 34651 -31032
tri 34651 -32164 35783 -31032 nw
tri 35783 -32164 36915 -31032 se
rect 36915 -32164 43399 -31032
rect -40146 -33296 -35783 -32164
tri -35783 -33296 -34651 -32164 sw
tri -34651 -33296 -33519 -32164 ne
rect -33519 -33296 -24752 -32164
tri -24752 -33296 -23620 -32164 sw
tri -23620 -33296 -22488 -32164 ne
rect -22488 -33296 22488 -32164
tri 22488 -33296 23620 -32164 nw
tri 23620 -33296 24752 -32164 se
rect 24752 -32183 34632 -32164
tri 34632 -32183 34651 -32164 nw
tri 35764 -32183 35783 -32164 se
rect 35783 -32183 43399 -32164
rect 24752 -33296 33500 -32183
rect -40146 -34304 -34651 -33296
tri -34651 -34304 -33643 -33296 sw
tri -33519 -34304 -32511 -33296 ne
rect -32511 -33504 -23620 -33296
tri -23620 -33504 -23412 -33296 sw
tri -22488 -33504 -22280 -33296 ne
rect -22280 -33504 22280 -33296
tri 22280 -33504 22488 -33296 nw
tri 23412 -33504 23620 -33296 se
rect 23620 -33315 33500 -33296
tri 33500 -33315 34632 -32183 nw
tri 34632 -33315 35764 -32183 se
rect 35764 -33315 43399 -32183
rect 23620 -33504 32368 -33315
rect -32511 -34304 -23412 -33504
rect -40146 -35436 -33643 -34304
tri -33643 -35436 -32511 -34304 sw
tri -32511 -35436 -31379 -34304 ne
rect -31379 -34636 -23412 -34304
tri -23412 -34636 -22280 -33504 sw
tri -22280 -34636 -21148 -33504 ne
rect -21148 -34636 21148 -33504
tri 21148 -34636 22280 -33504 nw
tri 22280 -34636 23412 -33504 se
rect 23412 -34447 32368 -33504
tri 32368 -34447 33500 -33315 nw
tri 33500 -34447 34632 -33315 se
rect 34632 -34447 43399 -33315
tri 43399 -34447 49100 -28746 nw
rect 23412 -34636 31236 -34447
rect -31379 -35436 -22280 -34636
rect -40146 -36568 -32511 -35436
tri -32511 -36568 -31379 -35436 sw
tri -31379 -36568 -30247 -35436 ne
rect -30247 -35768 -22280 -35436
tri -22280 -35768 -21148 -34636 sw
tri -21148 -35768 -20016 -34636 ne
rect -20016 -35768 20016 -34636
tri 20016 -35768 21148 -34636 nw
tri 21148 -35768 22280 -34636 se
rect 22280 -35579 31236 -34636
tri 31236 -35579 32368 -34447 nw
tri 32368 -35579 33500 -34447 se
rect 33500 -35579 41300 -34447
rect 22280 -35768 30247 -35579
rect -30247 -36568 -21148 -35768
rect -40146 -37700 -31379 -36568
tri -31379 -37700 -30247 -36568 sw
tri -30247 -37700 -29115 -36568 ne
rect -29115 -36900 -21148 -36568
tri -21148 -36900 -20016 -35768 sw
tri -20016 -36900 -18884 -35768 ne
rect -18884 -36900 18884 -35768
tri 18884 -36900 20016 -35768 nw
tri 20016 -36900 21148 -35768 se
rect 21148 -36568 30247 -35768
tri 30247 -36568 31236 -35579 nw
tri 31379 -36568 32368 -35579 se
rect 32368 -36546 41300 -35579
tri 41300 -36546 43399 -34447 nw
rect 32368 -36568 35783 -36546
rect 21148 -36900 29115 -36568
rect -29115 -37700 -20016 -36900
tri -20016 -37700 -19216 -36900 sw
tri 19216 -37700 20016 -36900 se
rect 20016 -37700 29115 -36900
tri 29115 -37700 30247 -36568 nw
tri 30247 -37700 31379 -36568 se
rect 31379 -37700 35783 -36568
tri -40146 -45500 -32346 -37700 ne
rect -32346 -38832 -30247 -37700
tri -30247 -38832 -29115 -37700 sw
tri -29115 -38832 -27983 -37700 ne
rect -27983 -38832 27983 -37700
tri 27983 -38832 29115 -37700 nw
tri 29115 -38832 30247 -37700 se
rect 30247 -38832 35783 -37700
rect -32346 -39964 -29115 -38832
tri -29115 -39964 -27983 -38832 sw
tri -27983 -39964 -26851 -38832 ne
rect -26851 -39799 27016 -38832
tri 27016 -39799 27983 -38832 nw
tri 28148 -39799 29115 -38832 se
rect 29115 -39799 35783 -38832
rect -26851 -39964 25884 -39799
rect -32346 -41096 -27983 -39964
tri -27983 -41096 -26851 -39964 sw
tri -26851 -41096 -25719 -39964 ne
rect -25719 -40931 25884 -39964
tri 25884 -40931 27016 -39799 nw
tri 27016 -40931 28148 -39799 se
rect 28148 -40931 35783 -39799
rect -25719 -41096 24752 -40931
rect -32346 -41304 -26851 -41096
tri -26851 -41304 -26643 -41096 sw
tri -25719 -41304 -25511 -41096 ne
rect -25511 -41304 24752 -41096
rect -32346 -42436 -26643 -41304
tri -26643 -42436 -25511 -41304 sw
tri -25511 -42436 -24379 -41304 ne
rect -24379 -42063 24752 -41304
tri 24752 -42063 25884 -40931 nw
tri 25884 -42063 27016 -40931 se
rect 27016 -42063 35783 -40931
tri 35783 -42063 41300 -36546 nw
rect -24379 -42436 23620 -42063
rect -32346 -43568 -25511 -42436
tri -25511 -43568 -24379 -42436 sw
tri -24379 -43568 -23247 -42436 ne
rect -23247 -43195 23620 -42436
tri 23620 -43195 24752 -42063 nw
tri 24752 -43195 25884 -42063 se
rect 25884 -43195 33500 -42063
rect -23247 -43568 23247 -43195
tri 23247 -43568 23620 -43195 nw
tri 24379 -43568 24752 -43195 se
rect 24752 -43568 33500 -43195
rect -32346 -44700 -24379 -43568
tri -24379 -44700 -23247 -43568 sw
tri -23247 -44700 -22115 -43568 ne
rect -22115 -44700 22115 -43568
tri 22115 -44700 23247 -43568 nw
tri 23247 -44700 24379 -43568 se
rect 24379 -44346 33500 -43568
tri 33500 -44346 35783 -42063 nw
rect 24379 -44700 32346 -44346
rect -32346 -45500 -23247 -44700
tri -23247 -45500 -22447 -44700 sw
tri 22447 -45500 23247 -44700 se
rect 23247 -45500 32346 -44700
tri 32346 -45500 33500 -44346 nw
tri -32346 -51962 -25884 -45500 ne
rect -25884 -51962 25884 -45500
tri 25884 -51962 32346 -45500 nw
tri -25884 -52500 -25346 -51962 ne
rect -25346 -52500 25346 -51962
tri 25346 -52500 25884 -51962 nw
<< end >>
