magic
tech sky130B
timestamp 1663433502
<< pwell >>
rect -1087 -3129 1087 3129
<< mvnmos >>
rect -973 -3000 -923 3000
rect -894 -3000 -844 3000
rect -815 -3000 -765 3000
rect -736 -3000 -686 3000
rect -657 -3000 -607 3000
rect -578 -3000 -528 3000
rect -499 -3000 -449 3000
rect -420 -3000 -370 3000
rect -341 -3000 -291 3000
rect -262 -3000 -212 3000
rect -183 -3000 -133 3000
rect -104 -3000 -54 3000
rect -25 -3000 25 3000
rect 54 -3000 104 3000
rect 133 -3000 183 3000
rect 212 -3000 262 3000
rect 291 -3000 341 3000
rect 370 -3000 420 3000
rect 449 -3000 499 3000
rect 528 -3000 578 3000
rect 607 -3000 657 3000
rect 686 -3000 736 3000
rect 765 -3000 815 3000
rect 844 -3000 894 3000
rect 923 -3000 973 3000
<< mvndiff >>
rect -1002 2994 -973 3000
rect -1002 -2994 -996 2994
rect -979 -2994 -973 2994
rect -1002 -3000 -973 -2994
rect -923 2994 -894 3000
rect -923 -2994 -917 2994
rect -900 -2994 -894 2994
rect -923 -3000 -894 -2994
rect -844 2994 -815 3000
rect -844 -2994 -838 2994
rect -821 -2994 -815 2994
rect -844 -3000 -815 -2994
rect -765 2994 -736 3000
rect -765 -2994 -759 2994
rect -742 -2994 -736 2994
rect -765 -3000 -736 -2994
rect -686 2994 -657 3000
rect -686 -2994 -680 2994
rect -663 -2994 -657 2994
rect -686 -3000 -657 -2994
rect -607 2994 -578 3000
rect -607 -2994 -601 2994
rect -584 -2994 -578 2994
rect -607 -3000 -578 -2994
rect -528 2994 -499 3000
rect -528 -2994 -522 2994
rect -505 -2994 -499 2994
rect -528 -3000 -499 -2994
rect -449 2994 -420 3000
rect -449 -2994 -443 2994
rect -426 -2994 -420 2994
rect -449 -3000 -420 -2994
rect -370 2994 -341 3000
rect -370 -2994 -364 2994
rect -347 -2994 -341 2994
rect -370 -3000 -341 -2994
rect -291 2994 -262 3000
rect -291 -2994 -285 2994
rect -268 -2994 -262 2994
rect -291 -3000 -262 -2994
rect -212 2994 -183 3000
rect -212 -2994 -206 2994
rect -189 -2994 -183 2994
rect -212 -3000 -183 -2994
rect -133 2994 -104 3000
rect -133 -2994 -127 2994
rect -110 -2994 -104 2994
rect -133 -3000 -104 -2994
rect -54 2994 -25 3000
rect -54 -2994 -48 2994
rect -31 -2994 -25 2994
rect -54 -3000 -25 -2994
rect 25 2994 54 3000
rect 25 -2994 31 2994
rect 48 -2994 54 2994
rect 25 -3000 54 -2994
rect 104 2994 133 3000
rect 104 -2994 110 2994
rect 127 -2994 133 2994
rect 104 -3000 133 -2994
rect 183 2994 212 3000
rect 183 -2994 189 2994
rect 206 -2994 212 2994
rect 183 -3000 212 -2994
rect 262 2994 291 3000
rect 262 -2994 268 2994
rect 285 -2994 291 2994
rect 262 -3000 291 -2994
rect 341 2994 370 3000
rect 341 -2994 347 2994
rect 364 -2994 370 2994
rect 341 -3000 370 -2994
rect 420 2994 449 3000
rect 420 -2994 426 2994
rect 443 -2994 449 2994
rect 420 -3000 449 -2994
rect 499 2994 528 3000
rect 499 -2994 505 2994
rect 522 -2994 528 2994
rect 499 -3000 528 -2994
rect 578 2994 607 3000
rect 578 -2994 584 2994
rect 601 -2994 607 2994
rect 578 -3000 607 -2994
rect 657 2994 686 3000
rect 657 -2994 663 2994
rect 680 -2994 686 2994
rect 657 -3000 686 -2994
rect 736 2994 765 3000
rect 736 -2994 742 2994
rect 759 -2994 765 2994
rect 736 -3000 765 -2994
rect 815 2994 844 3000
rect 815 -2994 821 2994
rect 838 -2994 844 2994
rect 815 -3000 844 -2994
rect 894 2994 923 3000
rect 894 -2994 900 2994
rect 917 -2994 923 2994
rect 894 -3000 923 -2994
rect 973 2994 1002 3000
rect 973 -2994 979 2994
rect 996 -2994 1002 2994
rect 973 -3000 1002 -2994
<< mvndiffc >>
rect -996 -2994 -979 2994
rect -917 -2994 -900 2994
rect -838 -2994 -821 2994
rect -759 -2994 -742 2994
rect -680 -2994 -663 2994
rect -601 -2994 -584 2994
rect -522 -2994 -505 2994
rect -443 -2994 -426 2994
rect -364 -2994 -347 2994
rect -285 -2994 -268 2994
rect -206 -2994 -189 2994
rect -127 -2994 -110 2994
rect -48 -2994 -31 2994
rect 31 -2994 48 2994
rect 110 -2994 127 2994
rect 189 -2994 206 2994
rect 268 -2994 285 2994
rect 347 -2994 364 2994
rect 426 -2994 443 2994
rect 505 -2994 522 2994
rect 584 -2994 601 2994
rect 663 -2994 680 2994
rect 742 -2994 759 2994
rect 821 -2994 838 2994
rect 900 -2994 917 2994
rect 979 -2994 996 2994
<< mvpsubdiff >>
rect -1069 3105 1069 3111
rect -1069 3088 -1015 3105
rect 1015 3088 1069 3105
rect -1069 3082 1069 3088
rect -1069 3057 -1040 3082
rect -1069 -3057 -1063 3057
rect -1046 -3057 -1040 3057
rect 1040 3057 1069 3082
rect -1069 -3082 -1040 -3057
rect 1040 -3057 1046 3057
rect 1063 -3057 1069 3057
rect 1040 -3082 1069 -3057
rect -1069 -3088 1069 -3082
rect -1069 -3105 -1015 -3088
rect 1015 -3105 1069 -3088
rect -1069 -3111 1069 -3105
<< mvpsubdiffcont >>
rect -1015 3088 1015 3105
rect -1063 -3057 -1046 3057
rect 1046 -3057 1063 3057
rect -1015 -3105 1015 -3088
<< poly >>
rect -973 3036 -923 3044
rect -973 3019 -965 3036
rect -931 3019 -923 3036
rect -973 3000 -923 3019
rect -894 3036 -844 3044
rect -894 3019 -886 3036
rect -852 3019 -844 3036
rect -894 3000 -844 3019
rect -815 3036 -765 3044
rect -815 3019 -807 3036
rect -773 3019 -765 3036
rect -815 3000 -765 3019
rect -736 3036 -686 3044
rect -736 3019 -728 3036
rect -694 3019 -686 3036
rect -736 3000 -686 3019
rect -657 3036 -607 3044
rect -657 3019 -649 3036
rect -615 3019 -607 3036
rect -657 3000 -607 3019
rect -578 3036 -528 3044
rect -578 3019 -570 3036
rect -536 3019 -528 3036
rect -578 3000 -528 3019
rect -499 3036 -449 3044
rect -499 3019 -491 3036
rect -457 3019 -449 3036
rect -499 3000 -449 3019
rect -420 3036 -370 3044
rect -420 3019 -412 3036
rect -378 3019 -370 3036
rect -420 3000 -370 3019
rect -341 3036 -291 3044
rect -341 3019 -333 3036
rect -299 3019 -291 3036
rect -341 3000 -291 3019
rect -262 3036 -212 3044
rect -262 3019 -254 3036
rect -220 3019 -212 3036
rect -262 3000 -212 3019
rect -183 3036 -133 3044
rect -183 3019 -175 3036
rect -141 3019 -133 3036
rect -183 3000 -133 3019
rect -104 3036 -54 3044
rect -104 3019 -96 3036
rect -62 3019 -54 3036
rect -104 3000 -54 3019
rect -25 3036 25 3044
rect -25 3019 -17 3036
rect 17 3019 25 3036
rect -25 3000 25 3019
rect 54 3036 104 3044
rect 54 3019 62 3036
rect 96 3019 104 3036
rect 54 3000 104 3019
rect 133 3036 183 3044
rect 133 3019 141 3036
rect 175 3019 183 3036
rect 133 3000 183 3019
rect 212 3036 262 3044
rect 212 3019 220 3036
rect 254 3019 262 3036
rect 212 3000 262 3019
rect 291 3036 341 3044
rect 291 3019 299 3036
rect 333 3019 341 3036
rect 291 3000 341 3019
rect 370 3036 420 3044
rect 370 3019 378 3036
rect 412 3019 420 3036
rect 370 3000 420 3019
rect 449 3036 499 3044
rect 449 3019 457 3036
rect 491 3019 499 3036
rect 449 3000 499 3019
rect 528 3036 578 3044
rect 528 3019 536 3036
rect 570 3019 578 3036
rect 528 3000 578 3019
rect 607 3036 657 3044
rect 607 3019 615 3036
rect 649 3019 657 3036
rect 607 3000 657 3019
rect 686 3036 736 3044
rect 686 3019 694 3036
rect 728 3019 736 3036
rect 686 3000 736 3019
rect 765 3036 815 3044
rect 765 3019 773 3036
rect 807 3019 815 3036
rect 765 3000 815 3019
rect 844 3036 894 3044
rect 844 3019 852 3036
rect 886 3019 894 3036
rect 844 3000 894 3019
rect 923 3036 973 3044
rect 923 3019 931 3036
rect 965 3019 973 3036
rect 923 3000 973 3019
rect -973 -3019 -923 -3000
rect -973 -3036 -965 -3019
rect -931 -3036 -923 -3019
rect -973 -3044 -923 -3036
rect -894 -3019 -844 -3000
rect -894 -3036 -886 -3019
rect -852 -3036 -844 -3019
rect -894 -3044 -844 -3036
rect -815 -3019 -765 -3000
rect -815 -3036 -807 -3019
rect -773 -3036 -765 -3019
rect -815 -3044 -765 -3036
rect -736 -3019 -686 -3000
rect -736 -3036 -728 -3019
rect -694 -3036 -686 -3019
rect -736 -3044 -686 -3036
rect -657 -3019 -607 -3000
rect -657 -3036 -649 -3019
rect -615 -3036 -607 -3019
rect -657 -3044 -607 -3036
rect -578 -3019 -528 -3000
rect -578 -3036 -570 -3019
rect -536 -3036 -528 -3019
rect -578 -3044 -528 -3036
rect -499 -3019 -449 -3000
rect -499 -3036 -491 -3019
rect -457 -3036 -449 -3019
rect -499 -3044 -449 -3036
rect -420 -3019 -370 -3000
rect -420 -3036 -412 -3019
rect -378 -3036 -370 -3019
rect -420 -3044 -370 -3036
rect -341 -3019 -291 -3000
rect -341 -3036 -333 -3019
rect -299 -3036 -291 -3019
rect -341 -3044 -291 -3036
rect -262 -3019 -212 -3000
rect -262 -3036 -254 -3019
rect -220 -3036 -212 -3019
rect -262 -3044 -212 -3036
rect -183 -3019 -133 -3000
rect -183 -3036 -175 -3019
rect -141 -3036 -133 -3019
rect -183 -3044 -133 -3036
rect -104 -3019 -54 -3000
rect -104 -3036 -96 -3019
rect -62 -3036 -54 -3019
rect -104 -3044 -54 -3036
rect -25 -3019 25 -3000
rect -25 -3036 -17 -3019
rect 17 -3036 25 -3019
rect -25 -3044 25 -3036
rect 54 -3019 104 -3000
rect 54 -3036 62 -3019
rect 96 -3036 104 -3019
rect 54 -3044 104 -3036
rect 133 -3019 183 -3000
rect 133 -3036 141 -3019
rect 175 -3036 183 -3019
rect 133 -3044 183 -3036
rect 212 -3019 262 -3000
rect 212 -3036 220 -3019
rect 254 -3036 262 -3019
rect 212 -3044 262 -3036
rect 291 -3019 341 -3000
rect 291 -3036 299 -3019
rect 333 -3036 341 -3019
rect 291 -3044 341 -3036
rect 370 -3019 420 -3000
rect 370 -3036 378 -3019
rect 412 -3036 420 -3019
rect 370 -3044 420 -3036
rect 449 -3019 499 -3000
rect 449 -3036 457 -3019
rect 491 -3036 499 -3019
rect 449 -3044 499 -3036
rect 528 -3019 578 -3000
rect 528 -3036 536 -3019
rect 570 -3036 578 -3019
rect 528 -3044 578 -3036
rect 607 -3019 657 -3000
rect 607 -3036 615 -3019
rect 649 -3036 657 -3019
rect 607 -3044 657 -3036
rect 686 -3019 736 -3000
rect 686 -3036 694 -3019
rect 728 -3036 736 -3019
rect 686 -3044 736 -3036
rect 765 -3019 815 -3000
rect 765 -3036 773 -3019
rect 807 -3036 815 -3019
rect 765 -3044 815 -3036
rect 844 -3019 894 -3000
rect 844 -3036 852 -3019
rect 886 -3036 894 -3019
rect 844 -3044 894 -3036
rect 923 -3019 973 -3000
rect 923 -3036 931 -3019
rect 965 -3036 973 -3019
rect 923 -3044 973 -3036
<< polycont >>
rect -965 3019 -931 3036
rect -886 3019 -852 3036
rect -807 3019 -773 3036
rect -728 3019 -694 3036
rect -649 3019 -615 3036
rect -570 3019 -536 3036
rect -491 3019 -457 3036
rect -412 3019 -378 3036
rect -333 3019 -299 3036
rect -254 3019 -220 3036
rect -175 3019 -141 3036
rect -96 3019 -62 3036
rect -17 3019 17 3036
rect 62 3019 96 3036
rect 141 3019 175 3036
rect 220 3019 254 3036
rect 299 3019 333 3036
rect 378 3019 412 3036
rect 457 3019 491 3036
rect 536 3019 570 3036
rect 615 3019 649 3036
rect 694 3019 728 3036
rect 773 3019 807 3036
rect 852 3019 886 3036
rect 931 3019 965 3036
rect -965 -3036 -931 -3019
rect -886 -3036 -852 -3019
rect -807 -3036 -773 -3019
rect -728 -3036 -694 -3019
rect -649 -3036 -615 -3019
rect -570 -3036 -536 -3019
rect -491 -3036 -457 -3019
rect -412 -3036 -378 -3019
rect -333 -3036 -299 -3019
rect -254 -3036 -220 -3019
rect -175 -3036 -141 -3019
rect -96 -3036 -62 -3019
rect -17 -3036 17 -3019
rect 62 -3036 96 -3019
rect 141 -3036 175 -3019
rect 220 -3036 254 -3019
rect 299 -3036 333 -3019
rect 378 -3036 412 -3019
rect 457 -3036 491 -3019
rect 536 -3036 570 -3019
rect 615 -3036 649 -3019
rect 694 -3036 728 -3019
rect 773 -3036 807 -3019
rect 852 -3036 886 -3019
rect 931 -3036 965 -3019
<< locali >>
rect -1063 3088 -1015 3105
rect 1015 3088 1063 3105
rect -1063 3057 -1046 3088
rect 1046 3057 1063 3088
rect -973 3019 -965 3036
rect -931 3019 -923 3036
rect -894 3019 -886 3036
rect -852 3019 -844 3036
rect -815 3019 -807 3036
rect -773 3019 -765 3036
rect -736 3019 -728 3036
rect -694 3019 -686 3036
rect -657 3019 -649 3036
rect -615 3019 -607 3036
rect -578 3019 -570 3036
rect -536 3019 -528 3036
rect -499 3019 -491 3036
rect -457 3019 -449 3036
rect -420 3019 -412 3036
rect -378 3019 -370 3036
rect -341 3019 -333 3036
rect -299 3019 -291 3036
rect -262 3019 -254 3036
rect -220 3019 -212 3036
rect -183 3019 -175 3036
rect -141 3019 -133 3036
rect -104 3019 -96 3036
rect -62 3019 -54 3036
rect -25 3019 -17 3036
rect 17 3019 25 3036
rect 54 3019 62 3036
rect 96 3019 104 3036
rect 133 3019 141 3036
rect 175 3019 183 3036
rect 212 3019 220 3036
rect 254 3019 262 3036
rect 291 3019 299 3036
rect 333 3019 341 3036
rect 370 3019 378 3036
rect 412 3019 420 3036
rect 449 3019 457 3036
rect 491 3019 499 3036
rect 528 3019 536 3036
rect 570 3019 578 3036
rect 607 3019 615 3036
rect 649 3019 657 3036
rect 686 3019 694 3036
rect 728 3019 736 3036
rect 765 3019 773 3036
rect 807 3019 815 3036
rect 844 3019 852 3036
rect 886 3019 894 3036
rect 923 3019 931 3036
rect 965 3019 973 3036
rect -996 2994 -979 3002
rect -996 -3002 -979 -2994
rect -917 2994 -900 3002
rect -917 -3002 -900 -2994
rect -838 2994 -821 3002
rect -838 -3002 -821 -2994
rect -759 2994 -742 3002
rect -759 -3002 -742 -2994
rect -680 2994 -663 3002
rect -680 -3002 -663 -2994
rect -601 2994 -584 3002
rect -601 -3002 -584 -2994
rect -522 2994 -505 3002
rect -522 -3002 -505 -2994
rect -443 2994 -426 3002
rect -443 -3002 -426 -2994
rect -364 2994 -347 3002
rect -364 -3002 -347 -2994
rect -285 2994 -268 3002
rect -285 -3002 -268 -2994
rect -206 2994 -189 3002
rect -206 -3002 -189 -2994
rect -127 2994 -110 3002
rect -127 -3002 -110 -2994
rect -48 2994 -31 3002
rect -48 -3002 -31 -2994
rect 31 2994 48 3002
rect 31 -3002 48 -2994
rect 110 2994 127 3002
rect 110 -3002 127 -2994
rect 189 2994 206 3002
rect 189 -3002 206 -2994
rect 268 2994 285 3002
rect 268 -3002 285 -2994
rect 347 2994 364 3002
rect 347 -3002 364 -2994
rect 426 2994 443 3002
rect 426 -3002 443 -2994
rect 505 2994 522 3002
rect 505 -3002 522 -2994
rect 584 2994 601 3002
rect 584 -3002 601 -2994
rect 663 2994 680 3002
rect 663 -3002 680 -2994
rect 742 2994 759 3002
rect 742 -3002 759 -2994
rect 821 2994 838 3002
rect 821 -3002 838 -2994
rect 900 2994 917 3002
rect 900 -3002 917 -2994
rect 979 2994 996 3002
rect 979 -3002 996 -2994
rect -973 -3036 -965 -3019
rect -931 -3036 -923 -3019
rect -894 -3036 -886 -3019
rect -852 -3036 -844 -3019
rect -815 -3036 -807 -3019
rect -773 -3036 -765 -3019
rect -736 -3036 -728 -3019
rect -694 -3036 -686 -3019
rect -657 -3036 -649 -3019
rect -615 -3036 -607 -3019
rect -578 -3036 -570 -3019
rect -536 -3036 -528 -3019
rect -499 -3036 -491 -3019
rect -457 -3036 -449 -3019
rect -420 -3036 -412 -3019
rect -378 -3036 -370 -3019
rect -341 -3036 -333 -3019
rect -299 -3036 -291 -3019
rect -262 -3036 -254 -3019
rect -220 -3036 -212 -3019
rect -183 -3036 -175 -3019
rect -141 -3036 -133 -3019
rect -104 -3036 -96 -3019
rect -62 -3036 -54 -3019
rect -25 -3036 -17 -3019
rect 17 -3036 25 -3019
rect 54 -3036 62 -3019
rect 96 -3036 104 -3019
rect 133 -3036 141 -3019
rect 175 -3036 183 -3019
rect 212 -3036 220 -3019
rect 254 -3036 262 -3019
rect 291 -3036 299 -3019
rect 333 -3036 341 -3019
rect 370 -3036 378 -3019
rect 412 -3036 420 -3019
rect 449 -3036 457 -3019
rect 491 -3036 499 -3019
rect 528 -3036 536 -3019
rect 570 -3036 578 -3019
rect 607 -3036 615 -3019
rect 649 -3036 657 -3019
rect 686 -3036 694 -3019
rect 728 -3036 736 -3019
rect 765 -3036 773 -3019
rect 807 -3036 815 -3019
rect 844 -3036 852 -3019
rect 886 -3036 894 -3019
rect 923 -3036 931 -3019
rect 965 -3036 973 -3019
rect -1063 -3088 -1046 -3057
rect 1046 -3088 1063 -3057
rect -1063 -3105 -1015 -3088
rect 1015 -3105 1063 -3088
<< viali >>
rect -965 3019 -931 3036
rect -886 3019 -852 3036
rect -807 3019 -773 3036
rect -728 3019 -694 3036
rect -649 3019 -615 3036
rect -570 3019 -536 3036
rect -491 3019 -457 3036
rect -412 3019 -378 3036
rect -333 3019 -299 3036
rect -254 3019 -220 3036
rect -175 3019 -141 3036
rect -96 3019 -62 3036
rect -17 3019 17 3036
rect 62 3019 96 3036
rect 141 3019 175 3036
rect 220 3019 254 3036
rect 299 3019 333 3036
rect 378 3019 412 3036
rect 457 3019 491 3036
rect 536 3019 570 3036
rect 615 3019 649 3036
rect 694 3019 728 3036
rect 773 3019 807 3036
rect 852 3019 886 3036
rect 931 3019 965 3036
rect -996 -2994 -979 2994
rect -917 -2994 -900 2994
rect -838 -2994 -821 2994
rect -759 -2994 -742 2994
rect -680 -2994 -663 2994
rect -601 -2994 -584 2994
rect -522 -2994 -505 2994
rect -443 -2994 -426 2994
rect -364 -2994 -347 2994
rect -285 -2994 -268 2994
rect -206 -2994 -189 2994
rect -127 -2994 -110 2994
rect -48 -2994 -31 2994
rect 31 -2994 48 2994
rect 110 -2994 127 2994
rect 189 -2994 206 2994
rect 268 -2994 285 2994
rect 347 -2994 364 2994
rect 426 -2994 443 2994
rect 505 -2994 522 2994
rect 584 -2994 601 2994
rect 663 -2994 680 2994
rect 742 -2994 759 2994
rect 821 -2994 838 2994
rect 900 -2994 917 2994
rect 979 -2994 996 2994
rect -965 -3036 -931 -3019
rect -886 -3036 -852 -3019
rect -807 -3036 -773 -3019
rect -728 -3036 -694 -3019
rect -649 -3036 -615 -3019
rect -570 -3036 -536 -3019
rect -491 -3036 -457 -3019
rect -412 -3036 -378 -3019
rect -333 -3036 -299 -3019
rect -254 -3036 -220 -3019
rect -175 -3036 -141 -3019
rect -96 -3036 -62 -3019
rect -17 -3036 17 -3019
rect 62 -3036 96 -3019
rect 141 -3036 175 -3019
rect 220 -3036 254 -3019
rect 299 -3036 333 -3019
rect 378 -3036 412 -3019
rect 457 -3036 491 -3019
rect 536 -3036 570 -3019
rect 615 -3036 649 -3019
rect 694 -3036 728 -3019
rect 773 -3036 807 -3019
rect 852 -3036 886 -3019
rect 931 -3036 965 -3019
<< metal1 >>
rect -971 3036 -925 3039
rect -971 3019 -965 3036
rect -931 3019 -925 3036
rect -971 3016 -925 3019
rect -892 3036 -846 3039
rect -892 3019 -886 3036
rect -852 3019 -846 3036
rect -892 3016 -846 3019
rect -813 3036 -767 3039
rect -813 3019 -807 3036
rect -773 3019 -767 3036
rect -813 3016 -767 3019
rect -734 3036 -688 3039
rect -734 3019 -728 3036
rect -694 3019 -688 3036
rect -734 3016 -688 3019
rect -655 3036 -609 3039
rect -655 3019 -649 3036
rect -615 3019 -609 3036
rect -655 3016 -609 3019
rect -576 3036 -530 3039
rect -576 3019 -570 3036
rect -536 3019 -530 3036
rect -576 3016 -530 3019
rect -497 3036 -451 3039
rect -497 3019 -491 3036
rect -457 3019 -451 3036
rect -497 3016 -451 3019
rect -418 3036 -372 3039
rect -418 3019 -412 3036
rect -378 3019 -372 3036
rect -418 3016 -372 3019
rect -339 3036 -293 3039
rect -339 3019 -333 3036
rect -299 3019 -293 3036
rect -339 3016 -293 3019
rect -260 3036 -214 3039
rect -260 3019 -254 3036
rect -220 3019 -214 3036
rect -260 3016 -214 3019
rect -181 3036 -135 3039
rect -181 3019 -175 3036
rect -141 3019 -135 3036
rect -181 3016 -135 3019
rect -102 3036 -56 3039
rect -102 3019 -96 3036
rect -62 3019 -56 3036
rect -102 3016 -56 3019
rect -23 3036 23 3039
rect -23 3019 -17 3036
rect 17 3019 23 3036
rect -23 3016 23 3019
rect 56 3036 102 3039
rect 56 3019 62 3036
rect 96 3019 102 3036
rect 56 3016 102 3019
rect 135 3036 181 3039
rect 135 3019 141 3036
rect 175 3019 181 3036
rect 135 3016 181 3019
rect 214 3036 260 3039
rect 214 3019 220 3036
rect 254 3019 260 3036
rect 214 3016 260 3019
rect 293 3036 339 3039
rect 293 3019 299 3036
rect 333 3019 339 3036
rect 293 3016 339 3019
rect 372 3036 418 3039
rect 372 3019 378 3036
rect 412 3019 418 3036
rect 372 3016 418 3019
rect 451 3036 497 3039
rect 451 3019 457 3036
rect 491 3019 497 3036
rect 451 3016 497 3019
rect 530 3036 576 3039
rect 530 3019 536 3036
rect 570 3019 576 3036
rect 530 3016 576 3019
rect 609 3036 655 3039
rect 609 3019 615 3036
rect 649 3019 655 3036
rect 609 3016 655 3019
rect 688 3036 734 3039
rect 688 3019 694 3036
rect 728 3019 734 3036
rect 688 3016 734 3019
rect 767 3036 813 3039
rect 767 3019 773 3036
rect 807 3019 813 3036
rect 767 3016 813 3019
rect 846 3036 892 3039
rect 846 3019 852 3036
rect 886 3019 892 3036
rect 846 3016 892 3019
rect 925 3036 971 3039
rect 925 3019 931 3036
rect 965 3019 971 3036
rect 925 3016 971 3019
rect -999 2994 -976 3000
rect -999 -2994 -996 2994
rect -979 -2994 -976 2994
rect -999 -3000 -976 -2994
rect -920 2994 -897 3000
rect -920 -2994 -917 2994
rect -900 -2994 -897 2994
rect -920 -3000 -897 -2994
rect -841 2994 -818 3000
rect -841 -2994 -838 2994
rect -821 -2994 -818 2994
rect -841 -3000 -818 -2994
rect -762 2994 -739 3000
rect -762 -2994 -759 2994
rect -742 -2994 -739 2994
rect -762 -3000 -739 -2994
rect -683 2994 -660 3000
rect -683 -2994 -680 2994
rect -663 -2994 -660 2994
rect -683 -3000 -660 -2994
rect -604 2994 -581 3000
rect -604 -2994 -601 2994
rect -584 -2994 -581 2994
rect -604 -3000 -581 -2994
rect -525 2994 -502 3000
rect -525 -2994 -522 2994
rect -505 -2994 -502 2994
rect -525 -3000 -502 -2994
rect -446 2994 -423 3000
rect -446 -2994 -443 2994
rect -426 -2994 -423 2994
rect -446 -3000 -423 -2994
rect -367 2994 -344 3000
rect -367 -2994 -364 2994
rect -347 -2994 -344 2994
rect -367 -3000 -344 -2994
rect -288 2994 -265 3000
rect -288 -2994 -285 2994
rect -268 -2994 -265 2994
rect -288 -3000 -265 -2994
rect -209 2994 -186 3000
rect -209 -2994 -206 2994
rect -189 -2994 -186 2994
rect -209 -3000 -186 -2994
rect -130 2994 -107 3000
rect -130 -2994 -127 2994
rect -110 -2994 -107 2994
rect -130 -3000 -107 -2994
rect -51 2994 -28 3000
rect -51 -2994 -48 2994
rect -31 -2994 -28 2994
rect -51 -3000 -28 -2994
rect 28 2994 51 3000
rect 28 -2994 31 2994
rect 48 -2994 51 2994
rect 28 -3000 51 -2994
rect 107 2994 130 3000
rect 107 -2994 110 2994
rect 127 -2994 130 2994
rect 107 -3000 130 -2994
rect 186 2994 209 3000
rect 186 -2994 189 2994
rect 206 -2994 209 2994
rect 186 -3000 209 -2994
rect 265 2994 288 3000
rect 265 -2994 268 2994
rect 285 -2994 288 2994
rect 265 -3000 288 -2994
rect 344 2994 367 3000
rect 344 -2994 347 2994
rect 364 -2994 367 2994
rect 344 -3000 367 -2994
rect 423 2994 446 3000
rect 423 -2994 426 2994
rect 443 -2994 446 2994
rect 423 -3000 446 -2994
rect 502 2994 525 3000
rect 502 -2994 505 2994
rect 522 -2994 525 2994
rect 502 -3000 525 -2994
rect 581 2994 604 3000
rect 581 -2994 584 2994
rect 601 -2994 604 2994
rect 581 -3000 604 -2994
rect 660 2994 683 3000
rect 660 -2994 663 2994
rect 680 -2994 683 2994
rect 660 -3000 683 -2994
rect 739 2994 762 3000
rect 739 -2994 742 2994
rect 759 -2994 762 2994
rect 739 -3000 762 -2994
rect 818 2994 841 3000
rect 818 -2994 821 2994
rect 838 -2994 841 2994
rect 818 -3000 841 -2994
rect 897 2994 920 3000
rect 897 -2994 900 2994
rect 917 -2994 920 2994
rect 897 -3000 920 -2994
rect 976 2994 999 3000
rect 976 -2994 979 2994
rect 996 -2994 999 2994
rect 976 -3000 999 -2994
rect -971 -3019 -925 -3016
rect -971 -3036 -965 -3019
rect -931 -3036 -925 -3019
rect -971 -3039 -925 -3036
rect -892 -3019 -846 -3016
rect -892 -3036 -886 -3019
rect -852 -3036 -846 -3019
rect -892 -3039 -846 -3036
rect -813 -3019 -767 -3016
rect -813 -3036 -807 -3019
rect -773 -3036 -767 -3019
rect -813 -3039 -767 -3036
rect -734 -3019 -688 -3016
rect -734 -3036 -728 -3019
rect -694 -3036 -688 -3019
rect -734 -3039 -688 -3036
rect -655 -3019 -609 -3016
rect -655 -3036 -649 -3019
rect -615 -3036 -609 -3019
rect -655 -3039 -609 -3036
rect -576 -3019 -530 -3016
rect -576 -3036 -570 -3019
rect -536 -3036 -530 -3019
rect -576 -3039 -530 -3036
rect -497 -3019 -451 -3016
rect -497 -3036 -491 -3019
rect -457 -3036 -451 -3019
rect -497 -3039 -451 -3036
rect -418 -3019 -372 -3016
rect -418 -3036 -412 -3019
rect -378 -3036 -372 -3019
rect -418 -3039 -372 -3036
rect -339 -3019 -293 -3016
rect -339 -3036 -333 -3019
rect -299 -3036 -293 -3019
rect -339 -3039 -293 -3036
rect -260 -3019 -214 -3016
rect -260 -3036 -254 -3019
rect -220 -3036 -214 -3019
rect -260 -3039 -214 -3036
rect -181 -3019 -135 -3016
rect -181 -3036 -175 -3019
rect -141 -3036 -135 -3019
rect -181 -3039 -135 -3036
rect -102 -3019 -56 -3016
rect -102 -3036 -96 -3019
rect -62 -3036 -56 -3019
rect -102 -3039 -56 -3036
rect -23 -3019 23 -3016
rect -23 -3036 -17 -3019
rect 17 -3036 23 -3019
rect -23 -3039 23 -3036
rect 56 -3019 102 -3016
rect 56 -3036 62 -3019
rect 96 -3036 102 -3019
rect 56 -3039 102 -3036
rect 135 -3019 181 -3016
rect 135 -3036 141 -3019
rect 175 -3036 181 -3019
rect 135 -3039 181 -3036
rect 214 -3019 260 -3016
rect 214 -3036 220 -3019
rect 254 -3036 260 -3019
rect 214 -3039 260 -3036
rect 293 -3019 339 -3016
rect 293 -3036 299 -3019
rect 333 -3036 339 -3019
rect 293 -3039 339 -3036
rect 372 -3019 418 -3016
rect 372 -3036 378 -3019
rect 412 -3036 418 -3019
rect 372 -3039 418 -3036
rect 451 -3019 497 -3016
rect 451 -3036 457 -3019
rect 491 -3036 497 -3019
rect 451 -3039 497 -3036
rect 530 -3019 576 -3016
rect 530 -3036 536 -3019
rect 570 -3036 576 -3019
rect 530 -3039 576 -3036
rect 609 -3019 655 -3016
rect 609 -3036 615 -3019
rect 649 -3036 655 -3019
rect 609 -3039 655 -3036
rect 688 -3019 734 -3016
rect 688 -3036 694 -3019
rect 728 -3036 734 -3019
rect 688 -3039 734 -3036
rect 767 -3019 813 -3016
rect 767 -3036 773 -3019
rect 807 -3036 813 -3019
rect 767 -3039 813 -3036
rect 846 -3019 892 -3016
rect 846 -3036 852 -3019
rect 886 -3036 892 -3019
rect 846 -3039 892 -3036
rect 925 -3019 971 -3016
rect 925 -3036 931 -3019
rect 965 -3036 971 -3019
rect 925 -3039 971 -3036
<< properties >>
string FIXED_BBOX -1054 -3096 1054 3096
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 60 l 0.50 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
