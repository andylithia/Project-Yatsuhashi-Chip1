magic
tech sky130B
magscale 1 2
timestamp 1620310959
