magic
tech sky130B
magscale 1 2
timestamp 1662654558
<< metal1 >>
rect 580 3220 1400 3359
rect 2330 3300 2530 4860
rect 580 3120 610 3220
rect 1360 3120 1400 3220
rect 1480 3180 4260 3220
rect 1480 3080 1520 3180
rect 4240 3080 4260 3180
rect 1480 3040 4260 3080
rect 1480 100 4330 140
rect 650 -216 1419 98
rect 1480 0 1520 100
rect 4240 0 4330 100
rect 1480 -40 4330 0
rect 2309 -1750 2542 -182
<< via1 >>
rect 610 3120 1360 3220
rect 1520 3080 4240 3180
rect 1520 0 4240 100
<< metal2 >>
rect -600 4300 600 4800
rect 300 3300 600 4300
rect 2320 4139 2520 4860
rect 2323 4057 2522 4111
rect 4183 4057 4330 4111
rect -100 3250 600 3300
rect -100 3220 1390 3250
rect 1481 3220 1535 3300
rect 2400 3220 2470 4057
rect 3331 3220 3385 3300
rect 4260 3220 4330 4057
rect -100 3120 610 3220
rect 1360 3120 1390 3220
rect -100 3100 1390 3120
rect 1480 3180 4330 3220
rect -100 1400 100 3100
rect 1480 3080 1520 3180
rect 4240 3080 4330 3180
rect 1480 3040 4330 3080
rect 4260 2900 4330 3040
rect -380 440 0 470
rect -4000 420 -3600 440
rect -4000 380 -3980 420
rect -3620 380 -3600 420
rect -380 300 -360 440
rect -20 300 0 440
rect 4200 300 4400 2900
rect -380 280 0 300
rect 4250 260 4400 300
rect 4160 140 4400 260
rect 1480 100 4400 140
rect 0 39 211 76
rect 0 -219 677 39
rect 1480 0 1520 100
rect 4240 0 4400 100
rect 1480 -40 4400 0
rect 1481 -212 1535 -40
rect 9 -374 677 -219
rect 2398 -939 2468 -40
rect 3331 -237 3385 -40
rect 4250 -939 4400 -40
rect 2300 -993 2566 -939
rect 4145 -993 4400 -939
rect 4250 -995 4400 -993
rect 2309 -1750 2554 -1021
<< via2 >>
rect -3980 300 -3620 420
rect -2680 300 -2320 420
rect -1580 300 -1220 420
rect -360 300 -20 440
<< metal3 >>
rect -600 5700 500 5800
rect -600 4900 -500 5700
rect 400 4900 500 5700
rect -600 4400 500 4900
rect -250 1250 100 1300
rect -250 700 -200 1250
rect 50 700 100 1250
rect -250 650 100 700
rect -3500 480 -3220 580
rect -4000 420 -3600 460
rect -4000 300 -3980 420
rect -3620 300 -3600 420
rect -4000 200 -3600 300
rect -3400 -2140 -3220 480
rect -3040 480 -2760 580
rect -3040 -2140 -2860 480
rect -2700 420 -2300 440
rect -2700 300 -2680 420
rect -2320 300 -2300 420
rect -2700 200 -2300 300
rect -2200 -2140 -2020 580
rect -1840 -2140 -1660 580
rect -1600 420 -1200 440
rect -1600 300 -1580 420
rect -1220 300 -1200 420
rect -1600 200 -1200 300
rect -1100 -2140 -920 580
rect -400 440 60 460
rect -400 300 -360 440
rect -20 300 60 440
rect -400 200 60 300
<< via3 >>
rect -500 4900 400 5700
rect 1053 4117 1130 4642
rect 1328 4117 1405 4643
rect 1610 4117 1687 4643
rect 1886 4117 1963 4643
rect 2162 4117 2240 4643
rect 911 4051 2240 4117
rect 2626 4117 2704 4642
rect 2902 4117 2980 4642
rect 3178 4117 3256 4642
rect 3460 4117 3538 4642
rect 3736 4117 3814 4642
rect 2626 4051 3814 4117
rect 1300 1450 1400 2000
rect -200 700 50 1250
rect 1560 1200 1660 1760
rect -3980 300 -3620 420
rect -2680 300 -2320 420
rect -1580 300 -1220 420
rect -360 300 -20 440
rect 776 -995 2230 -933
rect 2626 -995 3813 -933
rect 776 -999 2240 -995
rect 776 -1524 854 -999
rect 1052 -1524 1130 -999
rect 1328 -1524 1406 -999
rect 1610 -1524 1688 -999
rect 1886 -1524 1964 -999
rect 2162 -1525 2240 -999
rect 2626 -999 3814 -995
rect 2626 -1525 2704 -999
rect 2902 -1525 2980 -999
rect 3178 -1525 3256 -999
rect 3460 -1525 3538 -999
rect 3736 -1525 3814 -999
<< metal4 >>
rect 1800 6400 2600 6800
rect -200 5800 2600 6400
rect -5900 5700 2600 5800
rect -5900 5600 -500 5700
rect -5800 4900 -500 5600
rect 400 5000 2600 5700
rect 400 4900 600 5000
rect -5800 4600 600 4900
rect 800 4700 4000 4800
rect -5800 3300 -4800 4600
rect 800 4300 900 4700
rect 3900 4300 4000 4700
rect 800 4117 1053 4300
rect 1130 4117 1328 4300
rect 1405 4117 1610 4300
rect 1687 4117 1886 4300
rect 1963 4117 2162 4300
rect 800 4051 911 4117
rect 2240 4051 2626 4300
rect 2704 4117 2902 4300
rect 2980 4117 3178 4300
rect 3256 4117 3460 4300
rect 3538 4117 3736 4300
rect 3814 4051 4000 4300
rect 800 4000 4000 4051
rect 4400 3600 5200 4100
rect -5800 1400 -5200 3300
rect 1200 3000 5200 3600
rect -4900 2400 -4500 3000
rect 1300 2800 5200 3000
rect 1300 2400 1900 2800
rect -4900 2100 -4400 2400
rect 200 2100 1900 2400
rect -4900 1700 -4500 2100
rect 1250 2000 1450 2100
rect 1250 1450 1300 2000
rect 1400 1450 1450 2000
rect 1250 1400 1450 1450
rect 1540 1760 1720 1800
rect -5800 -1400 -4800 1400
rect -250 1250 100 1300
rect -250 700 -200 1250
rect 50 1050 100 1250
rect 1540 1200 1560 1760
rect 1660 1200 1720 1760
rect 1540 1050 1720 1200
rect 50 750 1720 1050
rect 50 700 1900 750
rect -250 650 1900 700
rect -400 440 200 460
rect -4000 420 -3600 440
rect -4000 300 -3980 420
rect -3620 300 -3600 420
rect -4000 -1400 -3600 300
rect -2700 420 -2300 440
rect -2700 300 -2680 420
rect -2320 300 -2300 420
rect -2700 -1400 -2300 300
rect -1600 420 -1200 440
rect -1600 300 -1580 420
rect -1220 300 -1200 420
rect -1600 -1400 -1200 300
rect -400 300 -360 440
rect -20 300 200 440
rect -400 200 200 300
rect 1300 400 1900 650
rect 1300 200 5200 400
rect -400 -1400 400 200
rect 1200 -400 5200 200
rect 4400 -900 5200 -400
rect -5800 -1900 400 -1400
rect 600 -933 4000 -900
rect 600 -1200 776 -933
rect 2230 -995 2626 -933
rect 3813 -995 4000 -933
rect 854 -1200 1052 -999
rect 1130 -1200 1328 -999
rect 1406 -1200 1610 -999
rect 1688 -1200 1886 -999
rect 1964 -1200 2162 -999
rect 2240 -1200 2626 -995
rect 2704 -1200 2902 -999
rect 2980 -1200 3178 -999
rect 3256 -1200 3460 -999
rect 3538 -1200 3736 -999
rect 3814 -1200 4000 -995
rect 600 -1600 700 -1200
rect 3900 -1600 4000 -1200
rect 600 -1700 4000 -1600
rect -5800 -2000 2600 -1900
rect -400 -3200 2600 -2000
rect 1800 -3600 2600 -3200
<< via4 >>
rect 900 4643 3900 4700
rect 900 4642 1328 4643
rect 900 4300 1053 4642
rect 1053 4300 1130 4642
rect 1130 4300 1328 4642
rect 1328 4300 1405 4643
rect 1405 4300 1610 4643
rect 1610 4300 1687 4643
rect 1687 4300 1886 4643
rect 1886 4300 1963 4643
rect 1963 4300 2162 4643
rect 2162 4300 2240 4643
rect 2240 4642 3900 4643
rect 2240 4300 2626 4642
rect 2626 4300 2704 4642
rect 2704 4300 2902 4642
rect 2902 4300 2980 4642
rect 2980 4300 3178 4642
rect 3178 4300 3256 4642
rect 3256 4300 3460 4642
rect 3460 4300 3538 4642
rect 3538 4300 3736 4642
rect 3736 4300 3814 4642
rect 3814 4300 3900 4642
rect 700 -1524 776 -1200
rect 776 -1524 854 -1200
rect 854 -1524 1052 -1200
rect 1052 -1524 1130 -1200
rect 1130 -1524 1328 -1200
rect 1328 -1524 1406 -1200
rect 1406 -1524 1610 -1200
rect 1610 -1524 1688 -1200
rect 1688 -1524 1886 -1200
rect 1886 -1524 1964 -1200
rect 1964 -1524 2162 -1200
rect 700 -1525 2162 -1524
rect 2162 -1525 2240 -1200
rect 2240 -1525 2626 -1200
rect 2626 -1525 2704 -1200
rect 2704 -1525 2902 -1200
rect 2902 -1525 2980 -1200
rect 2980 -1525 3178 -1200
rect 3178 -1525 3256 -1200
rect 3256 -1525 3460 -1200
rect 3460 -1525 3538 -1200
rect 3538 -1525 3736 -1200
rect 3736 -1525 3814 -1200
rect 3814 -1525 3900 -1200
rect 700 -1600 3900 -1525
<< metal5 >>
rect -5900 5000 4000 5600
rect -5800 4700 4000 5000
rect -5800 4600 900 4700
rect -5800 200 -4800 4600
rect 700 4300 900 4600
rect 3900 4300 4000 4700
rect 700 4200 4000 4300
rect -5800 -200 400 200
rect -5800 -600 -4800 -200
rect -4000 -600 -3600 -200
rect -2800 -600 -2400 -200
rect -1600 -600 -1200 -200
rect -400 -600 400 -200
rect -5800 -1000 400 -600
rect -5800 -1400 -4800 -1000
rect -4000 -1400 -3600 -1000
rect -2800 -1400 -2400 -1000
rect -1600 -1400 -1200 -1000
rect -400 -1100 400 -1000
rect -400 -1200 4000 -1100
rect -400 -1400 700 -1200
rect -5800 -1600 700 -1400
rect 3900 -1600 4000 -1200
rect -5800 -1800 4000 -1600
rect -400 -2400 4000 -1800
use XCP_1  XCP_1_0
timestamp 1662654558
transform 1 0 1440 0 1 0
box -1440 0 2918 3190
use captuner_complete_2  captuner_complete_2_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659228637
transform 0 1 -2000 -1 0 3050
box -1150 -2500 2770 2500
use sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1653785680
transform 1 0 650 0 1 3300
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1_1
timestamp 1653785680
transform 1 0 2500 0 1 3300
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1_2
timestamp 1653785680
transform 1 0 650 0 1 -1750
box 0 0 1716 1568
use sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1  sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1_3
timestamp 1653785680
transform 1 0 2500 0 1 -1750
box 0 0 1716 1568
<< labels >>
rlabel metal5 -5900 5000 -5800 5600 1 VH
rlabel metal4 -5900 5600 -5800 5800 1 VL
rlabel metal4 4400 3000 5200 6000 1 I1
rlabel metal4 4400 -2800 5200 200 1 I2
rlabel metal3 -3400 -2140 -3220 -2080 1 G3
rlabel metal3 -3040 -2140 -2860 -2080 1 G2
rlabel metal3 -2200 -2140 -2020 -2080 1 G1
rlabel metal3 -1840 -2140 -1660 -2080 1 G0
rlabel metal3 -1100 -2140 -920 -2080 1 G4
<< end >>
