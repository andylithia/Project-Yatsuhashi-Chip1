magic
tech sky130B
timestamp 1662579390
<< nwell >>
rect -2318 -169 2318 169
<< pwell >>
rect -2387 169 2387 238
rect -2387 -169 -2318 169
rect 2318 -169 2387 169
rect -2387 -238 2387 -169
<< psubdiff >>
rect -2369 203 -2321 220
rect 2321 203 2369 220
rect -2369 172 -2352 203
rect 2352 172 2369 203
rect -2369 -203 -2352 -172
rect 2352 -203 2369 -172
rect -2369 -220 -2321 -203
rect 2321 -220 2369 -203
<< nsubdiff >>
rect -2300 134 -2252 151
rect -1246 134 -1198 151
rect -2300 103 -2283 134
rect -1215 103 -1198 134
rect -2300 -134 -2283 -103
rect -1215 -134 -1198 -103
rect -2300 -151 -2252 -134
rect -1246 -151 -1198 -134
rect -1134 134 -1086 151
rect -80 134 -32 151
rect -1134 103 -1117 134
rect -49 103 -32 134
rect -1134 -134 -1117 -103
rect -49 -134 -32 -103
rect -1134 -151 -1086 -134
rect -80 -151 -32 -134
rect 32 134 80 151
rect 1086 134 1134 151
rect 32 103 49 134
rect 1117 103 1134 134
rect 32 -134 49 -103
rect 1117 -134 1134 -103
rect 32 -151 80 -134
rect 1086 -151 1134 -134
rect 1198 134 1246 151
rect 2252 134 2300 151
rect 1198 103 1215 134
rect 2283 103 2300 134
rect 1198 -134 1215 -103
rect 2283 -134 2300 -103
rect 1198 -151 1246 -134
rect 2252 -151 2300 -134
<< psubdiffcont >>
rect -2321 203 2321 220
rect -2369 -172 -2352 172
rect 2352 -172 2369 172
rect -2321 -220 2321 -203
<< nsubdiffcont >>
rect -2252 134 -1246 151
rect -2300 -103 -2283 103
rect -1215 -103 -1198 103
rect -2252 -151 -1246 -134
rect -1086 134 -80 151
rect -1134 -103 -1117 103
rect -49 -103 -32 103
rect -1086 -151 -80 -134
rect 80 134 1086 151
rect 32 -103 49 103
rect 1117 -103 1134 103
rect 80 -151 1086 -134
rect 1246 134 2252 151
rect 1198 -103 1215 103
rect 2283 -103 2300 103
rect 1246 -151 2252 -134
<< pdiode >>
rect -2249 94 -1249 100
rect -2249 -94 -2243 94
rect -1255 -94 -1249 94
rect -2249 -100 -1249 -94
rect -1083 94 -83 100
rect -1083 -94 -1077 94
rect -89 -94 -83 94
rect -1083 -100 -83 -94
rect 83 94 1083 100
rect 83 -94 89 94
rect 1077 -94 1083 94
rect 83 -100 1083 -94
rect 1249 94 2249 100
rect 1249 -94 1255 94
rect 2243 -94 2249 94
rect 1249 -100 2249 -94
<< pdiodec >>
rect -2243 -94 -1255 94
rect -1077 -94 -89 94
rect 89 -94 1077 94
rect 1255 -94 2243 94
<< locali >>
rect -2369 203 -2321 220
rect 2321 203 2369 220
rect -2369 172 -2352 203
rect 2352 172 2369 203
rect -2300 134 -2252 151
rect -1246 134 -1198 151
rect -2300 103 -2283 134
rect -1215 103 -1198 134
rect -2251 -94 -2243 94
rect -1255 -94 -1247 94
rect -2300 -134 -2283 -103
rect -1215 -134 -1198 -103
rect -2300 -151 -2252 -134
rect -1246 -151 -1198 -134
rect -1134 134 -1086 151
rect -80 134 -32 151
rect -1134 103 -1117 134
rect -49 103 -32 134
rect -1085 -94 -1077 94
rect -89 -94 -81 94
rect -1134 -134 -1117 -103
rect -49 -134 -32 -103
rect -1134 -151 -1086 -134
rect -80 -151 -32 -134
rect 32 134 80 151
rect 1086 134 1134 151
rect 32 103 49 134
rect 1117 103 1134 134
rect 81 -94 89 94
rect 1077 -94 1085 94
rect 32 -134 49 -103
rect 1117 -134 1134 -103
rect 32 -151 80 -134
rect 1086 -151 1134 -134
rect 1198 134 1246 151
rect 2252 134 2300 151
rect 1198 103 1215 134
rect 2283 103 2300 134
rect 1247 -94 1255 94
rect 2243 -94 2251 94
rect 1198 -134 1215 -103
rect 2283 -134 2300 -103
rect 1198 -151 1246 -134
rect 2252 -151 2300 -134
rect -2369 -203 -2352 -172
rect 2352 -203 2369 -172
rect -2369 -220 -2321 -203
rect 2321 -220 2369 -203
<< viali >>
rect -2243 -94 -1255 94
rect -1077 -94 -89 94
rect 89 -94 1077 94
rect 1255 -94 2243 94
<< metal1 >>
rect -2249 94 -1249 97
rect -2249 -94 -2243 94
rect -1255 -94 -1249 94
rect -2249 -97 -1249 -94
rect -1083 94 -83 97
rect -1083 -94 -1077 94
rect -89 -94 -83 94
rect -1083 -97 -83 -94
rect 83 94 1083 97
rect 83 -94 89 94
rect 1077 -94 1083 94
rect 83 -97 1083 -94
rect 1249 94 2249 97
rect 1249 -94 1255 94
rect 2243 -94 2249 94
rect 1249 -97 2249 -94
<< properties >>
string FIXED_BBOX 1206 -142 2291 142
string gencell sky130_fd_pr__diode_pd2nw_05v5
string library sky130
string parameters w 10 l 2 area 20.0 peri 24.0 nx 4 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
