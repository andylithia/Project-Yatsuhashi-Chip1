magic
tech sky130B
magscale 1 2
timestamp 1662175719
<< error_p >>
rect -29 1049 29 1055
rect -29 1015 -17 1049
rect -29 1009 29 1015
rect -29 433 29 439
rect -29 399 -17 433
rect -29 393 29 399
rect -29 325 29 331
rect -29 291 -17 325
rect -29 285 29 291
rect -29 -291 29 -285
rect -29 -325 -17 -291
rect -29 -331 29 -325
rect -29 -399 29 -393
rect -29 -433 -17 -399
rect -29 -439 29 -433
rect -29 -1015 29 -1009
rect -29 -1049 -17 -1015
rect -29 -1055 29 -1049
<< pwell >>
rect -211 -1187 211 1187
<< nmos >>
rect -15 471 15 977
rect -15 -253 15 253
rect -15 -977 15 -471
<< ndiff >>
rect -73 965 -15 977
rect -73 483 -61 965
rect -27 483 -15 965
rect -73 471 -15 483
rect 15 965 73 977
rect 15 483 27 965
rect 61 483 73 965
rect 15 471 73 483
rect -73 241 -15 253
rect -73 -241 -61 241
rect -27 -241 -15 241
rect -73 -253 -15 -241
rect 15 241 73 253
rect 15 -241 27 241
rect 61 -241 73 241
rect 15 -253 73 -241
rect -73 -483 -15 -471
rect -73 -965 -61 -483
rect -27 -965 -15 -483
rect -73 -977 -15 -965
rect 15 -483 73 -471
rect 15 -965 27 -483
rect 61 -965 73 -483
rect 15 -977 73 -965
<< ndiffc >>
rect -61 483 -27 965
rect 27 483 61 965
rect -61 -241 -27 241
rect 27 -241 61 241
rect -61 -965 -27 -483
rect 27 -965 61 -483
<< psubdiff >>
rect -175 1117 -79 1151
rect 79 1117 175 1151
rect -175 1055 -141 1117
rect 141 1055 175 1117
rect -175 -1117 -141 -1055
rect 141 -1117 175 -1055
rect -175 -1151 -79 -1117
rect 79 -1151 175 -1117
<< psubdiffcont >>
rect -79 1117 79 1151
rect -175 -1055 -141 1055
rect 141 -1055 175 1055
rect -79 -1151 79 -1117
<< poly >>
rect -33 1049 33 1065
rect -33 1015 -17 1049
rect 17 1015 33 1049
rect -33 999 33 1015
rect -15 977 15 999
rect -15 449 15 471
rect -33 433 33 449
rect -33 399 -17 433
rect 17 399 33 433
rect -33 383 33 399
rect -33 325 33 341
rect -33 291 -17 325
rect 17 291 33 325
rect -33 275 33 291
rect -15 253 15 275
rect -15 -275 15 -253
rect -33 -291 33 -275
rect -33 -325 -17 -291
rect 17 -325 33 -291
rect -33 -341 33 -325
rect -33 -399 33 -383
rect -33 -433 -17 -399
rect 17 -433 33 -399
rect -33 -449 33 -433
rect -15 -471 15 -449
rect -15 -999 15 -977
rect -33 -1015 33 -999
rect -33 -1049 -17 -1015
rect 17 -1049 33 -1015
rect -33 -1065 33 -1049
<< polycont >>
rect -17 1015 17 1049
rect -17 399 17 433
rect -17 291 17 325
rect -17 -325 17 -291
rect -17 -433 17 -399
rect -17 -1049 17 -1015
<< locali >>
rect -175 1117 -79 1151
rect 79 1117 175 1151
rect -175 1055 -141 1117
rect 141 1055 175 1117
rect -33 1015 -17 1049
rect 17 1015 33 1049
rect -61 965 -27 981
rect -61 467 -27 483
rect 27 965 61 981
rect 27 467 61 483
rect -33 399 -17 433
rect 17 399 33 433
rect -33 291 -17 325
rect 17 291 33 325
rect -61 241 -27 257
rect -61 -257 -27 -241
rect 27 241 61 257
rect 27 -257 61 -241
rect -33 -325 -17 -291
rect 17 -325 33 -291
rect -33 -433 -17 -399
rect 17 -433 33 -399
rect -61 -483 -27 -467
rect -61 -981 -27 -965
rect 27 -483 61 -467
rect 27 -981 61 -965
rect -33 -1049 -17 -1015
rect 17 -1049 33 -1015
rect -175 -1117 -141 -1055
rect 141 -1117 175 -1055
rect -175 -1151 -79 -1117
rect 79 -1151 175 -1117
<< viali >>
rect -17 1015 17 1049
rect -61 483 -27 965
rect 27 483 61 965
rect -17 399 17 433
rect -17 291 17 325
rect -61 -241 -27 241
rect 27 -241 61 241
rect -17 -325 17 -291
rect -17 -433 17 -399
rect -61 -965 -27 -483
rect 27 -965 61 -483
rect -17 -1049 17 -1015
<< metal1 >>
rect -29 1049 29 1055
rect -29 1015 -17 1049
rect 17 1015 29 1049
rect -29 1009 29 1015
rect -67 965 -21 977
rect -67 483 -61 965
rect -27 483 -21 965
rect -67 471 -21 483
rect 21 965 67 977
rect 21 483 27 965
rect 61 483 67 965
rect 21 471 67 483
rect -29 433 29 439
rect -29 399 -17 433
rect 17 399 29 433
rect -29 393 29 399
rect -29 325 29 331
rect -29 291 -17 325
rect 17 291 29 325
rect -29 285 29 291
rect -67 241 -21 253
rect -67 -241 -61 241
rect -27 -241 -21 241
rect -67 -253 -21 -241
rect 21 241 67 253
rect 21 -241 27 241
rect 61 -241 67 241
rect 21 -253 67 -241
rect -29 -291 29 -285
rect -29 -325 -17 -291
rect 17 -325 29 -291
rect -29 -331 29 -325
rect -29 -399 29 -393
rect -29 -433 -17 -399
rect 17 -433 29 -399
rect -29 -439 29 -433
rect -67 -483 -21 -471
rect -67 -965 -61 -483
rect -27 -965 -21 -483
rect -67 -977 -21 -965
rect 21 -483 67 -471
rect 21 -965 27 -483
rect 61 -965 67 -483
rect 21 -977 67 -965
rect -29 -1015 29 -1009
rect -29 -1049 -17 -1015
rect 17 -1049 29 -1015
rect -29 -1055 29 -1049
<< properties >>
string FIXED_BBOX -158 -1134 158 1134
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.53 l 0.150 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
