magic
tech sky130A
timestamp 1659146707
<< metal1 >>
rect 1290 891 1340 900
rect 600 862 1340 891
rect 1120 800 1270 810
rect 1120 790 1240 800
rect 1230 770 1240 790
rect 1120 750 1240 770
rect 1230 730 1240 750
rect 1120 710 1240 730
rect 1230 690 1240 710
rect 1120 680 1240 690
rect 1120 670 1270 680
rect 1290 608 1340 862
rect 600 579 1340 608
rect 1114 520 1270 530
rect 1114 510 1240 520
rect 1230 490 1240 510
rect 1114 470 1240 490
rect 1230 450 1240 470
rect 1114 430 1240 450
rect 1230 410 1240 430
rect 1114 400 1240 410
rect 1114 390 1270 400
rect 1290 325 1340 579
rect 600 296 1340 325
rect 1114 230 1270 240
rect 1114 220 1240 230
rect 1230 200 1240 220
rect 1114 180 1240 200
rect 1230 160 1240 180
rect 1114 140 1240 160
rect 1230 120 1240 140
rect 1114 110 1240 120
rect 1114 100 1270 110
rect 1290 42 1340 296
rect 600 13 1340 42
rect 1114 -50 1270 -40
rect 1114 -60 1240 -50
rect 1230 -80 1240 -60
rect 1114 -100 1240 -80
rect 1230 -120 1240 -100
rect 1114 -140 1240 -120
rect 1230 -160 1240 -140
rect 1114 -170 1240 -160
rect 1114 -180 1270 -170
rect 1290 -241 1340 13
rect 600 -270 1340 -241
rect 1114 -340 1270 -330
rect 1114 -350 1240 -340
rect 1230 -370 1240 -350
rect 1114 -390 1240 -370
rect 1230 -410 1240 -390
rect 1114 -430 1240 -410
rect 1230 -450 1240 -430
rect 1114 -460 1240 -450
rect 1114 -470 1270 -460
rect 1290 -524 1340 -270
rect 600 -553 1340 -524
rect 1114 -620 1270 -610
rect 1114 -630 1240 -620
rect 1230 -650 1240 -630
rect 1114 -670 1240 -650
rect 1230 -690 1240 -670
rect 1114 -710 1240 -690
rect 1230 -730 1240 -710
rect 1114 -740 1240 -730
rect 1114 -750 1270 -740
rect 1290 -807 1340 -553
rect 600 -836 1340 -807
rect 1114 -900 1270 -890
rect 1114 -910 1240 -900
rect 1230 -930 1240 -910
rect 1114 -950 1240 -930
rect 1230 -970 1240 -950
rect 1114 -990 1240 -970
rect 1230 -1010 1240 -990
rect 1114 -1020 1240 -1010
rect 1114 -1030 1270 -1020
rect 1290 -1090 1340 -836
rect 600 -1119 1340 -1090
rect 1290 -1130 1340 -1119
<< via1 >>
rect 1240 680 1270 800
rect 1240 400 1270 520
rect 1240 110 1270 230
rect 1240 -170 1270 -50
rect 1240 -460 1270 -340
rect 1240 -740 1270 -620
rect 1240 -1020 1270 -900
<< metal2 >>
rect 1150 890 1200 900
rect 490 790 550 800
rect 490 390 500 790
rect 540 390 550 790
rect 490 380 550 390
rect 490 210 540 240
rect 490 120 500 210
rect 530 120 540 210
rect 490 100 540 120
rect 490 -60 540 -50
rect 490 -170 500 -60
rect 530 -170 540 -60
rect 490 -180 540 -170
rect 490 -340 540 -330
rect 490 -450 500 -340
rect 530 -450 540 -340
rect 490 -460 540 -450
rect 490 -710 540 -623
rect 490 -1020 500 -710
rect 530 -1020 540 -710
rect 1150 -1140 1160 890
rect 1190 -1140 1200 890
rect 1230 800 1290 810
rect 1230 680 1240 800
rect 1270 680 1290 800
rect 1230 675 1290 680
rect 1230 670 1375 675
rect 1250 600 1375 670
rect 1250 530 1290 600
rect 1230 520 1290 530
rect 1230 400 1240 520
rect 1270 400 1290 520
rect 1230 390 1290 400
rect 1230 230 1270 240
rect 1230 110 1240 230
rect 1270 150 1375 225
rect 1230 100 1270 110
rect 1230 -50 1270 -40
rect 1230 -170 1240 -50
rect 1270 -125 1375 -50
rect 1230 -180 1270 -170
rect 1230 -340 1270 -330
rect 1230 -460 1240 -340
rect 1270 -425 1375 -350
rect 1230 -470 1270 -460
rect 1230 -620 1290 -610
rect 1230 -740 1240 -620
rect 1270 -740 1290 -620
rect 1230 -750 1290 -740
rect 1250 -775 1290 -750
rect 1250 -850 1375 -775
rect 1250 -890 1290 -850
rect 1230 -900 1290 -890
rect 1230 -1020 1240 -900
rect 1270 -1020 1290 -900
rect 1230 -1030 1290 -1020
rect 1150 -1150 1200 -1140
<< via2 >>
rect 500 390 540 790
rect 500 120 530 210
rect 500 -170 530 -60
rect 500 -450 530 -340
rect 500 -1020 530 -710
rect 1160 -1140 1190 890
<< metal3 >>
rect -575 800 475 1200
rect 1050 890 1200 975
rect -575 790 550 800
rect -575 390 500 790
rect 540 390 550 790
rect -575 375 550 390
rect -575 350 475 375
rect -75 210 550 225
rect -75 120 500 210
rect 530 120 550 210
rect -75 100 550 120
rect -75 75 475 100
rect -575 -60 540 -50
rect -575 -170 500 -60
rect 530 -170 540 -60
rect -575 -180 540 -170
rect -575 -200 475 -180
rect -575 -330 475 -325
rect -575 -340 540 -330
rect -575 -450 500 -340
rect 530 -450 540 -340
rect -575 -460 540 -450
rect -575 -575 475 -460
rect -575 -710 540 -700
rect -575 -1020 500 -710
rect 530 -1020 540 -710
rect -575 -1040 540 -1020
rect -575 -1150 475 -1040
rect 1050 -1140 1160 890
rect 1190 -1140 1200 890
rect 1050 -1225 1200 -1140
<< mimcap >>
rect -550 1150 450 1175
rect -550 400 -525 1150
rect 425 400 450 1150
rect -550 375 450 400
rect -50 175 450 200
rect -50 125 -25 175
rect 425 125 450 175
rect -50 100 450 125
rect -550 -100 450 -75
rect -550 -150 -525 -100
rect 425 -150 450 -100
rect -550 -175 450 -150
rect -550 -375 450 -350
rect -550 -525 -525 -375
rect 425 -525 450 -375
rect -550 -550 450 -525
rect -550 -750 450 -725
rect -550 -1100 -525 -750
rect 425 -1100 450 -750
rect -550 -1125 450 -1100
<< mimcapcontact >>
rect -525 400 425 1150
rect -25 125 425 175
rect -525 -150 425 -100
rect -525 -525 425 -375
rect -525 -1100 425 -750
<< metal4 >>
rect 325 1200 475 1250
rect -575 1150 475 1200
rect -575 400 -525 1150
rect 425 400 475 1150
rect -575 350 475 400
rect 325 225 475 350
rect -75 175 475 225
rect -75 125 -25 175
rect 425 125 475 175
rect -75 75 475 125
rect 325 -50 475 75
rect -575 -100 475 -50
rect -575 -150 -525 -100
rect 425 -150 475 -100
rect -575 -200 475 -150
rect 325 -325 475 -200
rect -575 -375 475 -325
rect -575 -525 -525 -375
rect 425 -525 475 -375
rect -575 -575 475 -525
rect 325 -700 475 -575
rect -575 -750 475 -700
rect -575 -1100 -525 -750
rect 425 -1100 475 -750
rect -575 -1150 475 -1100
rect 325 -1250 475 -1150
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_0
timestamp 1659146707
transform 0 1 550 -1 0 338
box 0 -32 338 629
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_1
timestamp 1659146707
transform 0 1 550 -1 0 55
box 0 -32 338 629
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_2
timestamp 1659146707
transform 0 1 550 -1 0 -228
box 0 -32 338 629
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_3
timestamp 1659146707
transform 0 1 550 -1 0 -511
box 0 -32 338 629
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_4
timestamp 1659146707
transform 0 1 550 -1 0 -794
box 0 -32 338 629
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_5
timestamp 1659146707
transform 0 1 550 -1 0 621
box 0 -32 338 629
use sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered  sky130_fd_pr__rf_nfet_01v8_aM04W5p00L0p15_fingered_6
timestamp 1659146707
transform 0 1 550 -1 0 904
box 0 -32 338 629
<< labels >>
rlabel metal2 1350 600 1375 675 1 G4
rlabel metal2 1350 150 1375 225 1 G0
rlabel metal2 1350 -125 1375 -50 1 G1
rlabel metal2 1350 -425 1375 -350 1 G2
rlabel metal2 1350 -850 1375 -775 1 G3
rlabel metal3 1050 -1225 1200 -1150 1 BOT
rlabel metal4 325 -1250 475 -1200 1 TOP
rlabel metal1 1290 840 1340 900 1 SUB
<< end >>
