magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< error_s >>
rect 595 680 653 686
rect 595 646 607 680
rect 595 640 653 646
<< poly >>
rect 297 630 327 684
rect 297 28 327 54
<< locali >>
rect 80 1243 379 1277
rect 345 972 379 1243
rect 245 73 279 342
rect 245 39 558 73
<< metal1 >>
rect 80 1260 108 1316
rect 248 412 276 972
rect 544 832 572 1316
rect 80 384 276 412
rect 348 804 572 832
rect 80 0 108 384
rect 348 342 376 804
rect 610 649 638 677
rect 544 0 572 56
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 595 0 1 630
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 333 0 1 309
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_2
timestamp 1661296025
transform 1 0 233 0 1 939
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_3
timestamp 1661296025
transform 1 0 529 0 1 23
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_4
timestamp 1661296025
transform 1 0 65 0 1 1227
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_14  sky130_sram_1r1w_24x128_8_contact_14_0
timestamp 1661296025
transform 1 0 599 0 1 622
box -26 -26 76 108
use sky130_sram_1r1w_24x128_8_nmos_m1_w2_880_sli_dli  sky130_sram_1r1w_24x128_8_nmos_m1_w2_880_sli_dli_0
timestamp 1661296025
transform 1 0 237 0 1 684
box -26 -26 176 602
use sky130_sram_1r1w_24x128_8_nmos_m1_w2_880_sli_dli  sky130_sram_1r1w_24x128_8_nmos_m1_w2_880_sli_dli_1
timestamp 1661296025
transform 1 0 237 0 1 54
box -26 -26 176 602
<< labels >>
rlabel poly s 312 41 312 41 4 sel
port 1 nsew
rlabel metal1 s 80 1260 108 1316 4 bl
port 2 nsew
rlabel metal1 s 544 1260 572 1316 4 br
port 3 nsew
rlabel metal1 s 80 0 108 56 4 bl_out
port 4 nsew
rlabel metal1 s 544 0 572 56 4 br_out
port 5 nsew
rlabel metal1 s 610 649 638 677 4 gnd
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 624 1316
<< end >>
