magic
tech sky130A
magscale 1 2
timestamp 1658896172
<< metal1 >>
rect 0 8220 1200 8400
rect 0 7940 1400 8220
rect 4 7786 159 7940
rect 461 7880 856 7940
rect 461 7800 1460 7880
rect 780 7780 1460 7800
rect 760 7600 1440 7700
rect 760 7420 1440 7520
rect 740 7240 1420 7340
rect 740 7060 1420 7160
rect 740 6960 1420 6980
rect 740 6880 1640 6960
rect 1400 6800 1640 6880
rect 740 6700 1640 6800
rect 1400 6640 1640 6700
rect 780 6500 1460 6600
rect 740 6320 1420 6420
rect 740 6140 1420 6240
rect 740 5960 1420 6060
rect 740 5780 1420 5880
rect 0 5380 1400 5720
rect 0 5000 1200 5380
<< metal2 >>
rect 1686 6900 2159 8192
rect 1685 6692 2159 6900
rect 2720 6760 2840 8060
rect -460 5580 -80 5660
rect -460 5500 1260 5580
rect -460 5400 900 5500
rect 1000 5400 1100 5500
rect 1200 5400 1260 5500
rect -460 5300 1260 5400
rect 1686 5399 2159 6692
rect 2240 6640 2840 6760
rect -460 5200 900 5300
rect 1000 5200 1100 5300
rect 1200 5200 1260 5300
rect -460 5140 1260 5200
<< via2 >>
rect 2320 7140 2380 7200
rect 2420 7140 2480 7200
rect 2520 7140 2580 7200
rect 2320 7040 2380 7100
rect 2420 7040 2480 7100
rect 2520 7040 2580 7100
rect 900 5400 1000 5500
rect 1100 5400 1200 5500
rect 900 5200 1000 5300
rect 1100 5200 1200 5300
<< metal3 >>
rect 2200 7380 2600 8100
rect 11690 7404 12002 7406
rect 2300 7200 2600 7220
rect 2300 7140 2320 7200
rect 2380 7140 2420 7200
rect 2480 7140 2520 7200
rect 2580 7140 2600 7200
rect 2300 7100 2600 7140
rect 2300 7040 2320 7100
rect 2380 7040 2420 7100
rect 2480 7040 2520 7100
rect 2580 7040 2600 7100
rect 2300 7020 2600 7040
rect 11690 7140 12230 7404
rect 2300 6540 2640 7020
rect 2300 6280 2600 6540
rect 2200 5580 2600 6280
rect 11690 5802 12002 7140
rect 840 5560 2600 5580
rect 840 5500 2220 5560
rect 840 5400 900 5500
rect 1000 5400 1100 5500
rect 1200 5400 2220 5500
rect 840 5300 2220 5400
rect 840 5200 900 5300
rect 1000 5200 1100 5300
rect 1200 5200 2220 5300
rect 840 5140 2220 5200
<< metal4 >>
rect -340 7960 2120 8380
rect 1600 7940 2120 7960
use captuner_complete_1  captuner_complete_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1658896172
transform -1 0 -1920 0 1 4580
box -3300 1000 -300 3400
use general_purpose_current_mirror  general_purpose_current_mirror_0
timestamp 1658895968
transform 1 0 12234 0 1 4918
box -80 -180 6020 2500
use nfet_3x_2  nfet_3x_2_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/LNA
timestamp 1658896172
transform 0 -1 2780 -1 0 8192
box 0 -60 1292 1380
use nfet_3x_2  nfet_3x_2_1
timestamp 1658896172
transform 0 -1 2780 -1 0 6692
box 0 -60 1292 1380
use simsq_balun_0p1n_24GHz  simsq_balun_0p1n_24GHz_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1658891120
transform 1 0 2000 0 1 2800
box -2000 -2800 10000 9400
use sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1649977179
transform 1 0 12200 0 1 7670
box 0 0 4498 4610
use sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top_1
timestamp 1649977179
transform 1 0 12194 0 1 -118
box 0 0 4498 4610
use sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top_2
timestamp 1649977179
transform 1 0 -4614 0 1 332
box 0 0 4498 4610
use sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top  sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top_3
timestamp 1649977179
transform 1 0 -5162 0 1 8546
box 0 0 4498 4610
<< end >>
