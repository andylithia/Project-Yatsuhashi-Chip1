magic
tech sky130B
magscale 1 2
timestamp 1662175719
<< error_p >>
rect -29 1040 29 1046
rect -29 1006 -17 1040
rect -29 1000 29 1006
rect -29 430 29 436
rect -29 396 -17 430
rect -29 390 29 396
rect -29 322 29 328
rect -29 288 -17 322
rect -29 282 29 288
rect -29 -288 29 -282
rect -29 -322 -17 -288
rect -29 -328 29 -322
rect -29 -396 29 -390
rect -29 -430 -17 -396
rect -29 -436 29 -430
rect -29 -1006 29 -1000
rect -29 -1040 -17 -1006
rect -29 -1046 29 -1040
<< pwell >>
rect -211 -1178 211 1178
<< nmos >>
rect -15 468 15 968
rect -15 -250 15 250
rect -15 -968 15 -468
<< ndiff >>
rect -73 956 -15 968
rect -73 480 -61 956
rect -27 480 -15 956
rect -73 468 -15 480
rect 15 956 73 968
rect 15 480 27 956
rect 61 480 73 956
rect 15 468 73 480
rect -73 238 -15 250
rect -73 -238 -61 238
rect -27 -238 -15 238
rect -73 -250 -15 -238
rect 15 238 73 250
rect 15 -238 27 238
rect 61 -238 73 238
rect 15 -250 73 -238
rect -73 -480 -15 -468
rect -73 -956 -61 -480
rect -27 -956 -15 -480
rect -73 -968 -15 -956
rect 15 -480 73 -468
rect 15 -956 27 -480
rect 61 -956 73 -480
rect 15 -968 73 -956
<< ndiffc >>
rect -61 480 -27 956
rect 27 480 61 956
rect -61 -238 -27 238
rect 27 -238 61 238
rect -61 -956 -27 -480
rect 27 -956 61 -480
<< psubdiff >>
rect -175 1108 -79 1142
rect 79 1108 175 1142
rect -175 1046 -141 1108
rect 141 1046 175 1108
rect -175 -1108 -141 -1046
rect 141 -1108 175 -1046
rect -175 -1142 -79 -1108
rect 79 -1142 175 -1108
<< psubdiffcont >>
rect -79 1108 79 1142
rect -175 -1046 -141 1046
rect 141 -1046 175 1046
rect -79 -1142 79 -1108
<< poly >>
rect -33 1040 33 1056
rect -33 1006 -17 1040
rect 17 1006 33 1040
rect -33 990 33 1006
rect -15 968 15 990
rect -15 446 15 468
rect -33 430 33 446
rect -33 396 -17 430
rect 17 396 33 430
rect -33 380 33 396
rect -33 322 33 338
rect -33 288 -17 322
rect 17 288 33 322
rect -33 272 33 288
rect -15 250 15 272
rect -15 -272 15 -250
rect -33 -288 33 -272
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect -33 -338 33 -322
rect -33 -396 33 -380
rect -33 -430 -17 -396
rect 17 -430 33 -396
rect -33 -446 33 -430
rect -15 -468 15 -446
rect -15 -990 15 -968
rect -33 -1006 33 -990
rect -33 -1040 -17 -1006
rect 17 -1040 33 -1006
rect -33 -1056 33 -1040
<< polycont >>
rect -17 1006 17 1040
rect -17 396 17 430
rect -17 288 17 322
rect -17 -322 17 -288
rect -17 -430 17 -396
rect -17 -1040 17 -1006
<< locali >>
rect -175 1108 -79 1142
rect 79 1108 175 1142
rect -175 1046 -141 1108
rect 141 1046 175 1108
rect -33 1006 -17 1040
rect 17 1006 33 1040
rect -61 956 -27 972
rect -61 464 -27 480
rect 27 956 61 972
rect 27 464 61 480
rect -33 396 -17 430
rect 17 396 33 430
rect -33 288 -17 322
rect 17 288 33 322
rect -61 238 -27 254
rect -61 -254 -27 -238
rect 27 238 61 254
rect 27 -254 61 -238
rect -33 -322 -17 -288
rect 17 -322 33 -288
rect -33 -430 -17 -396
rect 17 -430 33 -396
rect -61 -480 -27 -464
rect -61 -972 -27 -956
rect 27 -480 61 -464
rect 27 -972 61 -956
rect -33 -1040 -17 -1006
rect 17 -1040 33 -1006
rect -175 -1108 -141 -1046
rect 141 -1108 175 -1046
rect -175 -1142 -79 -1108
rect 79 -1142 175 -1108
<< viali >>
rect -17 1006 17 1040
rect -61 480 -27 956
rect 27 480 61 956
rect -17 396 17 430
rect -17 288 17 322
rect -61 -238 -27 238
rect 27 -238 61 238
rect -17 -322 17 -288
rect -17 -430 17 -396
rect -61 -956 -27 -480
rect 27 -956 61 -480
rect -17 -1040 17 -1006
<< metal1 >>
rect -29 1040 29 1046
rect -29 1006 -17 1040
rect 17 1006 29 1040
rect -29 1000 29 1006
rect -67 956 -21 968
rect -67 480 -61 956
rect -27 480 -21 956
rect -67 468 -21 480
rect 21 956 67 968
rect 21 480 27 956
rect 61 480 67 956
rect 21 468 67 480
rect -29 430 29 436
rect -29 396 -17 430
rect 17 396 29 430
rect -29 390 29 396
rect -29 322 29 328
rect -29 288 -17 322
rect 17 288 29 322
rect -29 282 29 288
rect -67 238 -21 250
rect -67 -238 -61 238
rect -27 -238 -21 238
rect -67 -250 -21 -238
rect 21 238 67 250
rect 21 -238 27 238
rect 61 -238 67 238
rect 21 -250 67 -238
rect -29 -288 29 -282
rect -29 -322 -17 -288
rect 17 -322 29 -288
rect -29 -328 29 -322
rect -29 -396 29 -390
rect -29 -430 -17 -396
rect 17 -430 29 -396
rect -29 -436 29 -430
rect -67 -480 -21 -468
rect -67 -956 -61 -480
rect -27 -956 -21 -480
rect -67 -968 -21 -956
rect 21 -480 67 -468
rect 21 -956 27 -480
rect 61 -956 67 -480
rect 21 -968 67 -956
rect -29 -1006 29 -1000
rect -29 -1040 -17 -1006
rect 17 -1040 29 -1006
rect -29 -1046 29 -1040
<< properties >>
string FIXED_BBOX -158 -1125 158 1125
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.150 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
