magic
tech sky130B
timestamp 1658891120
<< metal1 >>
rect -1000 4600 4800 4700
rect -1000 4400 -800 4600
rect -600 4400 -500 4600
rect -300 4400 -200 4600
rect 0 4400 100 4600
rect 300 4400 400 4600
rect 600 4400 700 4600
rect 900 4400 1000 4600
rect 1200 4400 1300 4600
rect 1500 4400 1600 4600
rect 1800 4400 1900 4600
rect 2100 4400 2200 4600
rect 2400 4400 2500 4600
rect 2700 4400 2800 4600
rect 3000 4400 3100 4600
rect 3300 4400 3400 4600
rect 3600 4400 3700 4600
rect 3900 4400 4000 4600
rect 4200 4400 4300 4600
rect 4500 4400 4800 4600
rect -1000 4300 4800 4400
rect -1000 4100 -900 4300
rect -700 4200 4500 4300
rect -700 4100 -500 4200
rect -1000 4000 -500 4100
rect -400 4000 -200 4200
rect -1000 3800 -900 4000
rect -700 3900 -600 4000
rect -300 3900 -200 4000
rect -700 3800 -400 3900
rect -1000 3700 -300 3800
rect -100 3700 100 4200
rect -1000 3500 -900 3700
rect -700 3600 -600 3700
rect 0 3600 100 3700
rect -700 3500 -100 3600
rect -1000 3400 0 3500
rect 200 3400 400 4200
rect -1000 3200 -900 3400
rect -700 3300 -600 3400
rect 300 3300 400 3400
rect -700 3200 200 3300
rect -1000 3100 300 3200
rect 500 3100 700 4200
rect -1000 2900 -900 3100
rect -700 3000 -600 3100
rect 600 3000 700 3100
rect -700 2900 500 3000
rect -1000 2800 600 2900
rect 800 2800 1000 4200
rect 900 2700 1000 2800
rect 1100 2500 1300 4200
rect 1200 2400 1300 2500
rect 1400 2200 1600 4200
rect 1500 2100 1600 2200
rect 1700 1900 1800 4200
rect 1900 2200 2100 4200
rect 2200 2500 2400 4200
rect 2500 2800 2700 4200
rect 2800 3100 3000 4200
rect 3100 3400 3300 4200
rect 3400 3700 3600 4200
rect 3700 4000 3900 4200
rect 4000 4100 4500 4200
rect 4700 4100 4800 4300
rect 4000 4000 4800 4100
rect 3700 3900 3800 4000
rect 4300 3900 4500 4000
rect 3900 3800 4500 3900
rect 4700 3800 4800 4000
rect 3800 3700 4800 3800
rect 3400 3600 3500 3700
rect 4300 3600 4500 3700
rect 3600 3500 4500 3600
rect 4700 3500 4800 3700
rect 3500 3400 4800 3500
rect 3100 3300 3200 3400
rect 4300 3300 4500 3400
rect 3300 3200 4500 3300
rect 4700 3200 4800 3400
rect 3200 3100 4800 3200
rect 2800 3000 2900 3100
rect 4300 3000 4500 3100
rect 3000 2900 4500 3000
rect 4700 2900 4800 3100
rect 2900 2800 4800 2900
rect 2500 2700 2600 2800
rect 4300 2700 4500 2800
rect 2700 2600 4500 2700
rect 4700 2600 4800 2800
rect 2600 2500 4800 2600
rect 2200 2400 2300 2500
rect 4300 2400 4500 2500
rect 2400 2300 4500 2400
rect 4700 2300 4800 2500
rect 2300 2200 4800 2300
rect 1900 2100 2000 2200
rect 4300 2100 4500 2200
rect 2100 2000 4500 2100
rect 4700 2000 4800 2200
rect 2000 1900 4800 2000
rect 4300 1800 4500 1900
rect 2000 1700 4500 1800
rect 4700 1700 4800 1900
rect 1900 1600 4800 1700
rect 2000 1500 4500 1600
rect 4300 1400 4500 1500
rect 4700 1400 4800 1600
rect 1500 1100 1600 1200
rect -1000 1000 1200 1100
rect -1000 800 -900 1000
rect -700 900 1100 1000
rect -700 800 -600 900
rect 1200 800 1300 900
rect -1000 700 900 800
rect -1000 500 -900 700
rect -700 600 800 700
rect -700 500 -600 600
rect 900 500 1000 600
rect -1000 400 600 500
rect -1000 200 -900 400
rect -700 300 500 400
rect -700 200 -600 300
rect 600 200 700 300
rect -1000 100 300 200
rect -1000 -100 -900 100
rect -700 0 200 100
rect -700 -100 -600 0
rect 300 -100 400 0
rect -1000 -200 0 -100
rect -1000 -400 -900 -200
rect -700 -300 -100 -200
rect -700 -400 -600 -300
rect 0 -400 100 -300
rect -1000 -500 -300 -400
rect -1000 -700 -900 -500
rect -700 -600 -400 -500
rect -700 -700 -600 -600
rect -300 -700 -200 -600
rect -1000 -800 -500 -700
rect -1000 -1000 -900 -800
rect -700 -900 -500 -800
rect -400 -900 -200 -700
rect -100 -900 100 -400
rect 200 -900 400 -100
rect 500 -900 700 200
rect 800 -900 1000 500
rect 1100 -900 1300 800
rect 1400 -900 1600 1100
rect 1700 -900 1800 1400
rect 2000 1300 4800 1400
rect 2100 1200 4500 1300
rect 1900 1100 2000 1200
rect 4300 1100 4500 1200
rect 4700 1100 4800 1300
rect 1900 -900 2100 1100
rect 2300 1000 4800 1100
rect 2400 900 4500 1000
rect 2200 800 2300 900
rect 4300 800 4500 900
rect 4700 800 4800 1000
rect 2200 -900 2400 800
rect 2600 700 4800 800
rect 2700 600 4500 700
rect 2500 500 2600 600
rect 4300 500 4500 600
rect 4700 500 4800 700
rect 2500 -900 2700 500
rect 2900 400 4800 500
rect 3000 300 4500 400
rect 2800 200 2900 300
rect 4300 200 4500 300
rect 4700 200 4800 400
rect 2800 -900 3000 200
rect 3200 100 4800 200
rect 3300 0 4500 100
rect 3100 -100 3200 0
rect 4300 -100 4500 0
rect 4700 -100 4800 100
rect 3100 -900 3300 -100
rect 3500 -200 4800 -100
rect 3600 -300 4500 -200
rect 3400 -400 3500 -300
rect 4300 -400 4500 -300
rect 4700 -400 4800 -200
rect 3400 -900 3600 -400
rect 3800 -500 4800 -400
rect 3900 -600 4500 -500
rect 3700 -700 3800 -600
rect 4300 -700 4500 -600
rect 4700 -700 4800 -500
rect 3700 -900 3900 -700
rect 4000 -800 4800 -700
rect 4000 -900 4500 -800
rect -700 -1000 4500 -900
rect 4700 -1000 4800 -800
rect -1000 -1100 4800 -1000
rect -1000 -1300 -900 -1100
rect -700 -1300 -500 -1100
rect -300 -1300 -200 -1100
rect 0 -1300 100 -1100
rect 300 -1300 400 -1100
rect 600 -1300 700 -1100
rect 900 -1300 1000 -1100
rect 1200 -1300 1300 -1100
rect 1500 -1300 1600 -1100
rect 1800 -1300 1900 -1100
rect 2100 -1300 2200 -1100
rect 2400 -1300 2500 -1100
rect 2700 -1300 2800 -1100
rect 3000 -1300 3100 -1100
rect 3300 -1300 3400 -1100
rect 3600 -1300 3700 -1100
rect 3900 -1300 4000 -1100
rect 4200 -1300 4300 -1100
rect 4500 -1300 4800 -1100
rect -1000 -1400 4800 -1300
<< via1 >>
rect -800 4400 -600 4600
rect -500 4400 -300 4600
rect -200 4400 0 4600
rect 100 4400 300 4600
rect 400 4400 600 4600
rect 700 4400 900 4600
rect 1000 4400 1200 4600
rect 1300 4400 1500 4600
rect 1600 4400 1800 4600
rect 1900 4400 2100 4600
rect 2200 4400 2400 4600
rect 2500 4400 2700 4600
rect 2800 4400 3000 4600
rect 3100 4400 3300 4600
rect 3400 4400 3600 4600
rect 3700 4400 3900 4600
rect 4000 4400 4200 4600
rect 4300 4400 4500 4600
rect -900 4100 -700 4300
rect -900 3800 -700 4000
rect -900 3500 -700 3700
rect -900 3200 -700 3400
rect -900 2900 -700 3100
rect 4500 4100 4700 4300
rect 4500 3800 4700 4000
rect 4500 3500 4700 3700
rect 4500 3200 4700 3400
rect 4500 2900 4700 3100
rect 4500 2600 4700 2800
rect 4500 2300 4700 2500
rect 4500 2000 4700 2200
rect 4500 1700 4700 1900
rect 4500 1400 4700 1600
rect -900 800 -700 1000
rect -900 500 -700 700
rect -900 200 -700 400
rect -900 -100 -700 100
rect -900 -400 -700 -200
rect -900 -700 -700 -500
rect -900 -1000 -700 -800
rect 4500 1100 4700 1300
rect 4500 800 4700 1000
rect 4500 500 4700 700
rect 4500 200 4700 400
rect 4500 -100 4700 100
rect 4500 -400 4700 -200
rect 4500 -700 4700 -500
rect 4500 -1000 4700 -800
rect -900 -1300 -700 -1100
rect -500 -1300 -300 -1100
rect -200 -1300 0 -1100
rect 100 -1300 300 -1100
rect 400 -1300 600 -1100
rect 700 -1300 900 -1100
rect 1000 -1300 1200 -1100
rect 1300 -1300 1500 -1100
rect 1600 -1300 1800 -1100
rect 1900 -1300 2100 -1100
rect 2200 -1300 2400 -1100
rect 2500 -1300 2700 -1100
rect 2800 -1300 3000 -1100
rect 3100 -1300 3300 -1100
rect 3400 -1300 3600 -1100
rect 3700 -1300 3900 -1100
rect 4000 -1300 4200 -1100
rect 4300 -1300 4500 -1100
<< metal2 >>
rect -1000 4600 4800 4700
rect -1000 4400 -800 4600
rect -600 4400 -500 4600
rect -300 4400 -200 4600
rect 0 4400 100 4600
rect 300 4400 400 4600
rect 600 4400 700 4600
rect 900 4400 1000 4600
rect 1200 4400 1300 4600
rect 1500 4400 1600 4600
rect 1800 4400 1900 4600
rect 2100 4400 2200 4600
rect 2400 4400 2500 4600
rect 2700 4400 2800 4600
rect 3000 4400 3100 4600
rect 3300 4400 3400 4600
rect 3600 4400 3700 4600
rect 3900 4400 4000 4600
rect 4200 4400 4300 4600
rect 4500 4400 4800 4600
rect -1000 4300 4800 4400
rect -1000 4100 -900 4300
rect -700 4100 -500 4300
rect -1000 4000 -500 4100
rect -400 4000 -200 4300
rect -1000 3800 -900 4000
rect -700 3900 -600 4000
rect -300 3900 -200 4000
rect -700 3800 -400 3900
rect -1000 3700 -300 3800
rect -100 3700 100 4300
rect -1000 3500 -900 3700
rect -700 3600 -600 3700
rect 0 3600 100 3700
rect -700 3500 -100 3600
rect -1000 3400 0 3500
rect 200 3400 400 4300
rect -1000 3200 -900 3400
rect -700 3300 -600 3400
rect 300 3300 400 3400
rect -700 3200 200 3300
rect -1000 3100 300 3200
rect 500 3100 700 4300
rect -1000 2900 -900 3100
rect -700 3000 -600 3100
rect 600 3000 700 3100
rect -700 2900 500 3000
rect -1000 2800 600 2900
rect 800 2800 1000 4300
rect 900 2700 1000 2800
rect 1100 2500 1300 4300
rect 1200 2400 1300 2500
rect 1400 2200 1600 4300
rect 1500 2100 1600 2200
rect 1700 1900 1800 4300
rect 1900 2200 2100 4300
rect 2200 2500 2400 4300
rect 2500 2800 2700 4300
rect 2800 3100 3000 4300
rect 3100 3400 3300 4300
rect 3400 3700 3600 4300
rect 3700 4000 3900 4300
rect 4000 4100 4500 4300
rect 4700 4100 4800 4300
rect 4000 4000 4800 4100
rect 3700 3900 3800 4000
rect 4400 3900 4500 4000
rect 3900 3800 4500 3900
rect 4700 3800 4800 4000
rect 3800 3700 4800 3800
rect 3400 3600 3500 3700
rect 4400 3600 4500 3700
rect 3600 3500 4500 3600
rect 4700 3500 4800 3700
rect 3500 3400 4800 3500
rect 3100 3300 3200 3400
rect 4400 3300 4500 3400
rect 3300 3200 4500 3300
rect 4700 3200 4800 3400
rect 3200 3100 4800 3200
rect 2800 3000 2900 3100
rect 4400 3000 4500 3100
rect 3000 2900 4500 3000
rect 4700 2900 4800 3100
rect 2900 2800 4800 2900
rect 2500 2700 2600 2800
rect 4400 2700 4500 2800
rect 2700 2600 4500 2700
rect 4700 2600 4800 2800
rect 2600 2500 4800 2600
rect 2200 2400 2300 2500
rect 4400 2400 4500 2500
rect 2400 2300 4500 2400
rect 4700 2300 4800 2500
rect 2300 2200 4800 2300
rect 1900 2100 2000 2200
rect 4400 2100 4500 2200
rect 2100 2000 4500 2100
rect 4700 2000 4800 2200
rect 2000 1900 4800 2000
rect 4400 1800 4500 1900
rect 2000 1700 4500 1800
rect 4700 1700 4800 1900
rect 1900 1600 4800 1700
rect 2000 1500 4500 1600
rect 4400 1400 4500 1500
rect 4700 1400 4800 1600
rect 1500 1100 1600 1200
rect -1000 1000 1200 1100
rect -1000 800 -900 1000
rect -700 900 1100 1000
rect -700 800 -600 900
rect 1200 800 1300 900
rect -1000 700 900 800
rect -1000 500 -900 700
rect -700 600 800 700
rect -700 500 -600 600
rect 900 500 1000 600
rect -1000 400 600 500
rect -1000 200 -900 400
rect -700 300 500 400
rect -700 200 -600 300
rect 600 200 700 300
rect -1000 100 300 200
rect -1000 -100 -900 100
rect -700 0 200 100
rect -700 -100 -600 0
rect 300 -100 400 0
rect -1000 -200 0 -100
rect -1000 -400 -900 -200
rect -700 -300 -100 -200
rect -700 -400 -600 -300
rect 0 -400 100 -300
rect -1000 -500 -300 -400
rect -1000 -700 -900 -500
rect -700 -600 -400 -500
rect -700 -700 -600 -600
rect -300 -700 -200 -600
rect -1000 -800 -500 -700
rect -1000 -1000 -900 -800
rect -700 -1000 -500 -800
rect -400 -1000 -200 -700
rect -100 -1000 100 -400
rect 200 -1000 400 -100
rect 500 -1000 700 200
rect 800 -1000 1000 500
rect 1100 -1000 1300 800
rect 1400 -1000 1600 1100
rect 1700 -1000 1800 1400
rect 2000 1300 4800 1400
rect 2100 1200 4500 1300
rect 1900 1100 2000 1200
rect 4400 1100 4500 1200
rect 4700 1100 4800 1300
rect 1900 -1000 2100 1100
rect 2300 1000 4800 1100
rect 2400 900 4500 1000
rect 2200 800 2300 900
rect 4400 800 4500 900
rect 4700 800 4800 1000
rect 2200 -1000 2400 800
rect 2600 700 4800 800
rect 2700 600 4500 700
rect 2500 500 2600 600
rect 4400 500 4500 600
rect 4700 500 4800 700
rect 2500 -1000 2700 500
rect 2900 400 4800 500
rect 3000 300 4500 400
rect 2800 200 2900 300
rect 4400 200 4500 300
rect 4700 200 4800 400
rect 2800 -1000 3000 200
rect 3200 100 4800 200
rect 3300 0 4500 100
rect 3100 -100 3200 0
rect 4400 -100 4500 0
rect 4700 -100 4800 100
rect 3100 -1000 3300 -100
rect 3500 -200 4800 -100
rect 3600 -300 4500 -200
rect 3400 -400 3500 -300
rect 4400 -400 4500 -300
rect 4700 -400 4800 -200
rect 3400 -1000 3600 -400
rect 3800 -500 4800 -400
rect 3900 -600 4500 -500
rect 3700 -700 3800 -600
rect 4400 -700 4500 -600
rect 4700 -700 4800 -500
rect 3700 -1000 3900 -700
rect 4000 -800 4800 -700
rect 4000 -1000 4500 -800
rect 4700 -1000 4800 -800
rect -1000 -1100 4800 -1000
rect -1000 -1300 -900 -1100
rect -700 -1300 -500 -1100
rect -300 -1300 -200 -1100
rect 0 -1300 100 -1100
rect 300 -1300 400 -1100
rect 600 -1300 700 -1100
rect 900 -1300 1000 -1100
rect 1200 -1300 1300 -1100
rect 1500 -1300 1600 -1100
rect 1800 -1300 1900 -1100
rect 2100 -1300 2200 -1100
rect 2400 -1300 2500 -1100
rect 2700 -1300 2800 -1100
rect 3000 -1300 3100 -1100
rect 3300 -1300 3400 -1100
rect 3600 -1300 3700 -1100
rect 3900 -1300 4000 -1100
rect 4200 -1300 4300 -1100
rect 4500 -1300 4800 -1100
rect -1000 -1400 4800 -1300
<< via2 >>
rect -800 4400 -600 4600
rect -500 4400 -300 4600
rect -200 4400 0 4600
rect 100 4400 300 4600
rect 400 4400 600 4600
rect 700 4400 900 4600
rect 1000 4400 1200 4600
rect 1300 4400 1500 4600
rect 1600 4400 1800 4600
rect 1900 4400 2100 4600
rect 2200 4400 2400 4600
rect 2500 4400 2700 4600
rect 2800 4400 3000 4600
rect 3100 4400 3300 4600
rect 3400 4400 3600 4600
rect 3700 4400 3900 4600
rect 4000 4400 4200 4600
rect 4300 4400 4500 4600
rect -900 4100 -700 4300
rect -900 3800 -700 4000
rect -900 3500 -700 3700
rect -900 3200 -700 3400
rect -900 2900 -700 3100
rect 4500 4100 4700 4300
rect 4500 3800 4700 4000
rect 4500 3500 4700 3700
rect 4500 3200 4700 3400
rect 4500 2900 4700 3100
rect 4500 2600 4700 2800
rect 4500 2300 4700 2500
rect -900 800 -700 1000
rect -900 500 -700 700
rect -900 200 -700 400
rect -900 -100 -700 100
rect -900 -400 -700 -200
rect -900 -700 -700 -500
rect -900 -1000 -700 -800
rect 4500 800 4700 1000
rect 4500 500 4700 700
rect 4500 200 4700 400
rect 4500 -100 4700 100
rect 4500 -400 4700 -200
rect 4500 -700 4700 -500
rect 4500 -1000 4700 -800
rect -900 -1300 -700 -1100
rect -500 -1300 -300 -1100
rect -200 -1300 0 -1100
rect 100 -1300 300 -1100
rect 400 -1300 600 -1100
rect 700 -1300 900 -1100
rect 1000 -1300 1200 -1100
rect 1300 -1300 1500 -1100
rect 1600 -1300 1800 -1100
rect 1900 -1300 2100 -1100
rect 2200 -1300 2400 -1100
rect 2500 -1300 2700 -1100
rect 2800 -1300 3000 -1100
rect 3100 -1300 3300 -1100
rect 3400 -1300 3600 -1100
rect 3700 -1300 3900 -1100
rect 4000 -1300 4200 -1100
rect 4300 -1300 4500 -1100
<< metal3 >>
rect -1000 4600 4800 4700
rect -1000 4400 -800 4600
rect -600 4400 -500 4600
rect -300 4400 -200 4600
rect 0 4400 100 4600
rect 300 4400 400 4600
rect 600 4400 700 4600
rect 900 4400 1000 4600
rect 1200 4400 1300 4600
rect 1500 4400 1600 4600
rect 1800 4400 1900 4600
rect 2100 4400 2200 4600
rect 2400 4400 2500 4600
rect 2700 4400 2800 4600
rect 3000 4400 3100 4600
rect 3300 4400 3400 4600
rect 3600 4400 3700 4600
rect 3900 4400 4000 4600
rect 4200 4400 4300 4600
rect 4500 4400 4800 4600
rect -1000 4300 4800 4400
rect -1000 4100 -900 4300
rect -700 4100 -600 4300
rect -1000 4000 -600 4100
rect -1000 3800 -900 4000
rect -700 3800 -600 4000
rect -1000 3700 -600 3800
rect -1000 3500 -900 3700
rect -700 3500 -600 3700
rect -1000 3400 -600 3500
rect -1000 3200 -900 3400
rect -700 3200 -600 3400
rect -1000 3100 -600 3200
rect -1000 2900 -900 3100
rect -700 2900 -600 3100
rect -1000 2800 -600 2900
rect 4400 4100 4500 4300
rect 4700 4100 4800 4300
rect 4400 4000 4800 4100
rect 4400 3800 4500 4000
rect 4700 3800 4800 4000
rect 4400 3700 4800 3800
rect 4400 3500 4500 3700
rect 4700 3500 4800 3700
rect 4400 3400 4800 3500
rect 4400 3200 4500 3400
rect 4700 3200 4800 3400
rect 4400 3100 4800 3200
rect 4400 2900 4500 3100
rect 4700 2900 4800 3100
rect 4400 2800 4800 2900
rect -200 2600 300 2650
rect -200 2450 -150 2600
rect 0 2450 50 2600
rect 200 2450 300 2600
rect -200 2400 300 2450
rect 4400 2600 4500 2800
rect 4700 2600 4800 2800
rect 4400 2500 4800 2600
rect -150 2350 250 2400
rect 4400 2300 4500 2500
rect 4700 2300 4800 2500
rect 4400 2000 4800 2300
rect 1500 1850 2000 1900
rect 1500 1450 1550 1850
rect 1700 1450 1750 1850
rect 1900 1800 2000 1850
rect 1900 1500 5000 1800
rect 1900 1450 2000 1500
rect -150 1400 250 1450
rect 1500 1400 2000 1450
rect -200 1350 300 1400
rect -200 1200 -150 1350
rect 0 1200 50 1350
rect 200 1200 300 1350
rect -200 1150 300 1200
rect -1000 1000 -600 1100
rect -1000 800 -900 1000
rect -700 800 -600 1000
rect -1000 700 -600 800
rect -1000 500 -900 700
rect -700 500 -600 700
rect -1000 400 -600 500
rect -1000 200 -900 400
rect -700 200 -600 400
rect -1000 100 -600 200
rect -1000 -100 -900 100
rect -700 -100 -600 100
rect -1000 -200 -600 -100
rect -1000 -400 -900 -200
rect -700 -400 -600 -200
rect -1000 -500 -600 -400
rect -1000 -700 -900 -500
rect -700 -700 -600 -500
rect -1000 -800 -600 -700
rect -1000 -1000 -900 -800
rect -700 -1000 -600 -800
rect 4400 1000 4800 1300
rect 4400 800 4500 1000
rect 4700 800 4800 1000
rect 4400 700 4800 800
rect 4400 500 4500 700
rect 4700 500 4800 700
rect 4400 400 4800 500
rect 4400 200 4500 400
rect 4700 200 4800 400
rect 4400 100 4800 200
rect 4400 -100 4500 100
rect 4700 -100 4800 100
rect 4400 -200 4800 -100
rect 4400 -400 4500 -200
rect 4700 -400 4800 -200
rect 4400 -500 4800 -400
rect 4400 -700 4500 -500
rect 4700 -700 4800 -500
rect 4400 -800 4800 -700
rect 4400 -1000 4500 -800
rect 4700 -1000 4800 -800
rect -1000 -1100 4800 -1000
rect -1000 -1300 -900 -1100
rect -700 -1300 -500 -1100
rect -300 -1300 -200 -1100
rect 0 -1300 100 -1100
rect 300 -1300 400 -1100
rect 600 -1300 700 -1100
rect 900 -1300 1000 -1100
rect 1200 -1300 1300 -1100
rect 1500 -1300 1600 -1100
rect 1800 -1300 1900 -1100
rect 2100 -1300 2200 -1100
rect 2400 -1300 2500 -1100
rect 2700 -1300 2800 -1100
rect 3000 -1300 3100 -1100
rect 3300 -1300 3400 -1100
rect 3600 -1300 3700 -1100
rect 3900 -1300 4000 -1100
rect 4200 -1300 4300 -1100
rect 4500 -1300 4800 -1100
rect -1000 -1400 4800 -1300
<< via3 >>
rect -150 2450 0 2600
rect 50 2450 200 2600
rect 1550 1450 1700 1850
rect 1750 1450 1900 1850
rect -150 1200 0 1350
rect 50 1200 200 1350
<< metal4 >>
rect -200 2800 300 2850
rect -200 2650 -100 2800
rect 50 2650 100 2800
rect 250 2650 300 2800
rect -200 2600 300 2650
rect -200 2450 -150 2600
rect 0 2450 50 2600
rect 200 2450 300 2600
rect 3300 2800 3800 2850
rect 3300 2650 3400 2800
rect 3550 2650 3600 2800
rect 3750 2650 3800 2800
rect 3300 2600 3800 2650
rect 3300 2500 3350 2600
rect -200 2400 300 2450
rect 3250 2450 3350 2500
rect 3500 2450 3550 2600
rect 3700 2450 3800 2600
rect 3250 2400 3800 2450
rect 3200 2300 3750 2400
rect 3150 2200 3700 2300
rect 3100 2100 3650 2200
rect 3050 2000 3600 2100
rect 3000 1900 3550 2000
rect 600 1800 1100 1900
rect 1450 1850 1950 1900
rect 1450 1800 1550 1850
rect 600 1500 650 1800
rect 800 1500 900 1800
rect 1050 1500 1550 1800
rect 600 1400 1100 1500
rect 1450 1450 1550 1500
rect 1700 1450 1750 1850
rect 1900 1450 1950 1850
rect 2950 1800 3500 1900
rect 2900 1700 3450 1800
rect 2850 1600 3400 1700
rect 2800 1500 3350 1600
rect 1450 1400 1950 1450
rect 2750 1400 3300 1500
rect -200 1350 300 1400
rect -200 1200 -150 1350
rect 0 1200 50 1350
rect 200 1200 300 1350
rect 2700 1300 3250 1400
rect 2650 1200 3200 1300
rect -200 1150 300 1200
rect -200 1000 -100 1150
rect 50 1000 100 1150
rect 250 1000 300 1150
rect 2600 1100 3150 1200
rect 2550 1000 3100 1100
rect -200 950 300 1000
rect 2500 900 3050 1000
rect 2500 850 3000 900
rect 2500 700 2550 850
rect 2700 700 2750 850
rect 2900 700 3000 850
rect 2500 650 3000 700
rect 2500 500 2600 650
rect 2750 500 2800 650
rect 2950 500 3000 650
rect 2500 450 3000 500
<< via4 >>
rect -100 2650 50 2800
rect 100 2650 250 2800
rect -150 2450 0 2600
rect 50 2450 200 2600
rect 3400 2650 3550 2800
rect 3600 2650 3750 2800
rect 3350 2450 3500 2600
rect 3550 2450 3700 2600
rect 650 1500 800 1800
rect 900 1500 1050 1800
rect -150 1200 0 1350
rect 50 1200 200 1350
rect -100 1000 50 1150
rect 100 1000 250 1150
rect 2550 700 2700 850
rect 2750 700 2900 850
rect 2600 500 2750 650
rect 2800 500 2950 650
<< metal5 >>
rect -200 3400 3800 3900
rect -200 2800 300 3400
rect -200 2650 -100 2800
rect 50 2650 100 2800
rect 250 2650 300 2800
rect -200 2600 300 2650
rect -200 2450 -150 2600
rect 0 2450 50 2600
rect 200 2450 300 2600
rect -200 2400 300 2450
rect 600 2600 3000 3100
rect 600 1800 1100 2600
rect 2500 2500 3000 2600
rect 3300 2800 3800 3400
rect 3300 2650 3400 2800
rect 3550 2650 3600 2800
rect 3750 2650 3800 2800
rect 3300 2600 3800 2650
rect 2500 2400 3050 2500
rect 3300 2450 3350 2600
rect 3500 2450 3550 2600
rect 3700 2450 3800 2600
rect 3300 2400 3800 2450
rect 2550 2300 3100 2400
rect 2600 2200 3150 2300
rect 2650 2100 3200 2200
rect 2700 2000 3250 2100
rect 2750 1900 3300 2000
rect 2800 1800 3350 1900
rect 600 1500 650 1800
rect 800 1500 900 1800
rect 1050 1500 1100 1800
rect 2850 1700 3400 1800
rect 2900 1600 3450 1700
rect 2950 1500 3500 1600
rect -200 1350 300 1400
rect -200 1200 -150 1350
rect 0 1200 50 1350
rect 200 1200 300 1350
rect -200 1150 300 1200
rect -200 1000 -100 1150
rect 50 1000 100 1150
rect 250 1000 300 1150
rect -200 -100 300 1000
rect 600 700 1100 1500
rect 3000 1400 3550 1500
rect 3050 1300 3600 1400
rect 3100 1200 3650 1300
rect 3150 1100 3700 1200
rect 3200 1000 3800 1100
rect 3250 900 3800 1000
rect 2500 850 3000 900
rect 2500 700 2550 850
rect 2700 700 2750 850
rect 2900 700 3000 850
rect 600 650 3000 700
rect 600 500 2600 650
rect 2750 500 2800 650
rect 2950 500 3000 650
rect 600 200 3000 500
rect 3300 -100 3800 900
rect -200 -600 3800 -100
<< labels >>
rlabel metal3 -150 2350 250 2400 1 A
rlabel metal3 -150 1400 250 1450 1 B
rlabel metal3 4850 1500 5000 1800 1 C
rlabel metal3 4500 4350 4800 4700 1 G
<< end >>
