magic
tech sky130A
timestamp 1663980874
<< metal3 >>
rect 200 5200 2800 6200
rect 5600 5200 8200 6200
rect 8300 200 10900 1200
<< metal4 >>
rect 200 5200 900 8400
rect 400 -500 1100 4700
rect 1300 -1700 2000 2700
rect 2100 300 2800 9900
rect 3000 400 3700 8400
rect 4700 5200 5400 9900
rect 5600 5200 6300 8400
rect 3900 -1700 4600 4700
rect 4800 -500 5500 2700
rect 5800 -500 6500 4700
rect 6700 -1700 7400 2700
rect 7500 200 8200 9800
rect 8300 200 9000 8400
rect 10100 5200 10800 9800
rect 9200 -500 9900 2700
rect 10100 -1700 10800 4700
<< metal5 >>
rect 100 8400 1800 10200
rect 9100 9900 10800 10200
rect 2100 9200 10800 9900
rect 100 7700 9000 8400
rect -600 -500 9900 200
rect -600 -6400 1100 -500
rect 10800 -1000 12500 100
rect 1300 -1700 12500 -1000
rect 10800 -6500 12500 -1700
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_0
timestamp 1663721312
transform 1 0 200 0 1 -200
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_1
timestamp 1663721312
transform 1 0 2900 0 1 -200
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_2
timestamp 1663721312
transform 1 0 5600 0 1 -200
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_3
timestamp 1663721312
transform 1 0 8300 0 1 -200
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_4
timestamp 1663721312
transform 1 0 200 0 1 3300
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_5
timestamp 1663721312
transform 1 0 2900 0 1 3300
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_6
timestamp 1663721312
transform 1 0 5600 0 1 3300
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_7
timestamp 1663721312
transform 1 0 8300 0 1 3300
box 0 0 2569 3258
use octa_thick_1p5n_classe_flat  octa_thick_1p5n_classe_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1663980778
transform 1 0 55600 0 1 38400
box -33000 -30000 7750 10000
<< end >>
