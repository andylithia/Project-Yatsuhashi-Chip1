magic
tech sky130B
magscale 1 2
timestamp 1660708745
<< pwell >>
rect -5320 19520 -5280 19530
<< locali >>
rect -5330 20650 -4220 20660
rect -5330 20640 -5240 20650
rect -5330 19530 -5320 20640
rect -5286 20610 -5240 20640
rect -4310 20640 -4220 20650
rect -4310 20610 -4260 20640
rect -5286 20600 -4260 20610
rect -5286 19570 -5280 20600
rect -4270 19570 -4260 20600
rect -5286 19560 -4260 19570
rect -5286 19530 -5240 19560
rect -5330 19520 -5240 19530
rect -4310 19530 -4260 19560
rect -4226 19530 -4220 20640
rect -4310 19520 -4220 19530
rect -5330 19510 -4220 19520
<< viali >>
rect -5320 19530 -5286 20640
rect -5240 20610 -4310 20650
rect -5240 19520 -4310 19560
rect -4260 19530 -4226 20640
<< metal1 >>
rect -4226 20660 -4050 20700
rect -5330 20650 -4050 20660
rect -5330 20640 -5240 20650
rect -5330 19530 -5320 20640
rect -5286 20610 -5240 20640
rect -4310 20640 -4050 20650
rect -4310 20610 -4260 20640
rect -5286 20600 -4260 20610
rect -5286 20510 -5280 20600
rect -5090 20550 -5000 20560
rect -5286 20430 -5120 20510
rect -5090 20440 -5080 20550
rect -5010 20440 -5000 20550
rect -4550 20550 -4460 20560
rect -5090 20430 -5000 20440
rect -4971 20437 -4797 20509
rect -4755 20437 -4581 20509
rect -4550 20440 -4540 20550
rect -4470 20440 -4460 20550
rect -4270 20510 -4260 20600
rect -4550 20430 -4460 20440
rect -4430 20430 -4260 20510
rect -5286 19740 -5280 20430
rect -5286 19660 -5120 19740
rect -5079 19663 -4905 19735
rect -5286 19570 -5280 19660
rect -4870 19570 -4680 19750
rect -4270 19740 -4260 20430
rect -4650 19730 -4470 19740
rect -4650 19630 -4640 19730
rect -4480 19630 -4470 19730
rect -4440 19660 -4260 19740
rect -4270 19570 -4260 19660
rect -5286 19560 -4260 19570
rect -5286 19530 -5240 19560
rect -5330 19520 -5240 19530
rect -4310 19530 -4260 19560
rect -4226 20600 -4050 20640
rect -4226 20200 -3950 20600
rect -4226 20100 -4050 20200
rect -4226 19700 -3950 20100
rect -4226 19600 -4050 19700
rect -3950 19600 550 19700
rect -4226 19530 -4220 19600
rect -4310 19520 -4220 19530
rect -5330 19510 -4220 19520
rect -3950 19580 -3830 19600
rect -3570 19580 -3330 19600
rect -3070 19580 -2830 19600
rect -2570 19580 -2330 19600
rect -2070 19580 -1830 19600
rect -1570 19580 -1330 19600
rect -1070 19580 -830 19600
rect -570 19580 -330 19600
rect -70 19580 170 19600
rect 430 19580 550 19600
rect -3950 19320 -3850 19580
rect -3550 19320 -3350 19580
rect -3050 19320 -2850 19580
rect -2550 19320 -2350 19580
rect -2050 19320 -1850 19580
rect -1550 19320 -1350 19580
rect -1050 19320 -850 19580
rect -550 19320 -350 19580
rect -50 19320 150 19580
rect 450 19320 550 19580
rect -3950 19300 -3830 19320
rect -3570 19300 -3330 19320
rect -3070 19300 -2830 19320
rect -2570 19300 -2330 19320
rect -2070 19300 -1830 19320
rect -1570 19300 -1330 19320
rect -1070 19300 -830 19320
rect -570 19300 -330 19320
rect -70 19300 170 19320
rect 430 19300 550 19320
rect 3750 19600 5550 19700
rect 3750 19580 4170 19600
rect 4430 19580 4670 19600
rect 4930 19580 5170 19600
rect 5430 19580 5550 19600
rect 3750 19320 4150 19580
rect 4450 19320 4650 19580
rect 4950 19320 5150 19580
rect 5450 19320 5550 19580
rect 3750 19300 4170 19320
rect 4430 19300 4670 19320
rect 4930 19300 5170 19320
rect 5430 19300 5550 19320
rect -3950 19200 550 19300
rect -5950 19100 550 19200
rect -5950 19080 -5830 19100
rect -5570 19080 -5330 19100
rect -5070 19080 -4830 19100
rect -4570 19080 -4330 19100
rect -4070 19080 -3830 19100
rect -3570 19080 -3330 19100
rect -3070 19080 -2830 19100
rect -2570 19080 -2330 19100
rect -2070 19080 -1830 19100
rect -1570 19080 -1330 19100
rect -1070 19080 -830 19100
rect -570 19080 -330 19100
rect -70 19080 170 19100
rect 430 19080 550 19100
rect -5950 18820 -5850 19080
rect -5550 18820 -5350 19080
rect -5050 18820 -4850 19080
rect -4550 18820 -4350 19080
rect -4050 18820 -3850 19080
rect -3550 18820 -3350 19080
rect -3050 18820 -2850 19080
rect -2550 18820 -2350 19080
rect -2050 18820 -1850 19080
rect -1550 18820 -1350 19080
rect -1050 18820 -850 19080
rect -550 18820 -350 19080
rect -50 18820 150 19080
rect 450 18820 550 19080
rect -5950 18800 -5830 18820
rect -5570 18800 -5330 18820
rect -5070 18800 -4830 18820
rect -4570 18800 -4330 18820
rect -4070 18800 -3830 18820
rect -3570 18800 -3330 18820
rect -3070 18800 -2830 18820
rect -2570 18800 -2330 18820
rect -2070 18800 -1830 18820
rect -1570 18800 -1330 18820
rect -1070 18800 -830 18820
rect -570 18800 -330 18820
rect -70 18800 170 18820
rect 430 18800 550 18820
rect -5950 18600 550 18800
rect -5950 18580 -5830 18600
rect -5570 18580 -5330 18600
rect -5070 18580 -4830 18600
rect -4570 18580 -4330 18600
rect -4070 18580 -3830 18600
rect -3570 18580 -3330 18600
rect -3070 18580 -2830 18600
rect -2570 18580 -2330 18600
rect -2070 18580 -1830 18600
rect -1570 18580 -1330 18600
rect -1070 18580 -830 18600
rect -570 18580 -330 18600
rect -70 18580 170 18600
rect 430 18580 550 18600
rect -5950 18320 -5850 18580
rect -5550 18320 -5350 18580
rect -5050 18320 -4850 18580
rect -4550 18320 -4350 18580
rect -4050 18320 -3850 18580
rect -3550 18320 -3350 18580
rect -3050 18320 -2850 18580
rect -2550 18320 -2350 18580
rect -2050 18320 -1850 18580
rect -1550 18320 -1350 18580
rect -1050 18320 -850 18580
rect -550 18320 -350 18580
rect -50 18320 150 18580
rect 450 18320 550 18580
rect -5950 18300 -5830 18320
rect -5570 18300 -5330 18320
rect -5070 18300 -4830 18320
rect -4570 18300 -4330 18320
rect -4070 18300 -3830 18320
rect -3570 18300 -3330 18320
rect -3070 18300 -2830 18320
rect -2570 18300 -2330 18320
rect -2070 18300 -1830 18320
rect -1570 18300 -1330 18320
rect -1070 18300 -830 18320
rect -570 18300 -330 18320
rect -70 18300 170 18320
rect 430 18300 550 18320
rect -5950 18200 550 18300
rect -7950 18100 550 18200
rect -7950 18080 -7830 18100
rect -7570 18080 -7330 18100
rect -7070 18080 -6830 18100
rect -6570 18080 -6330 18100
rect -6070 18080 -5830 18100
rect -5570 18080 -5330 18100
rect -5070 18080 -4830 18100
rect -4570 18080 -4330 18100
rect -4070 18080 -3830 18100
rect -3570 18080 -3330 18100
rect -3070 18080 -2830 18100
rect -2570 18080 -2330 18100
rect -2070 18080 -1830 18100
rect -1570 18080 -1330 18100
rect -1070 18080 -830 18100
rect -570 18080 -330 18100
rect -70 18080 170 18100
rect 430 18080 550 18100
rect -7950 17820 -7850 18080
rect -7550 17820 -7350 18080
rect -7050 17820 -6850 18080
rect -6550 17820 -6350 18080
rect -6050 17820 -5850 18080
rect -5550 17820 -5350 18080
rect -5050 17820 -4850 18080
rect -4550 17820 -4350 18080
rect -4050 17820 -3850 18080
rect -3550 17820 -3350 18080
rect -3050 17820 -2850 18080
rect -2550 17820 -2350 18080
rect -2050 17820 -1850 18080
rect -1550 17820 -1350 18080
rect -1050 17820 -850 18080
rect -550 17820 -350 18080
rect -50 17820 150 18080
rect 450 18000 550 18080
rect 3700 19100 5550 19300
rect 3700 19080 4170 19100
rect 4430 19080 4670 19100
rect 4930 19080 5170 19100
rect 5430 19080 5550 19100
rect 3700 18820 4150 19080
rect 4450 18820 4650 19080
rect 4950 18820 5150 19080
rect 5450 18820 5550 19080
rect 3700 18800 4170 18820
rect 4430 18800 4670 18820
rect 4930 18800 5170 18820
rect 5430 18800 5550 18820
rect 3700 18600 5550 18800
rect 3700 18580 4170 18600
rect 4430 18580 4670 18600
rect 4930 18580 5170 18600
rect 5430 18580 5550 18600
rect 3700 18320 4150 18580
rect 4450 18320 4650 18580
rect 4950 18320 5150 18580
rect 5450 18320 5550 18580
rect 3700 18300 4170 18320
rect 4430 18300 4670 18320
rect 4930 18300 5170 18320
rect 5430 18300 5550 18320
rect 3700 18100 5550 18300
rect 3700 18080 4170 18100
rect 4430 18080 4670 18100
rect 4930 18080 5170 18100
rect 5430 18080 5550 18100
rect 3700 18000 4150 18080
rect 450 17820 4150 18000
rect 4450 17820 4650 18080
rect 4950 17820 5150 18080
rect 5450 17820 5550 18080
rect -7950 17800 -7830 17820
rect -7570 17800 -7330 17820
rect -7070 17800 -6830 17820
rect -6570 17800 -6330 17820
rect -6070 17800 -5830 17820
rect -5570 17800 -5330 17820
rect -5070 17800 -4830 17820
rect -4570 17800 -4330 17820
rect -4070 17800 -3830 17820
rect -3570 17800 -3330 17820
rect -3070 17800 -2830 17820
rect -2570 17800 -2330 17820
rect -2070 17800 -1830 17820
rect -1570 17800 -1330 17820
rect -1070 17800 -830 17820
rect -570 17800 -330 17820
rect -70 17800 170 17820
rect 430 17800 4170 17820
rect 4430 17800 4670 17820
rect 4930 17800 5170 17820
rect 5430 17800 5550 17820
rect -7950 17700 5550 17800
rect 50 17600 5550 17700
rect 50 17580 170 17600
rect 430 17580 670 17600
rect 930 17580 1170 17600
rect 1430 17580 1670 17600
rect 1930 17580 2170 17600
rect 2430 17580 2670 17600
rect 2930 17580 3170 17600
rect 3430 17580 3670 17600
rect 3930 17580 4170 17600
rect 4430 17580 4670 17600
rect 4930 17580 5170 17600
rect 5430 17580 5550 17600
rect 50 17320 150 17580
rect 450 17320 650 17580
rect 950 17320 1150 17580
rect 1450 17320 1650 17580
rect 1950 17320 2150 17580
rect 2450 17320 2650 17580
rect 2950 17320 3150 17580
rect 3450 17320 3650 17580
rect 3950 17320 4150 17580
rect 4450 17320 4650 17580
rect 4950 17320 5150 17580
rect 5450 17320 5550 17580
rect 50 17300 170 17320
rect 430 17300 670 17320
rect 930 17300 1170 17320
rect 1430 17300 1670 17320
rect 1930 17300 2170 17320
rect 2430 17300 2670 17320
rect 2930 17300 3170 17320
rect 3430 17300 3670 17320
rect 3930 17300 4170 17320
rect 4430 17300 4670 17320
rect 4930 17300 5170 17320
rect 5430 17300 5550 17320
rect 50 17200 5550 17300
rect -5950 -1900 50 -1800
rect -5950 -1920 -5830 -1900
rect -5570 -1920 -5330 -1900
rect -5070 -1920 -4830 -1900
rect -4570 -1920 -4330 -1900
rect -4070 -1920 -3830 -1900
rect -3570 -1920 -3330 -1900
rect -3070 -1920 -2830 -1900
rect -2570 -1920 -2330 -1900
rect -2070 -1920 -1830 -1900
rect -1570 -1920 -1330 -1900
rect -1070 -1920 -830 -1900
rect -570 -1920 -330 -1900
rect -70 -1920 50 -1900
rect -5950 -2180 -5850 -1920
rect -5550 -2180 -5350 -1920
rect -5050 -2180 -4850 -1920
rect -4550 -2180 -4350 -1920
rect -4050 -2180 -3850 -1920
rect -3550 -2180 -3350 -1920
rect -3050 -2180 -2850 -1920
rect -2550 -2180 -2350 -1920
rect -2050 -2180 -1850 -1920
rect -1550 -2180 -1350 -1920
rect -1050 -2180 -850 -1920
rect -550 -2180 -350 -1920
rect -50 -2180 50 -1920
rect -5950 -2200 -5830 -2180
rect -5570 -2200 -5330 -2180
rect -5070 -2200 -4830 -2180
rect -4570 -2200 -4330 -2180
rect -4070 -2200 -3830 -2180
rect -3570 -2200 -3330 -2180
rect -3070 -2200 -2830 -2180
rect -2570 -2200 -2330 -2180
rect -2070 -2200 -1830 -2180
rect -1570 -2200 -1330 -2180
rect -1070 -2200 -830 -2180
rect -570 -2200 -330 -2180
rect -70 -2200 50 -2180
rect -5950 -2300 50 -2200
rect -5950 -2400 4550 -2300
rect -5950 -2420 -5830 -2400
rect -5570 -2420 -5330 -2400
rect -5070 -2420 -4830 -2400
rect -4570 -2420 -4330 -2400
rect -4070 -2420 -3830 -2400
rect -3570 -2420 -3330 -2400
rect -3070 -2420 -2830 -2400
rect -2570 -2420 -2330 -2400
rect -2070 -2420 -1830 -2400
rect -1570 -2420 -1330 -2400
rect -1070 -2420 -830 -2400
rect -570 -2420 -330 -2400
rect -70 -2420 170 -2400
rect 430 -2420 670 -2400
rect 930 -2420 1170 -2400
rect 1430 -2420 1670 -2400
rect 1930 -2420 2170 -2400
rect 2430 -2420 2670 -2400
rect 2930 -2420 3170 -2400
rect 3430 -2420 3670 -2400
rect 3930 -2420 4170 -2400
rect 4430 -2420 4550 -2400
rect -5950 -2680 -5850 -2420
rect -5550 -2680 -5350 -2420
rect -5050 -2680 -4850 -2420
rect -4550 -2680 -4350 -2420
rect -4050 -2680 -3850 -2420
rect -3550 -2680 -3350 -2420
rect -3050 -2680 -2850 -2420
rect -2550 -2680 -2350 -2420
rect -2050 -2680 -1850 -2420
rect -1550 -2680 -1350 -2420
rect -1050 -2680 -850 -2420
rect -550 -2680 -350 -2420
rect -50 -2680 150 -2420
rect 450 -2680 650 -2420
rect 950 -2680 1150 -2420
rect 1450 -2680 1650 -2420
rect 1950 -2680 2150 -2420
rect 2450 -2680 2650 -2420
rect 2950 -2680 3150 -2420
rect 3450 -2680 3650 -2420
rect 3950 -2680 4150 -2420
rect 4450 -2680 4550 -2420
rect -5950 -2700 -5830 -2680
rect -5570 -2700 -5330 -2680
rect -5070 -2700 -4830 -2680
rect -4570 -2700 -4330 -2680
rect -4070 -2700 -3830 -2680
rect -3570 -2700 -3330 -2680
rect -3070 -2700 -2830 -2680
rect -2570 -2700 -2330 -2680
rect -2070 -2700 -1830 -2680
rect -1570 -2700 -1330 -2680
rect -1070 -2700 -830 -2680
rect -570 -2700 -330 -2680
rect -70 -2700 170 -2680
rect 430 -2700 670 -2680
rect 930 -2700 1170 -2680
rect 1430 -2700 1670 -2680
rect 1930 -2700 2170 -2680
rect 2430 -2700 2670 -2680
rect 2930 -2700 3170 -2680
rect 3430 -2700 3670 -2680
rect 3930 -2700 4170 -2680
rect 4430 -2700 4550 -2680
rect -5950 -2900 4550 -2700
rect -5950 -2920 -5830 -2900
rect -5570 -2920 -5330 -2900
rect -5070 -2920 -4830 -2900
rect -4570 -2920 -4330 -2900
rect -4070 -2920 -3830 -2900
rect -3570 -2920 -3330 -2900
rect -3070 -2920 -2830 -2900
rect -2570 -2920 -2330 -2900
rect -2070 -2920 -1830 -2900
rect -1570 -2920 -1330 -2900
rect -1070 -2920 -830 -2900
rect -570 -2920 -330 -2900
rect -70 -2920 170 -2900
rect 430 -2920 670 -2900
rect 930 -2920 1170 -2900
rect 1430 -2920 1670 -2900
rect 1930 -2920 2170 -2900
rect 2430 -2920 2670 -2900
rect 2930 -2920 3170 -2900
rect 3430 -2920 3670 -2900
rect 3930 -2920 4170 -2900
rect 4430 -2920 4550 -2900
rect -5950 -3180 -5850 -2920
rect -5550 -3180 -5350 -2920
rect -5050 -3180 -4850 -2920
rect -4550 -3180 -4350 -2920
rect -4050 -3180 -3850 -2920
rect -3550 -3180 -3350 -2920
rect -3050 -3180 -2850 -2920
rect -2550 -3180 -2350 -2920
rect -2050 -3180 -1850 -2920
rect -1550 -3180 -1350 -2920
rect -1050 -3180 -850 -2920
rect -550 -3180 -350 -2920
rect -50 -3180 150 -2920
rect 450 -3180 650 -2920
rect 950 -3180 1150 -2920
rect 1450 -3180 1650 -2920
rect 1950 -3180 2150 -2920
rect 2450 -3180 2650 -2920
rect 2950 -3180 3150 -2920
rect 3450 -3180 3650 -2920
rect 3950 -3180 4150 -2920
rect 4450 -3180 4550 -2920
rect -5950 -3200 -5830 -3180
rect -5570 -3200 -5330 -3180
rect -5070 -3200 -4830 -3180
rect -4570 -3200 -4330 -3180
rect -4070 -3200 -3830 -3180
rect -3570 -3200 -3330 -3180
rect -3070 -3200 -2830 -3180
rect -2570 -3200 -2330 -3180
rect -2070 -3200 -1830 -3180
rect -1570 -3200 -1330 -3180
rect -1070 -3200 -830 -3180
rect -570 -3200 -330 -3180
rect -70 -3200 170 -3180
rect 430 -3200 670 -3180
rect 930 -3200 1170 -3180
rect 1430 -3200 1670 -3180
rect 1930 -3200 2170 -3180
rect 2430 -3200 2670 -3180
rect 2930 -3200 3170 -3180
rect 3430 -3200 3670 -3180
rect 3930 -3200 4170 -3180
rect 4430 -3200 4550 -3180
rect -5950 -3400 4550 -3200
rect -5950 -3420 -5830 -3400
rect -5570 -3420 -5330 -3400
rect -5070 -3420 -4830 -3400
rect -4570 -3420 -4330 -3400
rect -4070 -3420 -3830 -3400
rect -3570 -3420 -3330 -3400
rect -3070 -3420 -2830 -3400
rect -2570 -3420 -2330 -3400
rect -2070 -3420 -1830 -3400
rect -1570 -3420 -1330 -3400
rect -1070 -3420 -830 -3400
rect -570 -3420 -330 -3400
rect -70 -3420 170 -3400
rect 430 -3420 670 -3400
rect 930 -3420 1170 -3400
rect 1430 -3420 1670 -3400
rect 1930 -3420 2170 -3400
rect 2430 -3420 2670 -3400
rect 2930 -3420 3170 -3400
rect 3430 -3420 3670 -3400
rect 3930 -3420 4170 -3400
rect 4430 -3420 4550 -3400
rect -5950 -3680 -5850 -3420
rect -5550 -3680 -5350 -3420
rect -5050 -3680 -4850 -3420
rect -4550 -3680 -4350 -3420
rect -4050 -3680 -3850 -3420
rect -3550 -3680 -3350 -3420
rect -3050 -3680 -2850 -3420
rect -2550 -3680 -2350 -3420
rect -2050 -3680 -1850 -3420
rect -1550 -3680 -1350 -3420
rect -1050 -3680 -850 -3420
rect -550 -3680 -350 -3420
rect -50 -3680 150 -3420
rect 450 -3680 650 -3420
rect 950 -3680 1150 -3420
rect 1450 -3680 1650 -3420
rect 1950 -3680 2150 -3420
rect 2450 -3680 2650 -3420
rect 2950 -3680 3150 -3420
rect 3450 -3680 3650 -3420
rect 3950 -3680 4150 -3420
rect 4450 -3680 4550 -3420
rect -5950 -3700 -5830 -3680
rect -5570 -3700 -5330 -3680
rect -5070 -3700 -4830 -3680
rect -4570 -3700 -4330 -3680
rect -4070 -3700 -3830 -3680
rect -3570 -3700 -3330 -3680
rect -3070 -3700 -2830 -3680
rect -2570 -3700 -2330 -3680
rect -2070 -3700 -1830 -3680
rect -1570 -3700 -1330 -3680
rect -1070 -3700 -830 -3680
rect -570 -3700 -330 -3680
rect -70 -3700 170 -3680
rect 430 -3700 670 -3680
rect 930 -3700 1170 -3680
rect 1430 -3700 1670 -3680
rect 1930 -3700 2170 -3680
rect 2430 -3700 2670 -3680
rect 2930 -3700 3170 -3680
rect 3430 -3700 3670 -3680
rect 3930 -3700 4170 -3680
rect 4430 -3700 4550 -3680
rect -5950 -3900 4550 -3700
rect -5950 -3920 -5830 -3900
rect -5570 -3920 -5330 -3900
rect -5070 -3920 -4830 -3900
rect -4570 -3920 -4330 -3900
rect -4070 -3920 -3830 -3900
rect -3570 -3920 -3330 -3900
rect -3070 -3920 -2830 -3900
rect -2570 -3920 -2330 -3900
rect -2070 -3920 -1830 -3900
rect -1570 -3920 -1330 -3900
rect -1070 -3920 -830 -3900
rect -570 -3920 -330 -3900
rect -70 -3920 170 -3900
rect 430 -3920 670 -3900
rect 930 -3920 1170 -3900
rect 1430 -3920 1670 -3900
rect 1930 -3920 2170 -3900
rect 2430 -3920 2670 -3900
rect 2930 -3920 3170 -3900
rect 3430 -3920 3670 -3900
rect 3930 -3920 4170 -3900
rect 4430 -3920 4550 -3900
rect -5950 -4180 -5850 -3920
rect -5550 -4180 -5350 -3920
rect -5050 -4180 -4850 -3920
rect -4550 -4180 -4350 -3920
rect -4050 -4180 -3850 -3920
rect -3550 -4180 -3350 -3920
rect -3050 -4180 -2850 -3920
rect -2550 -4180 -2350 -3920
rect -2050 -4180 -1850 -3920
rect -1550 -4180 -1350 -3920
rect -1050 -4180 -850 -3920
rect -550 -4180 -350 -3920
rect -50 -4180 150 -3920
rect 450 -4180 650 -3920
rect 950 -4180 1150 -3920
rect 1450 -4180 1650 -3920
rect 1950 -4180 2150 -3920
rect 2450 -4180 2650 -3920
rect 2950 -4180 3150 -3920
rect 3450 -4180 3650 -3920
rect 3950 -4180 4150 -3920
rect 4450 -4180 4550 -3920
rect -5950 -4200 -5830 -4180
rect -5570 -4200 -5330 -4180
rect -5070 -4200 -4830 -4180
rect -4570 -4200 -4330 -4180
rect -4070 -4200 -3830 -4180
rect -3570 -4200 -3330 -4180
rect -3070 -4200 -2830 -4180
rect -2570 -4200 -2330 -4180
rect -2070 -4200 -1830 -4180
rect -1570 -4200 -1330 -4180
rect -1070 -4200 -830 -4180
rect -570 -4200 -330 -4180
rect -70 -4200 170 -4180
rect 430 -4200 670 -4180
rect 930 -4200 1170 -4180
rect 1430 -4200 1670 -4180
rect 1930 -4200 2170 -4180
rect 2430 -4200 2670 -4180
rect 2930 -4200 3170 -4180
rect 3430 -4200 3670 -4180
rect 3930 -4200 4170 -4180
rect 4430 -4200 4550 -4180
rect -5950 -4400 4550 -4200
rect -5950 -4420 -5830 -4400
rect -5570 -4420 -5330 -4400
rect -5070 -4420 -4830 -4400
rect -4570 -4420 -4330 -4400
rect -4070 -4420 -3830 -4400
rect -3570 -4420 -3330 -4400
rect -3070 -4420 -2830 -4400
rect -2570 -4420 -2330 -4400
rect -2070 -4420 -1830 -4400
rect -1570 -4420 -1330 -4400
rect -1070 -4420 -830 -4400
rect -570 -4420 -330 -4400
rect -70 -4420 170 -4400
rect 430 -4420 670 -4400
rect 930 -4420 1170 -4400
rect 1430 -4420 1670 -4400
rect 1930 -4420 2170 -4400
rect 2430 -4420 2670 -4400
rect 2930 -4420 3170 -4400
rect 3430 -4420 3670 -4400
rect 3930 -4420 4170 -4400
rect 4430 -4420 4550 -4400
rect -5950 -4680 -5850 -4420
rect -5550 -4680 -5350 -4420
rect -5050 -4680 -4850 -4420
rect -4550 -4680 -4350 -4420
rect -4050 -4680 -3850 -4420
rect -3550 -4680 -3350 -4420
rect -3050 -4680 -2850 -4420
rect -2550 -4680 -2350 -4420
rect -2050 -4680 -1850 -4420
rect -1550 -4680 -1350 -4420
rect -1050 -4680 -850 -4420
rect -550 -4680 -350 -4420
rect -50 -4680 150 -4420
rect 450 -4680 650 -4420
rect 950 -4680 1150 -4420
rect 1450 -4680 1650 -4420
rect 1950 -4680 2150 -4420
rect 2450 -4680 2650 -4420
rect 2950 -4680 3150 -4420
rect 3450 -4680 3650 -4420
rect 3950 -4680 4150 -4420
rect 4450 -4680 4550 -4420
rect -5950 -4700 -5830 -4680
rect -5570 -4700 -5330 -4680
rect -5070 -4700 -4830 -4680
rect -4570 -4700 -4330 -4680
rect -4070 -4700 -3830 -4680
rect -3570 -4700 -3330 -4680
rect -3070 -4700 -2830 -4680
rect -2570 -4700 -2330 -4680
rect -2070 -4700 -1830 -4680
rect -1570 -4700 -1330 -4680
rect -1070 -4700 -830 -4680
rect -570 -4700 -330 -4680
rect -70 -4700 170 -4680
rect 430 -4700 670 -4680
rect 930 -4700 1170 -4680
rect 1430 -4700 1670 -4680
rect 1930 -4700 2170 -4680
rect 2430 -4700 2670 -4680
rect 2930 -4700 3170 -4680
rect 3430 -4700 3670 -4680
rect 3930 -4700 4170 -4680
rect 4430 -4700 4550 -4680
rect -5950 -4800 4550 -4700
<< via1 >>
rect -5080 20440 -5010 20550
rect -4540 20440 -4470 20550
rect -4640 19630 -4480 19730
<< metal2 >>
rect 7600 23560 8200 23600
rect 7600 23040 7640 23560
rect 8160 23040 8200 23560
rect 7600 23000 8200 23040
rect 7900 22300 8200 23000
rect 7900 22000 11000 22300
rect -5160 20840 -4960 20860
rect -5160 20580 -5140 20840
rect -4980 20580 -4960 20840
rect -5160 20560 -4960 20580
rect -4600 20840 -4400 20860
rect -4600 20580 -4580 20840
rect -4420 20580 -4400 20840
rect -4600 20560 -4400 20580
rect -5090 20550 -5000 20560
rect -5090 20440 -5080 20550
rect -5010 20440 -5000 20550
rect -5090 20430 -5000 20440
rect -4550 20550 -4460 20560
rect -4550 20440 -4540 20550
rect -4470 20440 -4460 20550
rect -4550 20430 -4460 20440
rect -4650 19730 -4470 19740
rect -4650 19540 -4640 19730
rect -4480 19540 -4470 19730
rect -4650 19530 -4470 19540
rect 10700 14900 11000 22000
rect 900 1600 2600 1650
rect 900 1250 950 1600
rect 2550 1250 2600 1600
rect 900 1200 2600 1250
rect 450 -2300 600 -2000
rect 750 -2300 900 -1990
rect 1050 -2300 1200 -1990
rect 1350 -2300 1500 -1990
rect 1650 -2300 1800 -1990
rect 1950 -2300 2100 -1990
rect 2250 -2300 2400 -1990
rect 2550 -2300 2700 -1990
rect 2850 -2300 3000 -1990
rect 3150 -2300 3300 -1990
rect 3450 -2300 3600 -1990
rect 3750 -2300 3900 -1990
rect 4050 -2300 4200 -1990
rect 4350 -2300 4500 -1990
rect 4650 -2300 4800 -1990
rect 400 -2350 4800 -2300
rect 400 -3050 450 -2350
rect 4750 -3050 4800 -2350
rect 400 -3100 4800 -3050
<< via2 >>
rect 7640 23040 8160 23560
rect -5140 20580 -4980 20840
rect -4580 20580 -4420 20840
rect -4640 19630 -4480 19730
rect -4640 19540 -4480 19630
rect 950 1250 2550 1600
rect 450 -3050 4750 -2350
<< metal3 >>
rect -5500 26200 -4400 26500
rect -4840 26100 -4400 26200
rect -5300 25420 -5000 25440
rect -5300 24180 -5280 25420
rect -5020 24180 -5000 25420
rect -5300 22380 -5000 24180
rect -5300 22300 -4920 22380
rect -5240 22220 -4860 22300
rect -5160 20860 -4860 22220
rect -4700 20860 -4400 26100
rect 7600 23560 8200 23600
rect 7600 23040 7640 23560
rect 8160 23040 8200 23560
rect 7600 23000 8200 23040
rect -5160 20840 -4960 20860
rect -5160 20580 -5140 20840
rect -4980 20580 -4960 20840
rect -5160 20560 -4960 20580
rect -4600 20840 -4400 20860
rect -4600 20580 -4580 20840
rect -4420 20580 -4400 20840
rect -4600 20560 -4400 20580
rect 6000 20500 11000 21400
rect -4650 19790 -4470 19800
rect -4650 19540 -4640 19790
rect -4480 19540 -4470 19790
rect -4650 19530 -4470 19540
rect -4850 19000 50 19450
rect -4850 18600 350 19000
rect -4850 18350 50 18600
rect 6000 16100 10400 20500
rect 10900 16100 11000 20500
rect 6000 16000 11000 16100
rect 650 1800 2850 1850
rect 650 1250 700 1800
rect 2800 1250 2850 1800
rect 650 1200 2850 1250
rect 3310 -470 3450 -460
rect 3310 -630 3320 -470
rect 3440 -630 3450 -470
rect 3310 -650 3450 -630
rect 400 -2350 4800 -2300
rect 400 -3050 450 -2350
rect 4750 -3050 4800 -2350
rect 400 -3100 4800 -3050
rect 400 -7600 4800 -3200
<< via3 >>
rect -5280 24180 -5020 25420
rect 7640 23040 8160 23560
rect -4640 19730 -4480 19790
rect -4640 19540 -4480 19730
rect 10400 16100 10900 20500
rect 700 1600 2800 1800
rect 700 1250 950 1600
rect 950 1250 2550 1600
rect 2550 1250 2800 1600
rect 3320 -630 3440 -470
rect 450 -3050 4750 -2350
<< mimcap >>
rect 6100 20400 10100 20500
rect -4800 19350 0 19400
rect -4800 18450 -4750 19350
rect -50 18450 0 19350
rect -4800 18400 0 18450
rect 6100 16200 6200 20400
rect 10000 16200 10100 20400
rect 6100 16100 10100 16200
rect 600 -3600 4600 -3400
rect 600 -7200 800 -3600
rect 4400 -7200 4600 -3600
rect 600 -7400 4600 -7200
<< mimcapcontact >>
rect -4750 18450 -50 19350
rect 6200 16200 10000 20400
rect 800 -7200 4400 -3600
<< metal4 >>
rect -1550 26100 -900 26700
rect -11040 20360 -10220 20920
rect -9620 20360 -8800 21360
rect -8260 20360 -7440 21360
rect -6940 20360 -6120 21480
rect -1550 20700 -1450 26100
rect 7600 23560 8200 23600
rect 7600 23040 7640 23560
rect 8160 23040 8200 23560
rect 7600 23000 8200 23040
rect -12880 20200 -6120 20360
rect 6000 20400 10200 20600
rect -4650 19790 -4470 19800
rect -4650 19540 -4640 19790
rect -4480 19540 -4470 19790
rect -4650 19400 -4470 19540
rect -4800 19350 0 19400
rect -4800 18450 -4750 19350
rect -50 18450 0 19350
rect -4800 18400 0 18450
rect 6000 18200 6200 20400
rect 4200 17400 6200 18200
rect 6000 16200 6200 17400
rect 10000 16200 10200 20400
rect 6000 16000 10200 16200
rect 10300 20500 11000 20600
rect 10300 16100 10400 20500
rect 10900 16100 11000 20500
rect 10300 16000 11000 16100
rect 3310 -434 3570 -430
rect 3310 -670 3320 -434
rect 3560 -670 3570 -434
rect 400 -2350 4800 -2200
rect 400 -3050 450 -2350
rect 4750 -3050 4800 -2350
rect 400 -3200 4800 -3050
rect 600 -3600 4600 -3200
rect 600 -7200 800 -3600
rect 4400 -7200 4600 -3600
rect 600 -7400 4600 -7200
<< via4 >>
rect 7640 23040 8160 23560
rect 10400 16100 10900 20500
rect 3320 -470 3560 -434
rect 3320 -630 3440 -470
rect 3440 -630 3560 -470
rect 3320 -670 3560 -630
<< mimcap2 >>
rect 6100 20400 10100 20500
rect 6100 16200 6200 20400
rect 10000 16200 10100 20400
rect 6100 16100 10100 16200
<< mimcap2contact >>
rect 6200 16200 10000 20400
<< metal5 >>
rect 7600 23560 8200 23600
rect 7600 23040 7640 23560
rect 8160 23040 8200 23560
rect 7600 23000 8200 23040
rect 6000 20500 11000 20600
rect 6000 20400 10400 20500
rect 6000 16200 6200 20400
rect 10000 16200 10400 20400
rect 6000 16100 10400 16200
rect 10900 16100 11000 20500
rect 6000 16000 11000 16100
rect 3200 -434 3800 -200
rect 3200 -670 3320 -434
rect 3560 -670 3800 -434
rect 3200 -1000 3800 -670
use OSC_5GHz_1  OSC_5GHz_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/OSC
timestamp 1660526289
transform -1 0 6096 0 -1 32150
box 10000 -14800 72400 31200
use PA_complete  PA_complete_0
timestamp 1660708745
transform 1 0 11200 0 1 15600
box -23000 -42000 71900 48000
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660275339
transform 1 0 -1050 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_1
timestamp 1660275339
transform 1 0 -1550 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_2
timestamp 1660275339
transform 1 0 -2050 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_3
timestamp 1660275339
transform 1 0 -2550 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_4
timestamp 1660275339
transform 1 0 -3050 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_5
timestamp 1660275339
transform 1 0 -3550 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_6
timestamp 1660275339
transform 1 0 -550 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_7
timestamp 1660275339
transform 1 0 -4050 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_8
timestamp 1660275339
transform 1 0 -4050 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_9
timestamp 1660275339
transform 1 0 -3550 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_10
timestamp 1660275339
transform 1 0 -3050 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_11
timestamp 1660275339
transform 1 0 -2550 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_12
timestamp 1660275339
transform 1 0 -2050 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_13
timestamp 1660275339
transform 1 0 -1550 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_14
timestamp 1660275339
transform 1 0 -1050 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_15
timestamp 1660275339
transform 1 0 -550 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_16
timestamp 1660275339
transform 1 0 -50 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_17
timestamp 1660275339
transform 1 0 450 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_18
timestamp 1660275339
transform 1 0 950 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_19
timestamp 1660275339
transform 1 0 1450 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_20
timestamp 1660275339
transform 1 0 1950 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_21
timestamp 1660275339
transform 1 0 2450 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_22
timestamp 1660275339
transform 1 0 2950 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_23
timestamp 1660275339
transform 1 0 3450 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_24
timestamp 1660275339
transform 1 0 3450 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_25
timestamp 1660275339
transform 1 0 3950 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_26
timestamp 1660275339
transform 1 0 4450 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_27
timestamp 1660275339
transform 1 0 4950 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_28
timestamp 1660275339
transform 1 0 3950 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_29
timestamp 1660275339
transform 1 0 4450 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_30
timestamp 1660275339
transform 1 0 4950 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_31
timestamp 1660275339
transform 1 0 3950 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_32
timestamp 1660275339
transform 1 0 4450 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_33
timestamp 1660275339
transform 1 0 4950 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_34
timestamp 1660275339
transform 1 0 3950 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_35
timestamp 1660275339
transform 1 0 4450 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_36
timestamp 1660275339
transform 1 0 4950 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_37
timestamp 1660275339
transform 1 0 3950 0 1 16800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_38
timestamp 1660275339
transform 1 0 4450 0 1 16800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_39
timestamp 1660275339
transform 1 0 4950 0 1 16800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_40
timestamp 1660275339
transform 1 0 3950 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_41
timestamp 1660275339
transform 1 0 4450 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_42
timestamp 1660275339
transform 1 0 4950 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_43
timestamp 1660275339
transform 1 0 3950 0 1 16300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_44
timestamp 1660275339
transform 1 0 4450 0 1 16300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_45
timestamp 1660275339
transform 1 0 4950 0 1 16300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_46
timestamp 1660275339
transform 1 0 3950 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_47
timestamp 1660275339
transform 1 0 4450 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_48
timestamp 1660275339
transform 1 0 4950 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501465
transform 1 0 -7950 0 1 19900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_1
timestamp 1659501465
transform 1 0 -9950 0 1 19900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_2
timestamp 1659501465
transform 1 0 -11950 0 1 19900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_3
timestamp 1659501465
transform 1 0 -11950 0 1 17900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_4
timestamp 1659501465
transform 1 0 -9950 0 1 17900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_5
timestamp 1659501465
transform 1 0 -11950 0 1 15900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_6
timestamp 1659501465
transform 1 0 -9950 0 1 15900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_7
timestamp 1659501465
transform 1 0 -11950 0 1 13900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_8
timestamp 1659501465
transform 1 0 -9950 0 1 13900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_9
timestamp 1659501465
transform 1 0 -11950 0 1 11900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_10
timestamp 1659501465
transform 1 0 -9950 0 1 9900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_11
timestamp 1659501465
transform 1 0 -11950 0 1 9900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_12
timestamp 1659501465
transform 1 0 -9950 0 1 11900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_13
timestamp 1659501465
transform 1 0 -11950 0 1 7900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_14
timestamp 1659501465
transform 1 0 -9950 0 1 7900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_15
timestamp 1659501465
transform 1 0 -11950 0 1 5900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_16
timestamp 1659501465
transform 1 0 -9950 0 1 5900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_17
timestamp 1659501465
transform 1 0 -11950 0 1 3900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_18
timestamp 1659501465
transform 1 0 -9950 0 1 1900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_19
timestamp 1659501465
transform 1 0 -11950 0 1 1900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_20
timestamp 1659501465
transform 1 0 -9950 0 1 3900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_21
timestamp 1659501465
transform 1 0 -11950 0 1 -100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_22
timestamp 1659501465
transform 1 0 -9950 0 1 -100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_23
timestamp 1659501465
transform 1 0 -1450 0 1 22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_26
timestamp 1659501465
transform 1 0 -1450 0 1 24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_27
timestamp 1659501465
transform 1 0 -7950 0 1 -100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_28
timestamp 1659501465
transform 1 0 -5950 0 1 -100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_31
timestamp 1659501465
transform 1 0 -3950 0 1 -100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_32
timestamp 1659501465
transform 1 0 -1950 0 1 -100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_33
timestamp 1659501465
transform 1 0 -1450 0 1 26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_36
timestamp 1659501465
transform 1 0 -15950 0 1 -100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_37
timestamp 1659501465
transform 1 0 -13950 0 1 -100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_38
timestamp 1659501465
transform 1 0 -15950 0 1 3900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_39
timestamp 1659501465
transform 1 0 -15950 0 1 1900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_40
timestamp 1659501465
transform 1 0 -13950 0 1 3900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_41
timestamp 1659501465
transform 1 0 -13950 0 1 1900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_42
timestamp 1659501465
transform 1 0 -15950 0 1 7900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_43
timestamp 1659501465
transform 1 0 -15950 0 1 5900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_44
timestamp 1659501465
transform 1 0 -13950 0 1 7900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_45
timestamp 1659501465
transform 1 0 -13950 0 1 5900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_46
timestamp 1659501465
transform 1 0 -15950 0 1 11900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_47
timestamp 1659501465
transform 1 0 -15950 0 1 9900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_48
timestamp 1659501465
transform 1 0 -13950 0 1 11900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_49
timestamp 1659501465
transform 1 0 -13950 0 1 9900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_51
timestamp 1659501465
transform 1 0 -15950 0 1 13900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_52
timestamp 1659501465
transform 1 0 -13950 0 1 15900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_53
timestamp 1659501465
transform 1 0 -13950 0 1 13900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_56
timestamp 1659501465
transform 1 0 -13950 0 1 19900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_57
timestamp 1659501465
transform 1 0 -13950 0 1 17900
box 0 -1700 2000 300
use pmirror_pfet_64x_complete  pmirror_pfet_64x_complete_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660185098
transform 1 0 400 0 1 -2100
box 0 0 4280 3344
use rfbcsa_1  rfbcsa_1_0
timestamp 1660307541
transform 1 0 650 0 1 18200
box -650 -18200 3840 2000
use sky130_fd_pr__res_generic_po_3TQ83P  sky130_fd_pr__res_generic_po_3TQ83P_0
timestamp 1659923628
transform 1 0 -4776 0 1 20086
box -577 -589 577 589
use spiral_ind_0p630nH_5GHz_to_gnd_noPGS  spiral_ind_0p630nH_5GHz_to_gnd_noPGS_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1659324110
transform 0 1 -4550 1 0 2200
box 0 -1600 15800 13000
<< labels >>
rlabel metal4 4200 17550 4500 18150 1 D
rlabel metal5 3200 -1000 3800 -200 1 IREF
<< end >>
