magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< locali >>
rect -43 652 81 686
<< metal1 >>
rect 336 12700 400 12752
rect 49 11955 113 12007
rect 164 11955 228 12007
rect 417 11955 481 12007
rect 785 11955 849 12007
rect 1153 11955 1217 12007
rect 1521 11955 1585 12007
rect 1440 11286 1504 11338
rect 49 10617 113 10669
rect 164 10617 228 10669
rect 417 10617 481 10669
rect 785 10617 849 10669
rect 1153 10617 1217 10669
rect 1521 10617 1585 10669
rect 336 9872 400 9924
rect 49 9127 113 9179
rect 164 9127 228 9179
rect 417 9127 481 9179
rect 785 9127 849 9179
rect 1153 9127 1217 9179
rect 1521 9127 1585 9179
rect 1440 8458 1504 8510
rect 49 7789 113 7841
rect 164 7789 228 7841
rect 417 7789 481 7841
rect 785 7789 849 7841
rect 1153 7789 1217 7841
rect 1521 7789 1585 7841
rect 336 7044 400 7096
rect 49 6299 113 6351
rect 164 6299 228 6351
rect 417 6299 481 6351
rect 785 6299 849 6351
rect 1153 6299 1217 6351
rect 1521 6299 1585 6351
rect 1440 5630 1504 5682
rect 49 4961 113 5013
rect 164 4961 228 5013
rect 417 4961 481 5013
rect 785 4961 849 5013
rect 1153 4961 1217 5013
rect 1521 4961 1585 5013
rect 336 4216 400 4268
rect 49 3471 113 3523
rect 164 3471 228 3523
rect 417 3471 481 3523
rect 785 3471 849 3523
rect 1153 3471 1217 3523
rect 1521 3471 1585 3523
rect 1440 2802 1504 2854
rect 49 2133 113 2185
rect 164 2133 228 2185
rect 417 2133 481 2185
rect 785 2133 849 2185
rect 1153 2133 1217 2185
rect 1521 2133 1585 2185
rect 336 1388 400 1440
rect -75 643 -11 695
rect 49 643 113 695
rect 164 643 228 695
rect 417 643 481 695
rect 785 643 849 695
rect 1153 643 1217 695
rect 1521 643 1585 695
rect 1440 -26 1504 26
<< metal2 >>
rect 340 12702 396 12750
rect 67 11326 95 11981
rect 168 11957 224 12005
rect 421 11957 477 12005
rect 789 11957 845 12005
rect 1157 11957 1213 12005
rect 1525 11957 1581 12005
rect 67 11298 210 11326
rect 182 10667 210 11298
rect 1444 11288 1500 11336
rect 67 9912 95 10643
rect 168 10619 224 10667
rect 421 10619 477 10667
rect 789 10619 845 10667
rect 1157 10619 1213 10667
rect 1525 10619 1581 10667
rect 67 9884 210 9912
rect 182 9177 210 9884
rect 340 9874 396 9922
rect 67 8498 95 9153
rect 168 9129 224 9177
rect 421 9129 477 9177
rect 789 9129 845 9177
rect 1157 9129 1213 9177
rect 1525 9129 1581 9177
rect 67 8470 210 8498
rect 182 7839 210 8470
rect 1444 8460 1500 8508
rect 67 7084 95 7815
rect 168 7791 224 7839
rect 421 7791 477 7839
rect 789 7791 845 7839
rect 1157 7791 1213 7839
rect 1525 7791 1581 7839
rect 67 7056 210 7084
rect 182 6349 210 7056
rect 340 7046 396 7094
rect 67 5670 95 6325
rect 168 6301 224 6349
rect 421 6301 477 6349
rect 789 6301 845 6349
rect 1157 6301 1213 6349
rect 1525 6301 1581 6349
rect 67 5642 210 5670
rect 182 5011 210 5642
rect 1444 5632 1500 5680
rect 67 4256 95 4987
rect 168 4963 224 5011
rect 421 4963 477 5011
rect 789 4963 845 5011
rect 1157 4963 1213 5011
rect 1525 4963 1581 5011
rect 67 4228 210 4256
rect 182 3521 210 4228
rect 340 4218 396 4266
rect 67 2842 95 3497
rect 168 3473 224 3521
rect 421 3473 477 3521
rect 789 3473 845 3521
rect 1157 3473 1213 3521
rect 1525 3473 1581 3521
rect 67 2814 210 2842
rect 182 2183 210 2814
rect 1444 2804 1500 2852
rect 67 1428 95 2159
rect 168 2135 224 2183
rect 421 2135 477 2183
rect 789 2135 845 2183
rect 1157 2135 1213 2183
rect 1525 2135 1581 2183
rect 67 1400 210 1428
rect 182 693 210 1400
rect 340 1390 396 1438
rect -57 655 -29 683
rect 168 645 224 693
rect 421 645 477 693
rect 789 645 845 693
rect 1157 645 1213 693
rect 1525 645 1581 693
rect 1444 -24 1500 24
<< metal3 >>
rect 293 12694 443 12758
rect 196 11951 1553 12011
rect 1397 11280 1547 11344
rect 196 10613 1553 10673
rect 293 9866 443 9930
rect 196 9123 1553 9183
rect 1397 8452 1547 8516
rect 196 7785 1553 7845
rect 293 7038 443 7102
rect 196 6295 1553 6355
rect 1397 5624 1547 5688
rect 196 4957 1553 5017
rect 293 4210 443 4274
rect 196 3467 1553 3527
rect 1397 2796 1547 2860
rect 196 2129 1553 2189
rect 293 1382 443 1446
rect 196 639 1553 699
rect 1397 -32 1547 32
<< metal4 >>
rect 335 -33 401 12776
rect 1439 -50 1505 12759
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 1524 0 1 11948
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 -72 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_2
timestamp 1661296025
transform 1 0 1443 0 1 11279
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_3
timestamp 1661296025
transform 1 0 1443 0 1 11279
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_4
timestamp 1661296025
transform 1 0 1443 0 1 8451
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_5
timestamp 1661296025
transform 1 0 1443 0 1 8451
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_6
timestamp 1661296025
transform 1 0 1443 0 1 5623
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_7
timestamp 1661296025
transform 1 0 1443 0 1 5623
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_8
timestamp 1661296025
transform 1 0 1443 0 1 2795
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_9
timestamp 1661296025
transform 1 0 1443 0 1 2795
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_10
timestamp 1661296025
transform 1 0 1443 0 1 -33
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_11
timestamp 1661296025
transform 1 0 339 0 1 12693
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_12
timestamp 1661296025
transform 1 0 339 0 1 9865
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_13
timestamp 1661296025
transform 1 0 339 0 1 9865
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_14
timestamp 1661296025
transform 1 0 339 0 1 7037
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_15
timestamp 1661296025
transform 1 0 339 0 1 7037
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_16
timestamp 1661296025
transform 1 0 339 0 1 4209
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_17
timestamp 1661296025
transform 1 0 339 0 1 4209
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_18
timestamp 1661296025
transform 1 0 339 0 1 1381
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_19
timestamp 1661296025
transform 1 0 339 0 1 1381
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_20
timestamp 1661296025
transform 1 0 167 0 1 11948
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_21
timestamp 1661296025
transform 1 0 52 0 1 11948
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_22
timestamp 1661296025
transform 1 0 1524 0 1 11948
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_23
timestamp 1661296025
transform 1 0 1156 0 1 11948
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_24
timestamp 1661296025
transform 1 0 788 0 1 11948
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_25
timestamp 1661296025
transform 1 0 420 0 1 11948
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_26
timestamp 1661296025
transform 1 0 167 0 1 10610
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_27
timestamp 1661296025
transform 1 0 52 0 1 10610
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_28
timestamp 1661296025
transform 1 0 1524 0 1 10610
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_29
timestamp 1661296025
transform 1 0 1156 0 1 10610
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_30
timestamp 1661296025
transform 1 0 788 0 1 10610
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_31
timestamp 1661296025
transform 1 0 420 0 1 10610
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_32
timestamp 1661296025
transform 1 0 167 0 1 9120
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_33
timestamp 1661296025
transform 1 0 52 0 1 9120
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_34
timestamp 1661296025
transform 1 0 1524 0 1 9120
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_35
timestamp 1661296025
transform 1 0 1156 0 1 9120
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_36
timestamp 1661296025
transform 1 0 788 0 1 9120
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_37
timestamp 1661296025
transform 1 0 420 0 1 9120
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_38
timestamp 1661296025
transform 1 0 167 0 1 7782
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_39
timestamp 1661296025
transform 1 0 52 0 1 7782
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_40
timestamp 1661296025
transform 1 0 1524 0 1 7782
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_41
timestamp 1661296025
transform 1 0 1156 0 1 7782
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_42
timestamp 1661296025
transform 1 0 788 0 1 7782
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_43
timestamp 1661296025
transform 1 0 420 0 1 7782
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_44
timestamp 1661296025
transform 1 0 167 0 1 6292
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_45
timestamp 1661296025
transform 1 0 52 0 1 6292
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_46
timestamp 1661296025
transform 1 0 1524 0 1 6292
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_47
timestamp 1661296025
transform 1 0 1156 0 1 6292
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_48
timestamp 1661296025
transform 1 0 788 0 1 6292
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_49
timestamp 1661296025
transform 1 0 420 0 1 6292
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_50
timestamp 1661296025
transform 1 0 167 0 1 4954
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_51
timestamp 1661296025
transform 1 0 52 0 1 4954
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_52
timestamp 1661296025
transform 1 0 1524 0 1 4954
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_53
timestamp 1661296025
transform 1 0 1156 0 1 4954
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_54
timestamp 1661296025
transform 1 0 788 0 1 4954
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_55
timestamp 1661296025
transform 1 0 420 0 1 4954
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_56
timestamp 1661296025
transform 1 0 167 0 1 3464
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_57
timestamp 1661296025
transform 1 0 52 0 1 3464
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_58
timestamp 1661296025
transform 1 0 1524 0 1 3464
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_59
timestamp 1661296025
transform 1 0 1156 0 1 3464
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_60
timestamp 1661296025
transform 1 0 788 0 1 3464
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_61
timestamp 1661296025
transform 1 0 420 0 1 3464
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_62
timestamp 1661296025
transform 1 0 167 0 1 2126
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_63
timestamp 1661296025
transform 1 0 52 0 1 2126
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_64
timestamp 1661296025
transform 1 0 1524 0 1 2126
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_65
timestamp 1661296025
transform 1 0 1156 0 1 2126
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_66
timestamp 1661296025
transform 1 0 788 0 1 2126
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_67
timestamp 1661296025
transform 1 0 420 0 1 2126
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_68
timestamp 1661296025
transform 1 0 167 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_69
timestamp 1661296025
transform 1 0 52 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_70
timestamp 1661296025
transform 1 0 1524 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_71
timestamp 1661296025
transform 1 0 1156 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_72
timestamp 1661296025
transform 1 0 788 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_73
timestamp 1661296025
transform 1 0 420 0 1 636
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_0
timestamp 1661296025
transform 1 0 -75 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_1
timestamp 1661296025
transform 1 0 1440 0 1 11280
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_2
timestamp 1661296025
transform 1 0 1440 0 1 11280
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_3
timestamp 1661296025
transform 1 0 1440 0 1 8452
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_4
timestamp 1661296025
transform 1 0 1440 0 1 8452
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_5
timestamp 1661296025
transform 1 0 1440 0 1 5624
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_6
timestamp 1661296025
transform 1 0 1440 0 1 5624
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_7
timestamp 1661296025
transform 1 0 1440 0 1 2796
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_8
timestamp 1661296025
transform 1 0 1440 0 1 2796
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_9
timestamp 1661296025
transform 1 0 1440 0 1 -32
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_10
timestamp 1661296025
transform 1 0 336 0 1 12694
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_11
timestamp 1661296025
transform 1 0 336 0 1 9866
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_12
timestamp 1661296025
transform 1 0 336 0 1 9866
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_13
timestamp 1661296025
transform 1 0 336 0 1 7038
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_14
timestamp 1661296025
transform 1 0 336 0 1 7038
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_15
timestamp 1661296025
transform 1 0 336 0 1 4210
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_16
timestamp 1661296025
transform 1 0 336 0 1 4210
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_17
timestamp 1661296025
transform 1 0 336 0 1 1382
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_18
timestamp 1661296025
transform 1 0 336 0 1 1382
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_19
timestamp 1661296025
transform 1 0 164 0 1 11949
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_20
timestamp 1661296025
transform 1 0 49 0 1 11949
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_21
timestamp 1661296025
transform 1 0 1521 0 1 11949
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_22
timestamp 1661296025
transform 1 0 1153 0 1 11949
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_23
timestamp 1661296025
transform 1 0 785 0 1 11949
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_24
timestamp 1661296025
transform 1 0 417 0 1 11949
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_25
timestamp 1661296025
transform 1 0 164 0 1 10611
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_26
timestamp 1661296025
transform 1 0 49 0 1 10611
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_27
timestamp 1661296025
transform 1 0 1521 0 1 10611
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_28
timestamp 1661296025
transform 1 0 1153 0 1 10611
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_29
timestamp 1661296025
transform 1 0 785 0 1 10611
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_30
timestamp 1661296025
transform 1 0 417 0 1 10611
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_31
timestamp 1661296025
transform 1 0 164 0 1 9121
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_32
timestamp 1661296025
transform 1 0 49 0 1 9121
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_33
timestamp 1661296025
transform 1 0 1521 0 1 9121
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_34
timestamp 1661296025
transform 1 0 1153 0 1 9121
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_35
timestamp 1661296025
transform 1 0 785 0 1 9121
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_36
timestamp 1661296025
transform 1 0 417 0 1 9121
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_37
timestamp 1661296025
transform 1 0 164 0 1 7783
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_38
timestamp 1661296025
transform 1 0 49 0 1 7783
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_39
timestamp 1661296025
transform 1 0 1521 0 1 7783
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_40
timestamp 1661296025
transform 1 0 1153 0 1 7783
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_41
timestamp 1661296025
transform 1 0 785 0 1 7783
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_42
timestamp 1661296025
transform 1 0 417 0 1 7783
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_43
timestamp 1661296025
transform 1 0 164 0 1 6293
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_44
timestamp 1661296025
transform 1 0 49 0 1 6293
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_45
timestamp 1661296025
transform 1 0 1521 0 1 6293
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_46
timestamp 1661296025
transform 1 0 1153 0 1 6293
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_47
timestamp 1661296025
transform 1 0 785 0 1 6293
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_48
timestamp 1661296025
transform 1 0 417 0 1 6293
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_49
timestamp 1661296025
transform 1 0 164 0 1 4955
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_50
timestamp 1661296025
transform 1 0 49 0 1 4955
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_51
timestamp 1661296025
transform 1 0 1521 0 1 4955
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_52
timestamp 1661296025
transform 1 0 1153 0 1 4955
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_53
timestamp 1661296025
transform 1 0 785 0 1 4955
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_54
timestamp 1661296025
transform 1 0 417 0 1 4955
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_55
timestamp 1661296025
transform 1 0 164 0 1 3465
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_56
timestamp 1661296025
transform 1 0 49 0 1 3465
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_57
timestamp 1661296025
transform 1 0 1521 0 1 3465
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_58
timestamp 1661296025
transform 1 0 1153 0 1 3465
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_59
timestamp 1661296025
transform 1 0 785 0 1 3465
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_60
timestamp 1661296025
transform 1 0 417 0 1 3465
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_61
timestamp 1661296025
transform 1 0 164 0 1 2127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_62
timestamp 1661296025
transform 1 0 49 0 1 2127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_63
timestamp 1661296025
transform 1 0 1521 0 1 2127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_64
timestamp 1661296025
transform 1 0 1153 0 1 2127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_65
timestamp 1661296025
transform 1 0 785 0 1 2127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_66
timestamp 1661296025
transform 1 0 417 0 1 2127
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_67
timestamp 1661296025
transform 1 0 164 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_68
timestamp 1661296025
transform 1 0 49 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_69
timestamp 1661296025
transform 1 0 1521 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_70
timestamp 1661296025
transform 1 0 1153 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_71
timestamp 1661296025
transform 1 0 785 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_72
timestamp 1661296025
transform 1 0 417 0 1 637
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_0
timestamp 1661296025
transform 1 0 1439 0 1 11275
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_1
timestamp 1661296025
transform 1 0 1439 0 1 11275
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_2
timestamp 1661296025
transform 1 0 1439 0 1 8447
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_3
timestamp 1661296025
transform 1 0 1439 0 1 8447
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_4
timestamp 1661296025
transform 1 0 1439 0 1 5619
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_5
timestamp 1661296025
transform 1 0 1439 0 1 5619
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_6
timestamp 1661296025
transform 1 0 1439 0 1 2791
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_7
timestamp 1661296025
transform 1 0 1439 0 1 2791
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_8
timestamp 1661296025
transform 1 0 1439 0 1 -37
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_9
timestamp 1661296025
transform 1 0 335 0 1 12689
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_10
timestamp 1661296025
transform 1 0 335 0 1 9861
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_11
timestamp 1661296025
transform 1 0 335 0 1 9861
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_12
timestamp 1661296025
transform 1 0 335 0 1 7033
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_13
timestamp 1661296025
transform 1 0 335 0 1 7033
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_14
timestamp 1661296025
transform 1 0 335 0 1 4205
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_15
timestamp 1661296025
transform 1 0 335 0 1 4205
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_16
timestamp 1661296025
transform 1 0 335 0 1 1377
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_17
timestamp 1661296025
transform 1 0 335 0 1 1377
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_18
timestamp 1661296025
transform 1 0 163 0 1 11944
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_19
timestamp 1661296025
transform 1 0 1520 0 1 11944
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_20
timestamp 1661296025
transform 1 0 1152 0 1 11944
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_21
timestamp 1661296025
transform 1 0 784 0 1 11944
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_22
timestamp 1661296025
transform 1 0 416 0 1 11944
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_23
timestamp 1661296025
transform 1 0 163 0 1 10606
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_24
timestamp 1661296025
transform 1 0 1520 0 1 10606
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_25
timestamp 1661296025
transform 1 0 1152 0 1 10606
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_26
timestamp 1661296025
transform 1 0 784 0 1 10606
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_27
timestamp 1661296025
transform 1 0 416 0 1 10606
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_28
timestamp 1661296025
transform 1 0 163 0 1 9116
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_29
timestamp 1661296025
transform 1 0 1520 0 1 9116
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_30
timestamp 1661296025
transform 1 0 1152 0 1 9116
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_31
timestamp 1661296025
transform 1 0 784 0 1 9116
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_32
timestamp 1661296025
transform 1 0 416 0 1 9116
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_33
timestamp 1661296025
transform 1 0 163 0 1 7778
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_34
timestamp 1661296025
transform 1 0 1520 0 1 7778
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_35
timestamp 1661296025
transform 1 0 1152 0 1 7778
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_36
timestamp 1661296025
transform 1 0 784 0 1 7778
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_37
timestamp 1661296025
transform 1 0 416 0 1 7778
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_38
timestamp 1661296025
transform 1 0 163 0 1 6288
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_39
timestamp 1661296025
transform 1 0 1520 0 1 6288
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_40
timestamp 1661296025
transform 1 0 1152 0 1 6288
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_41
timestamp 1661296025
transform 1 0 784 0 1 6288
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_42
timestamp 1661296025
transform 1 0 416 0 1 6288
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_43
timestamp 1661296025
transform 1 0 163 0 1 4950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_44
timestamp 1661296025
transform 1 0 1520 0 1 4950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_45
timestamp 1661296025
transform 1 0 1152 0 1 4950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_46
timestamp 1661296025
transform 1 0 784 0 1 4950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_47
timestamp 1661296025
transform 1 0 416 0 1 4950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_48
timestamp 1661296025
transform 1 0 163 0 1 3460
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_49
timestamp 1661296025
transform 1 0 1520 0 1 3460
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_50
timestamp 1661296025
transform 1 0 1152 0 1 3460
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_51
timestamp 1661296025
transform 1 0 784 0 1 3460
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_52
timestamp 1661296025
transform 1 0 416 0 1 3460
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_53
timestamp 1661296025
transform 1 0 163 0 1 2122
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_54
timestamp 1661296025
transform 1 0 1520 0 1 2122
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_55
timestamp 1661296025
transform 1 0 1152 0 1 2122
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_56
timestamp 1661296025
transform 1 0 784 0 1 2122
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_57
timestamp 1661296025
transform 1 0 416 0 1 2122
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_58
timestamp 1661296025
transform 1 0 163 0 1 632
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_59
timestamp 1661296025
transform 1 0 1520 0 1 632
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_60
timestamp 1661296025
transform 1 0 1152 0 1 632
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_61
timestamp 1661296025
transform 1 0 784 0 1 632
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_62
timestamp 1661296025
transform 1 0 416 0 1 632
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_0
timestamp 1661296025
transform 1 0 1434 0 1 11279
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_1
timestamp 1661296025
transform 1 0 1434 0 1 11279
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_2
timestamp 1661296025
transform 1 0 1434 0 1 8451
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_3
timestamp 1661296025
transform 1 0 1434 0 1 8451
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_4
timestamp 1661296025
transform 1 0 1434 0 1 5623
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_5
timestamp 1661296025
transform 1 0 1434 0 1 5623
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_6
timestamp 1661296025
transform 1 0 1434 0 1 2795
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_7
timestamp 1661296025
transform 1 0 1434 0 1 2795
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_8
timestamp 1661296025
transform 1 0 1434 0 1 -33
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_9
timestamp 1661296025
transform 1 0 330 0 1 12693
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_10
timestamp 1661296025
transform 1 0 330 0 1 9865
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_11
timestamp 1661296025
transform 1 0 330 0 1 9865
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_12
timestamp 1661296025
transform 1 0 330 0 1 7037
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_13
timestamp 1661296025
transform 1 0 330 0 1 7037
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_14
timestamp 1661296025
transform 1 0 330 0 1 4209
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_15
timestamp 1661296025
transform 1 0 330 0 1 4209
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_16
timestamp 1661296025
transform 1 0 330 0 1 1381
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_17
timestamp 1661296025
transform 1 0 330 0 1 1381
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_0
timestamp 1661296025
transform 1 0 1472 0 1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_1
timestamp 1661296025
transform 1 0 1104 0 1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_2
timestamp 1661296025
transform 1 0 736 0 1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_3
timestamp 1661296025
transform 1 0 368 0 1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_4
timestamp 1661296025
transform 1 0 0 0 1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_5
timestamp 1661296025
transform 1 0 1472 0 -1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_6
timestamp 1661296025
transform 1 0 1104 0 -1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_7
timestamp 1661296025
transform 1 0 736 0 -1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_8
timestamp 1661296025
transform 1 0 368 0 -1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_9
timestamp 1661296025
transform 1 0 0 0 -1 11312
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_10
timestamp 1661296025
transform 1 0 1472 0 1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_11
timestamp 1661296025
transform 1 0 1104 0 1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_12
timestamp 1661296025
transform 1 0 736 0 1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_13
timestamp 1661296025
transform 1 0 368 0 1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_14
timestamp 1661296025
transform 1 0 0 0 1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_15
timestamp 1661296025
transform 1 0 1472 0 -1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_16
timestamp 1661296025
transform 1 0 1104 0 -1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_17
timestamp 1661296025
transform 1 0 736 0 -1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_18
timestamp 1661296025
transform 1 0 368 0 -1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_19
timestamp 1661296025
transform 1 0 0 0 -1 8484
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_20
timestamp 1661296025
transform 1 0 1472 0 1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_21
timestamp 1661296025
transform 1 0 1104 0 1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_22
timestamp 1661296025
transform 1 0 736 0 1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_23
timestamp 1661296025
transform 1 0 368 0 1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_24
timestamp 1661296025
transform 1 0 0 0 1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_25
timestamp 1661296025
transform 1 0 1472 0 -1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_26
timestamp 1661296025
transform 1 0 1104 0 -1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_27
timestamp 1661296025
transform 1 0 736 0 -1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_28
timestamp 1661296025
transform 1 0 368 0 -1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_29
timestamp 1661296025
transform 1 0 0 0 -1 5656
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_30
timestamp 1661296025
transform 1 0 1472 0 1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_31
timestamp 1661296025
transform 1 0 1104 0 1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_32
timestamp 1661296025
transform 1 0 736 0 1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_33
timestamp 1661296025
transform 1 0 368 0 1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_34
timestamp 1661296025
transform 1 0 0 0 1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_35
timestamp 1661296025
transform 1 0 1472 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_36
timestamp 1661296025
transform 1 0 1104 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_37
timestamp 1661296025
transform 1 0 736 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_38
timestamp 1661296025
transform 1 0 368 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_39
timestamp 1661296025
transform 1 0 0 0 -1 2828
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_40
timestamp 1661296025
transform 1 0 1472 0 1 0
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_41
timestamp 1661296025
transform 1 0 1104 0 1 0
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_42
timestamp 1661296025
transform 1 0 736 0 1 0
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_43
timestamp 1661296025
transform 1 0 368 0 1 0
box -36 -17 404 1471
use sky130_sram_1r1w_24x128_8_pinv_16  sky130_sram_1r1w_24x128_8_pinv_16_44
timestamp 1661296025
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel metal4 s 335 -33 401 12776 4 vdd
port 1 nsew
rlabel metal4 s 1439 -50 1505 12759 4 gnd
port 2 nsew
rlabel metal2 s -57 655 -29 683 4 in
port 3 nsew
rlabel metal1 s 1539 11967 1567 11995 4 out
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1840 12726
<< end >>
