magic
tech sky130A
magscale 1 2
timestamp 1664895471
<< error_s >>
rect 1000 400 1024 1200
<< pwell >>
rect 30600 12500 31000 14016
<< psubdiff >>
rect 30634 13946 30730 13980
rect 30868 13946 30964 13980
rect 30634 13884 30668 13946
rect 30930 13884 30964 13946
rect 30634 12570 30668 12632
rect 30930 12570 30964 12632
rect 30634 12536 30730 12570
rect 30868 12536 30964 12570
<< psubdiffcont >>
rect 30730 13946 30868 13980
rect 30634 12632 30668 13884
rect 30930 12632 30964 13884
rect 30730 12536 30868 12570
<< xpolycontact >>
rect 30764 13418 30834 13850
rect 30764 12666 30834 13098
<< ppolyres >>
rect 30764 13098 30834 13418
<< locali >>
rect 30634 13946 30730 13980
rect 30868 13946 30964 13980
rect 30634 13884 30668 13946
rect 30930 13884 30964 13946
rect 30634 12570 30668 12632
rect 30930 12570 30964 12632
rect 30634 12536 30730 12570
rect 30868 12536 30964 12570
<< viali >>
rect 30780 13435 30818 13832
rect 30780 12684 30818 13081
<< metal1 >>
rect 26540 39190 26780 39200
rect 26540 39010 26550 39190
rect 26770 39010 26780 39190
rect 26540 39000 26780 39010
rect 28080 39190 28320 39200
rect 28080 39010 28090 39190
rect 28310 39010 28320 39190
rect 28080 39000 28320 39010
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect 30700 13900 30900 13910
rect 30700 13420 30710 13900
rect 30890 13420 30900 13900
rect 30700 13410 30900 13420
rect 30700 13090 30900 13100
rect 30700 12610 30710 13090
rect 30890 12610 30900 13090
rect 30700 12600 30900 12610
<< via1 >>
rect 26550 39010 26770 39190
rect 28090 39010 28310 39190
rect 30910 27030 31090 27250
rect 30910 25490 31090 25710
rect 30710 13832 30890 13900
rect 30710 13435 30780 13832
rect 30780 13435 30818 13832
rect 30818 13435 30890 13832
rect 30710 13420 30890 13435
rect 30710 13081 30890 13090
rect 30710 12684 30780 13081
rect 30780 12684 30818 13081
rect 30818 12684 30890 13081
rect 30710 12610 30890 12684
<< metal2 >>
rect 26540 39190 26780 39200
rect 26540 39010 26550 39190
rect 26770 39010 26780 39190
rect 26540 39000 26780 39010
rect 28080 39190 28320 39200
rect 28080 39010 28090 39190
rect 28310 39010 28320 39190
rect 28080 39000 28320 39010
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect 30700 13900 30900 13910
rect 30700 13420 30710 13900
rect 30890 13420 30900 13900
rect 30700 13410 30900 13420
rect 30700 13090 30900 13100
rect 30700 12610 30710 13090
rect 30890 12610 30900 13090
rect 30700 12600 30900 12610
<< via2 >>
rect 26550 39010 26770 39190
rect 28090 39010 28310 39190
rect 30910 27030 31090 27250
rect 30910 25490 31090 25710
rect 30710 13420 30890 13900
rect 30710 12610 30890 13090
<< metal3 >>
rect 26500 39280 26800 39300
rect 26500 38920 26520 39280
rect 26780 38920 26800 39280
rect 26500 38900 26800 38920
rect 28080 39290 28320 39300
rect 28080 38910 28090 39290
rect 28310 38910 28320 39290
rect 28080 38900 28320 38910
rect 1000 31700 2800 31800
rect 1000 31100 1400 31700
rect 2700 31100 2800 31700
rect 1000 31000 2800 31100
rect 24000 31700 31200 31800
rect 24000 31100 24100 31700
rect 25400 31100 31200 31700
rect 24000 31000 31200 31100
rect 30700 27250 31200 31000
rect 30700 27030 30910 27250
rect 31090 27030 31200 27250
rect 30700 27000 31200 27030
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25480 31200 25490
rect 30600 14000 31000 14010
rect 30600 13420 30610 14000
rect 30990 13420 31000 14000
rect 30600 13410 31000 13420
rect 30600 13090 31000 13100
rect 30600 12510 30610 13090
rect 30990 12510 31000 13090
rect 30600 12500 31000 12510
<< via3 >>
rect 26520 39190 26780 39280
rect 26520 39010 26550 39190
rect 26550 39010 26770 39190
rect 26770 39010 26780 39190
rect 26520 38920 26780 39010
rect 28090 39190 28310 39290
rect 28090 39010 28310 39190
rect 28090 38910 28310 39010
rect 1400 31100 2700 31700
rect 24100 31100 25400 31700
rect 30810 25490 30910 25710
rect 30910 25490 31090 25710
rect 31090 25490 31190 25710
rect 30610 13900 30990 14000
rect 30610 13420 30710 13900
rect 30710 13420 30890 13900
rect 30890 13420 30990 13900
rect 30610 12610 30710 13090
rect 30710 12610 30890 13090
rect 30890 12610 30990 13090
rect 30610 12510 30990 12610
<< metal4 >>
rect 26000 47500 27400 47600
rect 26000 46500 26100 47500
rect 27300 46500 27400 47500
rect 26000 46400 27400 46500
rect 26000 46000 27800 46400
rect 26000 40800 30200 46000
rect 26000 39280 27800 40800
rect 26000 38920 26520 39280
rect 26780 38920 27800 39280
rect 26000 38200 27800 38920
rect 28080 39290 28380 39300
rect 28080 38910 28090 39290
rect 28310 39270 28380 39290
rect 28350 38930 28380 39270
rect 28310 38910 28380 38930
rect 28080 38900 28380 38910
rect 26000 25500 26100 38200
rect 27400 25500 27800 38200
rect 26000 23200 27800 25500
rect 26000 16300 26100 23200
rect 27400 16300 27800 23200
rect 26000 15600 27800 16300
rect 26000 14400 26100 15600
rect 27700 14400 27800 15600
rect 26000 14300 27800 14400
rect 28400 38600 30200 38700
rect 28400 37600 28500 38600
rect 29700 37600 30200 38600
rect 28400 24900 30200 37600
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25450 30830 25490
rect 31170 25450 31200 25490
rect 30800 25430 31200 25450
rect 28400 14300 32900 24900
rect 28400 13800 30200 14300
rect 26000 13100 30200 13800
rect 30600 14000 31000 14010
rect 30600 13420 30610 14000
rect 30990 13420 31000 14000
rect 30600 13410 31000 13420
rect 26000 13090 31000 13100
rect 26000 12510 30610 13090
rect 30990 12510 31000 13090
rect 26000 12500 31000 12510
rect 26000 12400 28400 12500
rect 26000 11900 30200 12400
rect 26000 9200 26100 11900
rect 27400 11000 30200 11900
rect 26000 9100 26600 9200
rect 26500 8000 26600 9100
rect 27400 8000 27800 11000
rect 26500 7900 27800 8000
rect 26000 7400 27800 7900
rect 26000 3600 30200 7400
rect 1000 1200 2800 3600
rect 2600 400 2800 1200
rect 1000 200 2800 400
rect 24000 2200 30200 3600
rect 24000 1200 27800 2200
rect 24000 400 25800 1200
rect 27600 400 27800 1200
rect 24000 200 27800 400
<< via4 >>
rect 26100 46500 27300 47500
rect 28110 38930 28310 39270
rect 28310 38930 28350 39270
rect 26100 25500 27400 38200
rect 26100 16300 27400 23200
rect 26100 14400 27700 15600
rect 28500 37600 29700 38600
rect 30830 25490 31170 25690
rect 30830 25450 31170 25490
rect 30630 13440 30970 13980
rect 26100 9200 27400 11900
rect 26600 8000 27400 9200
rect 1000 400 2600 1200
rect 25800 400 27600 1200
<< mimcap2 >>
rect 26100 45800 30100 45900
rect 26100 41000 26200 45800
rect 30000 41000 30100 45800
rect 26100 40900 30100 41000
rect 28500 36900 30100 37000
rect 28500 26700 28600 36900
rect 30000 26700 30100 36900
rect 28500 26600 30100 26700
rect 28500 24700 32800 24800
rect 28500 14500 28600 24700
rect 32700 14500 32800 24700
rect 28500 14400 32800 14500
rect 26100 7200 30100 7300
rect 26100 2400 26200 7200
rect 30000 2400 30100 7200
rect 26100 2300 30100 2400
<< mimcap2contact >>
rect 26200 41000 30000 45800
rect 28600 26700 30000 36900
rect 28600 14500 32700 24700
rect 26200 2400 30000 7200
<< metal5 >>
rect 1300 48100 2800 48500
rect 24000 48100 25500 48500
rect 1000 46700 1300 47600
rect 25500 47500 27400 47600
rect 25500 46700 26100 47500
rect 26000 46500 26100 46700
rect 27300 46500 27400 47500
rect 26000 46400 27400 46500
rect 26000 45800 30200 46000
rect 26000 41000 26200 45800
rect 30000 41000 30200 45800
rect 26000 40800 30200 41000
rect 1000 39700 1200 40200
rect 25400 39270 29800 39300
rect 25400 38930 28110 39270
rect 28350 38930 29800 39270
rect 25400 38800 29800 38930
rect 28400 38600 29800 38800
rect 26000 38200 27500 38300
rect 26000 25500 26100 38200
rect 27400 25500 27500 38200
rect 28400 37600 28500 38600
rect 29700 37600 29800 38600
rect 28400 37500 29800 37600
rect 28400 36900 30200 37100
rect 28400 26700 28600 36900
rect 30000 26700 30200 36900
rect 28400 26500 30200 26700
rect 26000 25400 27500 25500
rect 30800 25690 31200 25720
rect 30800 25450 30830 25690
rect 31170 25450 31200 25690
rect 30800 24900 31200 25450
rect 1000 24700 1200 24900
rect 25400 24700 32900 24900
rect 1000 24000 2100 24700
rect 25400 24600 28600 24700
rect 1000 23800 1200 24000
rect 24500 23900 28600 24600
rect 25400 23800 28600 23900
rect 25400 23500 25600 23800
rect 26000 23200 27500 23300
rect 1000 16500 1300 17900
rect 26000 16300 26100 23200
rect 27400 16300 27500 23200
rect 26000 16200 27500 16300
rect 25500 15600 28000 15700
rect 25500 14400 26100 15600
rect 27700 14400 28000 15600
rect 25500 14300 28000 14400
rect 28400 14500 28600 23800
rect 32700 14500 32900 24700
rect 28400 14300 32900 14500
rect 26800 13800 28000 14300
rect 30600 13980 31000 14300
rect 26800 12500 30200 13800
rect 30600 13440 30630 13980
rect 30970 13440 31000 13980
rect 30600 13410 31000 13440
rect 26000 11900 27500 12000
rect 1000 9100 1200 9600
rect 26000 9200 26100 11900
rect 26000 9100 26600 9200
rect 25400 8200 26100 8700
rect 26500 8000 26600 9100
rect 27400 8000 27500 11900
rect 26500 7900 27500 8000
rect 28400 7400 30200 12500
rect 26000 7200 30200 7400
rect 24000 2200 25400 3600
rect 26000 2400 26200 7200
rect 30000 2400 30200 7200
rect 26000 2200 30200 2400
rect 24000 1700 25500 2200
rect 1000 1200 1400 1400
rect 24000 1200 27800 1400
rect 24000 400 25800 1200
rect 27600 400 27800 1200
rect 1000 200 2800 400
rect 1300 0 2800 200
rect 24000 200 27800 400
rect 24000 0 25500 200
use cascode_1  cascode_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/CLASSE
timestamp 1664506494
transform 1 0 14700 0 1 -3700
box -14700 3700 10800 52200
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_0 ./CLASSE
timestamp 1664814488
transform -1 0 31001 0 1 26369
box -199 -889 199 889
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_4
timestamp 1664814488
transform 0 -1 27431 -1 0 39101
box -199 -889 199 889
use sky130_fd_pr__res_high_po_0p35_FFWWQH  sky130_fd_pr__res_high_po_0p35_FFWWQH_1
timestamp 1664805031
transform -1 0 30799 0 1 13258
box -201 -758 201 758
<< labels >>
rlabel metal5 25800 8200 26100 8700 1 VINP
rlabel metal5 1300 0 2800 400 1 VSS
rlabel metal5 24000 0 25500 400 1 VSSH
rlabel metal5 1300 48100 2800 48500 1 VDN
rlabel metal5 24000 48100 25500 48500 1 VDP
rlabel metal5 900 39700 1200 40200 1 VGN
rlabel metal5 25600 38800 25900 39300 1 VGP
rlabel metal5 900 16500 1200 17900 1 N
rlabel metal5 25600 14300 25900 15700 1 P
rlabel metal3 25600 31000 25800 31800 1 P2
<< end >>
