magic
tech sky130B
magscale 1 2
timestamp 1660708695
<< metal1 >>
rect 1540 9540 2030 9620
rect 1670 9120 1750 9540
rect 1540 9040 2020 9120
rect 1670 8620 1750 9040
rect 1540 8540 2020 8620
rect 1670 8120 1750 8540
rect 1540 8040 2010 8120
rect 1670 7630 1750 8040
rect 0 7580 200 7600
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 10200 7580 10400 7600
rect 10200 7420 10220 7580
rect 10380 7420 10400 7580
rect 10200 7400 10400 7420
rect 0 7100 200 7120
rect 0 6480 200 6500
rect 0 6120 20 6480
rect 180 6120 200 6480
rect 0 6100 200 6120
rect 10200 380 10400 400
rect 10200 220 10220 380
rect 10380 220 10400 380
rect 10200 200 10400 220
<< via1 >>
rect 20 7120 180 7580
rect 10220 7420 10380 7580
rect 20 6120 180 6480
rect 10220 220 10380 380
<< metal2 >>
rect 0 7580 200 7600
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 10200 7580 10400 7600
rect 10200 7420 10220 7580
rect 10380 7420 10400 7580
rect 10200 7400 10400 7420
rect 0 7100 200 7120
rect 0 6480 200 6500
rect 0 6120 20 6480
rect 180 6120 200 6480
rect 0 6100 200 6120
rect 10200 380 10400 400
rect 10200 220 10220 380
rect 10380 220 10400 380
rect 10200 200 10400 220
<< via2 >>
rect 20 7120 180 7580
rect 10220 7420 10380 7580
rect 20 6120 180 6480
rect 10220 220 10380 380
<< metal3 >>
rect -4200 12400 1000 12600
rect -4200 11800 -1400 12400
rect 800 11800 1000 12400
rect -4200 11400 1000 11800
rect 6200 11600 11200 11700
rect -8000 8400 -5000 8600
rect -8000 6000 -7800 8400
rect -5200 7200 -5000 8400
rect -4200 8000 400 11400
rect -1600 7920 400 8000
rect -1600 7740 -1580 7920
rect -20 7740 400 7920
rect -1600 7720 200 7740
rect 0 7580 200 7720
rect 1540 7640 1900 9100
rect 1500 7600 1900 7640
rect 6200 8400 10700 11600
rect 11100 8400 11200 11600
rect 6200 8300 11200 8400
rect -5200 6400 -200 7200
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 0 7100 200 7120
rect 6200 6800 9000 8300
rect 10200 7580 11200 7600
rect 10200 7420 10220 7580
rect 10380 7420 11200 7580
rect 10200 7400 11200 7420
rect 5400 6700 9500 6800
rect -100 6480 200 6500
rect -100 6400 20 6480
rect -5200 6120 20 6400
rect 180 6120 200 6480
rect -5200 6000 200 6120
rect -8000 5800 200 6000
rect -1600 2400 200 5800
rect 5500 939 9000 1100
rect 5800 -400 9000 939
rect 11000 400 11200 7400
rect 10200 380 11200 400
rect 10200 220 10220 380
rect 10380 220 11200 380
rect 10200 200 11200 220
rect 11000 0 11200 200
rect 11000 -200 11600 0
rect 5800 -500 10800 -400
rect 5800 -3700 10300 -500
rect 10700 -3700 10800 -500
rect 5800 -3800 10800 -3700
rect 11400 -5500 11600 -200
<< via3 >>
rect -1400 11800 800 12400
rect -7800 6000 -5200 8400
rect -1580 7740 -20 7920
rect 10700 8400 11100 11600
rect 10300 -3700 10700 -500
<< mimcap >>
rect 6300 11500 10100 11600
rect -4150 11300 350 11350
rect -4150 8300 -4100 11300
rect 300 8300 350 11300
rect 6300 8500 6400 11500
rect 10000 8500 10100 11500
rect 6300 8400 10100 8500
rect -4150 8250 350 8300
rect 5900 -600 9700 -500
rect 5900 -3600 6000 -600
rect 9600 -3600 9700 -600
rect 5900 -3700 9700 -3600
<< mimcapcontact >>
rect -4100 8300 300 11300
rect 6400 8500 10000 11500
rect 6000 -3600 9600 -600
<< metal4 >>
rect -1000 18400 1000 20400
rect -1600 12400 1000 18400
rect -1600 11800 -1400 12400
rect 800 11800 1000 12400
rect -1600 11600 1000 11800
rect 6200 11500 10200 11700
rect 6200 11400 6400 11500
rect -4200 11300 6400 11400
rect -8000 8400 -5000 8600
rect -8000 6000 -7800 8400
rect -5200 6000 -5000 8400
rect -4200 8300 -4100 11300
rect 300 11200 6400 11300
rect 300 10000 2000 11200
rect 300 8300 400 10000
rect -4200 8200 400 8300
rect 1800 8200 2000 10000
rect 4200 8500 6400 11200
rect 10000 8500 10200 11500
rect 4200 8300 10200 8500
rect 10600 11600 11200 11700
rect 10600 8400 10700 11600
rect 11100 8400 11200 11600
rect 10600 8300 11200 8400
rect 4200 8200 4439 8300
rect 1800 8001 4439 8200
rect 1800 8000 4400 8001
rect -1600 7920 0 7940
rect -1600 7740 -1580 7920
rect -20 7740 0 7920
rect -1600 7580 -1560 7740
rect -40 7580 0 7740
rect -1600 7540 0 7580
rect -8000 5800 -5000 6000
rect 10200 1800 17800 6000
rect 3700 -400 4400 400
rect 3700 -600 9800 -400
rect 3700 -3600 6000 -600
rect 9600 -3600 9800 -600
rect 3700 -3800 9800 -3600
rect 10200 -500 10800 -400
rect 10200 -3700 10300 -500
rect 10700 -3700 10800 -500
rect 10200 -3800 10800 -3700
rect 11800 -17800 16400 1800
rect 11800 -41000 12000 -17800
rect 16200 -41000 16400 -17800
rect 11800 -41200 16400 -41000
<< via4 >>
rect -1400 11800 800 12400
rect -7800 6000 -5200 8400
rect 2000 8200 4200 11200
rect 10700 8400 11100 11600
rect -1560 7740 -40 7920
rect -1560 7580 -40 7740
rect 10300 -3700 10700 -500
rect 12000 -41000 16200 -17800
<< mimcap2 >>
rect 6300 11500 10100 11600
rect -4150 11300 350 11350
rect -4150 8300 -4100 11300
rect 300 8300 350 11300
rect 6300 8500 6400 11500
rect 10000 8500 10100 11500
rect 6300 8400 10100 8500
rect -4150 8250 350 8300
rect 5900 -600 9700 -500
rect 5900 -3600 6000 -600
rect 9600 -3600 9700 -600
rect 5900 -3700 9700 -3600
<< mimcap2contact >>
rect -4100 8300 300 11300
rect 6400 8500 10000 11500
rect 6000 -3600 9600 -600
<< metal5 >>
rect -23000 47000 17000 48000
rect -23000 16000 -22000 47000
rect 16000 33000 17000 47000
rect 16000 32000 71000 33000
rect -1000 18400 1000 20400
rect -4200 12400 1000 12600
rect -4200 11800 -1400 12400
rect 800 11800 1000 12400
rect -4200 11400 1000 11800
rect 6200 11600 11200 11700
rect 6200 11500 10700 11600
rect -4200 11300 400 11400
rect -8000 8400 -5000 10600
rect -8000 6000 -7800 8400
rect -5200 6000 -5000 8400
rect -4200 8300 -4100 11300
rect 300 8300 400 11300
rect -4200 8000 400 8300
rect 1800 11200 4400 11400
rect 1800 8200 2000 11200
rect 4200 8200 4400 11200
rect 6200 8500 6400 11500
rect 10000 8500 10700 11500
rect 6200 8400 10700 8500
rect 11100 8400 11200 11600
rect 6200 8300 11200 8400
rect 1800 8100 4400 8200
rect -3550 7500 -3100 8000
rect -1600 7920 0 8000
rect -1600 7580 -1560 7920
rect -40 7580 0 7920
rect 1800 7600 5900 8100
rect -1600 7540 0 7580
rect -8000 5800 -5000 6000
rect 27100 1900 31100 5850
rect 70000 5000 71000 32000
rect 5800 -500 10800 -400
rect 5800 -600 10300 -500
rect 5800 -3600 6000 -600
rect 9600 -3600 10300 -600
rect 5800 -3700 10300 -3600
rect 10700 -3700 10800 -500
rect 5800 -3800 10800 -3700
rect 66000 -9000 71000 5000
rect 64000 -11000 71000 -9000
rect 11800 -17800 16400 -17600
rect 7000 -42000 8000 -26000
rect 11800 -41000 12000 -17800
rect 16200 -41000 16400 -17800
rect 70000 -26000 71000 -11000
rect 11800 -41200 16400 -41000
rect 20000 -27000 71000 -26000
rect 20000 -42000 21000 -27000
use PA_core_1  PA_core_1_0
timestamp 1660307541
transform 0 -1 10000 1 0 700
box -700 -500 7196 10000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501637
transform 1 0 1900 0 1 7640
box 0 0 4000 4000
use nfet_diode_1  nfet_diode_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660705385
transform 1 0 40 0 1 0
box 340 7600 1560 9660
use sky130_fd_pr__res_high_po_0p35_ZE2H5K  sky130_fd_pr__res_high_po_0p35_ZE2H5K_0
timestamp 1660277336
transform 1 0 101 0 1 6798
box -201 -898 201 898
<< labels >>
rlabel metal5 -8000 8700 -5000 10600 1 INPUT
rlabel metal4 16400 1800 17800 6000 1 OUTPUT
rlabel metal5 1800 10000 4400 11400 1 GND
rlabel space -3560 7500 -3100 8000 1 IREF_L
rlabel metal5 9800 -2400 10800 -400 1 VGATE_CAS
rlabel metal5 10200 9700 11200 11700 1 VGATE_CAS
<< end >>
