magic
tech sky130A
magscale 1 2
timestamp 1665068237
<< pwell >>
rect -3400 38680 -3002 40458
rect 1300 39700 6438 46216
rect 7600 39700 12738 46216
rect 13900 39700 19038 46216
rect 20200 39700 25338 46216
rect 1300 32700 6438 39216
rect 7600 32700 12738 39216
rect 13900 32700 19038 39216
rect 20200 32700 25338 39216
rect 29802 38680 30200 40458
rect -4400 25480 -4002 27258
rect 1300 24400 6438 30916
rect 7600 24400 12738 30916
rect 13900 24400 19038 30916
rect 20200 24400 25338 30916
rect 30802 25480 31200 27258
rect 1300 17400 6438 23916
rect 7600 17400 12738 23916
rect 13900 17400 19038 23916
rect 20200 17400 25338 23916
rect -4400 12500 -3998 14016
rect 1300 9100 6438 15616
rect 7600 9100 12738 15616
rect 13900 9100 19038 15616
rect 20200 9100 25338 15616
rect 30798 12500 31200 14016
rect 1300 2100 6438 8616
rect 7600 2100 12738 8616
rect 13900 2100 19038 8616
rect 20200 2100 25338 8616
<< mvnmos >>
rect 1528 39958 1628 45958
rect 1686 39958 1786 45958
rect 1844 39958 1944 45958
rect 2002 39958 2102 45958
rect 2160 39958 2260 45958
rect 2318 39958 2418 45958
rect 2476 39958 2576 45958
rect 2634 39958 2734 45958
rect 2792 39958 2892 45958
rect 2950 39958 3050 45958
rect 3108 39958 3208 45958
rect 3266 39958 3366 45958
rect 3424 39958 3524 45958
rect 3582 39958 3682 45958
rect 3740 39958 3840 45958
rect 3898 39958 3998 45958
rect 4056 39958 4156 45958
rect 4214 39958 4314 45958
rect 4372 39958 4472 45958
rect 4530 39958 4630 45958
rect 4688 39958 4788 45958
rect 4846 39958 4946 45958
rect 5004 39958 5104 45958
rect 5162 39958 5262 45958
rect 5320 39958 5420 45958
rect 5478 39958 5578 45958
rect 5636 39958 5736 45958
rect 5794 39958 5894 45958
rect 5952 39958 6052 45958
rect 6110 39958 6210 45958
rect 7828 39958 7928 45958
rect 7986 39958 8086 45958
rect 8144 39958 8244 45958
rect 8302 39958 8402 45958
rect 8460 39958 8560 45958
rect 8618 39958 8718 45958
rect 8776 39958 8876 45958
rect 8934 39958 9034 45958
rect 9092 39958 9192 45958
rect 9250 39958 9350 45958
rect 9408 39958 9508 45958
rect 9566 39958 9666 45958
rect 9724 39958 9824 45958
rect 9882 39958 9982 45958
rect 10040 39958 10140 45958
rect 10198 39958 10298 45958
rect 10356 39958 10456 45958
rect 10514 39958 10614 45958
rect 10672 39958 10772 45958
rect 10830 39958 10930 45958
rect 10988 39958 11088 45958
rect 11146 39958 11246 45958
rect 11304 39958 11404 45958
rect 11462 39958 11562 45958
rect 11620 39958 11720 45958
rect 11778 39958 11878 45958
rect 11936 39958 12036 45958
rect 12094 39958 12194 45958
rect 12252 39958 12352 45958
rect 12410 39958 12510 45958
rect 14128 39958 14228 45958
rect 14286 39958 14386 45958
rect 14444 39958 14544 45958
rect 14602 39958 14702 45958
rect 14760 39958 14860 45958
rect 14918 39958 15018 45958
rect 15076 39958 15176 45958
rect 15234 39958 15334 45958
rect 15392 39958 15492 45958
rect 15550 39958 15650 45958
rect 15708 39958 15808 45958
rect 15866 39958 15966 45958
rect 16024 39958 16124 45958
rect 16182 39958 16282 45958
rect 16340 39958 16440 45958
rect 16498 39958 16598 45958
rect 16656 39958 16756 45958
rect 16814 39958 16914 45958
rect 16972 39958 17072 45958
rect 17130 39958 17230 45958
rect 17288 39958 17388 45958
rect 17446 39958 17546 45958
rect 17604 39958 17704 45958
rect 17762 39958 17862 45958
rect 17920 39958 18020 45958
rect 18078 39958 18178 45958
rect 18236 39958 18336 45958
rect 18394 39958 18494 45958
rect 18552 39958 18652 45958
rect 18710 39958 18810 45958
rect 20428 39958 20528 45958
rect 20586 39958 20686 45958
rect 20744 39958 20844 45958
rect 20902 39958 21002 45958
rect 21060 39958 21160 45958
rect 21218 39958 21318 45958
rect 21376 39958 21476 45958
rect 21534 39958 21634 45958
rect 21692 39958 21792 45958
rect 21850 39958 21950 45958
rect 22008 39958 22108 45958
rect 22166 39958 22266 45958
rect 22324 39958 22424 45958
rect 22482 39958 22582 45958
rect 22640 39958 22740 45958
rect 22798 39958 22898 45958
rect 22956 39958 23056 45958
rect 23114 39958 23214 45958
rect 23272 39958 23372 45958
rect 23430 39958 23530 45958
rect 23588 39958 23688 45958
rect 23746 39958 23846 45958
rect 23904 39958 24004 45958
rect 24062 39958 24162 45958
rect 24220 39958 24320 45958
rect 24378 39958 24478 45958
rect 24536 39958 24636 45958
rect 24694 39958 24794 45958
rect 24852 39958 24952 45958
rect 25010 39958 25110 45958
rect 1528 32958 1628 38958
rect 1686 32958 1786 38958
rect 1844 32958 1944 38958
rect 2002 32958 2102 38958
rect 2160 32958 2260 38958
rect 2318 32958 2418 38958
rect 2476 32958 2576 38958
rect 2634 32958 2734 38958
rect 2792 32958 2892 38958
rect 2950 32958 3050 38958
rect 3108 32958 3208 38958
rect 3266 32958 3366 38958
rect 3424 32958 3524 38958
rect 3582 32958 3682 38958
rect 3740 32958 3840 38958
rect 3898 32958 3998 38958
rect 4056 32958 4156 38958
rect 4214 32958 4314 38958
rect 4372 32958 4472 38958
rect 4530 32958 4630 38958
rect 4688 32958 4788 38958
rect 4846 32958 4946 38958
rect 5004 32958 5104 38958
rect 5162 32958 5262 38958
rect 5320 32958 5420 38958
rect 5478 32958 5578 38958
rect 5636 32958 5736 38958
rect 5794 32958 5894 38958
rect 5952 32958 6052 38958
rect 6110 32958 6210 38958
rect 7828 32958 7928 38958
rect 7986 32958 8086 38958
rect 8144 32958 8244 38958
rect 8302 32958 8402 38958
rect 8460 32958 8560 38958
rect 8618 32958 8718 38958
rect 8776 32958 8876 38958
rect 8934 32958 9034 38958
rect 9092 32958 9192 38958
rect 9250 32958 9350 38958
rect 9408 32958 9508 38958
rect 9566 32958 9666 38958
rect 9724 32958 9824 38958
rect 9882 32958 9982 38958
rect 10040 32958 10140 38958
rect 10198 32958 10298 38958
rect 10356 32958 10456 38958
rect 10514 32958 10614 38958
rect 10672 32958 10772 38958
rect 10830 32958 10930 38958
rect 10988 32958 11088 38958
rect 11146 32958 11246 38958
rect 11304 32958 11404 38958
rect 11462 32958 11562 38958
rect 11620 32958 11720 38958
rect 11778 32958 11878 38958
rect 11936 32958 12036 38958
rect 12094 32958 12194 38958
rect 12252 32958 12352 38958
rect 12410 32958 12510 38958
rect 14128 32958 14228 38958
rect 14286 32958 14386 38958
rect 14444 32958 14544 38958
rect 14602 32958 14702 38958
rect 14760 32958 14860 38958
rect 14918 32958 15018 38958
rect 15076 32958 15176 38958
rect 15234 32958 15334 38958
rect 15392 32958 15492 38958
rect 15550 32958 15650 38958
rect 15708 32958 15808 38958
rect 15866 32958 15966 38958
rect 16024 32958 16124 38958
rect 16182 32958 16282 38958
rect 16340 32958 16440 38958
rect 16498 32958 16598 38958
rect 16656 32958 16756 38958
rect 16814 32958 16914 38958
rect 16972 32958 17072 38958
rect 17130 32958 17230 38958
rect 17288 32958 17388 38958
rect 17446 32958 17546 38958
rect 17604 32958 17704 38958
rect 17762 32958 17862 38958
rect 17920 32958 18020 38958
rect 18078 32958 18178 38958
rect 18236 32958 18336 38958
rect 18394 32958 18494 38958
rect 18552 32958 18652 38958
rect 18710 32958 18810 38958
rect 20428 32958 20528 38958
rect 20586 32958 20686 38958
rect 20744 32958 20844 38958
rect 20902 32958 21002 38958
rect 21060 32958 21160 38958
rect 21218 32958 21318 38958
rect 21376 32958 21476 38958
rect 21534 32958 21634 38958
rect 21692 32958 21792 38958
rect 21850 32958 21950 38958
rect 22008 32958 22108 38958
rect 22166 32958 22266 38958
rect 22324 32958 22424 38958
rect 22482 32958 22582 38958
rect 22640 32958 22740 38958
rect 22798 32958 22898 38958
rect 22956 32958 23056 38958
rect 23114 32958 23214 38958
rect 23272 32958 23372 38958
rect 23430 32958 23530 38958
rect 23588 32958 23688 38958
rect 23746 32958 23846 38958
rect 23904 32958 24004 38958
rect 24062 32958 24162 38958
rect 24220 32958 24320 38958
rect 24378 32958 24478 38958
rect 24536 32958 24636 38958
rect 24694 32958 24794 38958
rect 24852 32958 24952 38958
rect 25010 32958 25110 38958
rect 1528 24658 1628 30658
rect 1686 24658 1786 30658
rect 1844 24658 1944 30658
rect 2002 24658 2102 30658
rect 2160 24658 2260 30658
rect 2318 24658 2418 30658
rect 2476 24658 2576 30658
rect 2634 24658 2734 30658
rect 2792 24658 2892 30658
rect 2950 24658 3050 30658
rect 3108 24658 3208 30658
rect 3266 24658 3366 30658
rect 3424 24658 3524 30658
rect 3582 24658 3682 30658
rect 3740 24658 3840 30658
rect 3898 24658 3998 30658
rect 4056 24658 4156 30658
rect 4214 24658 4314 30658
rect 4372 24658 4472 30658
rect 4530 24658 4630 30658
rect 4688 24658 4788 30658
rect 4846 24658 4946 30658
rect 5004 24658 5104 30658
rect 5162 24658 5262 30658
rect 5320 24658 5420 30658
rect 5478 24658 5578 30658
rect 5636 24658 5736 30658
rect 5794 24658 5894 30658
rect 5952 24658 6052 30658
rect 6110 24658 6210 30658
rect 7828 24658 7928 30658
rect 7986 24658 8086 30658
rect 8144 24658 8244 30658
rect 8302 24658 8402 30658
rect 8460 24658 8560 30658
rect 8618 24658 8718 30658
rect 8776 24658 8876 30658
rect 8934 24658 9034 30658
rect 9092 24658 9192 30658
rect 9250 24658 9350 30658
rect 9408 24658 9508 30658
rect 9566 24658 9666 30658
rect 9724 24658 9824 30658
rect 9882 24658 9982 30658
rect 10040 24658 10140 30658
rect 10198 24658 10298 30658
rect 10356 24658 10456 30658
rect 10514 24658 10614 30658
rect 10672 24658 10772 30658
rect 10830 24658 10930 30658
rect 10988 24658 11088 30658
rect 11146 24658 11246 30658
rect 11304 24658 11404 30658
rect 11462 24658 11562 30658
rect 11620 24658 11720 30658
rect 11778 24658 11878 30658
rect 11936 24658 12036 30658
rect 12094 24658 12194 30658
rect 12252 24658 12352 30658
rect 12410 24658 12510 30658
rect 14128 24658 14228 30658
rect 14286 24658 14386 30658
rect 14444 24658 14544 30658
rect 14602 24658 14702 30658
rect 14760 24658 14860 30658
rect 14918 24658 15018 30658
rect 15076 24658 15176 30658
rect 15234 24658 15334 30658
rect 15392 24658 15492 30658
rect 15550 24658 15650 30658
rect 15708 24658 15808 30658
rect 15866 24658 15966 30658
rect 16024 24658 16124 30658
rect 16182 24658 16282 30658
rect 16340 24658 16440 30658
rect 16498 24658 16598 30658
rect 16656 24658 16756 30658
rect 16814 24658 16914 30658
rect 16972 24658 17072 30658
rect 17130 24658 17230 30658
rect 17288 24658 17388 30658
rect 17446 24658 17546 30658
rect 17604 24658 17704 30658
rect 17762 24658 17862 30658
rect 17920 24658 18020 30658
rect 18078 24658 18178 30658
rect 18236 24658 18336 30658
rect 18394 24658 18494 30658
rect 18552 24658 18652 30658
rect 18710 24658 18810 30658
rect 20428 24658 20528 30658
rect 20586 24658 20686 30658
rect 20744 24658 20844 30658
rect 20902 24658 21002 30658
rect 21060 24658 21160 30658
rect 21218 24658 21318 30658
rect 21376 24658 21476 30658
rect 21534 24658 21634 30658
rect 21692 24658 21792 30658
rect 21850 24658 21950 30658
rect 22008 24658 22108 30658
rect 22166 24658 22266 30658
rect 22324 24658 22424 30658
rect 22482 24658 22582 30658
rect 22640 24658 22740 30658
rect 22798 24658 22898 30658
rect 22956 24658 23056 30658
rect 23114 24658 23214 30658
rect 23272 24658 23372 30658
rect 23430 24658 23530 30658
rect 23588 24658 23688 30658
rect 23746 24658 23846 30658
rect 23904 24658 24004 30658
rect 24062 24658 24162 30658
rect 24220 24658 24320 30658
rect 24378 24658 24478 30658
rect 24536 24658 24636 30658
rect 24694 24658 24794 30658
rect 24852 24658 24952 30658
rect 25010 24658 25110 30658
rect 1528 17658 1628 23658
rect 1686 17658 1786 23658
rect 1844 17658 1944 23658
rect 2002 17658 2102 23658
rect 2160 17658 2260 23658
rect 2318 17658 2418 23658
rect 2476 17658 2576 23658
rect 2634 17658 2734 23658
rect 2792 17658 2892 23658
rect 2950 17658 3050 23658
rect 3108 17658 3208 23658
rect 3266 17658 3366 23658
rect 3424 17658 3524 23658
rect 3582 17658 3682 23658
rect 3740 17658 3840 23658
rect 3898 17658 3998 23658
rect 4056 17658 4156 23658
rect 4214 17658 4314 23658
rect 4372 17658 4472 23658
rect 4530 17658 4630 23658
rect 4688 17658 4788 23658
rect 4846 17658 4946 23658
rect 5004 17658 5104 23658
rect 5162 17658 5262 23658
rect 5320 17658 5420 23658
rect 5478 17658 5578 23658
rect 5636 17658 5736 23658
rect 5794 17658 5894 23658
rect 5952 17658 6052 23658
rect 6110 17658 6210 23658
rect 7828 17658 7928 23658
rect 7986 17658 8086 23658
rect 8144 17658 8244 23658
rect 8302 17658 8402 23658
rect 8460 17658 8560 23658
rect 8618 17658 8718 23658
rect 8776 17658 8876 23658
rect 8934 17658 9034 23658
rect 9092 17658 9192 23658
rect 9250 17658 9350 23658
rect 9408 17658 9508 23658
rect 9566 17658 9666 23658
rect 9724 17658 9824 23658
rect 9882 17658 9982 23658
rect 10040 17658 10140 23658
rect 10198 17658 10298 23658
rect 10356 17658 10456 23658
rect 10514 17658 10614 23658
rect 10672 17658 10772 23658
rect 10830 17658 10930 23658
rect 10988 17658 11088 23658
rect 11146 17658 11246 23658
rect 11304 17658 11404 23658
rect 11462 17658 11562 23658
rect 11620 17658 11720 23658
rect 11778 17658 11878 23658
rect 11936 17658 12036 23658
rect 12094 17658 12194 23658
rect 12252 17658 12352 23658
rect 12410 17658 12510 23658
rect 14128 17658 14228 23658
rect 14286 17658 14386 23658
rect 14444 17658 14544 23658
rect 14602 17658 14702 23658
rect 14760 17658 14860 23658
rect 14918 17658 15018 23658
rect 15076 17658 15176 23658
rect 15234 17658 15334 23658
rect 15392 17658 15492 23658
rect 15550 17658 15650 23658
rect 15708 17658 15808 23658
rect 15866 17658 15966 23658
rect 16024 17658 16124 23658
rect 16182 17658 16282 23658
rect 16340 17658 16440 23658
rect 16498 17658 16598 23658
rect 16656 17658 16756 23658
rect 16814 17658 16914 23658
rect 16972 17658 17072 23658
rect 17130 17658 17230 23658
rect 17288 17658 17388 23658
rect 17446 17658 17546 23658
rect 17604 17658 17704 23658
rect 17762 17658 17862 23658
rect 17920 17658 18020 23658
rect 18078 17658 18178 23658
rect 18236 17658 18336 23658
rect 18394 17658 18494 23658
rect 18552 17658 18652 23658
rect 18710 17658 18810 23658
rect 20428 17658 20528 23658
rect 20586 17658 20686 23658
rect 20744 17658 20844 23658
rect 20902 17658 21002 23658
rect 21060 17658 21160 23658
rect 21218 17658 21318 23658
rect 21376 17658 21476 23658
rect 21534 17658 21634 23658
rect 21692 17658 21792 23658
rect 21850 17658 21950 23658
rect 22008 17658 22108 23658
rect 22166 17658 22266 23658
rect 22324 17658 22424 23658
rect 22482 17658 22582 23658
rect 22640 17658 22740 23658
rect 22798 17658 22898 23658
rect 22956 17658 23056 23658
rect 23114 17658 23214 23658
rect 23272 17658 23372 23658
rect 23430 17658 23530 23658
rect 23588 17658 23688 23658
rect 23746 17658 23846 23658
rect 23904 17658 24004 23658
rect 24062 17658 24162 23658
rect 24220 17658 24320 23658
rect 24378 17658 24478 23658
rect 24536 17658 24636 23658
rect 24694 17658 24794 23658
rect 24852 17658 24952 23658
rect 25010 17658 25110 23658
rect 1528 9358 1628 15358
rect 1686 9358 1786 15358
rect 1844 9358 1944 15358
rect 2002 9358 2102 15358
rect 2160 9358 2260 15358
rect 2318 9358 2418 15358
rect 2476 9358 2576 15358
rect 2634 9358 2734 15358
rect 2792 9358 2892 15358
rect 2950 9358 3050 15358
rect 3108 9358 3208 15358
rect 3266 9358 3366 15358
rect 3424 9358 3524 15358
rect 3582 9358 3682 15358
rect 3740 9358 3840 15358
rect 3898 9358 3998 15358
rect 4056 9358 4156 15358
rect 4214 9358 4314 15358
rect 4372 9358 4472 15358
rect 4530 9358 4630 15358
rect 4688 9358 4788 15358
rect 4846 9358 4946 15358
rect 5004 9358 5104 15358
rect 5162 9358 5262 15358
rect 5320 9358 5420 15358
rect 5478 9358 5578 15358
rect 5636 9358 5736 15358
rect 5794 9358 5894 15358
rect 5952 9358 6052 15358
rect 6110 9358 6210 15358
rect 7828 9358 7928 15358
rect 7986 9358 8086 15358
rect 8144 9358 8244 15358
rect 8302 9358 8402 15358
rect 8460 9358 8560 15358
rect 8618 9358 8718 15358
rect 8776 9358 8876 15358
rect 8934 9358 9034 15358
rect 9092 9358 9192 15358
rect 9250 9358 9350 15358
rect 9408 9358 9508 15358
rect 9566 9358 9666 15358
rect 9724 9358 9824 15358
rect 9882 9358 9982 15358
rect 10040 9358 10140 15358
rect 10198 9358 10298 15358
rect 10356 9358 10456 15358
rect 10514 9358 10614 15358
rect 10672 9358 10772 15358
rect 10830 9358 10930 15358
rect 10988 9358 11088 15358
rect 11146 9358 11246 15358
rect 11304 9358 11404 15358
rect 11462 9358 11562 15358
rect 11620 9358 11720 15358
rect 11778 9358 11878 15358
rect 11936 9358 12036 15358
rect 12094 9358 12194 15358
rect 12252 9358 12352 15358
rect 12410 9358 12510 15358
rect 14128 9358 14228 15358
rect 14286 9358 14386 15358
rect 14444 9358 14544 15358
rect 14602 9358 14702 15358
rect 14760 9358 14860 15358
rect 14918 9358 15018 15358
rect 15076 9358 15176 15358
rect 15234 9358 15334 15358
rect 15392 9358 15492 15358
rect 15550 9358 15650 15358
rect 15708 9358 15808 15358
rect 15866 9358 15966 15358
rect 16024 9358 16124 15358
rect 16182 9358 16282 15358
rect 16340 9358 16440 15358
rect 16498 9358 16598 15358
rect 16656 9358 16756 15358
rect 16814 9358 16914 15358
rect 16972 9358 17072 15358
rect 17130 9358 17230 15358
rect 17288 9358 17388 15358
rect 17446 9358 17546 15358
rect 17604 9358 17704 15358
rect 17762 9358 17862 15358
rect 17920 9358 18020 15358
rect 18078 9358 18178 15358
rect 18236 9358 18336 15358
rect 18394 9358 18494 15358
rect 18552 9358 18652 15358
rect 18710 9358 18810 15358
rect 20428 9358 20528 15358
rect 20586 9358 20686 15358
rect 20744 9358 20844 15358
rect 20902 9358 21002 15358
rect 21060 9358 21160 15358
rect 21218 9358 21318 15358
rect 21376 9358 21476 15358
rect 21534 9358 21634 15358
rect 21692 9358 21792 15358
rect 21850 9358 21950 15358
rect 22008 9358 22108 15358
rect 22166 9358 22266 15358
rect 22324 9358 22424 15358
rect 22482 9358 22582 15358
rect 22640 9358 22740 15358
rect 22798 9358 22898 15358
rect 22956 9358 23056 15358
rect 23114 9358 23214 15358
rect 23272 9358 23372 15358
rect 23430 9358 23530 15358
rect 23588 9358 23688 15358
rect 23746 9358 23846 15358
rect 23904 9358 24004 15358
rect 24062 9358 24162 15358
rect 24220 9358 24320 15358
rect 24378 9358 24478 15358
rect 24536 9358 24636 15358
rect 24694 9358 24794 15358
rect 24852 9358 24952 15358
rect 25010 9358 25110 15358
rect 1528 2358 1628 8358
rect 1686 2358 1786 8358
rect 1844 2358 1944 8358
rect 2002 2358 2102 8358
rect 2160 2358 2260 8358
rect 2318 2358 2418 8358
rect 2476 2358 2576 8358
rect 2634 2358 2734 8358
rect 2792 2358 2892 8358
rect 2950 2358 3050 8358
rect 3108 2358 3208 8358
rect 3266 2358 3366 8358
rect 3424 2358 3524 8358
rect 3582 2358 3682 8358
rect 3740 2358 3840 8358
rect 3898 2358 3998 8358
rect 4056 2358 4156 8358
rect 4214 2358 4314 8358
rect 4372 2358 4472 8358
rect 4530 2358 4630 8358
rect 4688 2358 4788 8358
rect 4846 2358 4946 8358
rect 5004 2358 5104 8358
rect 5162 2358 5262 8358
rect 5320 2358 5420 8358
rect 5478 2358 5578 8358
rect 5636 2358 5736 8358
rect 5794 2358 5894 8358
rect 5952 2358 6052 8358
rect 6110 2358 6210 8358
rect 7828 2358 7928 8358
rect 7986 2358 8086 8358
rect 8144 2358 8244 8358
rect 8302 2358 8402 8358
rect 8460 2358 8560 8358
rect 8618 2358 8718 8358
rect 8776 2358 8876 8358
rect 8934 2358 9034 8358
rect 9092 2358 9192 8358
rect 9250 2358 9350 8358
rect 9408 2358 9508 8358
rect 9566 2358 9666 8358
rect 9724 2358 9824 8358
rect 9882 2358 9982 8358
rect 10040 2358 10140 8358
rect 10198 2358 10298 8358
rect 10356 2358 10456 8358
rect 10514 2358 10614 8358
rect 10672 2358 10772 8358
rect 10830 2358 10930 8358
rect 10988 2358 11088 8358
rect 11146 2358 11246 8358
rect 11304 2358 11404 8358
rect 11462 2358 11562 8358
rect 11620 2358 11720 8358
rect 11778 2358 11878 8358
rect 11936 2358 12036 8358
rect 12094 2358 12194 8358
rect 12252 2358 12352 8358
rect 12410 2358 12510 8358
rect 14128 2358 14228 8358
rect 14286 2358 14386 8358
rect 14444 2358 14544 8358
rect 14602 2358 14702 8358
rect 14760 2358 14860 8358
rect 14918 2358 15018 8358
rect 15076 2358 15176 8358
rect 15234 2358 15334 8358
rect 15392 2358 15492 8358
rect 15550 2358 15650 8358
rect 15708 2358 15808 8358
rect 15866 2358 15966 8358
rect 16024 2358 16124 8358
rect 16182 2358 16282 8358
rect 16340 2358 16440 8358
rect 16498 2358 16598 8358
rect 16656 2358 16756 8358
rect 16814 2358 16914 8358
rect 16972 2358 17072 8358
rect 17130 2358 17230 8358
rect 17288 2358 17388 8358
rect 17446 2358 17546 8358
rect 17604 2358 17704 8358
rect 17762 2358 17862 8358
rect 17920 2358 18020 8358
rect 18078 2358 18178 8358
rect 18236 2358 18336 8358
rect 18394 2358 18494 8358
rect 18552 2358 18652 8358
rect 18710 2358 18810 8358
rect 20428 2358 20528 8358
rect 20586 2358 20686 8358
rect 20744 2358 20844 8358
rect 20902 2358 21002 8358
rect 21060 2358 21160 8358
rect 21218 2358 21318 8358
rect 21376 2358 21476 8358
rect 21534 2358 21634 8358
rect 21692 2358 21792 8358
rect 21850 2358 21950 8358
rect 22008 2358 22108 8358
rect 22166 2358 22266 8358
rect 22324 2358 22424 8358
rect 22482 2358 22582 8358
rect 22640 2358 22740 8358
rect 22798 2358 22898 8358
rect 22956 2358 23056 8358
rect 23114 2358 23214 8358
rect 23272 2358 23372 8358
rect 23430 2358 23530 8358
rect 23588 2358 23688 8358
rect 23746 2358 23846 8358
rect 23904 2358 24004 8358
rect 24062 2358 24162 8358
rect 24220 2358 24320 8358
rect 24378 2358 24478 8358
rect 24536 2358 24636 8358
rect 24694 2358 24794 8358
rect 24852 2358 24952 8358
rect 25010 2358 25110 8358
<< mvndiff >>
rect 1470 45946 1528 45958
rect 1470 39970 1482 45946
rect 1516 39970 1528 45946
rect 1470 39958 1528 39970
rect 1628 45946 1686 45958
rect 1628 39970 1640 45946
rect 1674 39970 1686 45946
rect 1628 39958 1686 39970
rect 1786 45946 1844 45958
rect 1786 39970 1798 45946
rect 1832 39970 1844 45946
rect 1786 39958 1844 39970
rect 1944 45946 2002 45958
rect 1944 39970 1956 45946
rect 1990 39970 2002 45946
rect 1944 39958 2002 39970
rect 2102 45946 2160 45958
rect 2102 39970 2114 45946
rect 2148 39970 2160 45946
rect 2102 39958 2160 39970
rect 2260 45946 2318 45958
rect 2260 39970 2272 45946
rect 2306 39970 2318 45946
rect 2260 39958 2318 39970
rect 2418 45946 2476 45958
rect 2418 39970 2430 45946
rect 2464 39970 2476 45946
rect 2418 39958 2476 39970
rect 2576 45946 2634 45958
rect 2576 39970 2588 45946
rect 2622 39970 2634 45946
rect 2576 39958 2634 39970
rect 2734 45946 2792 45958
rect 2734 39970 2746 45946
rect 2780 39970 2792 45946
rect 2734 39958 2792 39970
rect 2892 45946 2950 45958
rect 2892 39970 2904 45946
rect 2938 39970 2950 45946
rect 2892 39958 2950 39970
rect 3050 45946 3108 45958
rect 3050 39970 3062 45946
rect 3096 39970 3108 45946
rect 3050 39958 3108 39970
rect 3208 45946 3266 45958
rect 3208 39970 3220 45946
rect 3254 39970 3266 45946
rect 3208 39958 3266 39970
rect 3366 45946 3424 45958
rect 3366 39970 3378 45946
rect 3412 39970 3424 45946
rect 3366 39958 3424 39970
rect 3524 45946 3582 45958
rect 3524 39970 3536 45946
rect 3570 39970 3582 45946
rect 3524 39958 3582 39970
rect 3682 45946 3740 45958
rect 3682 39970 3694 45946
rect 3728 39970 3740 45946
rect 3682 39958 3740 39970
rect 3840 45946 3898 45958
rect 3840 39970 3852 45946
rect 3886 39970 3898 45946
rect 3840 39958 3898 39970
rect 3998 45946 4056 45958
rect 3998 39970 4010 45946
rect 4044 39970 4056 45946
rect 3998 39958 4056 39970
rect 4156 45946 4214 45958
rect 4156 39970 4168 45946
rect 4202 39970 4214 45946
rect 4156 39958 4214 39970
rect 4314 45946 4372 45958
rect 4314 39970 4326 45946
rect 4360 39970 4372 45946
rect 4314 39958 4372 39970
rect 4472 45946 4530 45958
rect 4472 39970 4484 45946
rect 4518 39970 4530 45946
rect 4472 39958 4530 39970
rect 4630 45946 4688 45958
rect 4630 39970 4642 45946
rect 4676 39970 4688 45946
rect 4630 39958 4688 39970
rect 4788 45946 4846 45958
rect 4788 39970 4800 45946
rect 4834 39970 4846 45946
rect 4788 39958 4846 39970
rect 4946 45946 5004 45958
rect 4946 39970 4958 45946
rect 4992 39970 5004 45946
rect 4946 39958 5004 39970
rect 5104 45946 5162 45958
rect 5104 39970 5116 45946
rect 5150 39970 5162 45946
rect 5104 39958 5162 39970
rect 5262 45946 5320 45958
rect 5262 39970 5274 45946
rect 5308 39970 5320 45946
rect 5262 39958 5320 39970
rect 5420 45946 5478 45958
rect 5420 39970 5432 45946
rect 5466 39970 5478 45946
rect 5420 39958 5478 39970
rect 5578 45946 5636 45958
rect 5578 39970 5590 45946
rect 5624 39970 5636 45946
rect 5578 39958 5636 39970
rect 5736 45946 5794 45958
rect 5736 39970 5748 45946
rect 5782 39970 5794 45946
rect 5736 39958 5794 39970
rect 5894 45946 5952 45958
rect 5894 39970 5906 45946
rect 5940 39970 5952 45946
rect 5894 39958 5952 39970
rect 6052 45946 6110 45958
rect 6052 39970 6064 45946
rect 6098 39970 6110 45946
rect 6052 39958 6110 39970
rect 6210 45946 6268 45958
rect 6210 39970 6222 45946
rect 6256 39970 6268 45946
rect 6210 39958 6268 39970
rect 7770 45946 7828 45958
rect 7770 39970 7782 45946
rect 7816 39970 7828 45946
rect 7770 39958 7828 39970
rect 7928 45946 7986 45958
rect 7928 39970 7940 45946
rect 7974 39970 7986 45946
rect 7928 39958 7986 39970
rect 8086 45946 8144 45958
rect 8086 39970 8098 45946
rect 8132 39970 8144 45946
rect 8086 39958 8144 39970
rect 8244 45946 8302 45958
rect 8244 39970 8256 45946
rect 8290 39970 8302 45946
rect 8244 39958 8302 39970
rect 8402 45946 8460 45958
rect 8402 39970 8414 45946
rect 8448 39970 8460 45946
rect 8402 39958 8460 39970
rect 8560 45946 8618 45958
rect 8560 39970 8572 45946
rect 8606 39970 8618 45946
rect 8560 39958 8618 39970
rect 8718 45946 8776 45958
rect 8718 39970 8730 45946
rect 8764 39970 8776 45946
rect 8718 39958 8776 39970
rect 8876 45946 8934 45958
rect 8876 39970 8888 45946
rect 8922 39970 8934 45946
rect 8876 39958 8934 39970
rect 9034 45946 9092 45958
rect 9034 39970 9046 45946
rect 9080 39970 9092 45946
rect 9034 39958 9092 39970
rect 9192 45946 9250 45958
rect 9192 39970 9204 45946
rect 9238 39970 9250 45946
rect 9192 39958 9250 39970
rect 9350 45946 9408 45958
rect 9350 39970 9362 45946
rect 9396 39970 9408 45946
rect 9350 39958 9408 39970
rect 9508 45946 9566 45958
rect 9508 39970 9520 45946
rect 9554 39970 9566 45946
rect 9508 39958 9566 39970
rect 9666 45946 9724 45958
rect 9666 39970 9678 45946
rect 9712 39970 9724 45946
rect 9666 39958 9724 39970
rect 9824 45946 9882 45958
rect 9824 39970 9836 45946
rect 9870 39970 9882 45946
rect 9824 39958 9882 39970
rect 9982 45946 10040 45958
rect 9982 39970 9994 45946
rect 10028 39970 10040 45946
rect 9982 39958 10040 39970
rect 10140 45946 10198 45958
rect 10140 39970 10152 45946
rect 10186 39970 10198 45946
rect 10140 39958 10198 39970
rect 10298 45946 10356 45958
rect 10298 39970 10310 45946
rect 10344 39970 10356 45946
rect 10298 39958 10356 39970
rect 10456 45946 10514 45958
rect 10456 39970 10468 45946
rect 10502 39970 10514 45946
rect 10456 39958 10514 39970
rect 10614 45946 10672 45958
rect 10614 39970 10626 45946
rect 10660 39970 10672 45946
rect 10614 39958 10672 39970
rect 10772 45946 10830 45958
rect 10772 39970 10784 45946
rect 10818 39970 10830 45946
rect 10772 39958 10830 39970
rect 10930 45946 10988 45958
rect 10930 39970 10942 45946
rect 10976 39970 10988 45946
rect 10930 39958 10988 39970
rect 11088 45946 11146 45958
rect 11088 39970 11100 45946
rect 11134 39970 11146 45946
rect 11088 39958 11146 39970
rect 11246 45946 11304 45958
rect 11246 39970 11258 45946
rect 11292 39970 11304 45946
rect 11246 39958 11304 39970
rect 11404 45946 11462 45958
rect 11404 39970 11416 45946
rect 11450 39970 11462 45946
rect 11404 39958 11462 39970
rect 11562 45946 11620 45958
rect 11562 39970 11574 45946
rect 11608 39970 11620 45946
rect 11562 39958 11620 39970
rect 11720 45946 11778 45958
rect 11720 39970 11732 45946
rect 11766 39970 11778 45946
rect 11720 39958 11778 39970
rect 11878 45946 11936 45958
rect 11878 39970 11890 45946
rect 11924 39970 11936 45946
rect 11878 39958 11936 39970
rect 12036 45946 12094 45958
rect 12036 39970 12048 45946
rect 12082 39970 12094 45946
rect 12036 39958 12094 39970
rect 12194 45946 12252 45958
rect 12194 39970 12206 45946
rect 12240 39970 12252 45946
rect 12194 39958 12252 39970
rect 12352 45946 12410 45958
rect 12352 39970 12364 45946
rect 12398 39970 12410 45946
rect 12352 39958 12410 39970
rect 12510 45946 12568 45958
rect 12510 39970 12522 45946
rect 12556 39970 12568 45946
rect 12510 39958 12568 39970
rect 14070 45946 14128 45958
rect 14070 39970 14082 45946
rect 14116 39970 14128 45946
rect 14070 39958 14128 39970
rect 14228 45946 14286 45958
rect 14228 39970 14240 45946
rect 14274 39970 14286 45946
rect 14228 39958 14286 39970
rect 14386 45946 14444 45958
rect 14386 39970 14398 45946
rect 14432 39970 14444 45946
rect 14386 39958 14444 39970
rect 14544 45946 14602 45958
rect 14544 39970 14556 45946
rect 14590 39970 14602 45946
rect 14544 39958 14602 39970
rect 14702 45946 14760 45958
rect 14702 39970 14714 45946
rect 14748 39970 14760 45946
rect 14702 39958 14760 39970
rect 14860 45946 14918 45958
rect 14860 39970 14872 45946
rect 14906 39970 14918 45946
rect 14860 39958 14918 39970
rect 15018 45946 15076 45958
rect 15018 39970 15030 45946
rect 15064 39970 15076 45946
rect 15018 39958 15076 39970
rect 15176 45946 15234 45958
rect 15176 39970 15188 45946
rect 15222 39970 15234 45946
rect 15176 39958 15234 39970
rect 15334 45946 15392 45958
rect 15334 39970 15346 45946
rect 15380 39970 15392 45946
rect 15334 39958 15392 39970
rect 15492 45946 15550 45958
rect 15492 39970 15504 45946
rect 15538 39970 15550 45946
rect 15492 39958 15550 39970
rect 15650 45946 15708 45958
rect 15650 39970 15662 45946
rect 15696 39970 15708 45946
rect 15650 39958 15708 39970
rect 15808 45946 15866 45958
rect 15808 39970 15820 45946
rect 15854 39970 15866 45946
rect 15808 39958 15866 39970
rect 15966 45946 16024 45958
rect 15966 39970 15978 45946
rect 16012 39970 16024 45946
rect 15966 39958 16024 39970
rect 16124 45946 16182 45958
rect 16124 39970 16136 45946
rect 16170 39970 16182 45946
rect 16124 39958 16182 39970
rect 16282 45946 16340 45958
rect 16282 39970 16294 45946
rect 16328 39970 16340 45946
rect 16282 39958 16340 39970
rect 16440 45946 16498 45958
rect 16440 39970 16452 45946
rect 16486 39970 16498 45946
rect 16440 39958 16498 39970
rect 16598 45946 16656 45958
rect 16598 39970 16610 45946
rect 16644 39970 16656 45946
rect 16598 39958 16656 39970
rect 16756 45946 16814 45958
rect 16756 39970 16768 45946
rect 16802 39970 16814 45946
rect 16756 39958 16814 39970
rect 16914 45946 16972 45958
rect 16914 39970 16926 45946
rect 16960 39970 16972 45946
rect 16914 39958 16972 39970
rect 17072 45946 17130 45958
rect 17072 39970 17084 45946
rect 17118 39970 17130 45946
rect 17072 39958 17130 39970
rect 17230 45946 17288 45958
rect 17230 39970 17242 45946
rect 17276 39970 17288 45946
rect 17230 39958 17288 39970
rect 17388 45946 17446 45958
rect 17388 39970 17400 45946
rect 17434 39970 17446 45946
rect 17388 39958 17446 39970
rect 17546 45946 17604 45958
rect 17546 39970 17558 45946
rect 17592 39970 17604 45946
rect 17546 39958 17604 39970
rect 17704 45946 17762 45958
rect 17704 39970 17716 45946
rect 17750 39970 17762 45946
rect 17704 39958 17762 39970
rect 17862 45946 17920 45958
rect 17862 39970 17874 45946
rect 17908 39970 17920 45946
rect 17862 39958 17920 39970
rect 18020 45946 18078 45958
rect 18020 39970 18032 45946
rect 18066 39970 18078 45946
rect 18020 39958 18078 39970
rect 18178 45946 18236 45958
rect 18178 39970 18190 45946
rect 18224 39970 18236 45946
rect 18178 39958 18236 39970
rect 18336 45946 18394 45958
rect 18336 39970 18348 45946
rect 18382 39970 18394 45946
rect 18336 39958 18394 39970
rect 18494 45946 18552 45958
rect 18494 39970 18506 45946
rect 18540 39970 18552 45946
rect 18494 39958 18552 39970
rect 18652 45946 18710 45958
rect 18652 39970 18664 45946
rect 18698 39970 18710 45946
rect 18652 39958 18710 39970
rect 18810 45946 18868 45958
rect 18810 39970 18822 45946
rect 18856 39970 18868 45946
rect 18810 39958 18868 39970
rect 20370 45946 20428 45958
rect 20370 39970 20382 45946
rect 20416 39970 20428 45946
rect 20370 39958 20428 39970
rect 20528 45946 20586 45958
rect 20528 39970 20540 45946
rect 20574 39970 20586 45946
rect 20528 39958 20586 39970
rect 20686 45946 20744 45958
rect 20686 39970 20698 45946
rect 20732 39970 20744 45946
rect 20686 39958 20744 39970
rect 20844 45946 20902 45958
rect 20844 39970 20856 45946
rect 20890 39970 20902 45946
rect 20844 39958 20902 39970
rect 21002 45946 21060 45958
rect 21002 39970 21014 45946
rect 21048 39970 21060 45946
rect 21002 39958 21060 39970
rect 21160 45946 21218 45958
rect 21160 39970 21172 45946
rect 21206 39970 21218 45946
rect 21160 39958 21218 39970
rect 21318 45946 21376 45958
rect 21318 39970 21330 45946
rect 21364 39970 21376 45946
rect 21318 39958 21376 39970
rect 21476 45946 21534 45958
rect 21476 39970 21488 45946
rect 21522 39970 21534 45946
rect 21476 39958 21534 39970
rect 21634 45946 21692 45958
rect 21634 39970 21646 45946
rect 21680 39970 21692 45946
rect 21634 39958 21692 39970
rect 21792 45946 21850 45958
rect 21792 39970 21804 45946
rect 21838 39970 21850 45946
rect 21792 39958 21850 39970
rect 21950 45946 22008 45958
rect 21950 39970 21962 45946
rect 21996 39970 22008 45946
rect 21950 39958 22008 39970
rect 22108 45946 22166 45958
rect 22108 39970 22120 45946
rect 22154 39970 22166 45946
rect 22108 39958 22166 39970
rect 22266 45946 22324 45958
rect 22266 39970 22278 45946
rect 22312 39970 22324 45946
rect 22266 39958 22324 39970
rect 22424 45946 22482 45958
rect 22424 39970 22436 45946
rect 22470 39970 22482 45946
rect 22424 39958 22482 39970
rect 22582 45946 22640 45958
rect 22582 39970 22594 45946
rect 22628 39970 22640 45946
rect 22582 39958 22640 39970
rect 22740 45946 22798 45958
rect 22740 39970 22752 45946
rect 22786 39970 22798 45946
rect 22740 39958 22798 39970
rect 22898 45946 22956 45958
rect 22898 39970 22910 45946
rect 22944 39970 22956 45946
rect 22898 39958 22956 39970
rect 23056 45946 23114 45958
rect 23056 39970 23068 45946
rect 23102 39970 23114 45946
rect 23056 39958 23114 39970
rect 23214 45946 23272 45958
rect 23214 39970 23226 45946
rect 23260 39970 23272 45946
rect 23214 39958 23272 39970
rect 23372 45946 23430 45958
rect 23372 39970 23384 45946
rect 23418 39970 23430 45946
rect 23372 39958 23430 39970
rect 23530 45946 23588 45958
rect 23530 39970 23542 45946
rect 23576 39970 23588 45946
rect 23530 39958 23588 39970
rect 23688 45946 23746 45958
rect 23688 39970 23700 45946
rect 23734 39970 23746 45946
rect 23688 39958 23746 39970
rect 23846 45946 23904 45958
rect 23846 39970 23858 45946
rect 23892 39970 23904 45946
rect 23846 39958 23904 39970
rect 24004 45946 24062 45958
rect 24004 39970 24016 45946
rect 24050 39970 24062 45946
rect 24004 39958 24062 39970
rect 24162 45946 24220 45958
rect 24162 39970 24174 45946
rect 24208 39970 24220 45946
rect 24162 39958 24220 39970
rect 24320 45946 24378 45958
rect 24320 39970 24332 45946
rect 24366 39970 24378 45946
rect 24320 39958 24378 39970
rect 24478 45946 24536 45958
rect 24478 39970 24490 45946
rect 24524 39970 24536 45946
rect 24478 39958 24536 39970
rect 24636 45946 24694 45958
rect 24636 39970 24648 45946
rect 24682 39970 24694 45946
rect 24636 39958 24694 39970
rect 24794 45946 24852 45958
rect 24794 39970 24806 45946
rect 24840 39970 24852 45946
rect 24794 39958 24852 39970
rect 24952 45946 25010 45958
rect 24952 39970 24964 45946
rect 24998 39970 25010 45946
rect 24952 39958 25010 39970
rect 25110 45946 25168 45958
rect 25110 39970 25122 45946
rect 25156 39970 25168 45946
rect 25110 39958 25168 39970
rect 1470 38946 1528 38958
rect 1470 32970 1482 38946
rect 1516 32970 1528 38946
rect 1470 32958 1528 32970
rect 1628 38946 1686 38958
rect 1628 32970 1640 38946
rect 1674 32970 1686 38946
rect 1628 32958 1686 32970
rect 1786 38946 1844 38958
rect 1786 32970 1798 38946
rect 1832 32970 1844 38946
rect 1786 32958 1844 32970
rect 1944 38946 2002 38958
rect 1944 32970 1956 38946
rect 1990 32970 2002 38946
rect 1944 32958 2002 32970
rect 2102 38946 2160 38958
rect 2102 32970 2114 38946
rect 2148 32970 2160 38946
rect 2102 32958 2160 32970
rect 2260 38946 2318 38958
rect 2260 32970 2272 38946
rect 2306 32970 2318 38946
rect 2260 32958 2318 32970
rect 2418 38946 2476 38958
rect 2418 32970 2430 38946
rect 2464 32970 2476 38946
rect 2418 32958 2476 32970
rect 2576 38946 2634 38958
rect 2576 32970 2588 38946
rect 2622 32970 2634 38946
rect 2576 32958 2634 32970
rect 2734 38946 2792 38958
rect 2734 32970 2746 38946
rect 2780 32970 2792 38946
rect 2734 32958 2792 32970
rect 2892 38946 2950 38958
rect 2892 32970 2904 38946
rect 2938 32970 2950 38946
rect 2892 32958 2950 32970
rect 3050 38946 3108 38958
rect 3050 32970 3062 38946
rect 3096 32970 3108 38946
rect 3050 32958 3108 32970
rect 3208 38946 3266 38958
rect 3208 32970 3220 38946
rect 3254 32970 3266 38946
rect 3208 32958 3266 32970
rect 3366 38946 3424 38958
rect 3366 32970 3378 38946
rect 3412 32970 3424 38946
rect 3366 32958 3424 32970
rect 3524 38946 3582 38958
rect 3524 32970 3536 38946
rect 3570 32970 3582 38946
rect 3524 32958 3582 32970
rect 3682 38946 3740 38958
rect 3682 32970 3694 38946
rect 3728 32970 3740 38946
rect 3682 32958 3740 32970
rect 3840 38946 3898 38958
rect 3840 32970 3852 38946
rect 3886 32970 3898 38946
rect 3840 32958 3898 32970
rect 3998 38946 4056 38958
rect 3998 32970 4010 38946
rect 4044 32970 4056 38946
rect 3998 32958 4056 32970
rect 4156 38946 4214 38958
rect 4156 32970 4168 38946
rect 4202 32970 4214 38946
rect 4156 32958 4214 32970
rect 4314 38946 4372 38958
rect 4314 32970 4326 38946
rect 4360 32970 4372 38946
rect 4314 32958 4372 32970
rect 4472 38946 4530 38958
rect 4472 32970 4484 38946
rect 4518 32970 4530 38946
rect 4472 32958 4530 32970
rect 4630 38946 4688 38958
rect 4630 32970 4642 38946
rect 4676 32970 4688 38946
rect 4630 32958 4688 32970
rect 4788 38946 4846 38958
rect 4788 32970 4800 38946
rect 4834 32970 4846 38946
rect 4788 32958 4846 32970
rect 4946 38946 5004 38958
rect 4946 32970 4958 38946
rect 4992 32970 5004 38946
rect 4946 32958 5004 32970
rect 5104 38946 5162 38958
rect 5104 32970 5116 38946
rect 5150 32970 5162 38946
rect 5104 32958 5162 32970
rect 5262 38946 5320 38958
rect 5262 32970 5274 38946
rect 5308 32970 5320 38946
rect 5262 32958 5320 32970
rect 5420 38946 5478 38958
rect 5420 32970 5432 38946
rect 5466 32970 5478 38946
rect 5420 32958 5478 32970
rect 5578 38946 5636 38958
rect 5578 32970 5590 38946
rect 5624 32970 5636 38946
rect 5578 32958 5636 32970
rect 5736 38946 5794 38958
rect 5736 32970 5748 38946
rect 5782 32970 5794 38946
rect 5736 32958 5794 32970
rect 5894 38946 5952 38958
rect 5894 32970 5906 38946
rect 5940 32970 5952 38946
rect 5894 32958 5952 32970
rect 6052 38946 6110 38958
rect 6052 32970 6064 38946
rect 6098 32970 6110 38946
rect 6052 32958 6110 32970
rect 6210 38946 6268 38958
rect 6210 32970 6222 38946
rect 6256 32970 6268 38946
rect 6210 32958 6268 32970
rect 7770 38946 7828 38958
rect 7770 32970 7782 38946
rect 7816 32970 7828 38946
rect 7770 32958 7828 32970
rect 7928 38946 7986 38958
rect 7928 32970 7940 38946
rect 7974 32970 7986 38946
rect 7928 32958 7986 32970
rect 8086 38946 8144 38958
rect 8086 32970 8098 38946
rect 8132 32970 8144 38946
rect 8086 32958 8144 32970
rect 8244 38946 8302 38958
rect 8244 32970 8256 38946
rect 8290 32970 8302 38946
rect 8244 32958 8302 32970
rect 8402 38946 8460 38958
rect 8402 32970 8414 38946
rect 8448 32970 8460 38946
rect 8402 32958 8460 32970
rect 8560 38946 8618 38958
rect 8560 32970 8572 38946
rect 8606 32970 8618 38946
rect 8560 32958 8618 32970
rect 8718 38946 8776 38958
rect 8718 32970 8730 38946
rect 8764 32970 8776 38946
rect 8718 32958 8776 32970
rect 8876 38946 8934 38958
rect 8876 32970 8888 38946
rect 8922 32970 8934 38946
rect 8876 32958 8934 32970
rect 9034 38946 9092 38958
rect 9034 32970 9046 38946
rect 9080 32970 9092 38946
rect 9034 32958 9092 32970
rect 9192 38946 9250 38958
rect 9192 32970 9204 38946
rect 9238 32970 9250 38946
rect 9192 32958 9250 32970
rect 9350 38946 9408 38958
rect 9350 32970 9362 38946
rect 9396 32970 9408 38946
rect 9350 32958 9408 32970
rect 9508 38946 9566 38958
rect 9508 32970 9520 38946
rect 9554 32970 9566 38946
rect 9508 32958 9566 32970
rect 9666 38946 9724 38958
rect 9666 32970 9678 38946
rect 9712 32970 9724 38946
rect 9666 32958 9724 32970
rect 9824 38946 9882 38958
rect 9824 32970 9836 38946
rect 9870 32970 9882 38946
rect 9824 32958 9882 32970
rect 9982 38946 10040 38958
rect 9982 32970 9994 38946
rect 10028 32970 10040 38946
rect 9982 32958 10040 32970
rect 10140 38946 10198 38958
rect 10140 32970 10152 38946
rect 10186 32970 10198 38946
rect 10140 32958 10198 32970
rect 10298 38946 10356 38958
rect 10298 32970 10310 38946
rect 10344 32970 10356 38946
rect 10298 32958 10356 32970
rect 10456 38946 10514 38958
rect 10456 32970 10468 38946
rect 10502 32970 10514 38946
rect 10456 32958 10514 32970
rect 10614 38946 10672 38958
rect 10614 32970 10626 38946
rect 10660 32970 10672 38946
rect 10614 32958 10672 32970
rect 10772 38946 10830 38958
rect 10772 32970 10784 38946
rect 10818 32970 10830 38946
rect 10772 32958 10830 32970
rect 10930 38946 10988 38958
rect 10930 32970 10942 38946
rect 10976 32970 10988 38946
rect 10930 32958 10988 32970
rect 11088 38946 11146 38958
rect 11088 32970 11100 38946
rect 11134 32970 11146 38946
rect 11088 32958 11146 32970
rect 11246 38946 11304 38958
rect 11246 32970 11258 38946
rect 11292 32970 11304 38946
rect 11246 32958 11304 32970
rect 11404 38946 11462 38958
rect 11404 32970 11416 38946
rect 11450 32970 11462 38946
rect 11404 32958 11462 32970
rect 11562 38946 11620 38958
rect 11562 32970 11574 38946
rect 11608 32970 11620 38946
rect 11562 32958 11620 32970
rect 11720 38946 11778 38958
rect 11720 32970 11732 38946
rect 11766 32970 11778 38946
rect 11720 32958 11778 32970
rect 11878 38946 11936 38958
rect 11878 32970 11890 38946
rect 11924 32970 11936 38946
rect 11878 32958 11936 32970
rect 12036 38946 12094 38958
rect 12036 32970 12048 38946
rect 12082 32970 12094 38946
rect 12036 32958 12094 32970
rect 12194 38946 12252 38958
rect 12194 32970 12206 38946
rect 12240 32970 12252 38946
rect 12194 32958 12252 32970
rect 12352 38946 12410 38958
rect 12352 32970 12364 38946
rect 12398 32970 12410 38946
rect 12352 32958 12410 32970
rect 12510 38946 12568 38958
rect 12510 32970 12522 38946
rect 12556 32970 12568 38946
rect 12510 32958 12568 32970
rect 14070 38946 14128 38958
rect 14070 32970 14082 38946
rect 14116 32970 14128 38946
rect 14070 32958 14128 32970
rect 14228 38946 14286 38958
rect 14228 32970 14240 38946
rect 14274 32970 14286 38946
rect 14228 32958 14286 32970
rect 14386 38946 14444 38958
rect 14386 32970 14398 38946
rect 14432 32970 14444 38946
rect 14386 32958 14444 32970
rect 14544 38946 14602 38958
rect 14544 32970 14556 38946
rect 14590 32970 14602 38946
rect 14544 32958 14602 32970
rect 14702 38946 14760 38958
rect 14702 32970 14714 38946
rect 14748 32970 14760 38946
rect 14702 32958 14760 32970
rect 14860 38946 14918 38958
rect 14860 32970 14872 38946
rect 14906 32970 14918 38946
rect 14860 32958 14918 32970
rect 15018 38946 15076 38958
rect 15018 32970 15030 38946
rect 15064 32970 15076 38946
rect 15018 32958 15076 32970
rect 15176 38946 15234 38958
rect 15176 32970 15188 38946
rect 15222 32970 15234 38946
rect 15176 32958 15234 32970
rect 15334 38946 15392 38958
rect 15334 32970 15346 38946
rect 15380 32970 15392 38946
rect 15334 32958 15392 32970
rect 15492 38946 15550 38958
rect 15492 32970 15504 38946
rect 15538 32970 15550 38946
rect 15492 32958 15550 32970
rect 15650 38946 15708 38958
rect 15650 32970 15662 38946
rect 15696 32970 15708 38946
rect 15650 32958 15708 32970
rect 15808 38946 15866 38958
rect 15808 32970 15820 38946
rect 15854 32970 15866 38946
rect 15808 32958 15866 32970
rect 15966 38946 16024 38958
rect 15966 32970 15978 38946
rect 16012 32970 16024 38946
rect 15966 32958 16024 32970
rect 16124 38946 16182 38958
rect 16124 32970 16136 38946
rect 16170 32970 16182 38946
rect 16124 32958 16182 32970
rect 16282 38946 16340 38958
rect 16282 32970 16294 38946
rect 16328 32970 16340 38946
rect 16282 32958 16340 32970
rect 16440 38946 16498 38958
rect 16440 32970 16452 38946
rect 16486 32970 16498 38946
rect 16440 32958 16498 32970
rect 16598 38946 16656 38958
rect 16598 32970 16610 38946
rect 16644 32970 16656 38946
rect 16598 32958 16656 32970
rect 16756 38946 16814 38958
rect 16756 32970 16768 38946
rect 16802 32970 16814 38946
rect 16756 32958 16814 32970
rect 16914 38946 16972 38958
rect 16914 32970 16926 38946
rect 16960 32970 16972 38946
rect 16914 32958 16972 32970
rect 17072 38946 17130 38958
rect 17072 32970 17084 38946
rect 17118 32970 17130 38946
rect 17072 32958 17130 32970
rect 17230 38946 17288 38958
rect 17230 32970 17242 38946
rect 17276 32970 17288 38946
rect 17230 32958 17288 32970
rect 17388 38946 17446 38958
rect 17388 32970 17400 38946
rect 17434 32970 17446 38946
rect 17388 32958 17446 32970
rect 17546 38946 17604 38958
rect 17546 32970 17558 38946
rect 17592 32970 17604 38946
rect 17546 32958 17604 32970
rect 17704 38946 17762 38958
rect 17704 32970 17716 38946
rect 17750 32970 17762 38946
rect 17704 32958 17762 32970
rect 17862 38946 17920 38958
rect 17862 32970 17874 38946
rect 17908 32970 17920 38946
rect 17862 32958 17920 32970
rect 18020 38946 18078 38958
rect 18020 32970 18032 38946
rect 18066 32970 18078 38946
rect 18020 32958 18078 32970
rect 18178 38946 18236 38958
rect 18178 32970 18190 38946
rect 18224 32970 18236 38946
rect 18178 32958 18236 32970
rect 18336 38946 18394 38958
rect 18336 32970 18348 38946
rect 18382 32970 18394 38946
rect 18336 32958 18394 32970
rect 18494 38946 18552 38958
rect 18494 32970 18506 38946
rect 18540 32970 18552 38946
rect 18494 32958 18552 32970
rect 18652 38946 18710 38958
rect 18652 32970 18664 38946
rect 18698 32970 18710 38946
rect 18652 32958 18710 32970
rect 18810 38946 18868 38958
rect 18810 32970 18822 38946
rect 18856 32970 18868 38946
rect 18810 32958 18868 32970
rect 20370 38946 20428 38958
rect 20370 32970 20382 38946
rect 20416 32970 20428 38946
rect 20370 32958 20428 32970
rect 20528 38946 20586 38958
rect 20528 32970 20540 38946
rect 20574 32970 20586 38946
rect 20528 32958 20586 32970
rect 20686 38946 20744 38958
rect 20686 32970 20698 38946
rect 20732 32970 20744 38946
rect 20686 32958 20744 32970
rect 20844 38946 20902 38958
rect 20844 32970 20856 38946
rect 20890 32970 20902 38946
rect 20844 32958 20902 32970
rect 21002 38946 21060 38958
rect 21002 32970 21014 38946
rect 21048 32970 21060 38946
rect 21002 32958 21060 32970
rect 21160 38946 21218 38958
rect 21160 32970 21172 38946
rect 21206 32970 21218 38946
rect 21160 32958 21218 32970
rect 21318 38946 21376 38958
rect 21318 32970 21330 38946
rect 21364 32970 21376 38946
rect 21318 32958 21376 32970
rect 21476 38946 21534 38958
rect 21476 32970 21488 38946
rect 21522 32970 21534 38946
rect 21476 32958 21534 32970
rect 21634 38946 21692 38958
rect 21634 32970 21646 38946
rect 21680 32970 21692 38946
rect 21634 32958 21692 32970
rect 21792 38946 21850 38958
rect 21792 32970 21804 38946
rect 21838 32970 21850 38946
rect 21792 32958 21850 32970
rect 21950 38946 22008 38958
rect 21950 32970 21962 38946
rect 21996 32970 22008 38946
rect 21950 32958 22008 32970
rect 22108 38946 22166 38958
rect 22108 32970 22120 38946
rect 22154 32970 22166 38946
rect 22108 32958 22166 32970
rect 22266 38946 22324 38958
rect 22266 32970 22278 38946
rect 22312 32970 22324 38946
rect 22266 32958 22324 32970
rect 22424 38946 22482 38958
rect 22424 32970 22436 38946
rect 22470 32970 22482 38946
rect 22424 32958 22482 32970
rect 22582 38946 22640 38958
rect 22582 32970 22594 38946
rect 22628 32970 22640 38946
rect 22582 32958 22640 32970
rect 22740 38946 22798 38958
rect 22740 32970 22752 38946
rect 22786 32970 22798 38946
rect 22740 32958 22798 32970
rect 22898 38946 22956 38958
rect 22898 32970 22910 38946
rect 22944 32970 22956 38946
rect 22898 32958 22956 32970
rect 23056 38946 23114 38958
rect 23056 32970 23068 38946
rect 23102 32970 23114 38946
rect 23056 32958 23114 32970
rect 23214 38946 23272 38958
rect 23214 32970 23226 38946
rect 23260 32970 23272 38946
rect 23214 32958 23272 32970
rect 23372 38946 23430 38958
rect 23372 32970 23384 38946
rect 23418 32970 23430 38946
rect 23372 32958 23430 32970
rect 23530 38946 23588 38958
rect 23530 32970 23542 38946
rect 23576 32970 23588 38946
rect 23530 32958 23588 32970
rect 23688 38946 23746 38958
rect 23688 32970 23700 38946
rect 23734 32970 23746 38946
rect 23688 32958 23746 32970
rect 23846 38946 23904 38958
rect 23846 32970 23858 38946
rect 23892 32970 23904 38946
rect 23846 32958 23904 32970
rect 24004 38946 24062 38958
rect 24004 32970 24016 38946
rect 24050 32970 24062 38946
rect 24004 32958 24062 32970
rect 24162 38946 24220 38958
rect 24162 32970 24174 38946
rect 24208 32970 24220 38946
rect 24162 32958 24220 32970
rect 24320 38946 24378 38958
rect 24320 32970 24332 38946
rect 24366 32970 24378 38946
rect 24320 32958 24378 32970
rect 24478 38946 24536 38958
rect 24478 32970 24490 38946
rect 24524 32970 24536 38946
rect 24478 32958 24536 32970
rect 24636 38946 24694 38958
rect 24636 32970 24648 38946
rect 24682 32970 24694 38946
rect 24636 32958 24694 32970
rect 24794 38946 24852 38958
rect 24794 32970 24806 38946
rect 24840 32970 24852 38946
rect 24794 32958 24852 32970
rect 24952 38946 25010 38958
rect 24952 32970 24964 38946
rect 24998 32970 25010 38946
rect 24952 32958 25010 32970
rect 25110 38946 25168 38958
rect 25110 32970 25122 38946
rect 25156 32970 25168 38946
rect 25110 32958 25168 32970
rect 1470 30646 1528 30658
rect 1470 24670 1482 30646
rect 1516 24670 1528 30646
rect 1470 24658 1528 24670
rect 1628 30646 1686 30658
rect 1628 24670 1640 30646
rect 1674 24670 1686 30646
rect 1628 24658 1686 24670
rect 1786 30646 1844 30658
rect 1786 24670 1798 30646
rect 1832 24670 1844 30646
rect 1786 24658 1844 24670
rect 1944 30646 2002 30658
rect 1944 24670 1956 30646
rect 1990 24670 2002 30646
rect 1944 24658 2002 24670
rect 2102 30646 2160 30658
rect 2102 24670 2114 30646
rect 2148 24670 2160 30646
rect 2102 24658 2160 24670
rect 2260 30646 2318 30658
rect 2260 24670 2272 30646
rect 2306 24670 2318 30646
rect 2260 24658 2318 24670
rect 2418 30646 2476 30658
rect 2418 24670 2430 30646
rect 2464 24670 2476 30646
rect 2418 24658 2476 24670
rect 2576 30646 2634 30658
rect 2576 24670 2588 30646
rect 2622 24670 2634 30646
rect 2576 24658 2634 24670
rect 2734 30646 2792 30658
rect 2734 24670 2746 30646
rect 2780 24670 2792 30646
rect 2734 24658 2792 24670
rect 2892 30646 2950 30658
rect 2892 24670 2904 30646
rect 2938 24670 2950 30646
rect 2892 24658 2950 24670
rect 3050 30646 3108 30658
rect 3050 24670 3062 30646
rect 3096 24670 3108 30646
rect 3050 24658 3108 24670
rect 3208 30646 3266 30658
rect 3208 24670 3220 30646
rect 3254 24670 3266 30646
rect 3208 24658 3266 24670
rect 3366 30646 3424 30658
rect 3366 24670 3378 30646
rect 3412 24670 3424 30646
rect 3366 24658 3424 24670
rect 3524 30646 3582 30658
rect 3524 24670 3536 30646
rect 3570 24670 3582 30646
rect 3524 24658 3582 24670
rect 3682 30646 3740 30658
rect 3682 24670 3694 30646
rect 3728 24670 3740 30646
rect 3682 24658 3740 24670
rect 3840 30646 3898 30658
rect 3840 24670 3852 30646
rect 3886 24670 3898 30646
rect 3840 24658 3898 24670
rect 3998 30646 4056 30658
rect 3998 24670 4010 30646
rect 4044 24670 4056 30646
rect 3998 24658 4056 24670
rect 4156 30646 4214 30658
rect 4156 24670 4168 30646
rect 4202 24670 4214 30646
rect 4156 24658 4214 24670
rect 4314 30646 4372 30658
rect 4314 24670 4326 30646
rect 4360 24670 4372 30646
rect 4314 24658 4372 24670
rect 4472 30646 4530 30658
rect 4472 24670 4484 30646
rect 4518 24670 4530 30646
rect 4472 24658 4530 24670
rect 4630 30646 4688 30658
rect 4630 24670 4642 30646
rect 4676 24670 4688 30646
rect 4630 24658 4688 24670
rect 4788 30646 4846 30658
rect 4788 24670 4800 30646
rect 4834 24670 4846 30646
rect 4788 24658 4846 24670
rect 4946 30646 5004 30658
rect 4946 24670 4958 30646
rect 4992 24670 5004 30646
rect 4946 24658 5004 24670
rect 5104 30646 5162 30658
rect 5104 24670 5116 30646
rect 5150 24670 5162 30646
rect 5104 24658 5162 24670
rect 5262 30646 5320 30658
rect 5262 24670 5274 30646
rect 5308 24670 5320 30646
rect 5262 24658 5320 24670
rect 5420 30646 5478 30658
rect 5420 24670 5432 30646
rect 5466 24670 5478 30646
rect 5420 24658 5478 24670
rect 5578 30646 5636 30658
rect 5578 24670 5590 30646
rect 5624 24670 5636 30646
rect 5578 24658 5636 24670
rect 5736 30646 5794 30658
rect 5736 24670 5748 30646
rect 5782 24670 5794 30646
rect 5736 24658 5794 24670
rect 5894 30646 5952 30658
rect 5894 24670 5906 30646
rect 5940 24670 5952 30646
rect 5894 24658 5952 24670
rect 6052 30646 6110 30658
rect 6052 24670 6064 30646
rect 6098 24670 6110 30646
rect 6052 24658 6110 24670
rect 6210 30646 6268 30658
rect 6210 24670 6222 30646
rect 6256 24670 6268 30646
rect 6210 24658 6268 24670
rect 7770 30646 7828 30658
rect 7770 24670 7782 30646
rect 7816 24670 7828 30646
rect 7770 24658 7828 24670
rect 7928 30646 7986 30658
rect 7928 24670 7940 30646
rect 7974 24670 7986 30646
rect 7928 24658 7986 24670
rect 8086 30646 8144 30658
rect 8086 24670 8098 30646
rect 8132 24670 8144 30646
rect 8086 24658 8144 24670
rect 8244 30646 8302 30658
rect 8244 24670 8256 30646
rect 8290 24670 8302 30646
rect 8244 24658 8302 24670
rect 8402 30646 8460 30658
rect 8402 24670 8414 30646
rect 8448 24670 8460 30646
rect 8402 24658 8460 24670
rect 8560 30646 8618 30658
rect 8560 24670 8572 30646
rect 8606 24670 8618 30646
rect 8560 24658 8618 24670
rect 8718 30646 8776 30658
rect 8718 24670 8730 30646
rect 8764 24670 8776 30646
rect 8718 24658 8776 24670
rect 8876 30646 8934 30658
rect 8876 24670 8888 30646
rect 8922 24670 8934 30646
rect 8876 24658 8934 24670
rect 9034 30646 9092 30658
rect 9034 24670 9046 30646
rect 9080 24670 9092 30646
rect 9034 24658 9092 24670
rect 9192 30646 9250 30658
rect 9192 24670 9204 30646
rect 9238 24670 9250 30646
rect 9192 24658 9250 24670
rect 9350 30646 9408 30658
rect 9350 24670 9362 30646
rect 9396 24670 9408 30646
rect 9350 24658 9408 24670
rect 9508 30646 9566 30658
rect 9508 24670 9520 30646
rect 9554 24670 9566 30646
rect 9508 24658 9566 24670
rect 9666 30646 9724 30658
rect 9666 24670 9678 30646
rect 9712 24670 9724 30646
rect 9666 24658 9724 24670
rect 9824 30646 9882 30658
rect 9824 24670 9836 30646
rect 9870 24670 9882 30646
rect 9824 24658 9882 24670
rect 9982 30646 10040 30658
rect 9982 24670 9994 30646
rect 10028 24670 10040 30646
rect 9982 24658 10040 24670
rect 10140 30646 10198 30658
rect 10140 24670 10152 30646
rect 10186 24670 10198 30646
rect 10140 24658 10198 24670
rect 10298 30646 10356 30658
rect 10298 24670 10310 30646
rect 10344 24670 10356 30646
rect 10298 24658 10356 24670
rect 10456 30646 10514 30658
rect 10456 24670 10468 30646
rect 10502 24670 10514 30646
rect 10456 24658 10514 24670
rect 10614 30646 10672 30658
rect 10614 24670 10626 30646
rect 10660 24670 10672 30646
rect 10614 24658 10672 24670
rect 10772 30646 10830 30658
rect 10772 24670 10784 30646
rect 10818 24670 10830 30646
rect 10772 24658 10830 24670
rect 10930 30646 10988 30658
rect 10930 24670 10942 30646
rect 10976 24670 10988 30646
rect 10930 24658 10988 24670
rect 11088 30646 11146 30658
rect 11088 24670 11100 30646
rect 11134 24670 11146 30646
rect 11088 24658 11146 24670
rect 11246 30646 11304 30658
rect 11246 24670 11258 30646
rect 11292 24670 11304 30646
rect 11246 24658 11304 24670
rect 11404 30646 11462 30658
rect 11404 24670 11416 30646
rect 11450 24670 11462 30646
rect 11404 24658 11462 24670
rect 11562 30646 11620 30658
rect 11562 24670 11574 30646
rect 11608 24670 11620 30646
rect 11562 24658 11620 24670
rect 11720 30646 11778 30658
rect 11720 24670 11732 30646
rect 11766 24670 11778 30646
rect 11720 24658 11778 24670
rect 11878 30646 11936 30658
rect 11878 24670 11890 30646
rect 11924 24670 11936 30646
rect 11878 24658 11936 24670
rect 12036 30646 12094 30658
rect 12036 24670 12048 30646
rect 12082 24670 12094 30646
rect 12036 24658 12094 24670
rect 12194 30646 12252 30658
rect 12194 24670 12206 30646
rect 12240 24670 12252 30646
rect 12194 24658 12252 24670
rect 12352 30646 12410 30658
rect 12352 24670 12364 30646
rect 12398 24670 12410 30646
rect 12352 24658 12410 24670
rect 12510 30646 12568 30658
rect 12510 24670 12522 30646
rect 12556 24670 12568 30646
rect 12510 24658 12568 24670
rect 14070 30646 14128 30658
rect 14070 24670 14082 30646
rect 14116 24670 14128 30646
rect 14070 24658 14128 24670
rect 14228 30646 14286 30658
rect 14228 24670 14240 30646
rect 14274 24670 14286 30646
rect 14228 24658 14286 24670
rect 14386 30646 14444 30658
rect 14386 24670 14398 30646
rect 14432 24670 14444 30646
rect 14386 24658 14444 24670
rect 14544 30646 14602 30658
rect 14544 24670 14556 30646
rect 14590 24670 14602 30646
rect 14544 24658 14602 24670
rect 14702 30646 14760 30658
rect 14702 24670 14714 30646
rect 14748 24670 14760 30646
rect 14702 24658 14760 24670
rect 14860 30646 14918 30658
rect 14860 24670 14872 30646
rect 14906 24670 14918 30646
rect 14860 24658 14918 24670
rect 15018 30646 15076 30658
rect 15018 24670 15030 30646
rect 15064 24670 15076 30646
rect 15018 24658 15076 24670
rect 15176 30646 15234 30658
rect 15176 24670 15188 30646
rect 15222 24670 15234 30646
rect 15176 24658 15234 24670
rect 15334 30646 15392 30658
rect 15334 24670 15346 30646
rect 15380 24670 15392 30646
rect 15334 24658 15392 24670
rect 15492 30646 15550 30658
rect 15492 24670 15504 30646
rect 15538 24670 15550 30646
rect 15492 24658 15550 24670
rect 15650 30646 15708 30658
rect 15650 24670 15662 30646
rect 15696 24670 15708 30646
rect 15650 24658 15708 24670
rect 15808 30646 15866 30658
rect 15808 24670 15820 30646
rect 15854 24670 15866 30646
rect 15808 24658 15866 24670
rect 15966 30646 16024 30658
rect 15966 24670 15978 30646
rect 16012 24670 16024 30646
rect 15966 24658 16024 24670
rect 16124 30646 16182 30658
rect 16124 24670 16136 30646
rect 16170 24670 16182 30646
rect 16124 24658 16182 24670
rect 16282 30646 16340 30658
rect 16282 24670 16294 30646
rect 16328 24670 16340 30646
rect 16282 24658 16340 24670
rect 16440 30646 16498 30658
rect 16440 24670 16452 30646
rect 16486 24670 16498 30646
rect 16440 24658 16498 24670
rect 16598 30646 16656 30658
rect 16598 24670 16610 30646
rect 16644 24670 16656 30646
rect 16598 24658 16656 24670
rect 16756 30646 16814 30658
rect 16756 24670 16768 30646
rect 16802 24670 16814 30646
rect 16756 24658 16814 24670
rect 16914 30646 16972 30658
rect 16914 24670 16926 30646
rect 16960 24670 16972 30646
rect 16914 24658 16972 24670
rect 17072 30646 17130 30658
rect 17072 24670 17084 30646
rect 17118 24670 17130 30646
rect 17072 24658 17130 24670
rect 17230 30646 17288 30658
rect 17230 24670 17242 30646
rect 17276 24670 17288 30646
rect 17230 24658 17288 24670
rect 17388 30646 17446 30658
rect 17388 24670 17400 30646
rect 17434 24670 17446 30646
rect 17388 24658 17446 24670
rect 17546 30646 17604 30658
rect 17546 24670 17558 30646
rect 17592 24670 17604 30646
rect 17546 24658 17604 24670
rect 17704 30646 17762 30658
rect 17704 24670 17716 30646
rect 17750 24670 17762 30646
rect 17704 24658 17762 24670
rect 17862 30646 17920 30658
rect 17862 24670 17874 30646
rect 17908 24670 17920 30646
rect 17862 24658 17920 24670
rect 18020 30646 18078 30658
rect 18020 24670 18032 30646
rect 18066 24670 18078 30646
rect 18020 24658 18078 24670
rect 18178 30646 18236 30658
rect 18178 24670 18190 30646
rect 18224 24670 18236 30646
rect 18178 24658 18236 24670
rect 18336 30646 18394 30658
rect 18336 24670 18348 30646
rect 18382 24670 18394 30646
rect 18336 24658 18394 24670
rect 18494 30646 18552 30658
rect 18494 24670 18506 30646
rect 18540 24670 18552 30646
rect 18494 24658 18552 24670
rect 18652 30646 18710 30658
rect 18652 24670 18664 30646
rect 18698 24670 18710 30646
rect 18652 24658 18710 24670
rect 18810 30646 18868 30658
rect 18810 24670 18822 30646
rect 18856 24670 18868 30646
rect 18810 24658 18868 24670
rect 20370 30646 20428 30658
rect 20370 24670 20382 30646
rect 20416 24670 20428 30646
rect 20370 24658 20428 24670
rect 20528 30646 20586 30658
rect 20528 24670 20540 30646
rect 20574 24670 20586 30646
rect 20528 24658 20586 24670
rect 20686 30646 20744 30658
rect 20686 24670 20698 30646
rect 20732 24670 20744 30646
rect 20686 24658 20744 24670
rect 20844 30646 20902 30658
rect 20844 24670 20856 30646
rect 20890 24670 20902 30646
rect 20844 24658 20902 24670
rect 21002 30646 21060 30658
rect 21002 24670 21014 30646
rect 21048 24670 21060 30646
rect 21002 24658 21060 24670
rect 21160 30646 21218 30658
rect 21160 24670 21172 30646
rect 21206 24670 21218 30646
rect 21160 24658 21218 24670
rect 21318 30646 21376 30658
rect 21318 24670 21330 30646
rect 21364 24670 21376 30646
rect 21318 24658 21376 24670
rect 21476 30646 21534 30658
rect 21476 24670 21488 30646
rect 21522 24670 21534 30646
rect 21476 24658 21534 24670
rect 21634 30646 21692 30658
rect 21634 24670 21646 30646
rect 21680 24670 21692 30646
rect 21634 24658 21692 24670
rect 21792 30646 21850 30658
rect 21792 24670 21804 30646
rect 21838 24670 21850 30646
rect 21792 24658 21850 24670
rect 21950 30646 22008 30658
rect 21950 24670 21962 30646
rect 21996 24670 22008 30646
rect 21950 24658 22008 24670
rect 22108 30646 22166 30658
rect 22108 24670 22120 30646
rect 22154 24670 22166 30646
rect 22108 24658 22166 24670
rect 22266 30646 22324 30658
rect 22266 24670 22278 30646
rect 22312 24670 22324 30646
rect 22266 24658 22324 24670
rect 22424 30646 22482 30658
rect 22424 24670 22436 30646
rect 22470 24670 22482 30646
rect 22424 24658 22482 24670
rect 22582 30646 22640 30658
rect 22582 24670 22594 30646
rect 22628 24670 22640 30646
rect 22582 24658 22640 24670
rect 22740 30646 22798 30658
rect 22740 24670 22752 30646
rect 22786 24670 22798 30646
rect 22740 24658 22798 24670
rect 22898 30646 22956 30658
rect 22898 24670 22910 30646
rect 22944 24670 22956 30646
rect 22898 24658 22956 24670
rect 23056 30646 23114 30658
rect 23056 24670 23068 30646
rect 23102 24670 23114 30646
rect 23056 24658 23114 24670
rect 23214 30646 23272 30658
rect 23214 24670 23226 30646
rect 23260 24670 23272 30646
rect 23214 24658 23272 24670
rect 23372 30646 23430 30658
rect 23372 24670 23384 30646
rect 23418 24670 23430 30646
rect 23372 24658 23430 24670
rect 23530 30646 23588 30658
rect 23530 24670 23542 30646
rect 23576 24670 23588 30646
rect 23530 24658 23588 24670
rect 23688 30646 23746 30658
rect 23688 24670 23700 30646
rect 23734 24670 23746 30646
rect 23688 24658 23746 24670
rect 23846 30646 23904 30658
rect 23846 24670 23858 30646
rect 23892 24670 23904 30646
rect 23846 24658 23904 24670
rect 24004 30646 24062 30658
rect 24004 24670 24016 30646
rect 24050 24670 24062 30646
rect 24004 24658 24062 24670
rect 24162 30646 24220 30658
rect 24162 24670 24174 30646
rect 24208 24670 24220 30646
rect 24162 24658 24220 24670
rect 24320 30646 24378 30658
rect 24320 24670 24332 30646
rect 24366 24670 24378 30646
rect 24320 24658 24378 24670
rect 24478 30646 24536 30658
rect 24478 24670 24490 30646
rect 24524 24670 24536 30646
rect 24478 24658 24536 24670
rect 24636 30646 24694 30658
rect 24636 24670 24648 30646
rect 24682 24670 24694 30646
rect 24636 24658 24694 24670
rect 24794 30646 24852 30658
rect 24794 24670 24806 30646
rect 24840 24670 24852 30646
rect 24794 24658 24852 24670
rect 24952 30646 25010 30658
rect 24952 24670 24964 30646
rect 24998 24670 25010 30646
rect 24952 24658 25010 24670
rect 25110 30646 25168 30658
rect 25110 24670 25122 30646
rect 25156 24670 25168 30646
rect 25110 24658 25168 24670
rect 1470 23646 1528 23658
rect 1470 17670 1482 23646
rect 1516 17670 1528 23646
rect 1470 17658 1528 17670
rect 1628 23646 1686 23658
rect 1628 17670 1640 23646
rect 1674 17670 1686 23646
rect 1628 17658 1686 17670
rect 1786 23646 1844 23658
rect 1786 17670 1798 23646
rect 1832 17670 1844 23646
rect 1786 17658 1844 17670
rect 1944 23646 2002 23658
rect 1944 17670 1956 23646
rect 1990 17670 2002 23646
rect 1944 17658 2002 17670
rect 2102 23646 2160 23658
rect 2102 17670 2114 23646
rect 2148 17670 2160 23646
rect 2102 17658 2160 17670
rect 2260 23646 2318 23658
rect 2260 17670 2272 23646
rect 2306 17670 2318 23646
rect 2260 17658 2318 17670
rect 2418 23646 2476 23658
rect 2418 17670 2430 23646
rect 2464 17670 2476 23646
rect 2418 17658 2476 17670
rect 2576 23646 2634 23658
rect 2576 17670 2588 23646
rect 2622 17670 2634 23646
rect 2576 17658 2634 17670
rect 2734 23646 2792 23658
rect 2734 17670 2746 23646
rect 2780 17670 2792 23646
rect 2734 17658 2792 17670
rect 2892 23646 2950 23658
rect 2892 17670 2904 23646
rect 2938 17670 2950 23646
rect 2892 17658 2950 17670
rect 3050 23646 3108 23658
rect 3050 17670 3062 23646
rect 3096 17670 3108 23646
rect 3050 17658 3108 17670
rect 3208 23646 3266 23658
rect 3208 17670 3220 23646
rect 3254 17670 3266 23646
rect 3208 17658 3266 17670
rect 3366 23646 3424 23658
rect 3366 17670 3378 23646
rect 3412 17670 3424 23646
rect 3366 17658 3424 17670
rect 3524 23646 3582 23658
rect 3524 17670 3536 23646
rect 3570 17670 3582 23646
rect 3524 17658 3582 17670
rect 3682 23646 3740 23658
rect 3682 17670 3694 23646
rect 3728 17670 3740 23646
rect 3682 17658 3740 17670
rect 3840 23646 3898 23658
rect 3840 17670 3852 23646
rect 3886 17670 3898 23646
rect 3840 17658 3898 17670
rect 3998 23646 4056 23658
rect 3998 17670 4010 23646
rect 4044 17670 4056 23646
rect 3998 17658 4056 17670
rect 4156 23646 4214 23658
rect 4156 17670 4168 23646
rect 4202 17670 4214 23646
rect 4156 17658 4214 17670
rect 4314 23646 4372 23658
rect 4314 17670 4326 23646
rect 4360 17670 4372 23646
rect 4314 17658 4372 17670
rect 4472 23646 4530 23658
rect 4472 17670 4484 23646
rect 4518 17670 4530 23646
rect 4472 17658 4530 17670
rect 4630 23646 4688 23658
rect 4630 17670 4642 23646
rect 4676 17670 4688 23646
rect 4630 17658 4688 17670
rect 4788 23646 4846 23658
rect 4788 17670 4800 23646
rect 4834 17670 4846 23646
rect 4788 17658 4846 17670
rect 4946 23646 5004 23658
rect 4946 17670 4958 23646
rect 4992 17670 5004 23646
rect 4946 17658 5004 17670
rect 5104 23646 5162 23658
rect 5104 17670 5116 23646
rect 5150 17670 5162 23646
rect 5104 17658 5162 17670
rect 5262 23646 5320 23658
rect 5262 17670 5274 23646
rect 5308 17670 5320 23646
rect 5262 17658 5320 17670
rect 5420 23646 5478 23658
rect 5420 17670 5432 23646
rect 5466 17670 5478 23646
rect 5420 17658 5478 17670
rect 5578 23646 5636 23658
rect 5578 17670 5590 23646
rect 5624 17670 5636 23646
rect 5578 17658 5636 17670
rect 5736 23646 5794 23658
rect 5736 17670 5748 23646
rect 5782 17670 5794 23646
rect 5736 17658 5794 17670
rect 5894 23646 5952 23658
rect 5894 17670 5906 23646
rect 5940 17670 5952 23646
rect 5894 17658 5952 17670
rect 6052 23646 6110 23658
rect 6052 17670 6064 23646
rect 6098 17670 6110 23646
rect 6052 17658 6110 17670
rect 6210 23646 6268 23658
rect 6210 17670 6222 23646
rect 6256 17670 6268 23646
rect 6210 17658 6268 17670
rect 7770 23646 7828 23658
rect 7770 17670 7782 23646
rect 7816 17670 7828 23646
rect 7770 17658 7828 17670
rect 7928 23646 7986 23658
rect 7928 17670 7940 23646
rect 7974 17670 7986 23646
rect 7928 17658 7986 17670
rect 8086 23646 8144 23658
rect 8086 17670 8098 23646
rect 8132 17670 8144 23646
rect 8086 17658 8144 17670
rect 8244 23646 8302 23658
rect 8244 17670 8256 23646
rect 8290 17670 8302 23646
rect 8244 17658 8302 17670
rect 8402 23646 8460 23658
rect 8402 17670 8414 23646
rect 8448 17670 8460 23646
rect 8402 17658 8460 17670
rect 8560 23646 8618 23658
rect 8560 17670 8572 23646
rect 8606 17670 8618 23646
rect 8560 17658 8618 17670
rect 8718 23646 8776 23658
rect 8718 17670 8730 23646
rect 8764 17670 8776 23646
rect 8718 17658 8776 17670
rect 8876 23646 8934 23658
rect 8876 17670 8888 23646
rect 8922 17670 8934 23646
rect 8876 17658 8934 17670
rect 9034 23646 9092 23658
rect 9034 17670 9046 23646
rect 9080 17670 9092 23646
rect 9034 17658 9092 17670
rect 9192 23646 9250 23658
rect 9192 17670 9204 23646
rect 9238 17670 9250 23646
rect 9192 17658 9250 17670
rect 9350 23646 9408 23658
rect 9350 17670 9362 23646
rect 9396 17670 9408 23646
rect 9350 17658 9408 17670
rect 9508 23646 9566 23658
rect 9508 17670 9520 23646
rect 9554 17670 9566 23646
rect 9508 17658 9566 17670
rect 9666 23646 9724 23658
rect 9666 17670 9678 23646
rect 9712 17670 9724 23646
rect 9666 17658 9724 17670
rect 9824 23646 9882 23658
rect 9824 17670 9836 23646
rect 9870 17670 9882 23646
rect 9824 17658 9882 17670
rect 9982 23646 10040 23658
rect 9982 17670 9994 23646
rect 10028 17670 10040 23646
rect 9982 17658 10040 17670
rect 10140 23646 10198 23658
rect 10140 17670 10152 23646
rect 10186 17670 10198 23646
rect 10140 17658 10198 17670
rect 10298 23646 10356 23658
rect 10298 17670 10310 23646
rect 10344 17670 10356 23646
rect 10298 17658 10356 17670
rect 10456 23646 10514 23658
rect 10456 17670 10468 23646
rect 10502 17670 10514 23646
rect 10456 17658 10514 17670
rect 10614 23646 10672 23658
rect 10614 17670 10626 23646
rect 10660 17670 10672 23646
rect 10614 17658 10672 17670
rect 10772 23646 10830 23658
rect 10772 17670 10784 23646
rect 10818 17670 10830 23646
rect 10772 17658 10830 17670
rect 10930 23646 10988 23658
rect 10930 17670 10942 23646
rect 10976 17670 10988 23646
rect 10930 17658 10988 17670
rect 11088 23646 11146 23658
rect 11088 17670 11100 23646
rect 11134 17670 11146 23646
rect 11088 17658 11146 17670
rect 11246 23646 11304 23658
rect 11246 17670 11258 23646
rect 11292 17670 11304 23646
rect 11246 17658 11304 17670
rect 11404 23646 11462 23658
rect 11404 17670 11416 23646
rect 11450 17670 11462 23646
rect 11404 17658 11462 17670
rect 11562 23646 11620 23658
rect 11562 17670 11574 23646
rect 11608 17670 11620 23646
rect 11562 17658 11620 17670
rect 11720 23646 11778 23658
rect 11720 17670 11732 23646
rect 11766 17670 11778 23646
rect 11720 17658 11778 17670
rect 11878 23646 11936 23658
rect 11878 17670 11890 23646
rect 11924 17670 11936 23646
rect 11878 17658 11936 17670
rect 12036 23646 12094 23658
rect 12036 17670 12048 23646
rect 12082 17670 12094 23646
rect 12036 17658 12094 17670
rect 12194 23646 12252 23658
rect 12194 17670 12206 23646
rect 12240 17670 12252 23646
rect 12194 17658 12252 17670
rect 12352 23646 12410 23658
rect 12352 17670 12364 23646
rect 12398 17670 12410 23646
rect 12352 17658 12410 17670
rect 12510 23646 12568 23658
rect 12510 17670 12522 23646
rect 12556 17670 12568 23646
rect 12510 17658 12568 17670
rect 14070 23646 14128 23658
rect 14070 17670 14082 23646
rect 14116 17670 14128 23646
rect 14070 17658 14128 17670
rect 14228 23646 14286 23658
rect 14228 17670 14240 23646
rect 14274 17670 14286 23646
rect 14228 17658 14286 17670
rect 14386 23646 14444 23658
rect 14386 17670 14398 23646
rect 14432 17670 14444 23646
rect 14386 17658 14444 17670
rect 14544 23646 14602 23658
rect 14544 17670 14556 23646
rect 14590 17670 14602 23646
rect 14544 17658 14602 17670
rect 14702 23646 14760 23658
rect 14702 17670 14714 23646
rect 14748 17670 14760 23646
rect 14702 17658 14760 17670
rect 14860 23646 14918 23658
rect 14860 17670 14872 23646
rect 14906 17670 14918 23646
rect 14860 17658 14918 17670
rect 15018 23646 15076 23658
rect 15018 17670 15030 23646
rect 15064 17670 15076 23646
rect 15018 17658 15076 17670
rect 15176 23646 15234 23658
rect 15176 17670 15188 23646
rect 15222 17670 15234 23646
rect 15176 17658 15234 17670
rect 15334 23646 15392 23658
rect 15334 17670 15346 23646
rect 15380 17670 15392 23646
rect 15334 17658 15392 17670
rect 15492 23646 15550 23658
rect 15492 17670 15504 23646
rect 15538 17670 15550 23646
rect 15492 17658 15550 17670
rect 15650 23646 15708 23658
rect 15650 17670 15662 23646
rect 15696 17670 15708 23646
rect 15650 17658 15708 17670
rect 15808 23646 15866 23658
rect 15808 17670 15820 23646
rect 15854 17670 15866 23646
rect 15808 17658 15866 17670
rect 15966 23646 16024 23658
rect 15966 17670 15978 23646
rect 16012 17670 16024 23646
rect 15966 17658 16024 17670
rect 16124 23646 16182 23658
rect 16124 17670 16136 23646
rect 16170 17670 16182 23646
rect 16124 17658 16182 17670
rect 16282 23646 16340 23658
rect 16282 17670 16294 23646
rect 16328 17670 16340 23646
rect 16282 17658 16340 17670
rect 16440 23646 16498 23658
rect 16440 17670 16452 23646
rect 16486 17670 16498 23646
rect 16440 17658 16498 17670
rect 16598 23646 16656 23658
rect 16598 17670 16610 23646
rect 16644 17670 16656 23646
rect 16598 17658 16656 17670
rect 16756 23646 16814 23658
rect 16756 17670 16768 23646
rect 16802 17670 16814 23646
rect 16756 17658 16814 17670
rect 16914 23646 16972 23658
rect 16914 17670 16926 23646
rect 16960 17670 16972 23646
rect 16914 17658 16972 17670
rect 17072 23646 17130 23658
rect 17072 17670 17084 23646
rect 17118 17670 17130 23646
rect 17072 17658 17130 17670
rect 17230 23646 17288 23658
rect 17230 17670 17242 23646
rect 17276 17670 17288 23646
rect 17230 17658 17288 17670
rect 17388 23646 17446 23658
rect 17388 17670 17400 23646
rect 17434 17670 17446 23646
rect 17388 17658 17446 17670
rect 17546 23646 17604 23658
rect 17546 17670 17558 23646
rect 17592 17670 17604 23646
rect 17546 17658 17604 17670
rect 17704 23646 17762 23658
rect 17704 17670 17716 23646
rect 17750 17670 17762 23646
rect 17704 17658 17762 17670
rect 17862 23646 17920 23658
rect 17862 17670 17874 23646
rect 17908 17670 17920 23646
rect 17862 17658 17920 17670
rect 18020 23646 18078 23658
rect 18020 17670 18032 23646
rect 18066 17670 18078 23646
rect 18020 17658 18078 17670
rect 18178 23646 18236 23658
rect 18178 17670 18190 23646
rect 18224 17670 18236 23646
rect 18178 17658 18236 17670
rect 18336 23646 18394 23658
rect 18336 17670 18348 23646
rect 18382 17670 18394 23646
rect 18336 17658 18394 17670
rect 18494 23646 18552 23658
rect 18494 17670 18506 23646
rect 18540 17670 18552 23646
rect 18494 17658 18552 17670
rect 18652 23646 18710 23658
rect 18652 17670 18664 23646
rect 18698 17670 18710 23646
rect 18652 17658 18710 17670
rect 18810 23646 18868 23658
rect 18810 17670 18822 23646
rect 18856 17670 18868 23646
rect 18810 17658 18868 17670
rect 20370 23646 20428 23658
rect 20370 17670 20382 23646
rect 20416 17670 20428 23646
rect 20370 17658 20428 17670
rect 20528 23646 20586 23658
rect 20528 17670 20540 23646
rect 20574 17670 20586 23646
rect 20528 17658 20586 17670
rect 20686 23646 20744 23658
rect 20686 17670 20698 23646
rect 20732 17670 20744 23646
rect 20686 17658 20744 17670
rect 20844 23646 20902 23658
rect 20844 17670 20856 23646
rect 20890 17670 20902 23646
rect 20844 17658 20902 17670
rect 21002 23646 21060 23658
rect 21002 17670 21014 23646
rect 21048 17670 21060 23646
rect 21002 17658 21060 17670
rect 21160 23646 21218 23658
rect 21160 17670 21172 23646
rect 21206 17670 21218 23646
rect 21160 17658 21218 17670
rect 21318 23646 21376 23658
rect 21318 17670 21330 23646
rect 21364 17670 21376 23646
rect 21318 17658 21376 17670
rect 21476 23646 21534 23658
rect 21476 17670 21488 23646
rect 21522 17670 21534 23646
rect 21476 17658 21534 17670
rect 21634 23646 21692 23658
rect 21634 17670 21646 23646
rect 21680 17670 21692 23646
rect 21634 17658 21692 17670
rect 21792 23646 21850 23658
rect 21792 17670 21804 23646
rect 21838 17670 21850 23646
rect 21792 17658 21850 17670
rect 21950 23646 22008 23658
rect 21950 17670 21962 23646
rect 21996 17670 22008 23646
rect 21950 17658 22008 17670
rect 22108 23646 22166 23658
rect 22108 17670 22120 23646
rect 22154 17670 22166 23646
rect 22108 17658 22166 17670
rect 22266 23646 22324 23658
rect 22266 17670 22278 23646
rect 22312 17670 22324 23646
rect 22266 17658 22324 17670
rect 22424 23646 22482 23658
rect 22424 17670 22436 23646
rect 22470 17670 22482 23646
rect 22424 17658 22482 17670
rect 22582 23646 22640 23658
rect 22582 17670 22594 23646
rect 22628 17670 22640 23646
rect 22582 17658 22640 17670
rect 22740 23646 22798 23658
rect 22740 17670 22752 23646
rect 22786 17670 22798 23646
rect 22740 17658 22798 17670
rect 22898 23646 22956 23658
rect 22898 17670 22910 23646
rect 22944 17670 22956 23646
rect 22898 17658 22956 17670
rect 23056 23646 23114 23658
rect 23056 17670 23068 23646
rect 23102 17670 23114 23646
rect 23056 17658 23114 17670
rect 23214 23646 23272 23658
rect 23214 17670 23226 23646
rect 23260 17670 23272 23646
rect 23214 17658 23272 17670
rect 23372 23646 23430 23658
rect 23372 17670 23384 23646
rect 23418 17670 23430 23646
rect 23372 17658 23430 17670
rect 23530 23646 23588 23658
rect 23530 17670 23542 23646
rect 23576 17670 23588 23646
rect 23530 17658 23588 17670
rect 23688 23646 23746 23658
rect 23688 17670 23700 23646
rect 23734 17670 23746 23646
rect 23688 17658 23746 17670
rect 23846 23646 23904 23658
rect 23846 17670 23858 23646
rect 23892 17670 23904 23646
rect 23846 17658 23904 17670
rect 24004 23646 24062 23658
rect 24004 17670 24016 23646
rect 24050 17670 24062 23646
rect 24004 17658 24062 17670
rect 24162 23646 24220 23658
rect 24162 17670 24174 23646
rect 24208 17670 24220 23646
rect 24162 17658 24220 17670
rect 24320 23646 24378 23658
rect 24320 17670 24332 23646
rect 24366 17670 24378 23646
rect 24320 17658 24378 17670
rect 24478 23646 24536 23658
rect 24478 17670 24490 23646
rect 24524 17670 24536 23646
rect 24478 17658 24536 17670
rect 24636 23646 24694 23658
rect 24636 17670 24648 23646
rect 24682 17670 24694 23646
rect 24636 17658 24694 17670
rect 24794 23646 24852 23658
rect 24794 17670 24806 23646
rect 24840 17670 24852 23646
rect 24794 17658 24852 17670
rect 24952 23646 25010 23658
rect 24952 17670 24964 23646
rect 24998 17670 25010 23646
rect 24952 17658 25010 17670
rect 25110 23646 25168 23658
rect 25110 17670 25122 23646
rect 25156 17670 25168 23646
rect 25110 17658 25168 17670
rect 1470 15346 1528 15358
rect 1470 9370 1482 15346
rect 1516 9370 1528 15346
rect 1470 9358 1528 9370
rect 1628 15346 1686 15358
rect 1628 9370 1640 15346
rect 1674 9370 1686 15346
rect 1628 9358 1686 9370
rect 1786 15346 1844 15358
rect 1786 9370 1798 15346
rect 1832 9370 1844 15346
rect 1786 9358 1844 9370
rect 1944 15346 2002 15358
rect 1944 9370 1956 15346
rect 1990 9370 2002 15346
rect 1944 9358 2002 9370
rect 2102 15346 2160 15358
rect 2102 9370 2114 15346
rect 2148 9370 2160 15346
rect 2102 9358 2160 9370
rect 2260 15346 2318 15358
rect 2260 9370 2272 15346
rect 2306 9370 2318 15346
rect 2260 9358 2318 9370
rect 2418 15346 2476 15358
rect 2418 9370 2430 15346
rect 2464 9370 2476 15346
rect 2418 9358 2476 9370
rect 2576 15346 2634 15358
rect 2576 9370 2588 15346
rect 2622 9370 2634 15346
rect 2576 9358 2634 9370
rect 2734 15346 2792 15358
rect 2734 9370 2746 15346
rect 2780 9370 2792 15346
rect 2734 9358 2792 9370
rect 2892 15346 2950 15358
rect 2892 9370 2904 15346
rect 2938 9370 2950 15346
rect 2892 9358 2950 9370
rect 3050 15346 3108 15358
rect 3050 9370 3062 15346
rect 3096 9370 3108 15346
rect 3050 9358 3108 9370
rect 3208 15346 3266 15358
rect 3208 9370 3220 15346
rect 3254 9370 3266 15346
rect 3208 9358 3266 9370
rect 3366 15346 3424 15358
rect 3366 9370 3378 15346
rect 3412 9370 3424 15346
rect 3366 9358 3424 9370
rect 3524 15346 3582 15358
rect 3524 9370 3536 15346
rect 3570 9370 3582 15346
rect 3524 9358 3582 9370
rect 3682 15346 3740 15358
rect 3682 9370 3694 15346
rect 3728 9370 3740 15346
rect 3682 9358 3740 9370
rect 3840 15346 3898 15358
rect 3840 9370 3852 15346
rect 3886 9370 3898 15346
rect 3840 9358 3898 9370
rect 3998 15346 4056 15358
rect 3998 9370 4010 15346
rect 4044 9370 4056 15346
rect 3998 9358 4056 9370
rect 4156 15346 4214 15358
rect 4156 9370 4168 15346
rect 4202 9370 4214 15346
rect 4156 9358 4214 9370
rect 4314 15346 4372 15358
rect 4314 9370 4326 15346
rect 4360 9370 4372 15346
rect 4314 9358 4372 9370
rect 4472 15346 4530 15358
rect 4472 9370 4484 15346
rect 4518 9370 4530 15346
rect 4472 9358 4530 9370
rect 4630 15346 4688 15358
rect 4630 9370 4642 15346
rect 4676 9370 4688 15346
rect 4630 9358 4688 9370
rect 4788 15346 4846 15358
rect 4788 9370 4800 15346
rect 4834 9370 4846 15346
rect 4788 9358 4846 9370
rect 4946 15346 5004 15358
rect 4946 9370 4958 15346
rect 4992 9370 5004 15346
rect 4946 9358 5004 9370
rect 5104 15346 5162 15358
rect 5104 9370 5116 15346
rect 5150 9370 5162 15346
rect 5104 9358 5162 9370
rect 5262 15346 5320 15358
rect 5262 9370 5274 15346
rect 5308 9370 5320 15346
rect 5262 9358 5320 9370
rect 5420 15346 5478 15358
rect 5420 9370 5432 15346
rect 5466 9370 5478 15346
rect 5420 9358 5478 9370
rect 5578 15346 5636 15358
rect 5578 9370 5590 15346
rect 5624 9370 5636 15346
rect 5578 9358 5636 9370
rect 5736 15346 5794 15358
rect 5736 9370 5748 15346
rect 5782 9370 5794 15346
rect 5736 9358 5794 9370
rect 5894 15346 5952 15358
rect 5894 9370 5906 15346
rect 5940 9370 5952 15346
rect 5894 9358 5952 9370
rect 6052 15346 6110 15358
rect 6052 9370 6064 15346
rect 6098 9370 6110 15346
rect 6052 9358 6110 9370
rect 6210 15346 6268 15358
rect 6210 9370 6222 15346
rect 6256 9370 6268 15346
rect 6210 9358 6268 9370
rect 7770 15346 7828 15358
rect 7770 9370 7782 15346
rect 7816 9370 7828 15346
rect 7770 9358 7828 9370
rect 7928 15346 7986 15358
rect 7928 9370 7940 15346
rect 7974 9370 7986 15346
rect 7928 9358 7986 9370
rect 8086 15346 8144 15358
rect 8086 9370 8098 15346
rect 8132 9370 8144 15346
rect 8086 9358 8144 9370
rect 8244 15346 8302 15358
rect 8244 9370 8256 15346
rect 8290 9370 8302 15346
rect 8244 9358 8302 9370
rect 8402 15346 8460 15358
rect 8402 9370 8414 15346
rect 8448 9370 8460 15346
rect 8402 9358 8460 9370
rect 8560 15346 8618 15358
rect 8560 9370 8572 15346
rect 8606 9370 8618 15346
rect 8560 9358 8618 9370
rect 8718 15346 8776 15358
rect 8718 9370 8730 15346
rect 8764 9370 8776 15346
rect 8718 9358 8776 9370
rect 8876 15346 8934 15358
rect 8876 9370 8888 15346
rect 8922 9370 8934 15346
rect 8876 9358 8934 9370
rect 9034 15346 9092 15358
rect 9034 9370 9046 15346
rect 9080 9370 9092 15346
rect 9034 9358 9092 9370
rect 9192 15346 9250 15358
rect 9192 9370 9204 15346
rect 9238 9370 9250 15346
rect 9192 9358 9250 9370
rect 9350 15346 9408 15358
rect 9350 9370 9362 15346
rect 9396 9370 9408 15346
rect 9350 9358 9408 9370
rect 9508 15346 9566 15358
rect 9508 9370 9520 15346
rect 9554 9370 9566 15346
rect 9508 9358 9566 9370
rect 9666 15346 9724 15358
rect 9666 9370 9678 15346
rect 9712 9370 9724 15346
rect 9666 9358 9724 9370
rect 9824 15346 9882 15358
rect 9824 9370 9836 15346
rect 9870 9370 9882 15346
rect 9824 9358 9882 9370
rect 9982 15346 10040 15358
rect 9982 9370 9994 15346
rect 10028 9370 10040 15346
rect 9982 9358 10040 9370
rect 10140 15346 10198 15358
rect 10140 9370 10152 15346
rect 10186 9370 10198 15346
rect 10140 9358 10198 9370
rect 10298 15346 10356 15358
rect 10298 9370 10310 15346
rect 10344 9370 10356 15346
rect 10298 9358 10356 9370
rect 10456 15346 10514 15358
rect 10456 9370 10468 15346
rect 10502 9370 10514 15346
rect 10456 9358 10514 9370
rect 10614 15346 10672 15358
rect 10614 9370 10626 15346
rect 10660 9370 10672 15346
rect 10614 9358 10672 9370
rect 10772 15346 10830 15358
rect 10772 9370 10784 15346
rect 10818 9370 10830 15346
rect 10772 9358 10830 9370
rect 10930 15346 10988 15358
rect 10930 9370 10942 15346
rect 10976 9370 10988 15346
rect 10930 9358 10988 9370
rect 11088 15346 11146 15358
rect 11088 9370 11100 15346
rect 11134 9370 11146 15346
rect 11088 9358 11146 9370
rect 11246 15346 11304 15358
rect 11246 9370 11258 15346
rect 11292 9370 11304 15346
rect 11246 9358 11304 9370
rect 11404 15346 11462 15358
rect 11404 9370 11416 15346
rect 11450 9370 11462 15346
rect 11404 9358 11462 9370
rect 11562 15346 11620 15358
rect 11562 9370 11574 15346
rect 11608 9370 11620 15346
rect 11562 9358 11620 9370
rect 11720 15346 11778 15358
rect 11720 9370 11732 15346
rect 11766 9370 11778 15346
rect 11720 9358 11778 9370
rect 11878 15346 11936 15358
rect 11878 9370 11890 15346
rect 11924 9370 11936 15346
rect 11878 9358 11936 9370
rect 12036 15346 12094 15358
rect 12036 9370 12048 15346
rect 12082 9370 12094 15346
rect 12036 9358 12094 9370
rect 12194 15346 12252 15358
rect 12194 9370 12206 15346
rect 12240 9370 12252 15346
rect 12194 9358 12252 9370
rect 12352 15346 12410 15358
rect 12352 9370 12364 15346
rect 12398 9370 12410 15346
rect 12352 9358 12410 9370
rect 12510 15346 12568 15358
rect 12510 9370 12522 15346
rect 12556 9370 12568 15346
rect 12510 9358 12568 9370
rect 14070 15346 14128 15358
rect 14070 9370 14082 15346
rect 14116 9370 14128 15346
rect 14070 9358 14128 9370
rect 14228 15346 14286 15358
rect 14228 9370 14240 15346
rect 14274 9370 14286 15346
rect 14228 9358 14286 9370
rect 14386 15346 14444 15358
rect 14386 9370 14398 15346
rect 14432 9370 14444 15346
rect 14386 9358 14444 9370
rect 14544 15346 14602 15358
rect 14544 9370 14556 15346
rect 14590 9370 14602 15346
rect 14544 9358 14602 9370
rect 14702 15346 14760 15358
rect 14702 9370 14714 15346
rect 14748 9370 14760 15346
rect 14702 9358 14760 9370
rect 14860 15346 14918 15358
rect 14860 9370 14872 15346
rect 14906 9370 14918 15346
rect 14860 9358 14918 9370
rect 15018 15346 15076 15358
rect 15018 9370 15030 15346
rect 15064 9370 15076 15346
rect 15018 9358 15076 9370
rect 15176 15346 15234 15358
rect 15176 9370 15188 15346
rect 15222 9370 15234 15346
rect 15176 9358 15234 9370
rect 15334 15346 15392 15358
rect 15334 9370 15346 15346
rect 15380 9370 15392 15346
rect 15334 9358 15392 9370
rect 15492 15346 15550 15358
rect 15492 9370 15504 15346
rect 15538 9370 15550 15346
rect 15492 9358 15550 9370
rect 15650 15346 15708 15358
rect 15650 9370 15662 15346
rect 15696 9370 15708 15346
rect 15650 9358 15708 9370
rect 15808 15346 15866 15358
rect 15808 9370 15820 15346
rect 15854 9370 15866 15346
rect 15808 9358 15866 9370
rect 15966 15346 16024 15358
rect 15966 9370 15978 15346
rect 16012 9370 16024 15346
rect 15966 9358 16024 9370
rect 16124 15346 16182 15358
rect 16124 9370 16136 15346
rect 16170 9370 16182 15346
rect 16124 9358 16182 9370
rect 16282 15346 16340 15358
rect 16282 9370 16294 15346
rect 16328 9370 16340 15346
rect 16282 9358 16340 9370
rect 16440 15346 16498 15358
rect 16440 9370 16452 15346
rect 16486 9370 16498 15346
rect 16440 9358 16498 9370
rect 16598 15346 16656 15358
rect 16598 9370 16610 15346
rect 16644 9370 16656 15346
rect 16598 9358 16656 9370
rect 16756 15346 16814 15358
rect 16756 9370 16768 15346
rect 16802 9370 16814 15346
rect 16756 9358 16814 9370
rect 16914 15346 16972 15358
rect 16914 9370 16926 15346
rect 16960 9370 16972 15346
rect 16914 9358 16972 9370
rect 17072 15346 17130 15358
rect 17072 9370 17084 15346
rect 17118 9370 17130 15346
rect 17072 9358 17130 9370
rect 17230 15346 17288 15358
rect 17230 9370 17242 15346
rect 17276 9370 17288 15346
rect 17230 9358 17288 9370
rect 17388 15346 17446 15358
rect 17388 9370 17400 15346
rect 17434 9370 17446 15346
rect 17388 9358 17446 9370
rect 17546 15346 17604 15358
rect 17546 9370 17558 15346
rect 17592 9370 17604 15346
rect 17546 9358 17604 9370
rect 17704 15346 17762 15358
rect 17704 9370 17716 15346
rect 17750 9370 17762 15346
rect 17704 9358 17762 9370
rect 17862 15346 17920 15358
rect 17862 9370 17874 15346
rect 17908 9370 17920 15346
rect 17862 9358 17920 9370
rect 18020 15346 18078 15358
rect 18020 9370 18032 15346
rect 18066 9370 18078 15346
rect 18020 9358 18078 9370
rect 18178 15346 18236 15358
rect 18178 9370 18190 15346
rect 18224 9370 18236 15346
rect 18178 9358 18236 9370
rect 18336 15346 18394 15358
rect 18336 9370 18348 15346
rect 18382 9370 18394 15346
rect 18336 9358 18394 9370
rect 18494 15346 18552 15358
rect 18494 9370 18506 15346
rect 18540 9370 18552 15346
rect 18494 9358 18552 9370
rect 18652 15346 18710 15358
rect 18652 9370 18664 15346
rect 18698 9370 18710 15346
rect 18652 9358 18710 9370
rect 18810 15346 18868 15358
rect 18810 9370 18822 15346
rect 18856 9370 18868 15346
rect 18810 9358 18868 9370
rect 20370 15346 20428 15358
rect 20370 9370 20382 15346
rect 20416 9370 20428 15346
rect 20370 9358 20428 9370
rect 20528 15346 20586 15358
rect 20528 9370 20540 15346
rect 20574 9370 20586 15346
rect 20528 9358 20586 9370
rect 20686 15346 20744 15358
rect 20686 9370 20698 15346
rect 20732 9370 20744 15346
rect 20686 9358 20744 9370
rect 20844 15346 20902 15358
rect 20844 9370 20856 15346
rect 20890 9370 20902 15346
rect 20844 9358 20902 9370
rect 21002 15346 21060 15358
rect 21002 9370 21014 15346
rect 21048 9370 21060 15346
rect 21002 9358 21060 9370
rect 21160 15346 21218 15358
rect 21160 9370 21172 15346
rect 21206 9370 21218 15346
rect 21160 9358 21218 9370
rect 21318 15346 21376 15358
rect 21318 9370 21330 15346
rect 21364 9370 21376 15346
rect 21318 9358 21376 9370
rect 21476 15346 21534 15358
rect 21476 9370 21488 15346
rect 21522 9370 21534 15346
rect 21476 9358 21534 9370
rect 21634 15346 21692 15358
rect 21634 9370 21646 15346
rect 21680 9370 21692 15346
rect 21634 9358 21692 9370
rect 21792 15346 21850 15358
rect 21792 9370 21804 15346
rect 21838 9370 21850 15346
rect 21792 9358 21850 9370
rect 21950 15346 22008 15358
rect 21950 9370 21962 15346
rect 21996 9370 22008 15346
rect 21950 9358 22008 9370
rect 22108 15346 22166 15358
rect 22108 9370 22120 15346
rect 22154 9370 22166 15346
rect 22108 9358 22166 9370
rect 22266 15346 22324 15358
rect 22266 9370 22278 15346
rect 22312 9370 22324 15346
rect 22266 9358 22324 9370
rect 22424 15346 22482 15358
rect 22424 9370 22436 15346
rect 22470 9370 22482 15346
rect 22424 9358 22482 9370
rect 22582 15346 22640 15358
rect 22582 9370 22594 15346
rect 22628 9370 22640 15346
rect 22582 9358 22640 9370
rect 22740 15346 22798 15358
rect 22740 9370 22752 15346
rect 22786 9370 22798 15346
rect 22740 9358 22798 9370
rect 22898 15346 22956 15358
rect 22898 9370 22910 15346
rect 22944 9370 22956 15346
rect 22898 9358 22956 9370
rect 23056 15346 23114 15358
rect 23056 9370 23068 15346
rect 23102 9370 23114 15346
rect 23056 9358 23114 9370
rect 23214 15346 23272 15358
rect 23214 9370 23226 15346
rect 23260 9370 23272 15346
rect 23214 9358 23272 9370
rect 23372 15346 23430 15358
rect 23372 9370 23384 15346
rect 23418 9370 23430 15346
rect 23372 9358 23430 9370
rect 23530 15346 23588 15358
rect 23530 9370 23542 15346
rect 23576 9370 23588 15346
rect 23530 9358 23588 9370
rect 23688 15346 23746 15358
rect 23688 9370 23700 15346
rect 23734 9370 23746 15346
rect 23688 9358 23746 9370
rect 23846 15346 23904 15358
rect 23846 9370 23858 15346
rect 23892 9370 23904 15346
rect 23846 9358 23904 9370
rect 24004 15346 24062 15358
rect 24004 9370 24016 15346
rect 24050 9370 24062 15346
rect 24004 9358 24062 9370
rect 24162 15346 24220 15358
rect 24162 9370 24174 15346
rect 24208 9370 24220 15346
rect 24162 9358 24220 9370
rect 24320 15346 24378 15358
rect 24320 9370 24332 15346
rect 24366 9370 24378 15346
rect 24320 9358 24378 9370
rect 24478 15346 24536 15358
rect 24478 9370 24490 15346
rect 24524 9370 24536 15346
rect 24478 9358 24536 9370
rect 24636 15346 24694 15358
rect 24636 9370 24648 15346
rect 24682 9370 24694 15346
rect 24636 9358 24694 9370
rect 24794 15346 24852 15358
rect 24794 9370 24806 15346
rect 24840 9370 24852 15346
rect 24794 9358 24852 9370
rect 24952 15346 25010 15358
rect 24952 9370 24964 15346
rect 24998 9370 25010 15346
rect 24952 9358 25010 9370
rect 25110 15346 25168 15358
rect 25110 9370 25122 15346
rect 25156 9370 25168 15346
rect 25110 9358 25168 9370
rect 1470 8346 1528 8358
rect 1470 2370 1482 8346
rect 1516 2370 1528 8346
rect 1470 2358 1528 2370
rect 1628 8346 1686 8358
rect 1628 2370 1640 8346
rect 1674 2370 1686 8346
rect 1628 2358 1686 2370
rect 1786 8346 1844 8358
rect 1786 2370 1798 8346
rect 1832 2370 1844 8346
rect 1786 2358 1844 2370
rect 1944 8346 2002 8358
rect 1944 2370 1956 8346
rect 1990 2370 2002 8346
rect 1944 2358 2002 2370
rect 2102 8346 2160 8358
rect 2102 2370 2114 8346
rect 2148 2370 2160 8346
rect 2102 2358 2160 2370
rect 2260 8346 2318 8358
rect 2260 2370 2272 8346
rect 2306 2370 2318 8346
rect 2260 2358 2318 2370
rect 2418 8346 2476 8358
rect 2418 2370 2430 8346
rect 2464 2370 2476 8346
rect 2418 2358 2476 2370
rect 2576 8346 2634 8358
rect 2576 2370 2588 8346
rect 2622 2370 2634 8346
rect 2576 2358 2634 2370
rect 2734 8346 2792 8358
rect 2734 2370 2746 8346
rect 2780 2370 2792 8346
rect 2734 2358 2792 2370
rect 2892 8346 2950 8358
rect 2892 2370 2904 8346
rect 2938 2370 2950 8346
rect 2892 2358 2950 2370
rect 3050 8346 3108 8358
rect 3050 2370 3062 8346
rect 3096 2370 3108 8346
rect 3050 2358 3108 2370
rect 3208 8346 3266 8358
rect 3208 2370 3220 8346
rect 3254 2370 3266 8346
rect 3208 2358 3266 2370
rect 3366 8346 3424 8358
rect 3366 2370 3378 8346
rect 3412 2370 3424 8346
rect 3366 2358 3424 2370
rect 3524 8346 3582 8358
rect 3524 2370 3536 8346
rect 3570 2370 3582 8346
rect 3524 2358 3582 2370
rect 3682 8346 3740 8358
rect 3682 2370 3694 8346
rect 3728 2370 3740 8346
rect 3682 2358 3740 2370
rect 3840 8346 3898 8358
rect 3840 2370 3852 8346
rect 3886 2370 3898 8346
rect 3840 2358 3898 2370
rect 3998 8346 4056 8358
rect 3998 2370 4010 8346
rect 4044 2370 4056 8346
rect 3998 2358 4056 2370
rect 4156 8346 4214 8358
rect 4156 2370 4168 8346
rect 4202 2370 4214 8346
rect 4156 2358 4214 2370
rect 4314 8346 4372 8358
rect 4314 2370 4326 8346
rect 4360 2370 4372 8346
rect 4314 2358 4372 2370
rect 4472 8346 4530 8358
rect 4472 2370 4484 8346
rect 4518 2370 4530 8346
rect 4472 2358 4530 2370
rect 4630 8346 4688 8358
rect 4630 2370 4642 8346
rect 4676 2370 4688 8346
rect 4630 2358 4688 2370
rect 4788 8346 4846 8358
rect 4788 2370 4800 8346
rect 4834 2370 4846 8346
rect 4788 2358 4846 2370
rect 4946 8346 5004 8358
rect 4946 2370 4958 8346
rect 4992 2370 5004 8346
rect 4946 2358 5004 2370
rect 5104 8346 5162 8358
rect 5104 2370 5116 8346
rect 5150 2370 5162 8346
rect 5104 2358 5162 2370
rect 5262 8346 5320 8358
rect 5262 2370 5274 8346
rect 5308 2370 5320 8346
rect 5262 2358 5320 2370
rect 5420 8346 5478 8358
rect 5420 2370 5432 8346
rect 5466 2370 5478 8346
rect 5420 2358 5478 2370
rect 5578 8346 5636 8358
rect 5578 2370 5590 8346
rect 5624 2370 5636 8346
rect 5578 2358 5636 2370
rect 5736 8346 5794 8358
rect 5736 2370 5748 8346
rect 5782 2370 5794 8346
rect 5736 2358 5794 2370
rect 5894 8346 5952 8358
rect 5894 2370 5906 8346
rect 5940 2370 5952 8346
rect 5894 2358 5952 2370
rect 6052 8346 6110 8358
rect 6052 2370 6064 8346
rect 6098 2370 6110 8346
rect 6052 2358 6110 2370
rect 6210 8346 6268 8358
rect 6210 2370 6222 8346
rect 6256 2370 6268 8346
rect 6210 2358 6268 2370
rect 7770 8346 7828 8358
rect 7770 2370 7782 8346
rect 7816 2370 7828 8346
rect 7770 2358 7828 2370
rect 7928 8346 7986 8358
rect 7928 2370 7940 8346
rect 7974 2370 7986 8346
rect 7928 2358 7986 2370
rect 8086 8346 8144 8358
rect 8086 2370 8098 8346
rect 8132 2370 8144 8346
rect 8086 2358 8144 2370
rect 8244 8346 8302 8358
rect 8244 2370 8256 8346
rect 8290 2370 8302 8346
rect 8244 2358 8302 2370
rect 8402 8346 8460 8358
rect 8402 2370 8414 8346
rect 8448 2370 8460 8346
rect 8402 2358 8460 2370
rect 8560 8346 8618 8358
rect 8560 2370 8572 8346
rect 8606 2370 8618 8346
rect 8560 2358 8618 2370
rect 8718 8346 8776 8358
rect 8718 2370 8730 8346
rect 8764 2370 8776 8346
rect 8718 2358 8776 2370
rect 8876 8346 8934 8358
rect 8876 2370 8888 8346
rect 8922 2370 8934 8346
rect 8876 2358 8934 2370
rect 9034 8346 9092 8358
rect 9034 2370 9046 8346
rect 9080 2370 9092 8346
rect 9034 2358 9092 2370
rect 9192 8346 9250 8358
rect 9192 2370 9204 8346
rect 9238 2370 9250 8346
rect 9192 2358 9250 2370
rect 9350 8346 9408 8358
rect 9350 2370 9362 8346
rect 9396 2370 9408 8346
rect 9350 2358 9408 2370
rect 9508 8346 9566 8358
rect 9508 2370 9520 8346
rect 9554 2370 9566 8346
rect 9508 2358 9566 2370
rect 9666 8346 9724 8358
rect 9666 2370 9678 8346
rect 9712 2370 9724 8346
rect 9666 2358 9724 2370
rect 9824 8346 9882 8358
rect 9824 2370 9836 8346
rect 9870 2370 9882 8346
rect 9824 2358 9882 2370
rect 9982 8346 10040 8358
rect 9982 2370 9994 8346
rect 10028 2370 10040 8346
rect 9982 2358 10040 2370
rect 10140 8346 10198 8358
rect 10140 2370 10152 8346
rect 10186 2370 10198 8346
rect 10140 2358 10198 2370
rect 10298 8346 10356 8358
rect 10298 2370 10310 8346
rect 10344 2370 10356 8346
rect 10298 2358 10356 2370
rect 10456 8346 10514 8358
rect 10456 2370 10468 8346
rect 10502 2370 10514 8346
rect 10456 2358 10514 2370
rect 10614 8346 10672 8358
rect 10614 2370 10626 8346
rect 10660 2370 10672 8346
rect 10614 2358 10672 2370
rect 10772 8346 10830 8358
rect 10772 2370 10784 8346
rect 10818 2370 10830 8346
rect 10772 2358 10830 2370
rect 10930 8346 10988 8358
rect 10930 2370 10942 8346
rect 10976 2370 10988 8346
rect 10930 2358 10988 2370
rect 11088 8346 11146 8358
rect 11088 2370 11100 8346
rect 11134 2370 11146 8346
rect 11088 2358 11146 2370
rect 11246 8346 11304 8358
rect 11246 2370 11258 8346
rect 11292 2370 11304 8346
rect 11246 2358 11304 2370
rect 11404 8346 11462 8358
rect 11404 2370 11416 8346
rect 11450 2370 11462 8346
rect 11404 2358 11462 2370
rect 11562 8346 11620 8358
rect 11562 2370 11574 8346
rect 11608 2370 11620 8346
rect 11562 2358 11620 2370
rect 11720 8346 11778 8358
rect 11720 2370 11732 8346
rect 11766 2370 11778 8346
rect 11720 2358 11778 2370
rect 11878 8346 11936 8358
rect 11878 2370 11890 8346
rect 11924 2370 11936 8346
rect 11878 2358 11936 2370
rect 12036 8346 12094 8358
rect 12036 2370 12048 8346
rect 12082 2370 12094 8346
rect 12036 2358 12094 2370
rect 12194 8346 12252 8358
rect 12194 2370 12206 8346
rect 12240 2370 12252 8346
rect 12194 2358 12252 2370
rect 12352 8346 12410 8358
rect 12352 2370 12364 8346
rect 12398 2370 12410 8346
rect 12352 2358 12410 2370
rect 12510 8346 12568 8358
rect 12510 2370 12522 8346
rect 12556 2370 12568 8346
rect 12510 2358 12568 2370
rect 14070 8346 14128 8358
rect 14070 2370 14082 8346
rect 14116 2370 14128 8346
rect 14070 2358 14128 2370
rect 14228 8346 14286 8358
rect 14228 2370 14240 8346
rect 14274 2370 14286 8346
rect 14228 2358 14286 2370
rect 14386 8346 14444 8358
rect 14386 2370 14398 8346
rect 14432 2370 14444 8346
rect 14386 2358 14444 2370
rect 14544 8346 14602 8358
rect 14544 2370 14556 8346
rect 14590 2370 14602 8346
rect 14544 2358 14602 2370
rect 14702 8346 14760 8358
rect 14702 2370 14714 8346
rect 14748 2370 14760 8346
rect 14702 2358 14760 2370
rect 14860 8346 14918 8358
rect 14860 2370 14872 8346
rect 14906 2370 14918 8346
rect 14860 2358 14918 2370
rect 15018 8346 15076 8358
rect 15018 2370 15030 8346
rect 15064 2370 15076 8346
rect 15018 2358 15076 2370
rect 15176 8346 15234 8358
rect 15176 2370 15188 8346
rect 15222 2370 15234 8346
rect 15176 2358 15234 2370
rect 15334 8346 15392 8358
rect 15334 2370 15346 8346
rect 15380 2370 15392 8346
rect 15334 2358 15392 2370
rect 15492 8346 15550 8358
rect 15492 2370 15504 8346
rect 15538 2370 15550 8346
rect 15492 2358 15550 2370
rect 15650 8346 15708 8358
rect 15650 2370 15662 8346
rect 15696 2370 15708 8346
rect 15650 2358 15708 2370
rect 15808 8346 15866 8358
rect 15808 2370 15820 8346
rect 15854 2370 15866 8346
rect 15808 2358 15866 2370
rect 15966 8346 16024 8358
rect 15966 2370 15978 8346
rect 16012 2370 16024 8346
rect 15966 2358 16024 2370
rect 16124 8346 16182 8358
rect 16124 2370 16136 8346
rect 16170 2370 16182 8346
rect 16124 2358 16182 2370
rect 16282 8346 16340 8358
rect 16282 2370 16294 8346
rect 16328 2370 16340 8346
rect 16282 2358 16340 2370
rect 16440 8346 16498 8358
rect 16440 2370 16452 8346
rect 16486 2370 16498 8346
rect 16440 2358 16498 2370
rect 16598 8346 16656 8358
rect 16598 2370 16610 8346
rect 16644 2370 16656 8346
rect 16598 2358 16656 2370
rect 16756 8346 16814 8358
rect 16756 2370 16768 8346
rect 16802 2370 16814 8346
rect 16756 2358 16814 2370
rect 16914 8346 16972 8358
rect 16914 2370 16926 8346
rect 16960 2370 16972 8346
rect 16914 2358 16972 2370
rect 17072 8346 17130 8358
rect 17072 2370 17084 8346
rect 17118 2370 17130 8346
rect 17072 2358 17130 2370
rect 17230 8346 17288 8358
rect 17230 2370 17242 8346
rect 17276 2370 17288 8346
rect 17230 2358 17288 2370
rect 17388 8346 17446 8358
rect 17388 2370 17400 8346
rect 17434 2370 17446 8346
rect 17388 2358 17446 2370
rect 17546 8346 17604 8358
rect 17546 2370 17558 8346
rect 17592 2370 17604 8346
rect 17546 2358 17604 2370
rect 17704 8346 17762 8358
rect 17704 2370 17716 8346
rect 17750 2370 17762 8346
rect 17704 2358 17762 2370
rect 17862 8346 17920 8358
rect 17862 2370 17874 8346
rect 17908 2370 17920 8346
rect 17862 2358 17920 2370
rect 18020 8346 18078 8358
rect 18020 2370 18032 8346
rect 18066 2370 18078 8346
rect 18020 2358 18078 2370
rect 18178 8346 18236 8358
rect 18178 2370 18190 8346
rect 18224 2370 18236 8346
rect 18178 2358 18236 2370
rect 18336 8346 18394 8358
rect 18336 2370 18348 8346
rect 18382 2370 18394 8346
rect 18336 2358 18394 2370
rect 18494 8346 18552 8358
rect 18494 2370 18506 8346
rect 18540 2370 18552 8346
rect 18494 2358 18552 2370
rect 18652 8346 18710 8358
rect 18652 2370 18664 8346
rect 18698 2370 18710 8346
rect 18652 2358 18710 2370
rect 18810 8346 18868 8358
rect 18810 2370 18822 8346
rect 18856 2370 18868 8346
rect 18810 2358 18868 2370
rect 20370 8346 20428 8358
rect 20370 2370 20382 8346
rect 20416 2370 20428 8346
rect 20370 2358 20428 2370
rect 20528 8346 20586 8358
rect 20528 2370 20540 8346
rect 20574 2370 20586 8346
rect 20528 2358 20586 2370
rect 20686 8346 20744 8358
rect 20686 2370 20698 8346
rect 20732 2370 20744 8346
rect 20686 2358 20744 2370
rect 20844 8346 20902 8358
rect 20844 2370 20856 8346
rect 20890 2370 20902 8346
rect 20844 2358 20902 2370
rect 21002 8346 21060 8358
rect 21002 2370 21014 8346
rect 21048 2370 21060 8346
rect 21002 2358 21060 2370
rect 21160 8346 21218 8358
rect 21160 2370 21172 8346
rect 21206 2370 21218 8346
rect 21160 2358 21218 2370
rect 21318 8346 21376 8358
rect 21318 2370 21330 8346
rect 21364 2370 21376 8346
rect 21318 2358 21376 2370
rect 21476 8346 21534 8358
rect 21476 2370 21488 8346
rect 21522 2370 21534 8346
rect 21476 2358 21534 2370
rect 21634 8346 21692 8358
rect 21634 2370 21646 8346
rect 21680 2370 21692 8346
rect 21634 2358 21692 2370
rect 21792 8346 21850 8358
rect 21792 2370 21804 8346
rect 21838 2370 21850 8346
rect 21792 2358 21850 2370
rect 21950 8346 22008 8358
rect 21950 2370 21962 8346
rect 21996 2370 22008 8346
rect 21950 2358 22008 2370
rect 22108 8346 22166 8358
rect 22108 2370 22120 8346
rect 22154 2370 22166 8346
rect 22108 2358 22166 2370
rect 22266 8346 22324 8358
rect 22266 2370 22278 8346
rect 22312 2370 22324 8346
rect 22266 2358 22324 2370
rect 22424 8346 22482 8358
rect 22424 2370 22436 8346
rect 22470 2370 22482 8346
rect 22424 2358 22482 2370
rect 22582 8346 22640 8358
rect 22582 2370 22594 8346
rect 22628 2370 22640 8346
rect 22582 2358 22640 2370
rect 22740 8346 22798 8358
rect 22740 2370 22752 8346
rect 22786 2370 22798 8346
rect 22740 2358 22798 2370
rect 22898 8346 22956 8358
rect 22898 2370 22910 8346
rect 22944 2370 22956 8346
rect 22898 2358 22956 2370
rect 23056 8346 23114 8358
rect 23056 2370 23068 8346
rect 23102 2370 23114 8346
rect 23056 2358 23114 2370
rect 23214 8346 23272 8358
rect 23214 2370 23226 8346
rect 23260 2370 23272 8346
rect 23214 2358 23272 2370
rect 23372 8346 23430 8358
rect 23372 2370 23384 8346
rect 23418 2370 23430 8346
rect 23372 2358 23430 2370
rect 23530 8346 23588 8358
rect 23530 2370 23542 8346
rect 23576 2370 23588 8346
rect 23530 2358 23588 2370
rect 23688 8346 23746 8358
rect 23688 2370 23700 8346
rect 23734 2370 23746 8346
rect 23688 2358 23746 2370
rect 23846 8346 23904 8358
rect 23846 2370 23858 8346
rect 23892 2370 23904 8346
rect 23846 2358 23904 2370
rect 24004 8346 24062 8358
rect 24004 2370 24016 8346
rect 24050 2370 24062 8346
rect 24004 2358 24062 2370
rect 24162 8346 24220 8358
rect 24162 2370 24174 8346
rect 24208 2370 24220 8346
rect 24162 2358 24220 2370
rect 24320 8346 24378 8358
rect 24320 2370 24332 8346
rect 24366 2370 24378 8346
rect 24320 2358 24378 2370
rect 24478 8346 24536 8358
rect 24478 2370 24490 8346
rect 24524 2370 24536 8346
rect 24478 2358 24536 2370
rect 24636 8346 24694 8358
rect 24636 2370 24648 8346
rect 24682 2370 24694 8346
rect 24636 2358 24694 2370
rect 24794 8346 24852 8358
rect 24794 2370 24806 8346
rect 24840 2370 24852 8346
rect 24794 2358 24852 2370
rect 24952 8346 25010 8358
rect 24952 2370 24964 8346
rect 24998 2370 25010 8346
rect 24952 2358 25010 2370
rect 25110 8346 25168 8358
rect 25110 2370 25122 8346
rect 25156 2370 25168 8346
rect 25110 2358 25168 2370
<< mvndiffc >>
rect 1482 39970 1516 45946
rect 1640 39970 1674 45946
rect 1798 39970 1832 45946
rect 1956 39970 1990 45946
rect 2114 39970 2148 45946
rect 2272 39970 2306 45946
rect 2430 39970 2464 45946
rect 2588 39970 2622 45946
rect 2746 39970 2780 45946
rect 2904 39970 2938 45946
rect 3062 39970 3096 45946
rect 3220 39970 3254 45946
rect 3378 39970 3412 45946
rect 3536 39970 3570 45946
rect 3694 39970 3728 45946
rect 3852 39970 3886 45946
rect 4010 39970 4044 45946
rect 4168 39970 4202 45946
rect 4326 39970 4360 45946
rect 4484 39970 4518 45946
rect 4642 39970 4676 45946
rect 4800 39970 4834 45946
rect 4958 39970 4992 45946
rect 5116 39970 5150 45946
rect 5274 39970 5308 45946
rect 5432 39970 5466 45946
rect 5590 39970 5624 45946
rect 5748 39970 5782 45946
rect 5906 39970 5940 45946
rect 6064 39970 6098 45946
rect 6222 39970 6256 45946
rect 7782 39970 7816 45946
rect 7940 39970 7974 45946
rect 8098 39970 8132 45946
rect 8256 39970 8290 45946
rect 8414 39970 8448 45946
rect 8572 39970 8606 45946
rect 8730 39970 8764 45946
rect 8888 39970 8922 45946
rect 9046 39970 9080 45946
rect 9204 39970 9238 45946
rect 9362 39970 9396 45946
rect 9520 39970 9554 45946
rect 9678 39970 9712 45946
rect 9836 39970 9870 45946
rect 9994 39970 10028 45946
rect 10152 39970 10186 45946
rect 10310 39970 10344 45946
rect 10468 39970 10502 45946
rect 10626 39970 10660 45946
rect 10784 39970 10818 45946
rect 10942 39970 10976 45946
rect 11100 39970 11134 45946
rect 11258 39970 11292 45946
rect 11416 39970 11450 45946
rect 11574 39970 11608 45946
rect 11732 39970 11766 45946
rect 11890 39970 11924 45946
rect 12048 39970 12082 45946
rect 12206 39970 12240 45946
rect 12364 39970 12398 45946
rect 12522 39970 12556 45946
rect 14082 39970 14116 45946
rect 14240 39970 14274 45946
rect 14398 39970 14432 45946
rect 14556 39970 14590 45946
rect 14714 39970 14748 45946
rect 14872 39970 14906 45946
rect 15030 39970 15064 45946
rect 15188 39970 15222 45946
rect 15346 39970 15380 45946
rect 15504 39970 15538 45946
rect 15662 39970 15696 45946
rect 15820 39970 15854 45946
rect 15978 39970 16012 45946
rect 16136 39970 16170 45946
rect 16294 39970 16328 45946
rect 16452 39970 16486 45946
rect 16610 39970 16644 45946
rect 16768 39970 16802 45946
rect 16926 39970 16960 45946
rect 17084 39970 17118 45946
rect 17242 39970 17276 45946
rect 17400 39970 17434 45946
rect 17558 39970 17592 45946
rect 17716 39970 17750 45946
rect 17874 39970 17908 45946
rect 18032 39970 18066 45946
rect 18190 39970 18224 45946
rect 18348 39970 18382 45946
rect 18506 39970 18540 45946
rect 18664 39970 18698 45946
rect 18822 39970 18856 45946
rect 20382 39970 20416 45946
rect 20540 39970 20574 45946
rect 20698 39970 20732 45946
rect 20856 39970 20890 45946
rect 21014 39970 21048 45946
rect 21172 39970 21206 45946
rect 21330 39970 21364 45946
rect 21488 39970 21522 45946
rect 21646 39970 21680 45946
rect 21804 39970 21838 45946
rect 21962 39970 21996 45946
rect 22120 39970 22154 45946
rect 22278 39970 22312 45946
rect 22436 39970 22470 45946
rect 22594 39970 22628 45946
rect 22752 39970 22786 45946
rect 22910 39970 22944 45946
rect 23068 39970 23102 45946
rect 23226 39970 23260 45946
rect 23384 39970 23418 45946
rect 23542 39970 23576 45946
rect 23700 39970 23734 45946
rect 23858 39970 23892 45946
rect 24016 39970 24050 45946
rect 24174 39970 24208 45946
rect 24332 39970 24366 45946
rect 24490 39970 24524 45946
rect 24648 39970 24682 45946
rect 24806 39970 24840 45946
rect 24964 39970 24998 45946
rect 25122 39970 25156 45946
rect 1482 32970 1516 38946
rect 1640 32970 1674 38946
rect 1798 32970 1832 38946
rect 1956 32970 1990 38946
rect 2114 32970 2148 38946
rect 2272 32970 2306 38946
rect 2430 32970 2464 38946
rect 2588 32970 2622 38946
rect 2746 32970 2780 38946
rect 2904 32970 2938 38946
rect 3062 32970 3096 38946
rect 3220 32970 3254 38946
rect 3378 32970 3412 38946
rect 3536 32970 3570 38946
rect 3694 32970 3728 38946
rect 3852 32970 3886 38946
rect 4010 32970 4044 38946
rect 4168 32970 4202 38946
rect 4326 32970 4360 38946
rect 4484 32970 4518 38946
rect 4642 32970 4676 38946
rect 4800 32970 4834 38946
rect 4958 32970 4992 38946
rect 5116 32970 5150 38946
rect 5274 32970 5308 38946
rect 5432 32970 5466 38946
rect 5590 32970 5624 38946
rect 5748 32970 5782 38946
rect 5906 32970 5940 38946
rect 6064 32970 6098 38946
rect 6222 32970 6256 38946
rect 7782 32970 7816 38946
rect 7940 32970 7974 38946
rect 8098 32970 8132 38946
rect 8256 32970 8290 38946
rect 8414 32970 8448 38946
rect 8572 32970 8606 38946
rect 8730 32970 8764 38946
rect 8888 32970 8922 38946
rect 9046 32970 9080 38946
rect 9204 32970 9238 38946
rect 9362 32970 9396 38946
rect 9520 32970 9554 38946
rect 9678 32970 9712 38946
rect 9836 32970 9870 38946
rect 9994 32970 10028 38946
rect 10152 32970 10186 38946
rect 10310 32970 10344 38946
rect 10468 32970 10502 38946
rect 10626 32970 10660 38946
rect 10784 32970 10818 38946
rect 10942 32970 10976 38946
rect 11100 32970 11134 38946
rect 11258 32970 11292 38946
rect 11416 32970 11450 38946
rect 11574 32970 11608 38946
rect 11732 32970 11766 38946
rect 11890 32970 11924 38946
rect 12048 32970 12082 38946
rect 12206 32970 12240 38946
rect 12364 32970 12398 38946
rect 12522 32970 12556 38946
rect 14082 32970 14116 38946
rect 14240 32970 14274 38946
rect 14398 32970 14432 38946
rect 14556 32970 14590 38946
rect 14714 32970 14748 38946
rect 14872 32970 14906 38946
rect 15030 32970 15064 38946
rect 15188 32970 15222 38946
rect 15346 32970 15380 38946
rect 15504 32970 15538 38946
rect 15662 32970 15696 38946
rect 15820 32970 15854 38946
rect 15978 32970 16012 38946
rect 16136 32970 16170 38946
rect 16294 32970 16328 38946
rect 16452 32970 16486 38946
rect 16610 32970 16644 38946
rect 16768 32970 16802 38946
rect 16926 32970 16960 38946
rect 17084 32970 17118 38946
rect 17242 32970 17276 38946
rect 17400 32970 17434 38946
rect 17558 32970 17592 38946
rect 17716 32970 17750 38946
rect 17874 32970 17908 38946
rect 18032 32970 18066 38946
rect 18190 32970 18224 38946
rect 18348 32970 18382 38946
rect 18506 32970 18540 38946
rect 18664 32970 18698 38946
rect 18822 32970 18856 38946
rect 20382 32970 20416 38946
rect 20540 32970 20574 38946
rect 20698 32970 20732 38946
rect 20856 32970 20890 38946
rect 21014 32970 21048 38946
rect 21172 32970 21206 38946
rect 21330 32970 21364 38946
rect 21488 32970 21522 38946
rect 21646 32970 21680 38946
rect 21804 32970 21838 38946
rect 21962 32970 21996 38946
rect 22120 32970 22154 38946
rect 22278 32970 22312 38946
rect 22436 32970 22470 38946
rect 22594 32970 22628 38946
rect 22752 32970 22786 38946
rect 22910 32970 22944 38946
rect 23068 32970 23102 38946
rect 23226 32970 23260 38946
rect 23384 32970 23418 38946
rect 23542 32970 23576 38946
rect 23700 32970 23734 38946
rect 23858 32970 23892 38946
rect 24016 32970 24050 38946
rect 24174 32970 24208 38946
rect 24332 32970 24366 38946
rect 24490 32970 24524 38946
rect 24648 32970 24682 38946
rect 24806 32970 24840 38946
rect 24964 32970 24998 38946
rect 25122 32970 25156 38946
rect 1482 24670 1516 30646
rect 1640 24670 1674 30646
rect 1798 24670 1832 30646
rect 1956 24670 1990 30646
rect 2114 24670 2148 30646
rect 2272 24670 2306 30646
rect 2430 24670 2464 30646
rect 2588 24670 2622 30646
rect 2746 24670 2780 30646
rect 2904 24670 2938 30646
rect 3062 24670 3096 30646
rect 3220 24670 3254 30646
rect 3378 24670 3412 30646
rect 3536 24670 3570 30646
rect 3694 24670 3728 30646
rect 3852 24670 3886 30646
rect 4010 24670 4044 30646
rect 4168 24670 4202 30646
rect 4326 24670 4360 30646
rect 4484 24670 4518 30646
rect 4642 24670 4676 30646
rect 4800 24670 4834 30646
rect 4958 24670 4992 30646
rect 5116 24670 5150 30646
rect 5274 24670 5308 30646
rect 5432 24670 5466 30646
rect 5590 24670 5624 30646
rect 5748 24670 5782 30646
rect 5906 24670 5940 30646
rect 6064 24670 6098 30646
rect 6222 24670 6256 30646
rect 7782 24670 7816 30646
rect 7940 24670 7974 30646
rect 8098 24670 8132 30646
rect 8256 24670 8290 30646
rect 8414 24670 8448 30646
rect 8572 24670 8606 30646
rect 8730 24670 8764 30646
rect 8888 24670 8922 30646
rect 9046 24670 9080 30646
rect 9204 24670 9238 30646
rect 9362 24670 9396 30646
rect 9520 24670 9554 30646
rect 9678 24670 9712 30646
rect 9836 24670 9870 30646
rect 9994 24670 10028 30646
rect 10152 24670 10186 30646
rect 10310 24670 10344 30646
rect 10468 24670 10502 30646
rect 10626 24670 10660 30646
rect 10784 24670 10818 30646
rect 10942 24670 10976 30646
rect 11100 24670 11134 30646
rect 11258 24670 11292 30646
rect 11416 24670 11450 30646
rect 11574 24670 11608 30646
rect 11732 24670 11766 30646
rect 11890 24670 11924 30646
rect 12048 24670 12082 30646
rect 12206 24670 12240 30646
rect 12364 24670 12398 30646
rect 12522 24670 12556 30646
rect 14082 24670 14116 30646
rect 14240 24670 14274 30646
rect 14398 24670 14432 30646
rect 14556 24670 14590 30646
rect 14714 24670 14748 30646
rect 14872 24670 14906 30646
rect 15030 24670 15064 30646
rect 15188 24670 15222 30646
rect 15346 24670 15380 30646
rect 15504 24670 15538 30646
rect 15662 24670 15696 30646
rect 15820 24670 15854 30646
rect 15978 24670 16012 30646
rect 16136 24670 16170 30646
rect 16294 24670 16328 30646
rect 16452 24670 16486 30646
rect 16610 24670 16644 30646
rect 16768 24670 16802 30646
rect 16926 24670 16960 30646
rect 17084 24670 17118 30646
rect 17242 24670 17276 30646
rect 17400 24670 17434 30646
rect 17558 24670 17592 30646
rect 17716 24670 17750 30646
rect 17874 24670 17908 30646
rect 18032 24670 18066 30646
rect 18190 24670 18224 30646
rect 18348 24670 18382 30646
rect 18506 24670 18540 30646
rect 18664 24670 18698 30646
rect 18822 24670 18856 30646
rect 20382 24670 20416 30646
rect 20540 24670 20574 30646
rect 20698 24670 20732 30646
rect 20856 24670 20890 30646
rect 21014 24670 21048 30646
rect 21172 24670 21206 30646
rect 21330 24670 21364 30646
rect 21488 24670 21522 30646
rect 21646 24670 21680 30646
rect 21804 24670 21838 30646
rect 21962 24670 21996 30646
rect 22120 24670 22154 30646
rect 22278 24670 22312 30646
rect 22436 24670 22470 30646
rect 22594 24670 22628 30646
rect 22752 24670 22786 30646
rect 22910 24670 22944 30646
rect 23068 24670 23102 30646
rect 23226 24670 23260 30646
rect 23384 24670 23418 30646
rect 23542 24670 23576 30646
rect 23700 24670 23734 30646
rect 23858 24670 23892 30646
rect 24016 24670 24050 30646
rect 24174 24670 24208 30646
rect 24332 24670 24366 30646
rect 24490 24670 24524 30646
rect 24648 24670 24682 30646
rect 24806 24670 24840 30646
rect 24964 24670 24998 30646
rect 25122 24670 25156 30646
rect 1482 17670 1516 23646
rect 1640 17670 1674 23646
rect 1798 17670 1832 23646
rect 1956 17670 1990 23646
rect 2114 17670 2148 23646
rect 2272 17670 2306 23646
rect 2430 17670 2464 23646
rect 2588 17670 2622 23646
rect 2746 17670 2780 23646
rect 2904 17670 2938 23646
rect 3062 17670 3096 23646
rect 3220 17670 3254 23646
rect 3378 17670 3412 23646
rect 3536 17670 3570 23646
rect 3694 17670 3728 23646
rect 3852 17670 3886 23646
rect 4010 17670 4044 23646
rect 4168 17670 4202 23646
rect 4326 17670 4360 23646
rect 4484 17670 4518 23646
rect 4642 17670 4676 23646
rect 4800 17670 4834 23646
rect 4958 17670 4992 23646
rect 5116 17670 5150 23646
rect 5274 17670 5308 23646
rect 5432 17670 5466 23646
rect 5590 17670 5624 23646
rect 5748 17670 5782 23646
rect 5906 17670 5940 23646
rect 6064 17670 6098 23646
rect 6222 17670 6256 23646
rect 7782 17670 7816 23646
rect 7940 17670 7974 23646
rect 8098 17670 8132 23646
rect 8256 17670 8290 23646
rect 8414 17670 8448 23646
rect 8572 17670 8606 23646
rect 8730 17670 8764 23646
rect 8888 17670 8922 23646
rect 9046 17670 9080 23646
rect 9204 17670 9238 23646
rect 9362 17670 9396 23646
rect 9520 17670 9554 23646
rect 9678 17670 9712 23646
rect 9836 17670 9870 23646
rect 9994 17670 10028 23646
rect 10152 17670 10186 23646
rect 10310 17670 10344 23646
rect 10468 17670 10502 23646
rect 10626 17670 10660 23646
rect 10784 17670 10818 23646
rect 10942 17670 10976 23646
rect 11100 17670 11134 23646
rect 11258 17670 11292 23646
rect 11416 17670 11450 23646
rect 11574 17670 11608 23646
rect 11732 17670 11766 23646
rect 11890 17670 11924 23646
rect 12048 17670 12082 23646
rect 12206 17670 12240 23646
rect 12364 17670 12398 23646
rect 12522 17670 12556 23646
rect 14082 17670 14116 23646
rect 14240 17670 14274 23646
rect 14398 17670 14432 23646
rect 14556 17670 14590 23646
rect 14714 17670 14748 23646
rect 14872 17670 14906 23646
rect 15030 17670 15064 23646
rect 15188 17670 15222 23646
rect 15346 17670 15380 23646
rect 15504 17670 15538 23646
rect 15662 17670 15696 23646
rect 15820 17670 15854 23646
rect 15978 17670 16012 23646
rect 16136 17670 16170 23646
rect 16294 17670 16328 23646
rect 16452 17670 16486 23646
rect 16610 17670 16644 23646
rect 16768 17670 16802 23646
rect 16926 17670 16960 23646
rect 17084 17670 17118 23646
rect 17242 17670 17276 23646
rect 17400 17670 17434 23646
rect 17558 17670 17592 23646
rect 17716 17670 17750 23646
rect 17874 17670 17908 23646
rect 18032 17670 18066 23646
rect 18190 17670 18224 23646
rect 18348 17670 18382 23646
rect 18506 17670 18540 23646
rect 18664 17670 18698 23646
rect 18822 17670 18856 23646
rect 20382 17670 20416 23646
rect 20540 17670 20574 23646
rect 20698 17670 20732 23646
rect 20856 17670 20890 23646
rect 21014 17670 21048 23646
rect 21172 17670 21206 23646
rect 21330 17670 21364 23646
rect 21488 17670 21522 23646
rect 21646 17670 21680 23646
rect 21804 17670 21838 23646
rect 21962 17670 21996 23646
rect 22120 17670 22154 23646
rect 22278 17670 22312 23646
rect 22436 17670 22470 23646
rect 22594 17670 22628 23646
rect 22752 17670 22786 23646
rect 22910 17670 22944 23646
rect 23068 17670 23102 23646
rect 23226 17670 23260 23646
rect 23384 17670 23418 23646
rect 23542 17670 23576 23646
rect 23700 17670 23734 23646
rect 23858 17670 23892 23646
rect 24016 17670 24050 23646
rect 24174 17670 24208 23646
rect 24332 17670 24366 23646
rect 24490 17670 24524 23646
rect 24648 17670 24682 23646
rect 24806 17670 24840 23646
rect 24964 17670 24998 23646
rect 25122 17670 25156 23646
rect 1482 9370 1516 15346
rect 1640 9370 1674 15346
rect 1798 9370 1832 15346
rect 1956 9370 1990 15346
rect 2114 9370 2148 15346
rect 2272 9370 2306 15346
rect 2430 9370 2464 15346
rect 2588 9370 2622 15346
rect 2746 9370 2780 15346
rect 2904 9370 2938 15346
rect 3062 9370 3096 15346
rect 3220 9370 3254 15346
rect 3378 9370 3412 15346
rect 3536 9370 3570 15346
rect 3694 9370 3728 15346
rect 3852 9370 3886 15346
rect 4010 9370 4044 15346
rect 4168 9370 4202 15346
rect 4326 9370 4360 15346
rect 4484 9370 4518 15346
rect 4642 9370 4676 15346
rect 4800 9370 4834 15346
rect 4958 9370 4992 15346
rect 5116 9370 5150 15346
rect 5274 9370 5308 15346
rect 5432 9370 5466 15346
rect 5590 9370 5624 15346
rect 5748 9370 5782 15346
rect 5906 9370 5940 15346
rect 6064 9370 6098 15346
rect 6222 9370 6256 15346
rect 7782 9370 7816 15346
rect 7940 9370 7974 15346
rect 8098 9370 8132 15346
rect 8256 9370 8290 15346
rect 8414 9370 8448 15346
rect 8572 9370 8606 15346
rect 8730 9370 8764 15346
rect 8888 9370 8922 15346
rect 9046 9370 9080 15346
rect 9204 9370 9238 15346
rect 9362 9370 9396 15346
rect 9520 9370 9554 15346
rect 9678 9370 9712 15346
rect 9836 9370 9870 15346
rect 9994 9370 10028 15346
rect 10152 9370 10186 15346
rect 10310 9370 10344 15346
rect 10468 9370 10502 15346
rect 10626 9370 10660 15346
rect 10784 9370 10818 15346
rect 10942 9370 10976 15346
rect 11100 9370 11134 15346
rect 11258 9370 11292 15346
rect 11416 9370 11450 15346
rect 11574 9370 11608 15346
rect 11732 9370 11766 15346
rect 11890 9370 11924 15346
rect 12048 9370 12082 15346
rect 12206 9370 12240 15346
rect 12364 9370 12398 15346
rect 12522 9370 12556 15346
rect 14082 9370 14116 15346
rect 14240 9370 14274 15346
rect 14398 9370 14432 15346
rect 14556 9370 14590 15346
rect 14714 9370 14748 15346
rect 14872 9370 14906 15346
rect 15030 9370 15064 15346
rect 15188 9370 15222 15346
rect 15346 9370 15380 15346
rect 15504 9370 15538 15346
rect 15662 9370 15696 15346
rect 15820 9370 15854 15346
rect 15978 9370 16012 15346
rect 16136 9370 16170 15346
rect 16294 9370 16328 15346
rect 16452 9370 16486 15346
rect 16610 9370 16644 15346
rect 16768 9370 16802 15346
rect 16926 9370 16960 15346
rect 17084 9370 17118 15346
rect 17242 9370 17276 15346
rect 17400 9370 17434 15346
rect 17558 9370 17592 15346
rect 17716 9370 17750 15346
rect 17874 9370 17908 15346
rect 18032 9370 18066 15346
rect 18190 9370 18224 15346
rect 18348 9370 18382 15346
rect 18506 9370 18540 15346
rect 18664 9370 18698 15346
rect 18822 9370 18856 15346
rect 20382 9370 20416 15346
rect 20540 9370 20574 15346
rect 20698 9370 20732 15346
rect 20856 9370 20890 15346
rect 21014 9370 21048 15346
rect 21172 9370 21206 15346
rect 21330 9370 21364 15346
rect 21488 9370 21522 15346
rect 21646 9370 21680 15346
rect 21804 9370 21838 15346
rect 21962 9370 21996 15346
rect 22120 9370 22154 15346
rect 22278 9370 22312 15346
rect 22436 9370 22470 15346
rect 22594 9370 22628 15346
rect 22752 9370 22786 15346
rect 22910 9370 22944 15346
rect 23068 9370 23102 15346
rect 23226 9370 23260 15346
rect 23384 9370 23418 15346
rect 23542 9370 23576 15346
rect 23700 9370 23734 15346
rect 23858 9370 23892 15346
rect 24016 9370 24050 15346
rect 24174 9370 24208 15346
rect 24332 9370 24366 15346
rect 24490 9370 24524 15346
rect 24648 9370 24682 15346
rect 24806 9370 24840 15346
rect 24964 9370 24998 15346
rect 25122 9370 25156 15346
rect 1482 2370 1516 8346
rect 1640 2370 1674 8346
rect 1798 2370 1832 8346
rect 1956 2370 1990 8346
rect 2114 2370 2148 8346
rect 2272 2370 2306 8346
rect 2430 2370 2464 8346
rect 2588 2370 2622 8346
rect 2746 2370 2780 8346
rect 2904 2370 2938 8346
rect 3062 2370 3096 8346
rect 3220 2370 3254 8346
rect 3378 2370 3412 8346
rect 3536 2370 3570 8346
rect 3694 2370 3728 8346
rect 3852 2370 3886 8346
rect 4010 2370 4044 8346
rect 4168 2370 4202 8346
rect 4326 2370 4360 8346
rect 4484 2370 4518 8346
rect 4642 2370 4676 8346
rect 4800 2370 4834 8346
rect 4958 2370 4992 8346
rect 5116 2370 5150 8346
rect 5274 2370 5308 8346
rect 5432 2370 5466 8346
rect 5590 2370 5624 8346
rect 5748 2370 5782 8346
rect 5906 2370 5940 8346
rect 6064 2370 6098 8346
rect 6222 2370 6256 8346
rect 7782 2370 7816 8346
rect 7940 2370 7974 8346
rect 8098 2370 8132 8346
rect 8256 2370 8290 8346
rect 8414 2370 8448 8346
rect 8572 2370 8606 8346
rect 8730 2370 8764 8346
rect 8888 2370 8922 8346
rect 9046 2370 9080 8346
rect 9204 2370 9238 8346
rect 9362 2370 9396 8346
rect 9520 2370 9554 8346
rect 9678 2370 9712 8346
rect 9836 2370 9870 8346
rect 9994 2370 10028 8346
rect 10152 2370 10186 8346
rect 10310 2370 10344 8346
rect 10468 2370 10502 8346
rect 10626 2370 10660 8346
rect 10784 2370 10818 8346
rect 10942 2370 10976 8346
rect 11100 2370 11134 8346
rect 11258 2370 11292 8346
rect 11416 2370 11450 8346
rect 11574 2370 11608 8346
rect 11732 2370 11766 8346
rect 11890 2370 11924 8346
rect 12048 2370 12082 8346
rect 12206 2370 12240 8346
rect 12364 2370 12398 8346
rect 12522 2370 12556 8346
rect 14082 2370 14116 8346
rect 14240 2370 14274 8346
rect 14398 2370 14432 8346
rect 14556 2370 14590 8346
rect 14714 2370 14748 8346
rect 14872 2370 14906 8346
rect 15030 2370 15064 8346
rect 15188 2370 15222 8346
rect 15346 2370 15380 8346
rect 15504 2370 15538 8346
rect 15662 2370 15696 8346
rect 15820 2370 15854 8346
rect 15978 2370 16012 8346
rect 16136 2370 16170 8346
rect 16294 2370 16328 8346
rect 16452 2370 16486 8346
rect 16610 2370 16644 8346
rect 16768 2370 16802 8346
rect 16926 2370 16960 8346
rect 17084 2370 17118 8346
rect 17242 2370 17276 8346
rect 17400 2370 17434 8346
rect 17558 2370 17592 8346
rect 17716 2370 17750 8346
rect 17874 2370 17908 8346
rect 18032 2370 18066 8346
rect 18190 2370 18224 8346
rect 18348 2370 18382 8346
rect 18506 2370 18540 8346
rect 18664 2370 18698 8346
rect 18822 2370 18856 8346
rect 20382 2370 20416 8346
rect 20540 2370 20574 8346
rect 20698 2370 20732 8346
rect 20856 2370 20890 8346
rect 21014 2370 21048 8346
rect 21172 2370 21206 8346
rect 21330 2370 21364 8346
rect 21488 2370 21522 8346
rect 21646 2370 21680 8346
rect 21804 2370 21838 8346
rect 21962 2370 21996 8346
rect 22120 2370 22154 8346
rect 22278 2370 22312 8346
rect 22436 2370 22470 8346
rect 22594 2370 22628 8346
rect 22752 2370 22786 8346
rect 22910 2370 22944 8346
rect 23068 2370 23102 8346
rect 23226 2370 23260 8346
rect 23384 2370 23418 8346
rect 23542 2370 23576 8346
rect 23700 2370 23734 8346
rect 23858 2370 23892 8346
rect 24016 2370 24050 8346
rect 24174 2370 24208 8346
rect 24332 2370 24366 8346
rect 24490 2370 24524 8346
rect 24648 2370 24682 8346
rect 24806 2370 24840 8346
rect 24964 2370 24998 8346
rect 25122 2370 25156 8346
<< psubdiff >>
rect -3364 40388 -3268 40422
rect -3134 40388 -3038 40422
rect -3364 40326 -3330 40388
rect -3072 40326 -3038 40388
rect -3364 38750 -3330 38812
rect 29838 40388 29934 40422
rect 30068 40388 30164 40422
rect 29838 40326 29872 40388
rect -3072 38750 -3038 38812
rect -3364 38716 -3268 38750
rect -3134 38716 -3038 38750
rect 30130 40326 30164 40388
rect 29838 38750 29872 38812
rect 30130 38750 30164 38812
rect 29838 38716 29934 38750
rect 30068 38716 30164 38750
rect -4364 27188 -4268 27222
rect -4134 27188 -4038 27222
rect -4364 27126 -4330 27188
rect -4072 27126 -4038 27188
rect -4364 25550 -4330 25612
rect -4072 25550 -4038 25612
rect -4364 25516 -4268 25550
rect -4134 25516 -4038 25550
rect 30838 27188 30934 27222
rect 31068 27188 31164 27222
rect 30838 27126 30872 27188
rect 31130 27126 31164 27188
rect 30838 25550 30872 25612
rect 31130 25550 31164 25612
rect 30838 25516 30934 25550
rect 31068 25516 31164 25550
rect -4364 13946 -4268 13980
rect -4130 13946 -4034 13980
rect -4364 13884 -4330 13946
rect -4068 13884 -4034 13946
rect -4364 12570 -4330 12632
rect -4068 12570 -4034 12632
rect -4364 12536 -4268 12570
rect -4130 12536 -4034 12570
rect 30834 13946 30930 13980
rect 31068 13946 31164 13980
rect 30834 13884 30868 13946
rect 31130 13884 31164 13946
rect 30834 12570 30868 12632
rect 31130 12570 31164 12632
rect 30834 12536 30930 12570
rect 31068 12536 31164 12570
<< mvpsubdiff >>
rect 1336 46168 6402 46180
rect 1336 46134 1444 46168
rect 6294 46134 6402 46168
rect 1336 46122 6402 46134
rect 1336 46072 1394 46122
rect 1336 39844 1348 46072
rect 1382 39844 1394 46072
rect 6344 46072 6402 46122
rect 1336 39794 1394 39844
rect 6344 39844 6356 46072
rect 6390 39844 6402 46072
rect 6344 39794 6402 39844
rect 1336 39782 6402 39794
rect 1336 39748 1444 39782
rect 6294 39748 6402 39782
rect 1336 39736 6402 39748
rect 7636 46168 12702 46180
rect 7636 46134 7744 46168
rect 12594 46134 12702 46168
rect 7636 46122 12702 46134
rect 7636 46072 7694 46122
rect 7636 39844 7648 46072
rect 7682 39844 7694 46072
rect 12644 46072 12702 46122
rect 7636 39794 7694 39844
rect 12644 39844 12656 46072
rect 12690 39844 12702 46072
rect 12644 39794 12702 39844
rect 7636 39782 12702 39794
rect 7636 39748 7744 39782
rect 12594 39748 12702 39782
rect 7636 39736 12702 39748
rect 13936 46168 19002 46180
rect 13936 46134 14044 46168
rect 18894 46134 19002 46168
rect 13936 46122 19002 46134
rect 13936 46072 13994 46122
rect 13936 39844 13948 46072
rect 13982 39844 13994 46072
rect 18944 46072 19002 46122
rect 13936 39794 13994 39844
rect 18944 39844 18956 46072
rect 18990 39844 19002 46072
rect 18944 39794 19002 39844
rect 13936 39782 19002 39794
rect 13936 39748 14044 39782
rect 18894 39748 19002 39782
rect 13936 39736 19002 39748
rect 20236 46168 25302 46180
rect 20236 46134 20344 46168
rect 25194 46134 25302 46168
rect 20236 46122 25302 46134
rect 20236 46072 20294 46122
rect 20236 39844 20248 46072
rect 20282 39844 20294 46072
rect 25244 46072 25302 46122
rect 20236 39794 20294 39844
rect 25244 39844 25256 46072
rect 25290 39844 25302 46072
rect 25244 39794 25302 39844
rect 20236 39782 25302 39794
rect 20236 39748 20344 39782
rect 25194 39748 25302 39782
rect 20236 39736 25302 39748
rect 1336 39168 6402 39180
rect 1336 39134 1444 39168
rect 6294 39134 6402 39168
rect 1336 39122 6402 39134
rect 1336 39072 1394 39122
rect 1336 32844 1348 39072
rect 1382 32844 1394 39072
rect 6344 39072 6402 39122
rect 1336 32794 1394 32844
rect 6344 32844 6356 39072
rect 6390 32844 6402 39072
rect 6344 32794 6402 32844
rect 1336 32782 6402 32794
rect 1336 32748 1444 32782
rect 6294 32748 6402 32782
rect 1336 32736 6402 32748
rect 7636 39168 12702 39180
rect 7636 39134 7744 39168
rect 12594 39134 12702 39168
rect 7636 39122 12702 39134
rect 7636 39072 7694 39122
rect 7636 32844 7648 39072
rect 7682 32844 7694 39072
rect 12644 39072 12702 39122
rect 7636 32794 7694 32844
rect 12644 32844 12656 39072
rect 12690 32844 12702 39072
rect 12644 32794 12702 32844
rect 7636 32782 12702 32794
rect 7636 32748 7744 32782
rect 12594 32748 12702 32782
rect 7636 32736 12702 32748
rect 13936 39168 19002 39180
rect 13936 39134 14044 39168
rect 18894 39134 19002 39168
rect 13936 39122 19002 39134
rect 13936 39072 13994 39122
rect 13936 32844 13948 39072
rect 13982 32844 13994 39072
rect 18944 39072 19002 39122
rect 13936 32794 13994 32844
rect 18944 32844 18956 39072
rect 18990 32844 19002 39072
rect 18944 32794 19002 32844
rect 13936 32782 19002 32794
rect 13936 32748 14044 32782
rect 18894 32748 19002 32782
rect 13936 32736 19002 32748
rect 20236 39168 25302 39180
rect 20236 39134 20344 39168
rect 25194 39134 25302 39168
rect 20236 39122 25302 39134
rect 20236 39072 20294 39122
rect 20236 32844 20248 39072
rect 20282 32844 20294 39072
rect 25244 39072 25302 39122
rect 20236 32794 20294 32844
rect 25244 32844 25256 39072
rect 25290 32844 25302 39072
rect 25244 32794 25302 32844
rect 20236 32782 25302 32794
rect 20236 32748 20344 32782
rect 25194 32748 25302 32782
rect 20236 32736 25302 32748
rect 1336 30868 6402 30880
rect 1336 30834 1444 30868
rect 6294 30834 6402 30868
rect 1336 30822 6402 30834
rect 1336 30772 1394 30822
rect 1336 24544 1348 30772
rect 1382 24544 1394 30772
rect 6344 30772 6402 30822
rect 1336 24494 1394 24544
rect 6344 24544 6356 30772
rect 6390 24544 6402 30772
rect 6344 24494 6402 24544
rect 1336 24482 6402 24494
rect 1336 24448 1444 24482
rect 6294 24448 6402 24482
rect 1336 24436 6402 24448
rect 7636 30868 12702 30880
rect 7636 30834 7744 30868
rect 12594 30834 12702 30868
rect 7636 30822 12702 30834
rect 7636 30772 7694 30822
rect 7636 24544 7648 30772
rect 7682 24544 7694 30772
rect 12644 30772 12702 30822
rect 7636 24494 7694 24544
rect 12644 24544 12656 30772
rect 12690 24544 12702 30772
rect 12644 24494 12702 24544
rect 7636 24482 12702 24494
rect 7636 24448 7744 24482
rect 12594 24448 12702 24482
rect 7636 24436 12702 24448
rect 13936 30868 19002 30880
rect 13936 30834 14044 30868
rect 18894 30834 19002 30868
rect 13936 30822 19002 30834
rect 13936 30772 13994 30822
rect 13936 24544 13948 30772
rect 13982 24544 13994 30772
rect 18944 30772 19002 30822
rect 13936 24494 13994 24544
rect 18944 24544 18956 30772
rect 18990 24544 19002 30772
rect 18944 24494 19002 24544
rect 13936 24482 19002 24494
rect 13936 24448 14044 24482
rect 18894 24448 19002 24482
rect 13936 24436 19002 24448
rect 20236 30868 25302 30880
rect 20236 30834 20344 30868
rect 25194 30834 25302 30868
rect 20236 30822 25302 30834
rect 20236 30772 20294 30822
rect 20236 24544 20248 30772
rect 20282 24544 20294 30772
rect 25244 30772 25302 30822
rect 20236 24494 20294 24544
rect 25244 24544 25256 30772
rect 25290 24544 25302 30772
rect 25244 24494 25302 24544
rect 20236 24482 25302 24494
rect 20236 24448 20344 24482
rect 25194 24448 25302 24482
rect 20236 24436 25302 24448
rect 1336 23868 6402 23880
rect 1336 23834 1444 23868
rect 6294 23834 6402 23868
rect 1336 23822 6402 23834
rect 1336 23772 1394 23822
rect 1336 17544 1348 23772
rect 1382 17544 1394 23772
rect 6344 23772 6402 23822
rect 1336 17494 1394 17544
rect 6344 17544 6356 23772
rect 6390 17544 6402 23772
rect 6344 17494 6402 17544
rect 1336 17482 6402 17494
rect 1336 17448 1444 17482
rect 6294 17448 6402 17482
rect 1336 17436 6402 17448
rect 7636 23868 12702 23880
rect 7636 23834 7744 23868
rect 12594 23834 12702 23868
rect 7636 23822 12702 23834
rect 7636 23772 7694 23822
rect 7636 17544 7648 23772
rect 7682 17544 7694 23772
rect 12644 23772 12702 23822
rect 7636 17494 7694 17544
rect 12644 17544 12656 23772
rect 12690 17544 12702 23772
rect 12644 17494 12702 17544
rect 7636 17482 12702 17494
rect 7636 17448 7744 17482
rect 12594 17448 12702 17482
rect 7636 17436 12702 17448
rect 13936 23868 19002 23880
rect 13936 23834 14044 23868
rect 18894 23834 19002 23868
rect 13936 23822 19002 23834
rect 13936 23772 13994 23822
rect 13936 17544 13948 23772
rect 13982 17544 13994 23772
rect 18944 23772 19002 23822
rect 13936 17494 13994 17544
rect 18944 17544 18956 23772
rect 18990 17544 19002 23772
rect 18944 17494 19002 17544
rect 13936 17482 19002 17494
rect 13936 17448 14044 17482
rect 18894 17448 19002 17482
rect 13936 17436 19002 17448
rect 20236 23868 25302 23880
rect 20236 23834 20344 23868
rect 25194 23834 25302 23868
rect 20236 23822 25302 23834
rect 20236 23772 20294 23822
rect 20236 17544 20248 23772
rect 20282 17544 20294 23772
rect 25244 23772 25302 23822
rect 20236 17494 20294 17544
rect 25244 17544 25256 23772
rect 25290 17544 25302 23772
rect 25244 17494 25302 17544
rect 20236 17482 25302 17494
rect 20236 17448 20344 17482
rect 25194 17448 25302 17482
rect 20236 17436 25302 17448
rect 1336 15568 6402 15580
rect 1336 15534 1444 15568
rect 6294 15534 6402 15568
rect 1336 15522 6402 15534
rect 1336 15472 1394 15522
rect 1336 9244 1348 15472
rect 1382 9244 1394 15472
rect 6344 15472 6402 15522
rect 1336 9194 1394 9244
rect 6344 9244 6356 15472
rect 6390 9244 6402 15472
rect 6344 9194 6402 9244
rect 1336 9182 6402 9194
rect 1336 9148 1444 9182
rect 6294 9148 6402 9182
rect 1336 9136 6402 9148
rect 7636 15568 12702 15580
rect 7636 15534 7744 15568
rect 12594 15534 12702 15568
rect 7636 15522 12702 15534
rect 7636 15472 7694 15522
rect 7636 9244 7648 15472
rect 7682 9244 7694 15472
rect 12644 15472 12702 15522
rect 7636 9194 7694 9244
rect 12644 9244 12656 15472
rect 12690 9244 12702 15472
rect 12644 9194 12702 9244
rect 7636 9182 12702 9194
rect 7636 9148 7744 9182
rect 12594 9148 12702 9182
rect 7636 9136 12702 9148
rect 13936 15568 19002 15580
rect 13936 15534 14044 15568
rect 18894 15534 19002 15568
rect 13936 15522 19002 15534
rect 13936 15472 13994 15522
rect 13936 9244 13948 15472
rect 13982 9244 13994 15472
rect 18944 15472 19002 15522
rect 13936 9194 13994 9244
rect 18944 9244 18956 15472
rect 18990 9244 19002 15472
rect 18944 9194 19002 9244
rect 13936 9182 19002 9194
rect 13936 9148 14044 9182
rect 18894 9148 19002 9182
rect 13936 9136 19002 9148
rect 20236 15568 25302 15580
rect 20236 15534 20344 15568
rect 25194 15534 25302 15568
rect 20236 15522 25302 15534
rect 20236 15472 20294 15522
rect 20236 9244 20248 15472
rect 20282 9244 20294 15472
rect 25244 15472 25302 15522
rect 20236 9194 20294 9244
rect 25244 9244 25256 15472
rect 25290 9244 25302 15472
rect 25244 9194 25302 9244
rect 20236 9182 25302 9194
rect 20236 9148 20344 9182
rect 25194 9148 25302 9182
rect 20236 9136 25302 9148
rect 1336 8568 6402 8580
rect 1336 8534 1444 8568
rect 6294 8534 6402 8568
rect 1336 8522 6402 8534
rect 1336 8472 1394 8522
rect 1336 2244 1348 8472
rect 1382 2244 1394 8472
rect 6344 8472 6402 8522
rect 1336 2194 1394 2244
rect 6344 2244 6356 8472
rect 6390 2244 6402 8472
rect 6344 2194 6402 2244
rect 1336 2182 6402 2194
rect 1336 2148 1444 2182
rect 6294 2148 6402 2182
rect 1336 2136 6402 2148
rect 7636 8568 12702 8580
rect 7636 8534 7744 8568
rect 12594 8534 12702 8568
rect 7636 8522 12702 8534
rect 7636 8472 7694 8522
rect 7636 2244 7648 8472
rect 7682 2244 7694 8472
rect 12644 8472 12702 8522
rect 7636 2194 7694 2244
rect 12644 2244 12656 8472
rect 12690 2244 12702 8472
rect 12644 2194 12702 2244
rect 7636 2182 12702 2194
rect 7636 2148 7744 2182
rect 12594 2148 12702 2182
rect 7636 2136 12702 2148
rect 13936 8568 19002 8580
rect 13936 8534 14044 8568
rect 18894 8534 19002 8568
rect 13936 8522 19002 8534
rect 13936 8472 13994 8522
rect 13936 2244 13948 8472
rect 13982 2244 13994 8472
rect 18944 8472 19002 8522
rect 13936 2194 13994 2244
rect 18944 2244 18956 8472
rect 18990 2244 19002 8472
rect 18944 2194 19002 2244
rect 13936 2182 19002 2194
rect 13936 2148 14044 2182
rect 18894 2148 19002 2182
rect 13936 2136 19002 2148
rect 20236 8568 25302 8580
rect 20236 8534 20344 8568
rect 25194 8534 25302 8568
rect 20236 8522 25302 8534
rect 20236 8472 20294 8522
rect 20236 2244 20248 8472
rect 20282 2244 20294 8472
rect 25244 8472 25302 8522
rect 20236 2194 20294 2244
rect 25244 2244 25256 8472
rect 25290 2244 25302 8472
rect 25244 2194 25302 2244
rect 20236 2182 25302 2194
rect 20236 2148 20344 2182
rect 25194 2148 25302 2182
rect 20236 2136 25302 2148
<< psubdiffcont >>
rect -3268 40388 -3134 40422
rect -3364 38812 -3330 40326
rect -3072 38812 -3038 40326
rect 29934 40388 30068 40422
rect -3268 38716 -3134 38750
rect 29838 38812 29872 40326
rect 30130 38812 30164 40326
rect 29934 38716 30068 38750
rect -4268 27188 -4134 27222
rect -4364 25612 -4330 27126
rect -4072 25612 -4038 27126
rect -4268 25516 -4134 25550
rect 30934 27188 31068 27222
rect 30838 25612 30872 27126
rect 31130 25612 31164 27126
rect 30934 25516 31068 25550
rect -4268 13946 -4130 13980
rect -4364 12632 -4330 13884
rect -4068 12632 -4034 13884
rect -4268 12536 -4130 12570
rect 30930 13946 31068 13980
rect 30834 12632 30868 13884
rect 31130 12632 31164 13884
rect 30930 12536 31068 12570
<< mvpsubdiffcont >>
rect 1444 46134 6294 46168
rect 1348 39844 1382 46072
rect 6356 39844 6390 46072
rect 1444 39748 6294 39782
rect 7744 46134 12594 46168
rect 7648 39844 7682 46072
rect 12656 39844 12690 46072
rect 7744 39748 12594 39782
rect 14044 46134 18894 46168
rect 13948 39844 13982 46072
rect 18956 39844 18990 46072
rect 14044 39748 18894 39782
rect 20344 46134 25194 46168
rect 20248 39844 20282 46072
rect 25256 39844 25290 46072
rect 20344 39748 25194 39782
rect 1444 39134 6294 39168
rect 1348 32844 1382 39072
rect 6356 32844 6390 39072
rect 1444 32748 6294 32782
rect 7744 39134 12594 39168
rect 7648 32844 7682 39072
rect 12656 32844 12690 39072
rect 7744 32748 12594 32782
rect 14044 39134 18894 39168
rect 13948 32844 13982 39072
rect 18956 32844 18990 39072
rect 14044 32748 18894 32782
rect 20344 39134 25194 39168
rect 20248 32844 20282 39072
rect 25256 32844 25290 39072
rect 20344 32748 25194 32782
rect 1444 30834 6294 30868
rect 1348 24544 1382 30772
rect 6356 24544 6390 30772
rect 1444 24448 6294 24482
rect 7744 30834 12594 30868
rect 7648 24544 7682 30772
rect 12656 24544 12690 30772
rect 7744 24448 12594 24482
rect 14044 30834 18894 30868
rect 13948 24544 13982 30772
rect 18956 24544 18990 30772
rect 14044 24448 18894 24482
rect 20344 30834 25194 30868
rect 20248 24544 20282 30772
rect 25256 24544 25290 30772
rect 20344 24448 25194 24482
rect 1444 23834 6294 23868
rect 1348 17544 1382 23772
rect 6356 17544 6390 23772
rect 1444 17448 6294 17482
rect 7744 23834 12594 23868
rect 7648 17544 7682 23772
rect 12656 17544 12690 23772
rect 7744 17448 12594 17482
rect 14044 23834 18894 23868
rect 13948 17544 13982 23772
rect 18956 17544 18990 23772
rect 14044 17448 18894 17482
rect 20344 23834 25194 23868
rect 20248 17544 20282 23772
rect 25256 17544 25290 23772
rect 20344 17448 25194 17482
rect 1444 15534 6294 15568
rect 1348 9244 1382 15472
rect 6356 9244 6390 15472
rect 1444 9148 6294 9182
rect 7744 15534 12594 15568
rect 7648 9244 7682 15472
rect 12656 9244 12690 15472
rect 7744 9148 12594 9182
rect 14044 15534 18894 15568
rect 13948 9244 13982 15472
rect 18956 9244 18990 15472
rect 14044 9148 18894 9182
rect 20344 15534 25194 15568
rect 20248 9244 20282 15472
rect 25256 9244 25290 15472
rect 20344 9148 25194 9182
rect 1444 8534 6294 8568
rect 1348 2244 1382 8472
rect 6356 2244 6390 8472
rect 1444 2148 6294 2182
rect 7744 8534 12594 8568
rect 7648 2244 7682 8472
rect 12656 2244 12690 8472
rect 7744 2148 12594 2182
rect 14044 8534 18894 8568
rect 13948 2244 13982 8472
rect 18956 2244 18990 8472
rect 14044 2148 18894 2182
rect 20344 8534 25194 8568
rect 20248 2244 20282 8472
rect 25256 2244 25290 8472
rect 20344 2148 25194 2182
<< poly >>
rect -3234 40276 -3168 40292
rect -3234 40242 -3218 40276
rect -3184 40242 -3168 40276
rect -3234 40219 -3168 40242
rect -3234 38896 -3168 38919
rect -3234 38862 -3218 38896
rect -3184 38862 -3168 38896
rect -3234 38846 -3168 38862
rect 1528 46030 1628 46046
rect 1528 45996 1544 46030
rect 1612 45996 1628 46030
rect 1528 45958 1628 45996
rect 1686 46030 1786 46046
rect 1686 45996 1702 46030
rect 1770 45996 1786 46030
rect 1686 45958 1786 45996
rect 1844 46030 1944 46046
rect 1844 45996 1860 46030
rect 1928 45996 1944 46030
rect 1844 45958 1944 45996
rect 2002 46030 2102 46046
rect 2002 45996 2018 46030
rect 2086 45996 2102 46030
rect 2002 45958 2102 45996
rect 2160 46030 2260 46046
rect 2160 45996 2176 46030
rect 2244 45996 2260 46030
rect 2160 45958 2260 45996
rect 2318 46030 2418 46046
rect 2318 45996 2334 46030
rect 2402 45996 2418 46030
rect 2318 45958 2418 45996
rect 2476 46030 2576 46046
rect 2476 45996 2492 46030
rect 2560 45996 2576 46030
rect 2476 45958 2576 45996
rect 2634 46030 2734 46046
rect 2634 45996 2650 46030
rect 2718 45996 2734 46030
rect 2634 45958 2734 45996
rect 2792 46030 2892 46046
rect 2792 45996 2808 46030
rect 2876 45996 2892 46030
rect 2792 45958 2892 45996
rect 2950 46030 3050 46046
rect 2950 45996 2966 46030
rect 3034 45996 3050 46030
rect 2950 45958 3050 45996
rect 3108 46030 3208 46046
rect 3108 45996 3124 46030
rect 3192 45996 3208 46030
rect 3108 45958 3208 45996
rect 3266 46030 3366 46046
rect 3266 45996 3282 46030
rect 3350 45996 3366 46030
rect 3266 45958 3366 45996
rect 3424 46030 3524 46046
rect 3424 45996 3440 46030
rect 3508 45996 3524 46030
rect 3424 45958 3524 45996
rect 3582 46030 3682 46046
rect 3582 45996 3598 46030
rect 3666 45996 3682 46030
rect 3582 45958 3682 45996
rect 3740 46030 3840 46046
rect 3740 45996 3756 46030
rect 3824 45996 3840 46030
rect 3740 45958 3840 45996
rect 3898 46030 3998 46046
rect 3898 45996 3914 46030
rect 3982 45996 3998 46030
rect 3898 45958 3998 45996
rect 4056 46030 4156 46046
rect 4056 45996 4072 46030
rect 4140 45996 4156 46030
rect 4056 45958 4156 45996
rect 4214 46030 4314 46046
rect 4214 45996 4230 46030
rect 4298 45996 4314 46030
rect 4214 45958 4314 45996
rect 4372 46030 4472 46046
rect 4372 45996 4388 46030
rect 4456 45996 4472 46030
rect 4372 45958 4472 45996
rect 4530 46030 4630 46046
rect 4530 45996 4546 46030
rect 4614 45996 4630 46030
rect 4530 45958 4630 45996
rect 4688 46030 4788 46046
rect 4688 45996 4704 46030
rect 4772 45996 4788 46030
rect 4688 45958 4788 45996
rect 4846 46030 4946 46046
rect 4846 45996 4862 46030
rect 4930 45996 4946 46030
rect 4846 45958 4946 45996
rect 5004 46030 5104 46046
rect 5004 45996 5020 46030
rect 5088 45996 5104 46030
rect 5004 45958 5104 45996
rect 5162 46030 5262 46046
rect 5162 45996 5178 46030
rect 5246 45996 5262 46030
rect 5162 45958 5262 45996
rect 5320 46030 5420 46046
rect 5320 45996 5336 46030
rect 5404 45996 5420 46030
rect 5320 45958 5420 45996
rect 5478 46030 5578 46046
rect 5478 45996 5494 46030
rect 5562 45996 5578 46030
rect 5478 45958 5578 45996
rect 5636 46030 5736 46046
rect 5636 45996 5652 46030
rect 5720 45996 5736 46030
rect 5636 45958 5736 45996
rect 5794 46030 5894 46046
rect 5794 45996 5810 46030
rect 5878 45996 5894 46030
rect 5794 45958 5894 45996
rect 5952 46030 6052 46046
rect 5952 45996 5968 46030
rect 6036 45996 6052 46030
rect 5952 45958 6052 45996
rect 6110 46030 6210 46046
rect 6110 45996 6126 46030
rect 6194 45996 6210 46030
rect 6110 45958 6210 45996
rect 1528 39920 1628 39958
rect 1528 39886 1544 39920
rect 1612 39886 1628 39920
rect 1528 39870 1628 39886
rect 1686 39920 1786 39958
rect 1686 39886 1702 39920
rect 1770 39886 1786 39920
rect 1686 39870 1786 39886
rect 1844 39920 1944 39958
rect 1844 39886 1860 39920
rect 1928 39886 1944 39920
rect 1844 39870 1944 39886
rect 2002 39920 2102 39958
rect 2002 39886 2018 39920
rect 2086 39886 2102 39920
rect 2002 39870 2102 39886
rect 2160 39920 2260 39958
rect 2160 39886 2176 39920
rect 2244 39886 2260 39920
rect 2160 39870 2260 39886
rect 2318 39920 2418 39958
rect 2318 39886 2334 39920
rect 2402 39886 2418 39920
rect 2318 39870 2418 39886
rect 2476 39920 2576 39958
rect 2476 39886 2492 39920
rect 2560 39886 2576 39920
rect 2476 39870 2576 39886
rect 2634 39920 2734 39958
rect 2634 39886 2650 39920
rect 2718 39886 2734 39920
rect 2634 39870 2734 39886
rect 2792 39920 2892 39958
rect 2792 39886 2808 39920
rect 2876 39886 2892 39920
rect 2792 39870 2892 39886
rect 2950 39920 3050 39958
rect 2950 39886 2966 39920
rect 3034 39886 3050 39920
rect 2950 39870 3050 39886
rect 3108 39920 3208 39958
rect 3108 39886 3124 39920
rect 3192 39886 3208 39920
rect 3108 39870 3208 39886
rect 3266 39920 3366 39958
rect 3266 39886 3282 39920
rect 3350 39886 3366 39920
rect 3266 39870 3366 39886
rect 3424 39920 3524 39958
rect 3424 39886 3440 39920
rect 3508 39886 3524 39920
rect 3424 39870 3524 39886
rect 3582 39920 3682 39958
rect 3582 39886 3598 39920
rect 3666 39886 3682 39920
rect 3582 39870 3682 39886
rect 3740 39920 3840 39958
rect 3740 39886 3756 39920
rect 3824 39886 3840 39920
rect 3740 39870 3840 39886
rect 3898 39920 3998 39958
rect 3898 39886 3914 39920
rect 3982 39886 3998 39920
rect 3898 39870 3998 39886
rect 4056 39920 4156 39958
rect 4056 39886 4072 39920
rect 4140 39886 4156 39920
rect 4056 39870 4156 39886
rect 4214 39920 4314 39958
rect 4214 39886 4230 39920
rect 4298 39886 4314 39920
rect 4214 39870 4314 39886
rect 4372 39920 4472 39958
rect 4372 39886 4388 39920
rect 4456 39886 4472 39920
rect 4372 39870 4472 39886
rect 4530 39920 4630 39958
rect 4530 39886 4546 39920
rect 4614 39886 4630 39920
rect 4530 39870 4630 39886
rect 4688 39920 4788 39958
rect 4688 39886 4704 39920
rect 4772 39886 4788 39920
rect 4688 39870 4788 39886
rect 4846 39920 4946 39958
rect 4846 39886 4862 39920
rect 4930 39886 4946 39920
rect 4846 39870 4946 39886
rect 5004 39920 5104 39958
rect 5004 39886 5020 39920
rect 5088 39886 5104 39920
rect 5004 39870 5104 39886
rect 5162 39920 5262 39958
rect 5162 39886 5178 39920
rect 5246 39886 5262 39920
rect 5162 39870 5262 39886
rect 5320 39920 5420 39958
rect 5320 39886 5336 39920
rect 5404 39886 5420 39920
rect 5320 39870 5420 39886
rect 5478 39920 5578 39958
rect 5478 39886 5494 39920
rect 5562 39886 5578 39920
rect 5478 39870 5578 39886
rect 5636 39920 5736 39958
rect 5636 39886 5652 39920
rect 5720 39886 5736 39920
rect 5636 39870 5736 39886
rect 5794 39920 5894 39958
rect 5794 39886 5810 39920
rect 5878 39886 5894 39920
rect 5794 39870 5894 39886
rect 5952 39920 6052 39958
rect 5952 39886 5968 39920
rect 6036 39886 6052 39920
rect 5952 39870 6052 39886
rect 6110 39920 6210 39958
rect 6110 39886 6126 39920
rect 6194 39886 6210 39920
rect 6110 39870 6210 39886
rect 7828 46030 7928 46046
rect 7828 45996 7844 46030
rect 7912 45996 7928 46030
rect 7828 45958 7928 45996
rect 7986 46030 8086 46046
rect 7986 45996 8002 46030
rect 8070 45996 8086 46030
rect 7986 45958 8086 45996
rect 8144 46030 8244 46046
rect 8144 45996 8160 46030
rect 8228 45996 8244 46030
rect 8144 45958 8244 45996
rect 8302 46030 8402 46046
rect 8302 45996 8318 46030
rect 8386 45996 8402 46030
rect 8302 45958 8402 45996
rect 8460 46030 8560 46046
rect 8460 45996 8476 46030
rect 8544 45996 8560 46030
rect 8460 45958 8560 45996
rect 8618 46030 8718 46046
rect 8618 45996 8634 46030
rect 8702 45996 8718 46030
rect 8618 45958 8718 45996
rect 8776 46030 8876 46046
rect 8776 45996 8792 46030
rect 8860 45996 8876 46030
rect 8776 45958 8876 45996
rect 8934 46030 9034 46046
rect 8934 45996 8950 46030
rect 9018 45996 9034 46030
rect 8934 45958 9034 45996
rect 9092 46030 9192 46046
rect 9092 45996 9108 46030
rect 9176 45996 9192 46030
rect 9092 45958 9192 45996
rect 9250 46030 9350 46046
rect 9250 45996 9266 46030
rect 9334 45996 9350 46030
rect 9250 45958 9350 45996
rect 9408 46030 9508 46046
rect 9408 45996 9424 46030
rect 9492 45996 9508 46030
rect 9408 45958 9508 45996
rect 9566 46030 9666 46046
rect 9566 45996 9582 46030
rect 9650 45996 9666 46030
rect 9566 45958 9666 45996
rect 9724 46030 9824 46046
rect 9724 45996 9740 46030
rect 9808 45996 9824 46030
rect 9724 45958 9824 45996
rect 9882 46030 9982 46046
rect 9882 45996 9898 46030
rect 9966 45996 9982 46030
rect 9882 45958 9982 45996
rect 10040 46030 10140 46046
rect 10040 45996 10056 46030
rect 10124 45996 10140 46030
rect 10040 45958 10140 45996
rect 10198 46030 10298 46046
rect 10198 45996 10214 46030
rect 10282 45996 10298 46030
rect 10198 45958 10298 45996
rect 10356 46030 10456 46046
rect 10356 45996 10372 46030
rect 10440 45996 10456 46030
rect 10356 45958 10456 45996
rect 10514 46030 10614 46046
rect 10514 45996 10530 46030
rect 10598 45996 10614 46030
rect 10514 45958 10614 45996
rect 10672 46030 10772 46046
rect 10672 45996 10688 46030
rect 10756 45996 10772 46030
rect 10672 45958 10772 45996
rect 10830 46030 10930 46046
rect 10830 45996 10846 46030
rect 10914 45996 10930 46030
rect 10830 45958 10930 45996
rect 10988 46030 11088 46046
rect 10988 45996 11004 46030
rect 11072 45996 11088 46030
rect 10988 45958 11088 45996
rect 11146 46030 11246 46046
rect 11146 45996 11162 46030
rect 11230 45996 11246 46030
rect 11146 45958 11246 45996
rect 11304 46030 11404 46046
rect 11304 45996 11320 46030
rect 11388 45996 11404 46030
rect 11304 45958 11404 45996
rect 11462 46030 11562 46046
rect 11462 45996 11478 46030
rect 11546 45996 11562 46030
rect 11462 45958 11562 45996
rect 11620 46030 11720 46046
rect 11620 45996 11636 46030
rect 11704 45996 11720 46030
rect 11620 45958 11720 45996
rect 11778 46030 11878 46046
rect 11778 45996 11794 46030
rect 11862 45996 11878 46030
rect 11778 45958 11878 45996
rect 11936 46030 12036 46046
rect 11936 45996 11952 46030
rect 12020 45996 12036 46030
rect 11936 45958 12036 45996
rect 12094 46030 12194 46046
rect 12094 45996 12110 46030
rect 12178 45996 12194 46030
rect 12094 45958 12194 45996
rect 12252 46030 12352 46046
rect 12252 45996 12268 46030
rect 12336 45996 12352 46030
rect 12252 45958 12352 45996
rect 12410 46030 12510 46046
rect 12410 45996 12426 46030
rect 12494 45996 12510 46030
rect 12410 45958 12510 45996
rect 7828 39920 7928 39958
rect 7828 39886 7844 39920
rect 7912 39886 7928 39920
rect 7828 39870 7928 39886
rect 7986 39920 8086 39958
rect 7986 39886 8002 39920
rect 8070 39886 8086 39920
rect 7986 39870 8086 39886
rect 8144 39920 8244 39958
rect 8144 39886 8160 39920
rect 8228 39886 8244 39920
rect 8144 39870 8244 39886
rect 8302 39920 8402 39958
rect 8302 39886 8318 39920
rect 8386 39886 8402 39920
rect 8302 39870 8402 39886
rect 8460 39920 8560 39958
rect 8460 39886 8476 39920
rect 8544 39886 8560 39920
rect 8460 39870 8560 39886
rect 8618 39920 8718 39958
rect 8618 39886 8634 39920
rect 8702 39886 8718 39920
rect 8618 39870 8718 39886
rect 8776 39920 8876 39958
rect 8776 39886 8792 39920
rect 8860 39886 8876 39920
rect 8776 39870 8876 39886
rect 8934 39920 9034 39958
rect 8934 39886 8950 39920
rect 9018 39886 9034 39920
rect 8934 39870 9034 39886
rect 9092 39920 9192 39958
rect 9092 39886 9108 39920
rect 9176 39886 9192 39920
rect 9092 39870 9192 39886
rect 9250 39920 9350 39958
rect 9250 39886 9266 39920
rect 9334 39886 9350 39920
rect 9250 39870 9350 39886
rect 9408 39920 9508 39958
rect 9408 39886 9424 39920
rect 9492 39886 9508 39920
rect 9408 39870 9508 39886
rect 9566 39920 9666 39958
rect 9566 39886 9582 39920
rect 9650 39886 9666 39920
rect 9566 39870 9666 39886
rect 9724 39920 9824 39958
rect 9724 39886 9740 39920
rect 9808 39886 9824 39920
rect 9724 39870 9824 39886
rect 9882 39920 9982 39958
rect 9882 39886 9898 39920
rect 9966 39886 9982 39920
rect 9882 39870 9982 39886
rect 10040 39920 10140 39958
rect 10040 39886 10056 39920
rect 10124 39886 10140 39920
rect 10040 39870 10140 39886
rect 10198 39920 10298 39958
rect 10198 39886 10214 39920
rect 10282 39886 10298 39920
rect 10198 39870 10298 39886
rect 10356 39920 10456 39958
rect 10356 39886 10372 39920
rect 10440 39886 10456 39920
rect 10356 39870 10456 39886
rect 10514 39920 10614 39958
rect 10514 39886 10530 39920
rect 10598 39886 10614 39920
rect 10514 39870 10614 39886
rect 10672 39920 10772 39958
rect 10672 39886 10688 39920
rect 10756 39886 10772 39920
rect 10672 39870 10772 39886
rect 10830 39920 10930 39958
rect 10830 39886 10846 39920
rect 10914 39886 10930 39920
rect 10830 39870 10930 39886
rect 10988 39920 11088 39958
rect 10988 39886 11004 39920
rect 11072 39886 11088 39920
rect 10988 39870 11088 39886
rect 11146 39920 11246 39958
rect 11146 39886 11162 39920
rect 11230 39886 11246 39920
rect 11146 39870 11246 39886
rect 11304 39920 11404 39958
rect 11304 39886 11320 39920
rect 11388 39886 11404 39920
rect 11304 39870 11404 39886
rect 11462 39920 11562 39958
rect 11462 39886 11478 39920
rect 11546 39886 11562 39920
rect 11462 39870 11562 39886
rect 11620 39920 11720 39958
rect 11620 39886 11636 39920
rect 11704 39886 11720 39920
rect 11620 39870 11720 39886
rect 11778 39920 11878 39958
rect 11778 39886 11794 39920
rect 11862 39886 11878 39920
rect 11778 39870 11878 39886
rect 11936 39920 12036 39958
rect 11936 39886 11952 39920
rect 12020 39886 12036 39920
rect 11936 39870 12036 39886
rect 12094 39920 12194 39958
rect 12094 39886 12110 39920
rect 12178 39886 12194 39920
rect 12094 39870 12194 39886
rect 12252 39920 12352 39958
rect 12252 39886 12268 39920
rect 12336 39886 12352 39920
rect 12252 39870 12352 39886
rect 12410 39920 12510 39958
rect 12410 39886 12426 39920
rect 12494 39886 12510 39920
rect 12410 39870 12510 39886
rect 14128 46030 14228 46046
rect 14128 45996 14144 46030
rect 14212 45996 14228 46030
rect 14128 45958 14228 45996
rect 14286 46030 14386 46046
rect 14286 45996 14302 46030
rect 14370 45996 14386 46030
rect 14286 45958 14386 45996
rect 14444 46030 14544 46046
rect 14444 45996 14460 46030
rect 14528 45996 14544 46030
rect 14444 45958 14544 45996
rect 14602 46030 14702 46046
rect 14602 45996 14618 46030
rect 14686 45996 14702 46030
rect 14602 45958 14702 45996
rect 14760 46030 14860 46046
rect 14760 45996 14776 46030
rect 14844 45996 14860 46030
rect 14760 45958 14860 45996
rect 14918 46030 15018 46046
rect 14918 45996 14934 46030
rect 15002 45996 15018 46030
rect 14918 45958 15018 45996
rect 15076 46030 15176 46046
rect 15076 45996 15092 46030
rect 15160 45996 15176 46030
rect 15076 45958 15176 45996
rect 15234 46030 15334 46046
rect 15234 45996 15250 46030
rect 15318 45996 15334 46030
rect 15234 45958 15334 45996
rect 15392 46030 15492 46046
rect 15392 45996 15408 46030
rect 15476 45996 15492 46030
rect 15392 45958 15492 45996
rect 15550 46030 15650 46046
rect 15550 45996 15566 46030
rect 15634 45996 15650 46030
rect 15550 45958 15650 45996
rect 15708 46030 15808 46046
rect 15708 45996 15724 46030
rect 15792 45996 15808 46030
rect 15708 45958 15808 45996
rect 15866 46030 15966 46046
rect 15866 45996 15882 46030
rect 15950 45996 15966 46030
rect 15866 45958 15966 45996
rect 16024 46030 16124 46046
rect 16024 45996 16040 46030
rect 16108 45996 16124 46030
rect 16024 45958 16124 45996
rect 16182 46030 16282 46046
rect 16182 45996 16198 46030
rect 16266 45996 16282 46030
rect 16182 45958 16282 45996
rect 16340 46030 16440 46046
rect 16340 45996 16356 46030
rect 16424 45996 16440 46030
rect 16340 45958 16440 45996
rect 16498 46030 16598 46046
rect 16498 45996 16514 46030
rect 16582 45996 16598 46030
rect 16498 45958 16598 45996
rect 16656 46030 16756 46046
rect 16656 45996 16672 46030
rect 16740 45996 16756 46030
rect 16656 45958 16756 45996
rect 16814 46030 16914 46046
rect 16814 45996 16830 46030
rect 16898 45996 16914 46030
rect 16814 45958 16914 45996
rect 16972 46030 17072 46046
rect 16972 45996 16988 46030
rect 17056 45996 17072 46030
rect 16972 45958 17072 45996
rect 17130 46030 17230 46046
rect 17130 45996 17146 46030
rect 17214 45996 17230 46030
rect 17130 45958 17230 45996
rect 17288 46030 17388 46046
rect 17288 45996 17304 46030
rect 17372 45996 17388 46030
rect 17288 45958 17388 45996
rect 17446 46030 17546 46046
rect 17446 45996 17462 46030
rect 17530 45996 17546 46030
rect 17446 45958 17546 45996
rect 17604 46030 17704 46046
rect 17604 45996 17620 46030
rect 17688 45996 17704 46030
rect 17604 45958 17704 45996
rect 17762 46030 17862 46046
rect 17762 45996 17778 46030
rect 17846 45996 17862 46030
rect 17762 45958 17862 45996
rect 17920 46030 18020 46046
rect 17920 45996 17936 46030
rect 18004 45996 18020 46030
rect 17920 45958 18020 45996
rect 18078 46030 18178 46046
rect 18078 45996 18094 46030
rect 18162 45996 18178 46030
rect 18078 45958 18178 45996
rect 18236 46030 18336 46046
rect 18236 45996 18252 46030
rect 18320 45996 18336 46030
rect 18236 45958 18336 45996
rect 18394 46030 18494 46046
rect 18394 45996 18410 46030
rect 18478 45996 18494 46030
rect 18394 45958 18494 45996
rect 18552 46030 18652 46046
rect 18552 45996 18568 46030
rect 18636 45996 18652 46030
rect 18552 45958 18652 45996
rect 18710 46030 18810 46046
rect 18710 45996 18726 46030
rect 18794 45996 18810 46030
rect 18710 45958 18810 45996
rect 14128 39920 14228 39958
rect 14128 39886 14144 39920
rect 14212 39886 14228 39920
rect 14128 39870 14228 39886
rect 14286 39920 14386 39958
rect 14286 39886 14302 39920
rect 14370 39886 14386 39920
rect 14286 39870 14386 39886
rect 14444 39920 14544 39958
rect 14444 39886 14460 39920
rect 14528 39886 14544 39920
rect 14444 39870 14544 39886
rect 14602 39920 14702 39958
rect 14602 39886 14618 39920
rect 14686 39886 14702 39920
rect 14602 39870 14702 39886
rect 14760 39920 14860 39958
rect 14760 39886 14776 39920
rect 14844 39886 14860 39920
rect 14760 39870 14860 39886
rect 14918 39920 15018 39958
rect 14918 39886 14934 39920
rect 15002 39886 15018 39920
rect 14918 39870 15018 39886
rect 15076 39920 15176 39958
rect 15076 39886 15092 39920
rect 15160 39886 15176 39920
rect 15076 39870 15176 39886
rect 15234 39920 15334 39958
rect 15234 39886 15250 39920
rect 15318 39886 15334 39920
rect 15234 39870 15334 39886
rect 15392 39920 15492 39958
rect 15392 39886 15408 39920
rect 15476 39886 15492 39920
rect 15392 39870 15492 39886
rect 15550 39920 15650 39958
rect 15550 39886 15566 39920
rect 15634 39886 15650 39920
rect 15550 39870 15650 39886
rect 15708 39920 15808 39958
rect 15708 39886 15724 39920
rect 15792 39886 15808 39920
rect 15708 39870 15808 39886
rect 15866 39920 15966 39958
rect 15866 39886 15882 39920
rect 15950 39886 15966 39920
rect 15866 39870 15966 39886
rect 16024 39920 16124 39958
rect 16024 39886 16040 39920
rect 16108 39886 16124 39920
rect 16024 39870 16124 39886
rect 16182 39920 16282 39958
rect 16182 39886 16198 39920
rect 16266 39886 16282 39920
rect 16182 39870 16282 39886
rect 16340 39920 16440 39958
rect 16340 39886 16356 39920
rect 16424 39886 16440 39920
rect 16340 39870 16440 39886
rect 16498 39920 16598 39958
rect 16498 39886 16514 39920
rect 16582 39886 16598 39920
rect 16498 39870 16598 39886
rect 16656 39920 16756 39958
rect 16656 39886 16672 39920
rect 16740 39886 16756 39920
rect 16656 39870 16756 39886
rect 16814 39920 16914 39958
rect 16814 39886 16830 39920
rect 16898 39886 16914 39920
rect 16814 39870 16914 39886
rect 16972 39920 17072 39958
rect 16972 39886 16988 39920
rect 17056 39886 17072 39920
rect 16972 39870 17072 39886
rect 17130 39920 17230 39958
rect 17130 39886 17146 39920
rect 17214 39886 17230 39920
rect 17130 39870 17230 39886
rect 17288 39920 17388 39958
rect 17288 39886 17304 39920
rect 17372 39886 17388 39920
rect 17288 39870 17388 39886
rect 17446 39920 17546 39958
rect 17446 39886 17462 39920
rect 17530 39886 17546 39920
rect 17446 39870 17546 39886
rect 17604 39920 17704 39958
rect 17604 39886 17620 39920
rect 17688 39886 17704 39920
rect 17604 39870 17704 39886
rect 17762 39920 17862 39958
rect 17762 39886 17778 39920
rect 17846 39886 17862 39920
rect 17762 39870 17862 39886
rect 17920 39920 18020 39958
rect 17920 39886 17936 39920
rect 18004 39886 18020 39920
rect 17920 39870 18020 39886
rect 18078 39920 18178 39958
rect 18078 39886 18094 39920
rect 18162 39886 18178 39920
rect 18078 39870 18178 39886
rect 18236 39920 18336 39958
rect 18236 39886 18252 39920
rect 18320 39886 18336 39920
rect 18236 39870 18336 39886
rect 18394 39920 18494 39958
rect 18394 39886 18410 39920
rect 18478 39886 18494 39920
rect 18394 39870 18494 39886
rect 18552 39920 18652 39958
rect 18552 39886 18568 39920
rect 18636 39886 18652 39920
rect 18552 39870 18652 39886
rect 18710 39920 18810 39958
rect 18710 39886 18726 39920
rect 18794 39886 18810 39920
rect 18710 39870 18810 39886
rect 20428 46030 20528 46046
rect 20428 45996 20444 46030
rect 20512 45996 20528 46030
rect 20428 45958 20528 45996
rect 20586 46030 20686 46046
rect 20586 45996 20602 46030
rect 20670 45996 20686 46030
rect 20586 45958 20686 45996
rect 20744 46030 20844 46046
rect 20744 45996 20760 46030
rect 20828 45996 20844 46030
rect 20744 45958 20844 45996
rect 20902 46030 21002 46046
rect 20902 45996 20918 46030
rect 20986 45996 21002 46030
rect 20902 45958 21002 45996
rect 21060 46030 21160 46046
rect 21060 45996 21076 46030
rect 21144 45996 21160 46030
rect 21060 45958 21160 45996
rect 21218 46030 21318 46046
rect 21218 45996 21234 46030
rect 21302 45996 21318 46030
rect 21218 45958 21318 45996
rect 21376 46030 21476 46046
rect 21376 45996 21392 46030
rect 21460 45996 21476 46030
rect 21376 45958 21476 45996
rect 21534 46030 21634 46046
rect 21534 45996 21550 46030
rect 21618 45996 21634 46030
rect 21534 45958 21634 45996
rect 21692 46030 21792 46046
rect 21692 45996 21708 46030
rect 21776 45996 21792 46030
rect 21692 45958 21792 45996
rect 21850 46030 21950 46046
rect 21850 45996 21866 46030
rect 21934 45996 21950 46030
rect 21850 45958 21950 45996
rect 22008 46030 22108 46046
rect 22008 45996 22024 46030
rect 22092 45996 22108 46030
rect 22008 45958 22108 45996
rect 22166 46030 22266 46046
rect 22166 45996 22182 46030
rect 22250 45996 22266 46030
rect 22166 45958 22266 45996
rect 22324 46030 22424 46046
rect 22324 45996 22340 46030
rect 22408 45996 22424 46030
rect 22324 45958 22424 45996
rect 22482 46030 22582 46046
rect 22482 45996 22498 46030
rect 22566 45996 22582 46030
rect 22482 45958 22582 45996
rect 22640 46030 22740 46046
rect 22640 45996 22656 46030
rect 22724 45996 22740 46030
rect 22640 45958 22740 45996
rect 22798 46030 22898 46046
rect 22798 45996 22814 46030
rect 22882 45996 22898 46030
rect 22798 45958 22898 45996
rect 22956 46030 23056 46046
rect 22956 45996 22972 46030
rect 23040 45996 23056 46030
rect 22956 45958 23056 45996
rect 23114 46030 23214 46046
rect 23114 45996 23130 46030
rect 23198 45996 23214 46030
rect 23114 45958 23214 45996
rect 23272 46030 23372 46046
rect 23272 45996 23288 46030
rect 23356 45996 23372 46030
rect 23272 45958 23372 45996
rect 23430 46030 23530 46046
rect 23430 45996 23446 46030
rect 23514 45996 23530 46030
rect 23430 45958 23530 45996
rect 23588 46030 23688 46046
rect 23588 45996 23604 46030
rect 23672 45996 23688 46030
rect 23588 45958 23688 45996
rect 23746 46030 23846 46046
rect 23746 45996 23762 46030
rect 23830 45996 23846 46030
rect 23746 45958 23846 45996
rect 23904 46030 24004 46046
rect 23904 45996 23920 46030
rect 23988 45996 24004 46030
rect 23904 45958 24004 45996
rect 24062 46030 24162 46046
rect 24062 45996 24078 46030
rect 24146 45996 24162 46030
rect 24062 45958 24162 45996
rect 24220 46030 24320 46046
rect 24220 45996 24236 46030
rect 24304 45996 24320 46030
rect 24220 45958 24320 45996
rect 24378 46030 24478 46046
rect 24378 45996 24394 46030
rect 24462 45996 24478 46030
rect 24378 45958 24478 45996
rect 24536 46030 24636 46046
rect 24536 45996 24552 46030
rect 24620 45996 24636 46030
rect 24536 45958 24636 45996
rect 24694 46030 24794 46046
rect 24694 45996 24710 46030
rect 24778 45996 24794 46030
rect 24694 45958 24794 45996
rect 24852 46030 24952 46046
rect 24852 45996 24868 46030
rect 24936 45996 24952 46030
rect 24852 45958 24952 45996
rect 25010 46030 25110 46046
rect 25010 45996 25026 46030
rect 25094 45996 25110 46030
rect 25010 45958 25110 45996
rect 20428 39920 20528 39958
rect 20428 39886 20444 39920
rect 20512 39886 20528 39920
rect 20428 39870 20528 39886
rect 20586 39920 20686 39958
rect 20586 39886 20602 39920
rect 20670 39886 20686 39920
rect 20586 39870 20686 39886
rect 20744 39920 20844 39958
rect 20744 39886 20760 39920
rect 20828 39886 20844 39920
rect 20744 39870 20844 39886
rect 20902 39920 21002 39958
rect 20902 39886 20918 39920
rect 20986 39886 21002 39920
rect 20902 39870 21002 39886
rect 21060 39920 21160 39958
rect 21060 39886 21076 39920
rect 21144 39886 21160 39920
rect 21060 39870 21160 39886
rect 21218 39920 21318 39958
rect 21218 39886 21234 39920
rect 21302 39886 21318 39920
rect 21218 39870 21318 39886
rect 21376 39920 21476 39958
rect 21376 39886 21392 39920
rect 21460 39886 21476 39920
rect 21376 39870 21476 39886
rect 21534 39920 21634 39958
rect 21534 39886 21550 39920
rect 21618 39886 21634 39920
rect 21534 39870 21634 39886
rect 21692 39920 21792 39958
rect 21692 39886 21708 39920
rect 21776 39886 21792 39920
rect 21692 39870 21792 39886
rect 21850 39920 21950 39958
rect 21850 39886 21866 39920
rect 21934 39886 21950 39920
rect 21850 39870 21950 39886
rect 22008 39920 22108 39958
rect 22008 39886 22024 39920
rect 22092 39886 22108 39920
rect 22008 39870 22108 39886
rect 22166 39920 22266 39958
rect 22166 39886 22182 39920
rect 22250 39886 22266 39920
rect 22166 39870 22266 39886
rect 22324 39920 22424 39958
rect 22324 39886 22340 39920
rect 22408 39886 22424 39920
rect 22324 39870 22424 39886
rect 22482 39920 22582 39958
rect 22482 39886 22498 39920
rect 22566 39886 22582 39920
rect 22482 39870 22582 39886
rect 22640 39920 22740 39958
rect 22640 39886 22656 39920
rect 22724 39886 22740 39920
rect 22640 39870 22740 39886
rect 22798 39920 22898 39958
rect 22798 39886 22814 39920
rect 22882 39886 22898 39920
rect 22798 39870 22898 39886
rect 22956 39920 23056 39958
rect 22956 39886 22972 39920
rect 23040 39886 23056 39920
rect 22956 39870 23056 39886
rect 23114 39920 23214 39958
rect 23114 39886 23130 39920
rect 23198 39886 23214 39920
rect 23114 39870 23214 39886
rect 23272 39920 23372 39958
rect 23272 39886 23288 39920
rect 23356 39886 23372 39920
rect 23272 39870 23372 39886
rect 23430 39920 23530 39958
rect 23430 39886 23446 39920
rect 23514 39886 23530 39920
rect 23430 39870 23530 39886
rect 23588 39920 23688 39958
rect 23588 39886 23604 39920
rect 23672 39886 23688 39920
rect 23588 39870 23688 39886
rect 23746 39920 23846 39958
rect 23746 39886 23762 39920
rect 23830 39886 23846 39920
rect 23746 39870 23846 39886
rect 23904 39920 24004 39958
rect 23904 39886 23920 39920
rect 23988 39886 24004 39920
rect 23904 39870 24004 39886
rect 24062 39920 24162 39958
rect 24062 39886 24078 39920
rect 24146 39886 24162 39920
rect 24062 39870 24162 39886
rect 24220 39920 24320 39958
rect 24220 39886 24236 39920
rect 24304 39886 24320 39920
rect 24220 39870 24320 39886
rect 24378 39920 24478 39958
rect 24378 39886 24394 39920
rect 24462 39886 24478 39920
rect 24378 39870 24478 39886
rect 24536 39920 24636 39958
rect 24536 39886 24552 39920
rect 24620 39886 24636 39920
rect 24536 39870 24636 39886
rect 24694 39920 24794 39958
rect 24694 39886 24710 39920
rect 24778 39886 24794 39920
rect 24694 39870 24794 39886
rect 24852 39920 24952 39958
rect 24852 39886 24868 39920
rect 24936 39886 24952 39920
rect 24852 39870 24952 39886
rect 25010 39920 25110 39958
rect 25010 39886 25026 39920
rect 25094 39886 25110 39920
rect 25010 39870 25110 39886
rect 1528 39030 1628 39046
rect 1528 38996 1544 39030
rect 1612 38996 1628 39030
rect 1528 38958 1628 38996
rect 1686 39030 1786 39046
rect 1686 38996 1702 39030
rect 1770 38996 1786 39030
rect 1686 38958 1786 38996
rect 1844 39030 1944 39046
rect 1844 38996 1860 39030
rect 1928 38996 1944 39030
rect 1844 38958 1944 38996
rect 2002 39030 2102 39046
rect 2002 38996 2018 39030
rect 2086 38996 2102 39030
rect 2002 38958 2102 38996
rect 2160 39030 2260 39046
rect 2160 38996 2176 39030
rect 2244 38996 2260 39030
rect 2160 38958 2260 38996
rect 2318 39030 2418 39046
rect 2318 38996 2334 39030
rect 2402 38996 2418 39030
rect 2318 38958 2418 38996
rect 2476 39030 2576 39046
rect 2476 38996 2492 39030
rect 2560 38996 2576 39030
rect 2476 38958 2576 38996
rect 2634 39030 2734 39046
rect 2634 38996 2650 39030
rect 2718 38996 2734 39030
rect 2634 38958 2734 38996
rect 2792 39030 2892 39046
rect 2792 38996 2808 39030
rect 2876 38996 2892 39030
rect 2792 38958 2892 38996
rect 2950 39030 3050 39046
rect 2950 38996 2966 39030
rect 3034 38996 3050 39030
rect 2950 38958 3050 38996
rect 3108 39030 3208 39046
rect 3108 38996 3124 39030
rect 3192 38996 3208 39030
rect 3108 38958 3208 38996
rect 3266 39030 3366 39046
rect 3266 38996 3282 39030
rect 3350 38996 3366 39030
rect 3266 38958 3366 38996
rect 3424 39030 3524 39046
rect 3424 38996 3440 39030
rect 3508 38996 3524 39030
rect 3424 38958 3524 38996
rect 3582 39030 3682 39046
rect 3582 38996 3598 39030
rect 3666 38996 3682 39030
rect 3582 38958 3682 38996
rect 3740 39030 3840 39046
rect 3740 38996 3756 39030
rect 3824 38996 3840 39030
rect 3740 38958 3840 38996
rect 3898 39030 3998 39046
rect 3898 38996 3914 39030
rect 3982 38996 3998 39030
rect 3898 38958 3998 38996
rect 4056 39030 4156 39046
rect 4056 38996 4072 39030
rect 4140 38996 4156 39030
rect 4056 38958 4156 38996
rect 4214 39030 4314 39046
rect 4214 38996 4230 39030
rect 4298 38996 4314 39030
rect 4214 38958 4314 38996
rect 4372 39030 4472 39046
rect 4372 38996 4388 39030
rect 4456 38996 4472 39030
rect 4372 38958 4472 38996
rect 4530 39030 4630 39046
rect 4530 38996 4546 39030
rect 4614 38996 4630 39030
rect 4530 38958 4630 38996
rect 4688 39030 4788 39046
rect 4688 38996 4704 39030
rect 4772 38996 4788 39030
rect 4688 38958 4788 38996
rect 4846 39030 4946 39046
rect 4846 38996 4862 39030
rect 4930 38996 4946 39030
rect 4846 38958 4946 38996
rect 5004 39030 5104 39046
rect 5004 38996 5020 39030
rect 5088 38996 5104 39030
rect 5004 38958 5104 38996
rect 5162 39030 5262 39046
rect 5162 38996 5178 39030
rect 5246 38996 5262 39030
rect 5162 38958 5262 38996
rect 5320 39030 5420 39046
rect 5320 38996 5336 39030
rect 5404 38996 5420 39030
rect 5320 38958 5420 38996
rect 5478 39030 5578 39046
rect 5478 38996 5494 39030
rect 5562 38996 5578 39030
rect 5478 38958 5578 38996
rect 5636 39030 5736 39046
rect 5636 38996 5652 39030
rect 5720 38996 5736 39030
rect 5636 38958 5736 38996
rect 5794 39030 5894 39046
rect 5794 38996 5810 39030
rect 5878 38996 5894 39030
rect 5794 38958 5894 38996
rect 5952 39030 6052 39046
rect 5952 38996 5968 39030
rect 6036 38996 6052 39030
rect 5952 38958 6052 38996
rect 6110 39030 6210 39046
rect 6110 38996 6126 39030
rect 6194 38996 6210 39030
rect 6110 38958 6210 38996
rect 1528 32920 1628 32958
rect 1528 32886 1544 32920
rect 1612 32886 1628 32920
rect 1528 32870 1628 32886
rect 1686 32920 1786 32958
rect 1686 32886 1702 32920
rect 1770 32886 1786 32920
rect 1686 32870 1786 32886
rect 1844 32920 1944 32958
rect 1844 32886 1860 32920
rect 1928 32886 1944 32920
rect 1844 32870 1944 32886
rect 2002 32920 2102 32958
rect 2002 32886 2018 32920
rect 2086 32886 2102 32920
rect 2002 32870 2102 32886
rect 2160 32920 2260 32958
rect 2160 32886 2176 32920
rect 2244 32886 2260 32920
rect 2160 32870 2260 32886
rect 2318 32920 2418 32958
rect 2318 32886 2334 32920
rect 2402 32886 2418 32920
rect 2318 32870 2418 32886
rect 2476 32920 2576 32958
rect 2476 32886 2492 32920
rect 2560 32886 2576 32920
rect 2476 32870 2576 32886
rect 2634 32920 2734 32958
rect 2634 32886 2650 32920
rect 2718 32886 2734 32920
rect 2634 32870 2734 32886
rect 2792 32920 2892 32958
rect 2792 32886 2808 32920
rect 2876 32886 2892 32920
rect 2792 32870 2892 32886
rect 2950 32920 3050 32958
rect 2950 32886 2966 32920
rect 3034 32886 3050 32920
rect 2950 32870 3050 32886
rect 3108 32920 3208 32958
rect 3108 32886 3124 32920
rect 3192 32886 3208 32920
rect 3108 32870 3208 32886
rect 3266 32920 3366 32958
rect 3266 32886 3282 32920
rect 3350 32886 3366 32920
rect 3266 32870 3366 32886
rect 3424 32920 3524 32958
rect 3424 32886 3440 32920
rect 3508 32886 3524 32920
rect 3424 32870 3524 32886
rect 3582 32920 3682 32958
rect 3582 32886 3598 32920
rect 3666 32886 3682 32920
rect 3582 32870 3682 32886
rect 3740 32920 3840 32958
rect 3740 32886 3756 32920
rect 3824 32886 3840 32920
rect 3740 32870 3840 32886
rect 3898 32920 3998 32958
rect 3898 32886 3914 32920
rect 3982 32886 3998 32920
rect 3898 32870 3998 32886
rect 4056 32920 4156 32958
rect 4056 32886 4072 32920
rect 4140 32886 4156 32920
rect 4056 32870 4156 32886
rect 4214 32920 4314 32958
rect 4214 32886 4230 32920
rect 4298 32886 4314 32920
rect 4214 32870 4314 32886
rect 4372 32920 4472 32958
rect 4372 32886 4388 32920
rect 4456 32886 4472 32920
rect 4372 32870 4472 32886
rect 4530 32920 4630 32958
rect 4530 32886 4546 32920
rect 4614 32886 4630 32920
rect 4530 32870 4630 32886
rect 4688 32920 4788 32958
rect 4688 32886 4704 32920
rect 4772 32886 4788 32920
rect 4688 32870 4788 32886
rect 4846 32920 4946 32958
rect 4846 32886 4862 32920
rect 4930 32886 4946 32920
rect 4846 32870 4946 32886
rect 5004 32920 5104 32958
rect 5004 32886 5020 32920
rect 5088 32886 5104 32920
rect 5004 32870 5104 32886
rect 5162 32920 5262 32958
rect 5162 32886 5178 32920
rect 5246 32886 5262 32920
rect 5162 32870 5262 32886
rect 5320 32920 5420 32958
rect 5320 32886 5336 32920
rect 5404 32886 5420 32920
rect 5320 32870 5420 32886
rect 5478 32920 5578 32958
rect 5478 32886 5494 32920
rect 5562 32886 5578 32920
rect 5478 32870 5578 32886
rect 5636 32920 5736 32958
rect 5636 32886 5652 32920
rect 5720 32886 5736 32920
rect 5636 32870 5736 32886
rect 5794 32920 5894 32958
rect 5794 32886 5810 32920
rect 5878 32886 5894 32920
rect 5794 32870 5894 32886
rect 5952 32920 6052 32958
rect 5952 32886 5968 32920
rect 6036 32886 6052 32920
rect 5952 32870 6052 32886
rect 6110 32920 6210 32958
rect 6110 32886 6126 32920
rect 6194 32886 6210 32920
rect 6110 32870 6210 32886
rect 7828 39030 7928 39046
rect 7828 38996 7844 39030
rect 7912 38996 7928 39030
rect 7828 38958 7928 38996
rect 7986 39030 8086 39046
rect 7986 38996 8002 39030
rect 8070 38996 8086 39030
rect 7986 38958 8086 38996
rect 8144 39030 8244 39046
rect 8144 38996 8160 39030
rect 8228 38996 8244 39030
rect 8144 38958 8244 38996
rect 8302 39030 8402 39046
rect 8302 38996 8318 39030
rect 8386 38996 8402 39030
rect 8302 38958 8402 38996
rect 8460 39030 8560 39046
rect 8460 38996 8476 39030
rect 8544 38996 8560 39030
rect 8460 38958 8560 38996
rect 8618 39030 8718 39046
rect 8618 38996 8634 39030
rect 8702 38996 8718 39030
rect 8618 38958 8718 38996
rect 8776 39030 8876 39046
rect 8776 38996 8792 39030
rect 8860 38996 8876 39030
rect 8776 38958 8876 38996
rect 8934 39030 9034 39046
rect 8934 38996 8950 39030
rect 9018 38996 9034 39030
rect 8934 38958 9034 38996
rect 9092 39030 9192 39046
rect 9092 38996 9108 39030
rect 9176 38996 9192 39030
rect 9092 38958 9192 38996
rect 9250 39030 9350 39046
rect 9250 38996 9266 39030
rect 9334 38996 9350 39030
rect 9250 38958 9350 38996
rect 9408 39030 9508 39046
rect 9408 38996 9424 39030
rect 9492 38996 9508 39030
rect 9408 38958 9508 38996
rect 9566 39030 9666 39046
rect 9566 38996 9582 39030
rect 9650 38996 9666 39030
rect 9566 38958 9666 38996
rect 9724 39030 9824 39046
rect 9724 38996 9740 39030
rect 9808 38996 9824 39030
rect 9724 38958 9824 38996
rect 9882 39030 9982 39046
rect 9882 38996 9898 39030
rect 9966 38996 9982 39030
rect 9882 38958 9982 38996
rect 10040 39030 10140 39046
rect 10040 38996 10056 39030
rect 10124 38996 10140 39030
rect 10040 38958 10140 38996
rect 10198 39030 10298 39046
rect 10198 38996 10214 39030
rect 10282 38996 10298 39030
rect 10198 38958 10298 38996
rect 10356 39030 10456 39046
rect 10356 38996 10372 39030
rect 10440 38996 10456 39030
rect 10356 38958 10456 38996
rect 10514 39030 10614 39046
rect 10514 38996 10530 39030
rect 10598 38996 10614 39030
rect 10514 38958 10614 38996
rect 10672 39030 10772 39046
rect 10672 38996 10688 39030
rect 10756 38996 10772 39030
rect 10672 38958 10772 38996
rect 10830 39030 10930 39046
rect 10830 38996 10846 39030
rect 10914 38996 10930 39030
rect 10830 38958 10930 38996
rect 10988 39030 11088 39046
rect 10988 38996 11004 39030
rect 11072 38996 11088 39030
rect 10988 38958 11088 38996
rect 11146 39030 11246 39046
rect 11146 38996 11162 39030
rect 11230 38996 11246 39030
rect 11146 38958 11246 38996
rect 11304 39030 11404 39046
rect 11304 38996 11320 39030
rect 11388 38996 11404 39030
rect 11304 38958 11404 38996
rect 11462 39030 11562 39046
rect 11462 38996 11478 39030
rect 11546 38996 11562 39030
rect 11462 38958 11562 38996
rect 11620 39030 11720 39046
rect 11620 38996 11636 39030
rect 11704 38996 11720 39030
rect 11620 38958 11720 38996
rect 11778 39030 11878 39046
rect 11778 38996 11794 39030
rect 11862 38996 11878 39030
rect 11778 38958 11878 38996
rect 11936 39030 12036 39046
rect 11936 38996 11952 39030
rect 12020 38996 12036 39030
rect 11936 38958 12036 38996
rect 12094 39030 12194 39046
rect 12094 38996 12110 39030
rect 12178 38996 12194 39030
rect 12094 38958 12194 38996
rect 12252 39030 12352 39046
rect 12252 38996 12268 39030
rect 12336 38996 12352 39030
rect 12252 38958 12352 38996
rect 12410 39030 12510 39046
rect 12410 38996 12426 39030
rect 12494 38996 12510 39030
rect 12410 38958 12510 38996
rect 7828 32920 7928 32958
rect 7828 32886 7844 32920
rect 7912 32886 7928 32920
rect 7828 32870 7928 32886
rect 7986 32920 8086 32958
rect 7986 32886 8002 32920
rect 8070 32886 8086 32920
rect 7986 32870 8086 32886
rect 8144 32920 8244 32958
rect 8144 32886 8160 32920
rect 8228 32886 8244 32920
rect 8144 32870 8244 32886
rect 8302 32920 8402 32958
rect 8302 32886 8318 32920
rect 8386 32886 8402 32920
rect 8302 32870 8402 32886
rect 8460 32920 8560 32958
rect 8460 32886 8476 32920
rect 8544 32886 8560 32920
rect 8460 32870 8560 32886
rect 8618 32920 8718 32958
rect 8618 32886 8634 32920
rect 8702 32886 8718 32920
rect 8618 32870 8718 32886
rect 8776 32920 8876 32958
rect 8776 32886 8792 32920
rect 8860 32886 8876 32920
rect 8776 32870 8876 32886
rect 8934 32920 9034 32958
rect 8934 32886 8950 32920
rect 9018 32886 9034 32920
rect 8934 32870 9034 32886
rect 9092 32920 9192 32958
rect 9092 32886 9108 32920
rect 9176 32886 9192 32920
rect 9092 32870 9192 32886
rect 9250 32920 9350 32958
rect 9250 32886 9266 32920
rect 9334 32886 9350 32920
rect 9250 32870 9350 32886
rect 9408 32920 9508 32958
rect 9408 32886 9424 32920
rect 9492 32886 9508 32920
rect 9408 32870 9508 32886
rect 9566 32920 9666 32958
rect 9566 32886 9582 32920
rect 9650 32886 9666 32920
rect 9566 32870 9666 32886
rect 9724 32920 9824 32958
rect 9724 32886 9740 32920
rect 9808 32886 9824 32920
rect 9724 32870 9824 32886
rect 9882 32920 9982 32958
rect 9882 32886 9898 32920
rect 9966 32886 9982 32920
rect 9882 32870 9982 32886
rect 10040 32920 10140 32958
rect 10040 32886 10056 32920
rect 10124 32886 10140 32920
rect 10040 32870 10140 32886
rect 10198 32920 10298 32958
rect 10198 32886 10214 32920
rect 10282 32886 10298 32920
rect 10198 32870 10298 32886
rect 10356 32920 10456 32958
rect 10356 32886 10372 32920
rect 10440 32886 10456 32920
rect 10356 32870 10456 32886
rect 10514 32920 10614 32958
rect 10514 32886 10530 32920
rect 10598 32886 10614 32920
rect 10514 32870 10614 32886
rect 10672 32920 10772 32958
rect 10672 32886 10688 32920
rect 10756 32886 10772 32920
rect 10672 32870 10772 32886
rect 10830 32920 10930 32958
rect 10830 32886 10846 32920
rect 10914 32886 10930 32920
rect 10830 32870 10930 32886
rect 10988 32920 11088 32958
rect 10988 32886 11004 32920
rect 11072 32886 11088 32920
rect 10988 32870 11088 32886
rect 11146 32920 11246 32958
rect 11146 32886 11162 32920
rect 11230 32886 11246 32920
rect 11146 32870 11246 32886
rect 11304 32920 11404 32958
rect 11304 32886 11320 32920
rect 11388 32886 11404 32920
rect 11304 32870 11404 32886
rect 11462 32920 11562 32958
rect 11462 32886 11478 32920
rect 11546 32886 11562 32920
rect 11462 32870 11562 32886
rect 11620 32920 11720 32958
rect 11620 32886 11636 32920
rect 11704 32886 11720 32920
rect 11620 32870 11720 32886
rect 11778 32920 11878 32958
rect 11778 32886 11794 32920
rect 11862 32886 11878 32920
rect 11778 32870 11878 32886
rect 11936 32920 12036 32958
rect 11936 32886 11952 32920
rect 12020 32886 12036 32920
rect 11936 32870 12036 32886
rect 12094 32920 12194 32958
rect 12094 32886 12110 32920
rect 12178 32886 12194 32920
rect 12094 32870 12194 32886
rect 12252 32920 12352 32958
rect 12252 32886 12268 32920
rect 12336 32886 12352 32920
rect 12252 32870 12352 32886
rect 12410 32920 12510 32958
rect 12410 32886 12426 32920
rect 12494 32886 12510 32920
rect 12410 32870 12510 32886
rect 14128 39030 14228 39046
rect 14128 38996 14144 39030
rect 14212 38996 14228 39030
rect 14128 38958 14228 38996
rect 14286 39030 14386 39046
rect 14286 38996 14302 39030
rect 14370 38996 14386 39030
rect 14286 38958 14386 38996
rect 14444 39030 14544 39046
rect 14444 38996 14460 39030
rect 14528 38996 14544 39030
rect 14444 38958 14544 38996
rect 14602 39030 14702 39046
rect 14602 38996 14618 39030
rect 14686 38996 14702 39030
rect 14602 38958 14702 38996
rect 14760 39030 14860 39046
rect 14760 38996 14776 39030
rect 14844 38996 14860 39030
rect 14760 38958 14860 38996
rect 14918 39030 15018 39046
rect 14918 38996 14934 39030
rect 15002 38996 15018 39030
rect 14918 38958 15018 38996
rect 15076 39030 15176 39046
rect 15076 38996 15092 39030
rect 15160 38996 15176 39030
rect 15076 38958 15176 38996
rect 15234 39030 15334 39046
rect 15234 38996 15250 39030
rect 15318 38996 15334 39030
rect 15234 38958 15334 38996
rect 15392 39030 15492 39046
rect 15392 38996 15408 39030
rect 15476 38996 15492 39030
rect 15392 38958 15492 38996
rect 15550 39030 15650 39046
rect 15550 38996 15566 39030
rect 15634 38996 15650 39030
rect 15550 38958 15650 38996
rect 15708 39030 15808 39046
rect 15708 38996 15724 39030
rect 15792 38996 15808 39030
rect 15708 38958 15808 38996
rect 15866 39030 15966 39046
rect 15866 38996 15882 39030
rect 15950 38996 15966 39030
rect 15866 38958 15966 38996
rect 16024 39030 16124 39046
rect 16024 38996 16040 39030
rect 16108 38996 16124 39030
rect 16024 38958 16124 38996
rect 16182 39030 16282 39046
rect 16182 38996 16198 39030
rect 16266 38996 16282 39030
rect 16182 38958 16282 38996
rect 16340 39030 16440 39046
rect 16340 38996 16356 39030
rect 16424 38996 16440 39030
rect 16340 38958 16440 38996
rect 16498 39030 16598 39046
rect 16498 38996 16514 39030
rect 16582 38996 16598 39030
rect 16498 38958 16598 38996
rect 16656 39030 16756 39046
rect 16656 38996 16672 39030
rect 16740 38996 16756 39030
rect 16656 38958 16756 38996
rect 16814 39030 16914 39046
rect 16814 38996 16830 39030
rect 16898 38996 16914 39030
rect 16814 38958 16914 38996
rect 16972 39030 17072 39046
rect 16972 38996 16988 39030
rect 17056 38996 17072 39030
rect 16972 38958 17072 38996
rect 17130 39030 17230 39046
rect 17130 38996 17146 39030
rect 17214 38996 17230 39030
rect 17130 38958 17230 38996
rect 17288 39030 17388 39046
rect 17288 38996 17304 39030
rect 17372 38996 17388 39030
rect 17288 38958 17388 38996
rect 17446 39030 17546 39046
rect 17446 38996 17462 39030
rect 17530 38996 17546 39030
rect 17446 38958 17546 38996
rect 17604 39030 17704 39046
rect 17604 38996 17620 39030
rect 17688 38996 17704 39030
rect 17604 38958 17704 38996
rect 17762 39030 17862 39046
rect 17762 38996 17778 39030
rect 17846 38996 17862 39030
rect 17762 38958 17862 38996
rect 17920 39030 18020 39046
rect 17920 38996 17936 39030
rect 18004 38996 18020 39030
rect 17920 38958 18020 38996
rect 18078 39030 18178 39046
rect 18078 38996 18094 39030
rect 18162 38996 18178 39030
rect 18078 38958 18178 38996
rect 18236 39030 18336 39046
rect 18236 38996 18252 39030
rect 18320 38996 18336 39030
rect 18236 38958 18336 38996
rect 18394 39030 18494 39046
rect 18394 38996 18410 39030
rect 18478 38996 18494 39030
rect 18394 38958 18494 38996
rect 18552 39030 18652 39046
rect 18552 38996 18568 39030
rect 18636 38996 18652 39030
rect 18552 38958 18652 38996
rect 18710 39030 18810 39046
rect 18710 38996 18726 39030
rect 18794 38996 18810 39030
rect 18710 38958 18810 38996
rect 14128 32920 14228 32958
rect 14128 32886 14144 32920
rect 14212 32886 14228 32920
rect 14128 32870 14228 32886
rect 14286 32920 14386 32958
rect 14286 32886 14302 32920
rect 14370 32886 14386 32920
rect 14286 32870 14386 32886
rect 14444 32920 14544 32958
rect 14444 32886 14460 32920
rect 14528 32886 14544 32920
rect 14444 32870 14544 32886
rect 14602 32920 14702 32958
rect 14602 32886 14618 32920
rect 14686 32886 14702 32920
rect 14602 32870 14702 32886
rect 14760 32920 14860 32958
rect 14760 32886 14776 32920
rect 14844 32886 14860 32920
rect 14760 32870 14860 32886
rect 14918 32920 15018 32958
rect 14918 32886 14934 32920
rect 15002 32886 15018 32920
rect 14918 32870 15018 32886
rect 15076 32920 15176 32958
rect 15076 32886 15092 32920
rect 15160 32886 15176 32920
rect 15076 32870 15176 32886
rect 15234 32920 15334 32958
rect 15234 32886 15250 32920
rect 15318 32886 15334 32920
rect 15234 32870 15334 32886
rect 15392 32920 15492 32958
rect 15392 32886 15408 32920
rect 15476 32886 15492 32920
rect 15392 32870 15492 32886
rect 15550 32920 15650 32958
rect 15550 32886 15566 32920
rect 15634 32886 15650 32920
rect 15550 32870 15650 32886
rect 15708 32920 15808 32958
rect 15708 32886 15724 32920
rect 15792 32886 15808 32920
rect 15708 32870 15808 32886
rect 15866 32920 15966 32958
rect 15866 32886 15882 32920
rect 15950 32886 15966 32920
rect 15866 32870 15966 32886
rect 16024 32920 16124 32958
rect 16024 32886 16040 32920
rect 16108 32886 16124 32920
rect 16024 32870 16124 32886
rect 16182 32920 16282 32958
rect 16182 32886 16198 32920
rect 16266 32886 16282 32920
rect 16182 32870 16282 32886
rect 16340 32920 16440 32958
rect 16340 32886 16356 32920
rect 16424 32886 16440 32920
rect 16340 32870 16440 32886
rect 16498 32920 16598 32958
rect 16498 32886 16514 32920
rect 16582 32886 16598 32920
rect 16498 32870 16598 32886
rect 16656 32920 16756 32958
rect 16656 32886 16672 32920
rect 16740 32886 16756 32920
rect 16656 32870 16756 32886
rect 16814 32920 16914 32958
rect 16814 32886 16830 32920
rect 16898 32886 16914 32920
rect 16814 32870 16914 32886
rect 16972 32920 17072 32958
rect 16972 32886 16988 32920
rect 17056 32886 17072 32920
rect 16972 32870 17072 32886
rect 17130 32920 17230 32958
rect 17130 32886 17146 32920
rect 17214 32886 17230 32920
rect 17130 32870 17230 32886
rect 17288 32920 17388 32958
rect 17288 32886 17304 32920
rect 17372 32886 17388 32920
rect 17288 32870 17388 32886
rect 17446 32920 17546 32958
rect 17446 32886 17462 32920
rect 17530 32886 17546 32920
rect 17446 32870 17546 32886
rect 17604 32920 17704 32958
rect 17604 32886 17620 32920
rect 17688 32886 17704 32920
rect 17604 32870 17704 32886
rect 17762 32920 17862 32958
rect 17762 32886 17778 32920
rect 17846 32886 17862 32920
rect 17762 32870 17862 32886
rect 17920 32920 18020 32958
rect 17920 32886 17936 32920
rect 18004 32886 18020 32920
rect 17920 32870 18020 32886
rect 18078 32920 18178 32958
rect 18078 32886 18094 32920
rect 18162 32886 18178 32920
rect 18078 32870 18178 32886
rect 18236 32920 18336 32958
rect 18236 32886 18252 32920
rect 18320 32886 18336 32920
rect 18236 32870 18336 32886
rect 18394 32920 18494 32958
rect 18394 32886 18410 32920
rect 18478 32886 18494 32920
rect 18394 32870 18494 32886
rect 18552 32920 18652 32958
rect 18552 32886 18568 32920
rect 18636 32886 18652 32920
rect 18552 32870 18652 32886
rect 18710 32920 18810 32958
rect 18710 32886 18726 32920
rect 18794 32886 18810 32920
rect 18710 32870 18810 32886
rect 20428 39030 20528 39046
rect 20428 38996 20444 39030
rect 20512 38996 20528 39030
rect 20428 38958 20528 38996
rect 20586 39030 20686 39046
rect 20586 38996 20602 39030
rect 20670 38996 20686 39030
rect 20586 38958 20686 38996
rect 20744 39030 20844 39046
rect 20744 38996 20760 39030
rect 20828 38996 20844 39030
rect 20744 38958 20844 38996
rect 20902 39030 21002 39046
rect 20902 38996 20918 39030
rect 20986 38996 21002 39030
rect 20902 38958 21002 38996
rect 21060 39030 21160 39046
rect 21060 38996 21076 39030
rect 21144 38996 21160 39030
rect 21060 38958 21160 38996
rect 21218 39030 21318 39046
rect 21218 38996 21234 39030
rect 21302 38996 21318 39030
rect 21218 38958 21318 38996
rect 21376 39030 21476 39046
rect 21376 38996 21392 39030
rect 21460 38996 21476 39030
rect 21376 38958 21476 38996
rect 21534 39030 21634 39046
rect 21534 38996 21550 39030
rect 21618 38996 21634 39030
rect 21534 38958 21634 38996
rect 21692 39030 21792 39046
rect 21692 38996 21708 39030
rect 21776 38996 21792 39030
rect 21692 38958 21792 38996
rect 21850 39030 21950 39046
rect 21850 38996 21866 39030
rect 21934 38996 21950 39030
rect 21850 38958 21950 38996
rect 22008 39030 22108 39046
rect 22008 38996 22024 39030
rect 22092 38996 22108 39030
rect 22008 38958 22108 38996
rect 22166 39030 22266 39046
rect 22166 38996 22182 39030
rect 22250 38996 22266 39030
rect 22166 38958 22266 38996
rect 22324 39030 22424 39046
rect 22324 38996 22340 39030
rect 22408 38996 22424 39030
rect 22324 38958 22424 38996
rect 22482 39030 22582 39046
rect 22482 38996 22498 39030
rect 22566 38996 22582 39030
rect 22482 38958 22582 38996
rect 22640 39030 22740 39046
rect 22640 38996 22656 39030
rect 22724 38996 22740 39030
rect 22640 38958 22740 38996
rect 22798 39030 22898 39046
rect 22798 38996 22814 39030
rect 22882 38996 22898 39030
rect 22798 38958 22898 38996
rect 22956 39030 23056 39046
rect 22956 38996 22972 39030
rect 23040 38996 23056 39030
rect 22956 38958 23056 38996
rect 23114 39030 23214 39046
rect 23114 38996 23130 39030
rect 23198 38996 23214 39030
rect 23114 38958 23214 38996
rect 23272 39030 23372 39046
rect 23272 38996 23288 39030
rect 23356 38996 23372 39030
rect 23272 38958 23372 38996
rect 23430 39030 23530 39046
rect 23430 38996 23446 39030
rect 23514 38996 23530 39030
rect 23430 38958 23530 38996
rect 23588 39030 23688 39046
rect 23588 38996 23604 39030
rect 23672 38996 23688 39030
rect 23588 38958 23688 38996
rect 23746 39030 23846 39046
rect 23746 38996 23762 39030
rect 23830 38996 23846 39030
rect 23746 38958 23846 38996
rect 23904 39030 24004 39046
rect 23904 38996 23920 39030
rect 23988 38996 24004 39030
rect 23904 38958 24004 38996
rect 24062 39030 24162 39046
rect 24062 38996 24078 39030
rect 24146 38996 24162 39030
rect 24062 38958 24162 38996
rect 24220 39030 24320 39046
rect 24220 38996 24236 39030
rect 24304 38996 24320 39030
rect 24220 38958 24320 38996
rect 24378 39030 24478 39046
rect 24378 38996 24394 39030
rect 24462 38996 24478 39030
rect 24378 38958 24478 38996
rect 24536 39030 24636 39046
rect 24536 38996 24552 39030
rect 24620 38996 24636 39030
rect 24536 38958 24636 38996
rect 24694 39030 24794 39046
rect 24694 38996 24710 39030
rect 24778 38996 24794 39030
rect 24694 38958 24794 38996
rect 24852 39030 24952 39046
rect 24852 38996 24868 39030
rect 24936 38996 24952 39030
rect 24852 38958 24952 38996
rect 25010 39030 25110 39046
rect 25010 38996 25026 39030
rect 25094 38996 25110 39030
rect 25010 38958 25110 38996
rect 20428 32920 20528 32958
rect 20428 32886 20444 32920
rect 20512 32886 20528 32920
rect 20428 32870 20528 32886
rect 20586 32920 20686 32958
rect 20586 32886 20602 32920
rect 20670 32886 20686 32920
rect 20586 32870 20686 32886
rect 20744 32920 20844 32958
rect 20744 32886 20760 32920
rect 20828 32886 20844 32920
rect 20744 32870 20844 32886
rect 20902 32920 21002 32958
rect 20902 32886 20918 32920
rect 20986 32886 21002 32920
rect 20902 32870 21002 32886
rect 21060 32920 21160 32958
rect 21060 32886 21076 32920
rect 21144 32886 21160 32920
rect 21060 32870 21160 32886
rect 21218 32920 21318 32958
rect 21218 32886 21234 32920
rect 21302 32886 21318 32920
rect 21218 32870 21318 32886
rect 21376 32920 21476 32958
rect 21376 32886 21392 32920
rect 21460 32886 21476 32920
rect 21376 32870 21476 32886
rect 21534 32920 21634 32958
rect 21534 32886 21550 32920
rect 21618 32886 21634 32920
rect 21534 32870 21634 32886
rect 21692 32920 21792 32958
rect 21692 32886 21708 32920
rect 21776 32886 21792 32920
rect 21692 32870 21792 32886
rect 21850 32920 21950 32958
rect 21850 32886 21866 32920
rect 21934 32886 21950 32920
rect 21850 32870 21950 32886
rect 22008 32920 22108 32958
rect 22008 32886 22024 32920
rect 22092 32886 22108 32920
rect 22008 32870 22108 32886
rect 22166 32920 22266 32958
rect 22166 32886 22182 32920
rect 22250 32886 22266 32920
rect 22166 32870 22266 32886
rect 22324 32920 22424 32958
rect 22324 32886 22340 32920
rect 22408 32886 22424 32920
rect 22324 32870 22424 32886
rect 22482 32920 22582 32958
rect 22482 32886 22498 32920
rect 22566 32886 22582 32920
rect 22482 32870 22582 32886
rect 22640 32920 22740 32958
rect 22640 32886 22656 32920
rect 22724 32886 22740 32920
rect 22640 32870 22740 32886
rect 22798 32920 22898 32958
rect 22798 32886 22814 32920
rect 22882 32886 22898 32920
rect 22798 32870 22898 32886
rect 22956 32920 23056 32958
rect 22956 32886 22972 32920
rect 23040 32886 23056 32920
rect 22956 32870 23056 32886
rect 23114 32920 23214 32958
rect 23114 32886 23130 32920
rect 23198 32886 23214 32920
rect 23114 32870 23214 32886
rect 23272 32920 23372 32958
rect 23272 32886 23288 32920
rect 23356 32886 23372 32920
rect 23272 32870 23372 32886
rect 23430 32920 23530 32958
rect 23430 32886 23446 32920
rect 23514 32886 23530 32920
rect 23430 32870 23530 32886
rect 23588 32920 23688 32958
rect 23588 32886 23604 32920
rect 23672 32886 23688 32920
rect 23588 32870 23688 32886
rect 23746 32920 23846 32958
rect 23746 32886 23762 32920
rect 23830 32886 23846 32920
rect 23746 32870 23846 32886
rect 23904 32920 24004 32958
rect 23904 32886 23920 32920
rect 23988 32886 24004 32920
rect 23904 32870 24004 32886
rect 24062 32920 24162 32958
rect 24062 32886 24078 32920
rect 24146 32886 24162 32920
rect 24062 32870 24162 32886
rect 24220 32920 24320 32958
rect 24220 32886 24236 32920
rect 24304 32886 24320 32920
rect 24220 32870 24320 32886
rect 24378 32920 24478 32958
rect 24378 32886 24394 32920
rect 24462 32886 24478 32920
rect 24378 32870 24478 32886
rect 24536 32920 24636 32958
rect 24536 32886 24552 32920
rect 24620 32886 24636 32920
rect 24536 32870 24636 32886
rect 24694 32920 24794 32958
rect 24694 32886 24710 32920
rect 24778 32886 24794 32920
rect 24694 32870 24794 32886
rect 24852 32920 24952 32958
rect 24852 32886 24868 32920
rect 24936 32886 24952 32920
rect 24852 32870 24952 32886
rect 25010 32920 25110 32958
rect 25010 32886 25026 32920
rect 25094 32886 25110 32920
rect 25010 32870 25110 32886
rect 29968 40276 30034 40292
rect 29968 40242 29984 40276
rect 30018 40242 30034 40276
rect 29968 40219 30034 40242
rect 29968 38896 30034 38919
rect 29968 38862 29984 38896
rect 30018 38862 30034 38896
rect 29968 38846 30034 38862
rect -4234 27076 -4168 27092
rect -4234 27042 -4218 27076
rect -4184 27042 -4168 27076
rect -4234 27019 -4168 27042
rect -4234 25696 -4168 25719
rect -4234 25662 -4218 25696
rect -4184 25662 -4168 25696
rect -4234 25646 -4168 25662
rect 1528 30730 1628 30746
rect 1528 30696 1544 30730
rect 1612 30696 1628 30730
rect 1528 30658 1628 30696
rect 1686 30730 1786 30746
rect 1686 30696 1702 30730
rect 1770 30696 1786 30730
rect 1686 30658 1786 30696
rect 1844 30730 1944 30746
rect 1844 30696 1860 30730
rect 1928 30696 1944 30730
rect 1844 30658 1944 30696
rect 2002 30730 2102 30746
rect 2002 30696 2018 30730
rect 2086 30696 2102 30730
rect 2002 30658 2102 30696
rect 2160 30730 2260 30746
rect 2160 30696 2176 30730
rect 2244 30696 2260 30730
rect 2160 30658 2260 30696
rect 2318 30730 2418 30746
rect 2318 30696 2334 30730
rect 2402 30696 2418 30730
rect 2318 30658 2418 30696
rect 2476 30730 2576 30746
rect 2476 30696 2492 30730
rect 2560 30696 2576 30730
rect 2476 30658 2576 30696
rect 2634 30730 2734 30746
rect 2634 30696 2650 30730
rect 2718 30696 2734 30730
rect 2634 30658 2734 30696
rect 2792 30730 2892 30746
rect 2792 30696 2808 30730
rect 2876 30696 2892 30730
rect 2792 30658 2892 30696
rect 2950 30730 3050 30746
rect 2950 30696 2966 30730
rect 3034 30696 3050 30730
rect 2950 30658 3050 30696
rect 3108 30730 3208 30746
rect 3108 30696 3124 30730
rect 3192 30696 3208 30730
rect 3108 30658 3208 30696
rect 3266 30730 3366 30746
rect 3266 30696 3282 30730
rect 3350 30696 3366 30730
rect 3266 30658 3366 30696
rect 3424 30730 3524 30746
rect 3424 30696 3440 30730
rect 3508 30696 3524 30730
rect 3424 30658 3524 30696
rect 3582 30730 3682 30746
rect 3582 30696 3598 30730
rect 3666 30696 3682 30730
rect 3582 30658 3682 30696
rect 3740 30730 3840 30746
rect 3740 30696 3756 30730
rect 3824 30696 3840 30730
rect 3740 30658 3840 30696
rect 3898 30730 3998 30746
rect 3898 30696 3914 30730
rect 3982 30696 3998 30730
rect 3898 30658 3998 30696
rect 4056 30730 4156 30746
rect 4056 30696 4072 30730
rect 4140 30696 4156 30730
rect 4056 30658 4156 30696
rect 4214 30730 4314 30746
rect 4214 30696 4230 30730
rect 4298 30696 4314 30730
rect 4214 30658 4314 30696
rect 4372 30730 4472 30746
rect 4372 30696 4388 30730
rect 4456 30696 4472 30730
rect 4372 30658 4472 30696
rect 4530 30730 4630 30746
rect 4530 30696 4546 30730
rect 4614 30696 4630 30730
rect 4530 30658 4630 30696
rect 4688 30730 4788 30746
rect 4688 30696 4704 30730
rect 4772 30696 4788 30730
rect 4688 30658 4788 30696
rect 4846 30730 4946 30746
rect 4846 30696 4862 30730
rect 4930 30696 4946 30730
rect 4846 30658 4946 30696
rect 5004 30730 5104 30746
rect 5004 30696 5020 30730
rect 5088 30696 5104 30730
rect 5004 30658 5104 30696
rect 5162 30730 5262 30746
rect 5162 30696 5178 30730
rect 5246 30696 5262 30730
rect 5162 30658 5262 30696
rect 5320 30730 5420 30746
rect 5320 30696 5336 30730
rect 5404 30696 5420 30730
rect 5320 30658 5420 30696
rect 5478 30730 5578 30746
rect 5478 30696 5494 30730
rect 5562 30696 5578 30730
rect 5478 30658 5578 30696
rect 5636 30730 5736 30746
rect 5636 30696 5652 30730
rect 5720 30696 5736 30730
rect 5636 30658 5736 30696
rect 5794 30730 5894 30746
rect 5794 30696 5810 30730
rect 5878 30696 5894 30730
rect 5794 30658 5894 30696
rect 5952 30730 6052 30746
rect 5952 30696 5968 30730
rect 6036 30696 6052 30730
rect 5952 30658 6052 30696
rect 6110 30730 6210 30746
rect 6110 30696 6126 30730
rect 6194 30696 6210 30730
rect 6110 30658 6210 30696
rect 1528 24620 1628 24658
rect 1528 24586 1544 24620
rect 1612 24586 1628 24620
rect 1528 24570 1628 24586
rect 1686 24620 1786 24658
rect 1686 24586 1702 24620
rect 1770 24586 1786 24620
rect 1686 24570 1786 24586
rect 1844 24620 1944 24658
rect 1844 24586 1860 24620
rect 1928 24586 1944 24620
rect 1844 24570 1944 24586
rect 2002 24620 2102 24658
rect 2002 24586 2018 24620
rect 2086 24586 2102 24620
rect 2002 24570 2102 24586
rect 2160 24620 2260 24658
rect 2160 24586 2176 24620
rect 2244 24586 2260 24620
rect 2160 24570 2260 24586
rect 2318 24620 2418 24658
rect 2318 24586 2334 24620
rect 2402 24586 2418 24620
rect 2318 24570 2418 24586
rect 2476 24620 2576 24658
rect 2476 24586 2492 24620
rect 2560 24586 2576 24620
rect 2476 24570 2576 24586
rect 2634 24620 2734 24658
rect 2634 24586 2650 24620
rect 2718 24586 2734 24620
rect 2634 24570 2734 24586
rect 2792 24620 2892 24658
rect 2792 24586 2808 24620
rect 2876 24586 2892 24620
rect 2792 24570 2892 24586
rect 2950 24620 3050 24658
rect 2950 24586 2966 24620
rect 3034 24586 3050 24620
rect 2950 24570 3050 24586
rect 3108 24620 3208 24658
rect 3108 24586 3124 24620
rect 3192 24586 3208 24620
rect 3108 24570 3208 24586
rect 3266 24620 3366 24658
rect 3266 24586 3282 24620
rect 3350 24586 3366 24620
rect 3266 24570 3366 24586
rect 3424 24620 3524 24658
rect 3424 24586 3440 24620
rect 3508 24586 3524 24620
rect 3424 24570 3524 24586
rect 3582 24620 3682 24658
rect 3582 24586 3598 24620
rect 3666 24586 3682 24620
rect 3582 24570 3682 24586
rect 3740 24620 3840 24658
rect 3740 24586 3756 24620
rect 3824 24586 3840 24620
rect 3740 24570 3840 24586
rect 3898 24620 3998 24658
rect 3898 24586 3914 24620
rect 3982 24586 3998 24620
rect 3898 24570 3998 24586
rect 4056 24620 4156 24658
rect 4056 24586 4072 24620
rect 4140 24586 4156 24620
rect 4056 24570 4156 24586
rect 4214 24620 4314 24658
rect 4214 24586 4230 24620
rect 4298 24586 4314 24620
rect 4214 24570 4314 24586
rect 4372 24620 4472 24658
rect 4372 24586 4388 24620
rect 4456 24586 4472 24620
rect 4372 24570 4472 24586
rect 4530 24620 4630 24658
rect 4530 24586 4546 24620
rect 4614 24586 4630 24620
rect 4530 24570 4630 24586
rect 4688 24620 4788 24658
rect 4688 24586 4704 24620
rect 4772 24586 4788 24620
rect 4688 24570 4788 24586
rect 4846 24620 4946 24658
rect 4846 24586 4862 24620
rect 4930 24586 4946 24620
rect 4846 24570 4946 24586
rect 5004 24620 5104 24658
rect 5004 24586 5020 24620
rect 5088 24586 5104 24620
rect 5004 24570 5104 24586
rect 5162 24620 5262 24658
rect 5162 24586 5178 24620
rect 5246 24586 5262 24620
rect 5162 24570 5262 24586
rect 5320 24620 5420 24658
rect 5320 24586 5336 24620
rect 5404 24586 5420 24620
rect 5320 24570 5420 24586
rect 5478 24620 5578 24658
rect 5478 24586 5494 24620
rect 5562 24586 5578 24620
rect 5478 24570 5578 24586
rect 5636 24620 5736 24658
rect 5636 24586 5652 24620
rect 5720 24586 5736 24620
rect 5636 24570 5736 24586
rect 5794 24620 5894 24658
rect 5794 24586 5810 24620
rect 5878 24586 5894 24620
rect 5794 24570 5894 24586
rect 5952 24620 6052 24658
rect 5952 24586 5968 24620
rect 6036 24586 6052 24620
rect 5952 24570 6052 24586
rect 6110 24620 6210 24658
rect 6110 24586 6126 24620
rect 6194 24586 6210 24620
rect 6110 24570 6210 24586
rect 7828 30730 7928 30746
rect 7828 30696 7844 30730
rect 7912 30696 7928 30730
rect 7828 30658 7928 30696
rect 7986 30730 8086 30746
rect 7986 30696 8002 30730
rect 8070 30696 8086 30730
rect 7986 30658 8086 30696
rect 8144 30730 8244 30746
rect 8144 30696 8160 30730
rect 8228 30696 8244 30730
rect 8144 30658 8244 30696
rect 8302 30730 8402 30746
rect 8302 30696 8318 30730
rect 8386 30696 8402 30730
rect 8302 30658 8402 30696
rect 8460 30730 8560 30746
rect 8460 30696 8476 30730
rect 8544 30696 8560 30730
rect 8460 30658 8560 30696
rect 8618 30730 8718 30746
rect 8618 30696 8634 30730
rect 8702 30696 8718 30730
rect 8618 30658 8718 30696
rect 8776 30730 8876 30746
rect 8776 30696 8792 30730
rect 8860 30696 8876 30730
rect 8776 30658 8876 30696
rect 8934 30730 9034 30746
rect 8934 30696 8950 30730
rect 9018 30696 9034 30730
rect 8934 30658 9034 30696
rect 9092 30730 9192 30746
rect 9092 30696 9108 30730
rect 9176 30696 9192 30730
rect 9092 30658 9192 30696
rect 9250 30730 9350 30746
rect 9250 30696 9266 30730
rect 9334 30696 9350 30730
rect 9250 30658 9350 30696
rect 9408 30730 9508 30746
rect 9408 30696 9424 30730
rect 9492 30696 9508 30730
rect 9408 30658 9508 30696
rect 9566 30730 9666 30746
rect 9566 30696 9582 30730
rect 9650 30696 9666 30730
rect 9566 30658 9666 30696
rect 9724 30730 9824 30746
rect 9724 30696 9740 30730
rect 9808 30696 9824 30730
rect 9724 30658 9824 30696
rect 9882 30730 9982 30746
rect 9882 30696 9898 30730
rect 9966 30696 9982 30730
rect 9882 30658 9982 30696
rect 10040 30730 10140 30746
rect 10040 30696 10056 30730
rect 10124 30696 10140 30730
rect 10040 30658 10140 30696
rect 10198 30730 10298 30746
rect 10198 30696 10214 30730
rect 10282 30696 10298 30730
rect 10198 30658 10298 30696
rect 10356 30730 10456 30746
rect 10356 30696 10372 30730
rect 10440 30696 10456 30730
rect 10356 30658 10456 30696
rect 10514 30730 10614 30746
rect 10514 30696 10530 30730
rect 10598 30696 10614 30730
rect 10514 30658 10614 30696
rect 10672 30730 10772 30746
rect 10672 30696 10688 30730
rect 10756 30696 10772 30730
rect 10672 30658 10772 30696
rect 10830 30730 10930 30746
rect 10830 30696 10846 30730
rect 10914 30696 10930 30730
rect 10830 30658 10930 30696
rect 10988 30730 11088 30746
rect 10988 30696 11004 30730
rect 11072 30696 11088 30730
rect 10988 30658 11088 30696
rect 11146 30730 11246 30746
rect 11146 30696 11162 30730
rect 11230 30696 11246 30730
rect 11146 30658 11246 30696
rect 11304 30730 11404 30746
rect 11304 30696 11320 30730
rect 11388 30696 11404 30730
rect 11304 30658 11404 30696
rect 11462 30730 11562 30746
rect 11462 30696 11478 30730
rect 11546 30696 11562 30730
rect 11462 30658 11562 30696
rect 11620 30730 11720 30746
rect 11620 30696 11636 30730
rect 11704 30696 11720 30730
rect 11620 30658 11720 30696
rect 11778 30730 11878 30746
rect 11778 30696 11794 30730
rect 11862 30696 11878 30730
rect 11778 30658 11878 30696
rect 11936 30730 12036 30746
rect 11936 30696 11952 30730
rect 12020 30696 12036 30730
rect 11936 30658 12036 30696
rect 12094 30730 12194 30746
rect 12094 30696 12110 30730
rect 12178 30696 12194 30730
rect 12094 30658 12194 30696
rect 12252 30730 12352 30746
rect 12252 30696 12268 30730
rect 12336 30696 12352 30730
rect 12252 30658 12352 30696
rect 12410 30730 12510 30746
rect 12410 30696 12426 30730
rect 12494 30696 12510 30730
rect 12410 30658 12510 30696
rect 7828 24620 7928 24658
rect 7828 24586 7844 24620
rect 7912 24586 7928 24620
rect 7828 24570 7928 24586
rect 7986 24620 8086 24658
rect 7986 24586 8002 24620
rect 8070 24586 8086 24620
rect 7986 24570 8086 24586
rect 8144 24620 8244 24658
rect 8144 24586 8160 24620
rect 8228 24586 8244 24620
rect 8144 24570 8244 24586
rect 8302 24620 8402 24658
rect 8302 24586 8318 24620
rect 8386 24586 8402 24620
rect 8302 24570 8402 24586
rect 8460 24620 8560 24658
rect 8460 24586 8476 24620
rect 8544 24586 8560 24620
rect 8460 24570 8560 24586
rect 8618 24620 8718 24658
rect 8618 24586 8634 24620
rect 8702 24586 8718 24620
rect 8618 24570 8718 24586
rect 8776 24620 8876 24658
rect 8776 24586 8792 24620
rect 8860 24586 8876 24620
rect 8776 24570 8876 24586
rect 8934 24620 9034 24658
rect 8934 24586 8950 24620
rect 9018 24586 9034 24620
rect 8934 24570 9034 24586
rect 9092 24620 9192 24658
rect 9092 24586 9108 24620
rect 9176 24586 9192 24620
rect 9092 24570 9192 24586
rect 9250 24620 9350 24658
rect 9250 24586 9266 24620
rect 9334 24586 9350 24620
rect 9250 24570 9350 24586
rect 9408 24620 9508 24658
rect 9408 24586 9424 24620
rect 9492 24586 9508 24620
rect 9408 24570 9508 24586
rect 9566 24620 9666 24658
rect 9566 24586 9582 24620
rect 9650 24586 9666 24620
rect 9566 24570 9666 24586
rect 9724 24620 9824 24658
rect 9724 24586 9740 24620
rect 9808 24586 9824 24620
rect 9724 24570 9824 24586
rect 9882 24620 9982 24658
rect 9882 24586 9898 24620
rect 9966 24586 9982 24620
rect 9882 24570 9982 24586
rect 10040 24620 10140 24658
rect 10040 24586 10056 24620
rect 10124 24586 10140 24620
rect 10040 24570 10140 24586
rect 10198 24620 10298 24658
rect 10198 24586 10214 24620
rect 10282 24586 10298 24620
rect 10198 24570 10298 24586
rect 10356 24620 10456 24658
rect 10356 24586 10372 24620
rect 10440 24586 10456 24620
rect 10356 24570 10456 24586
rect 10514 24620 10614 24658
rect 10514 24586 10530 24620
rect 10598 24586 10614 24620
rect 10514 24570 10614 24586
rect 10672 24620 10772 24658
rect 10672 24586 10688 24620
rect 10756 24586 10772 24620
rect 10672 24570 10772 24586
rect 10830 24620 10930 24658
rect 10830 24586 10846 24620
rect 10914 24586 10930 24620
rect 10830 24570 10930 24586
rect 10988 24620 11088 24658
rect 10988 24586 11004 24620
rect 11072 24586 11088 24620
rect 10988 24570 11088 24586
rect 11146 24620 11246 24658
rect 11146 24586 11162 24620
rect 11230 24586 11246 24620
rect 11146 24570 11246 24586
rect 11304 24620 11404 24658
rect 11304 24586 11320 24620
rect 11388 24586 11404 24620
rect 11304 24570 11404 24586
rect 11462 24620 11562 24658
rect 11462 24586 11478 24620
rect 11546 24586 11562 24620
rect 11462 24570 11562 24586
rect 11620 24620 11720 24658
rect 11620 24586 11636 24620
rect 11704 24586 11720 24620
rect 11620 24570 11720 24586
rect 11778 24620 11878 24658
rect 11778 24586 11794 24620
rect 11862 24586 11878 24620
rect 11778 24570 11878 24586
rect 11936 24620 12036 24658
rect 11936 24586 11952 24620
rect 12020 24586 12036 24620
rect 11936 24570 12036 24586
rect 12094 24620 12194 24658
rect 12094 24586 12110 24620
rect 12178 24586 12194 24620
rect 12094 24570 12194 24586
rect 12252 24620 12352 24658
rect 12252 24586 12268 24620
rect 12336 24586 12352 24620
rect 12252 24570 12352 24586
rect 12410 24620 12510 24658
rect 12410 24586 12426 24620
rect 12494 24586 12510 24620
rect 12410 24570 12510 24586
rect 14128 30730 14228 30746
rect 14128 30696 14144 30730
rect 14212 30696 14228 30730
rect 14128 30658 14228 30696
rect 14286 30730 14386 30746
rect 14286 30696 14302 30730
rect 14370 30696 14386 30730
rect 14286 30658 14386 30696
rect 14444 30730 14544 30746
rect 14444 30696 14460 30730
rect 14528 30696 14544 30730
rect 14444 30658 14544 30696
rect 14602 30730 14702 30746
rect 14602 30696 14618 30730
rect 14686 30696 14702 30730
rect 14602 30658 14702 30696
rect 14760 30730 14860 30746
rect 14760 30696 14776 30730
rect 14844 30696 14860 30730
rect 14760 30658 14860 30696
rect 14918 30730 15018 30746
rect 14918 30696 14934 30730
rect 15002 30696 15018 30730
rect 14918 30658 15018 30696
rect 15076 30730 15176 30746
rect 15076 30696 15092 30730
rect 15160 30696 15176 30730
rect 15076 30658 15176 30696
rect 15234 30730 15334 30746
rect 15234 30696 15250 30730
rect 15318 30696 15334 30730
rect 15234 30658 15334 30696
rect 15392 30730 15492 30746
rect 15392 30696 15408 30730
rect 15476 30696 15492 30730
rect 15392 30658 15492 30696
rect 15550 30730 15650 30746
rect 15550 30696 15566 30730
rect 15634 30696 15650 30730
rect 15550 30658 15650 30696
rect 15708 30730 15808 30746
rect 15708 30696 15724 30730
rect 15792 30696 15808 30730
rect 15708 30658 15808 30696
rect 15866 30730 15966 30746
rect 15866 30696 15882 30730
rect 15950 30696 15966 30730
rect 15866 30658 15966 30696
rect 16024 30730 16124 30746
rect 16024 30696 16040 30730
rect 16108 30696 16124 30730
rect 16024 30658 16124 30696
rect 16182 30730 16282 30746
rect 16182 30696 16198 30730
rect 16266 30696 16282 30730
rect 16182 30658 16282 30696
rect 16340 30730 16440 30746
rect 16340 30696 16356 30730
rect 16424 30696 16440 30730
rect 16340 30658 16440 30696
rect 16498 30730 16598 30746
rect 16498 30696 16514 30730
rect 16582 30696 16598 30730
rect 16498 30658 16598 30696
rect 16656 30730 16756 30746
rect 16656 30696 16672 30730
rect 16740 30696 16756 30730
rect 16656 30658 16756 30696
rect 16814 30730 16914 30746
rect 16814 30696 16830 30730
rect 16898 30696 16914 30730
rect 16814 30658 16914 30696
rect 16972 30730 17072 30746
rect 16972 30696 16988 30730
rect 17056 30696 17072 30730
rect 16972 30658 17072 30696
rect 17130 30730 17230 30746
rect 17130 30696 17146 30730
rect 17214 30696 17230 30730
rect 17130 30658 17230 30696
rect 17288 30730 17388 30746
rect 17288 30696 17304 30730
rect 17372 30696 17388 30730
rect 17288 30658 17388 30696
rect 17446 30730 17546 30746
rect 17446 30696 17462 30730
rect 17530 30696 17546 30730
rect 17446 30658 17546 30696
rect 17604 30730 17704 30746
rect 17604 30696 17620 30730
rect 17688 30696 17704 30730
rect 17604 30658 17704 30696
rect 17762 30730 17862 30746
rect 17762 30696 17778 30730
rect 17846 30696 17862 30730
rect 17762 30658 17862 30696
rect 17920 30730 18020 30746
rect 17920 30696 17936 30730
rect 18004 30696 18020 30730
rect 17920 30658 18020 30696
rect 18078 30730 18178 30746
rect 18078 30696 18094 30730
rect 18162 30696 18178 30730
rect 18078 30658 18178 30696
rect 18236 30730 18336 30746
rect 18236 30696 18252 30730
rect 18320 30696 18336 30730
rect 18236 30658 18336 30696
rect 18394 30730 18494 30746
rect 18394 30696 18410 30730
rect 18478 30696 18494 30730
rect 18394 30658 18494 30696
rect 18552 30730 18652 30746
rect 18552 30696 18568 30730
rect 18636 30696 18652 30730
rect 18552 30658 18652 30696
rect 18710 30730 18810 30746
rect 18710 30696 18726 30730
rect 18794 30696 18810 30730
rect 18710 30658 18810 30696
rect 14128 24620 14228 24658
rect 14128 24586 14144 24620
rect 14212 24586 14228 24620
rect 14128 24570 14228 24586
rect 14286 24620 14386 24658
rect 14286 24586 14302 24620
rect 14370 24586 14386 24620
rect 14286 24570 14386 24586
rect 14444 24620 14544 24658
rect 14444 24586 14460 24620
rect 14528 24586 14544 24620
rect 14444 24570 14544 24586
rect 14602 24620 14702 24658
rect 14602 24586 14618 24620
rect 14686 24586 14702 24620
rect 14602 24570 14702 24586
rect 14760 24620 14860 24658
rect 14760 24586 14776 24620
rect 14844 24586 14860 24620
rect 14760 24570 14860 24586
rect 14918 24620 15018 24658
rect 14918 24586 14934 24620
rect 15002 24586 15018 24620
rect 14918 24570 15018 24586
rect 15076 24620 15176 24658
rect 15076 24586 15092 24620
rect 15160 24586 15176 24620
rect 15076 24570 15176 24586
rect 15234 24620 15334 24658
rect 15234 24586 15250 24620
rect 15318 24586 15334 24620
rect 15234 24570 15334 24586
rect 15392 24620 15492 24658
rect 15392 24586 15408 24620
rect 15476 24586 15492 24620
rect 15392 24570 15492 24586
rect 15550 24620 15650 24658
rect 15550 24586 15566 24620
rect 15634 24586 15650 24620
rect 15550 24570 15650 24586
rect 15708 24620 15808 24658
rect 15708 24586 15724 24620
rect 15792 24586 15808 24620
rect 15708 24570 15808 24586
rect 15866 24620 15966 24658
rect 15866 24586 15882 24620
rect 15950 24586 15966 24620
rect 15866 24570 15966 24586
rect 16024 24620 16124 24658
rect 16024 24586 16040 24620
rect 16108 24586 16124 24620
rect 16024 24570 16124 24586
rect 16182 24620 16282 24658
rect 16182 24586 16198 24620
rect 16266 24586 16282 24620
rect 16182 24570 16282 24586
rect 16340 24620 16440 24658
rect 16340 24586 16356 24620
rect 16424 24586 16440 24620
rect 16340 24570 16440 24586
rect 16498 24620 16598 24658
rect 16498 24586 16514 24620
rect 16582 24586 16598 24620
rect 16498 24570 16598 24586
rect 16656 24620 16756 24658
rect 16656 24586 16672 24620
rect 16740 24586 16756 24620
rect 16656 24570 16756 24586
rect 16814 24620 16914 24658
rect 16814 24586 16830 24620
rect 16898 24586 16914 24620
rect 16814 24570 16914 24586
rect 16972 24620 17072 24658
rect 16972 24586 16988 24620
rect 17056 24586 17072 24620
rect 16972 24570 17072 24586
rect 17130 24620 17230 24658
rect 17130 24586 17146 24620
rect 17214 24586 17230 24620
rect 17130 24570 17230 24586
rect 17288 24620 17388 24658
rect 17288 24586 17304 24620
rect 17372 24586 17388 24620
rect 17288 24570 17388 24586
rect 17446 24620 17546 24658
rect 17446 24586 17462 24620
rect 17530 24586 17546 24620
rect 17446 24570 17546 24586
rect 17604 24620 17704 24658
rect 17604 24586 17620 24620
rect 17688 24586 17704 24620
rect 17604 24570 17704 24586
rect 17762 24620 17862 24658
rect 17762 24586 17778 24620
rect 17846 24586 17862 24620
rect 17762 24570 17862 24586
rect 17920 24620 18020 24658
rect 17920 24586 17936 24620
rect 18004 24586 18020 24620
rect 17920 24570 18020 24586
rect 18078 24620 18178 24658
rect 18078 24586 18094 24620
rect 18162 24586 18178 24620
rect 18078 24570 18178 24586
rect 18236 24620 18336 24658
rect 18236 24586 18252 24620
rect 18320 24586 18336 24620
rect 18236 24570 18336 24586
rect 18394 24620 18494 24658
rect 18394 24586 18410 24620
rect 18478 24586 18494 24620
rect 18394 24570 18494 24586
rect 18552 24620 18652 24658
rect 18552 24586 18568 24620
rect 18636 24586 18652 24620
rect 18552 24570 18652 24586
rect 18710 24620 18810 24658
rect 18710 24586 18726 24620
rect 18794 24586 18810 24620
rect 18710 24570 18810 24586
rect 20428 30730 20528 30746
rect 20428 30696 20444 30730
rect 20512 30696 20528 30730
rect 20428 30658 20528 30696
rect 20586 30730 20686 30746
rect 20586 30696 20602 30730
rect 20670 30696 20686 30730
rect 20586 30658 20686 30696
rect 20744 30730 20844 30746
rect 20744 30696 20760 30730
rect 20828 30696 20844 30730
rect 20744 30658 20844 30696
rect 20902 30730 21002 30746
rect 20902 30696 20918 30730
rect 20986 30696 21002 30730
rect 20902 30658 21002 30696
rect 21060 30730 21160 30746
rect 21060 30696 21076 30730
rect 21144 30696 21160 30730
rect 21060 30658 21160 30696
rect 21218 30730 21318 30746
rect 21218 30696 21234 30730
rect 21302 30696 21318 30730
rect 21218 30658 21318 30696
rect 21376 30730 21476 30746
rect 21376 30696 21392 30730
rect 21460 30696 21476 30730
rect 21376 30658 21476 30696
rect 21534 30730 21634 30746
rect 21534 30696 21550 30730
rect 21618 30696 21634 30730
rect 21534 30658 21634 30696
rect 21692 30730 21792 30746
rect 21692 30696 21708 30730
rect 21776 30696 21792 30730
rect 21692 30658 21792 30696
rect 21850 30730 21950 30746
rect 21850 30696 21866 30730
rect 21934 30696 21950 30730
rect 21850 30658 21950 30696
rect 22008 30730 22108 30746
rect 22008 30696 22024 30730
rect 22092 30696 22108 30730
rect 22008 30658 22108 30696
rect 22166 30730 22266 30746
rect 22166 30696 22182 30730
rect 22250 30696 22266 30730
rect 22166 30658 22266 30696
rect 22324 30730 22424 30746
rect 22324 30696 22340 30730
rect 22408 30696 22424 30730
rect 22324 30658 22424 30696
rect 22482 30730 22582 30746
rect 22482 30696 22498 30730
rect 22566 30696 22582 30730
rect 22482 30658 22582 30696
rect 22640 30730 22740 30746
rect 22640 30696 22656 30730
rect 22724 30696 22740 30730
rect 22640 30658 22740 30696
rect 22798 30730 22898 30746
rect 22798 30696 22814 30730
rect 22882 30696 22898 30730
rect 22798 30658 22898 30696
rect 22956 30730 23056 30746
rect 22956 30696 22972 30730
rect 23040 30696 23056 30730
rect 22956 30658 23056 30696
rect 23114 30730 23214 30746
rect 23114 30696 23130 30730
rect 23198 30696 23214 30730
rect 23114 30658 23214 30696
rect 23272 30730 23372 30746
rect 23272 30696 23288 30730
rect 23356 30696 23372 30730
rect 23272 30658 23372 30696
rect 23430 30730 23530 30746
rect 23430 30696 23446 30730
rect 23514 30696 23530 30730
rect 23430 30658 23530 30696
rect 23588 30730 23688 30746
rect 23588 30696 23604 30730
rect 23672 30696 23688 30730
rect 23588 30658 23688 30696
rect 23746 30730 23846 30746
rect 23746 30696 23762 30730
rect 23830 30696 23846 30730
rect 23746 30658 23846 30696
rect 23904 30730 24004 30746
rect 23904 30696 23920 30730
rect 23988 30696 24004 30730
rect 23904 30658 24004 30696
rect 24062 30730 24162 30746
rect 24062 30696 24078 30730
rect 24146 30696 24162 30730
rect 24062 30658 24162 30696
rect 24220 30730 24320 30746
rect 24220 30696 24236 30730
rect 24304 30696 24320 30730
rect 24220 30658 24320 30696
rect 24378 30730 24478 30746
rect 24378 30696 24394 30730
rect 24462 30696 24478 30730
rect 24378 30658 24478 30696
rect 24536 30730 24636 30746
rect 24536 30696 24552 30730
rect 24620 30696 24636 30730
rect 24536 30658 24636 30696
rect 24694 30730 24794 30746
rect 24694 30696 24710 30730
rect 24778 30696 24794 30730
rect 24694 30658 24794 30696
rect 24852 30730 24952 30746
rect 24852 30696 24868 30730
rect 24936 30696 24952 30730
rect 24852 30658 24952 30696
rect 25010 30730 25110 30746
rect 25010 30696 25026 30730
rect 25094 30696 25110 30730
rect 25010 30658 25110 30696
rect 20428 24620 20528 24658
rect 20428 24586 20444 24620
rect 20512 24586 20528 24620
rect 20428 24570 20528 24586
rect 20586 24620 20686 24658
rect 20586 24586 20602 24620
rect 20670 24586 20686 24620
rect 20586 24570 20686 24586
rect 20744 24620 20844 24658
rect 20744 24586 20760 24620
rect 20828 24586 20844 24620
rect 20744 24570 20844 24586
rect 20902 24620 21002 24658
rect 20902 24586 20918 24620
rect 20986 24586 21002 24620
rect 20902 24570 21002 24586
rect 21060 24620 21160 24658
rect 21060 24586 21076 24620
rect 21144 24586 21160 24620
rect 21060 24570 21160 24586
rect 21218 24620 21318 24658
rect 21218 24586 21234 24620
rect 21302 24586 21318 24620
rect 21218 24570 21318 24586
rect 21376 24620 21476 24658
rect 21376 24586 21392 24620
rect 21460 24586 21476 24620
rect 21376 24570 21476 24586
rect 21534 24620 21634 24658
rect 21534 24586 21550 24620
rect 21618 24586 21634 24620
rect 21534 24570 21634 24586
rect 21692 24620 21792 24658
rect 21692 24586 21708 24620
rect 21776 24586 21792 24620
rect 21692 24570 21792 24586
rect 21850 24620 21950 24658
rect 21850 24586 21866 24620
rect 21934 24586 21950 24620
rect 21850 24570 21950 24586
rect 22008 24620 22108 24658
rect 22008 24586 22024 24620
rect 22092 24586 22108 24620
rect 22008 24570 22108 24586
rect 22166 24620 22266 24658
rect 22166 24586 22182 24620
rect 22250 24586 22266 24620
rect 22166 24570 22266 24586
rect 22324 24620 22424 24658
rect 22324 24586 22340 24620
rect 22408 24586 22424 24620
rect 22324 24570 22424 24586
rect 22482 24620 22582 24658
rect 22482 24586 22498 24620
rect 22566 24586 22582 24620
rect 22482 24570 22582 24586
rect 22640 24620 22740 24658
rect 22640 24586 22656 24620
rect 22724 24586 22740 24620
rect 22640 24570 22740 24586
rect 22798 24620 22898 24658
rect 22798 24586 22814 24620
rect 22882 24586 22898 24620
rect 22798 24570 22898 24586
rect 22956 24620 23056 24658
rect 22956 24586 22972 24620
rect 23040 24586 23056 24620
rect 22956 24570 23056 24586
rect 23114 24620 23214 24658
rect 23114 24586 23130 24620
rect 23198 24586 23214 24620
rect 23114 24570 23214 24586
rect 23272 24620 23372 24658
rect 23272 24586 23288 24620
rect 23356 24586 23372 24620
rect 23272 24570 23372 24586
rect 23430 24620 23530 24658
rect 23430 24586 23446 24620
rect 23514 24586 23530 24620
rect 23430 24570 23530 24586
rect 23588 24620 23688 24658
rect 23588 24586 23604 24620
rect 23672 24586 23688 24620
rect 23588 24570 23688 24586
rect 23746 24620 23846 24658
rect 23746 24586 23762 24620
rect 23830 24586 23846 24620
rect 23746 24570 23846 24586
rect 23904 24620 24004 24658
rect 23904 24586 23920 24620
rect 23988 24586 24004 24620
rect 23904 24570 24004 24586
rect 24062 24620 24162 24658
rect 24062 24586 24078 24620
rect 24146 24586 24162 24620
rect 24062 24570 24162 24586
rect 24220 24620 24320 24658
rect 24220 24586 24236 24620
rect 24304 24586 24320 24620
rect 24220 24570 24320 24586
rect 24378 24620 24478 24658
rect 24378 24586 24394 24620
rect 24462 24586 24478 24620
rect 24378 24570 24478 24586
rect 24536 24620 24636 24658
rect 24536 24586 24552 24620
rect 24620 24586 24636 24620
rect 24536 24570 24636 24586
rect 24694 24620 24794 24658
rect 24694 24586 24710 24620
rect 24778 24586 24794 24620
rect 24694 24570 24794 24586
rect 24852 24620 24952 24658
rect 24852 24586 24868 24620
rect 24936 24586 24952 24620
rect 24852 24570 24952 24586
rect 25010 24620 25110 24658
rect 25010 24586 25026 24620
rect 25094 24586 25110 24620
rect 25010 24570 25110 24586
rect 30968 27076 31034 27092
rect 30968 27042 30984 27076
rect 31018 27042 31034 27076
rect 30968 27019 31034 27042
rect 30968 25696 31034 25719
rect 30968 25662 30984 25696
rect 31018 25662 31034 25696
rect 30968 25646 31034 25662
rect 1528 23730 1628 23746
rect 1528 23696 1544 23730
rect 1612 23696 1628 23730
rect 1528 23658 1628 23696
rect 1686 23730 1786 23746
rect 1686 23696 1702 23730
rect 1770 23696 1786 23730
rect 1686 23658 1786 23696
rect 1844 23730 1944 23746
rect 1844 23696 1860 23730
rect 1928 23696 1944 23730
rect 1844 23658 1944 23696
rect 2002 23730 2102 23746
rect 2002 23696 2018 23730
rect 2086 23696 2102 23730
rect 2002 23658 2102 23696
rect 2160 23730 2260 23746
rect 2160 23696 2176 23730
rect 2244 23696 2260 23730
rect 2160 23658 2260 23696
rect 2318 23730 2418 23746
rect 2318 23696 2334 23730
rect 2402 23696 2418 23730
rect 2318 23658 2418 23696
rect 2476 23730 2576 23746
rect 2476 23696 2492 23730
rect 2560 23696 2576 23730
rect 2476 23658 2576 23696
rect 2634 23730 2734 23746
rect 2634 23696 2650 23730
rect 2718 23696 2734 23730
rect 2634 23658 2734 23696
rect 2792 23730 2892 23746
rect 2792 23696 2808 23730
rect 2876 23696 2892 23730
rect 2792 23658 2892 23696
rect 2950 23730 3050 23746
rect 2950 23696 2966 23730
rect 3034 23696 3050 23730
rect 2950 23658 3050 23696
rect 3108 23730 3208 23746
rect 3108 23696 3124 23730
rect 3192 23696 3208 23730
rect 3108 23658 3208 23696
rect 3266 23730 3366 23746
rect 3266 23696 3282 23730
rect 3350 23696 3366 23730
rect 3266 23658 3366 23696
rect 3424 23730 3524 23746
rect 3424 23696 3440 23730
rect 3508 23696 3524 23730
rect 3424 23658 3524 23696
rect 3582 23730 3682 23746
rect 3582 23696 3598 23730
rect 3666 23696 3682 23730
rect 3582 23658 3682 23696
rect 3740 23730 3840 23746
rect 3740 23696 3756 23730
rect 3824 23696 3840 23730
rect 3740 23658 3840 23696
rect 3898 23730 3998 23746
rect 3898 23696 3914 23730
rect 3982 23696 3998 23730
rect 3898 23658 3998 23696
rect 4056 23730 4156 23746
rect 4056 23696 4072 23730
rect 4140 23696 4156 23730
rect 4056 23658 4156 23696
rect 4214 23730 4314 23746
rect 4214 23696 4230 23730
rect 4298 23696 4314 23730
rect 4214 23658 4314 23696
rect 4372 23730 4472 23746
rect 4372 23696 4388 23730
rect 4456 23696 4472 23730
rect 4372 23658 4472 23696
rect 4530 23730 4630 23746
rect 4530 23696 4546 23730
rect 4614 23696 4630 23730
rect 4530 23658 4630 23696
rect 4688 23730 4788 23746
rect 4688 23696 4704 23730
rect 4772 23696 4788 23730
rect 4688 23658 4788 23696
rect 4846 23730 4946 23746
rect 4846 23696 4862 23730
rect 4930 23696 4946 23730
rect 4846 23658 4946 23696
rect 5004 23730 5104 23746
rect 5004 23696 5020 23730
rect 5088 23696 5104 23730
rect 5004 23658 5104 23696
rect 5162 23730 5262 23746
rect 5162 23696 5178 23730
rect 5246 23696 5262 23730
rect 5162 23658 5262 23696
rect 5320 23730 5420 23746
rect 5320 23696 5336 23730
rect 5404 23696 5420 23730
rect 5320 23658 5420 23696
rect 5478 23730 5578 23746
rect 5478 23696 5494 23730
rect 5562 23696 5578 23730
rect 5478 23658 5578 23696
rect 5636 23730 5736 23746
rect 5636 23696 5652 23730
rect 5720 23696 5736 23730
rect 5636 23658 5736 23696
rect 5794 23730 5894 23746
rect 5794 23696 5810 23730
rect 5878 23696 5894 23730
rect 5794 23658 5894 23696
rect 5952 23730 6052 23746
rect 5952 23696 5968 23730
rect 6036 23696 6052 23730
rect 5952 23658 6052 23696
rect 6110 23730 6210 23746
rect 6110 23696 6126 23730
rect 6194 23696 6210 23730
rect 6110 23658 6210 23696
rect 1528 17620 1628 17658
rect 1528 17586 1544 17620
rect 1612 17586 1628 17620
rect 1528 17570 1628 17586
rect 1686 17620 1786 17658
rect 1686 17586 1702 17620
rect 1770 17586 1786 17620
rect 1686 17570 1786 17586
rect 1844 17620 1944 17658
rect 1844 17586 1860 17620
rect 1928 17586 1944 17620
rect 1844 17570 1944 17586
rect 2002 17620 2102 17658
rect 2002 17586 2018 17620
rect 2086 17586 2102 17620
rect 2002 17570 2102 17586
rect 2160 17620 2260 17658
rect 2160 17586 2176 17620
rect 2244 17586 2260 17620
rect 2160 17570 2260 17586
rect 2318 17620 2418 17658
rect 2318 17586 2334 17620
rect 2402 17586 2418 17620
rect 2318 17570 2418 17586
rect 2476 17620 2576 17658
rect 2476 17586 2492 17620
rect 2560 17586 2576 17620
rect 2476 17570 2576 17586
rect 2634 17620 2734 17658
rect 2634 17586 2650 17620
rect 2718 17586 2734 17620
rect 2634 17570 2734 17586
rect 2792 17620 2892 17658
rect 2792 17586 2808 17620
rect 2876 17586 2892 17620
rect 2792 17570 2892 17586
rect 2950 17620 3050 17658
rect 2950 17586 2966 17620
rect 3034 17586 3050 17620
rect 2950 17570 3050 17586
rect 3108 17620 3208 17658
rect 3108 17586 3124 17620
rect 3192 17586 3208 17620
rect 3108 17570 3208 17586
rect 3266 17620 3366 17658
rect 3266 17586 3282 17620
rect 3350 17586 3366 17620
rect 3266 17570 3366 17586
rect 3424 17620 3524 17658
rect 3424 17586 3440 17620
rect 3508 17586 3524 17620
rect 3424 17570 3524 17586
rect 3582 17620 3682 17658
rect 3582 17586 3598 17620
rect 3666 17586 3682 17620
rect 3582 17570 3682 17586
rect 3740 17620 3840 17658
rect 3740 17586 3756 17620
rect 3824 17586 3840 17620
rect 3740 17570 3840 17586
rect 3898 17620 3998 17658
rect 3898 17586 3914 17620
rect 3982 17586 3998 17620
rect 3898 17570 3998 17586
rect 4056 17620 4156 17658
rect 4056 17586 4072 17620
rect 4140 17586 4156 17620
rect 4056 17570 4156 17586
rect 4214 17620 4314 17658
rect 4214 17586 4230 17620
rect 4298 17586 4314 17620
rect 4214 17570 4314 17586
rect 4372 17620 4472 17658
rect 4372 17586 4388 17620
rect 4456 17586 4472 17620
rect 4372 17570 4472 17586
rect 4530 17620 4630 17658
rect 4530 17586 4546 17620
rect 4614 17586 4630 17620
rect 4530 17570 4630 17586
rect 4688 17620 4788 17658
rect 4688 17586 4704 17620
rect 4772 17586 4788 17620
rect 4688 17570 4788 17586
rect 4846 17620 4946 17658
rect 4846 17586 4862 17620
rect 4930 17586 4946 17620
rect 4846 17570 4946 17586
rect 5004 17620 5104 17658
rect 5004 17586 5020 17620
rect 5088 17586 5104 17620
rect 5004 17570 5104 17586
rect 5162 17620 5262 17658
rect 5162 17586 5178 17620
rect 5246 17586 5262 17620
rect 5162 17570 5262 17586
rect 5320 17620 5420 17658
rect 5320 17586 5336 17620
rect 5404 17586 5420 17620
rect 5320 17570 5420 17586
rect 5478 17620 5578 17658
rect 5478 17586 5494 17620
rect 5562 17586 5578 17620
rect 5478 17570 5578 17586
rect 5636 17620 5736 17658
rect 5636 17586 5652 17620
rect 5720 17586 5736 17620
rect 5636 17570 5736 17586
rect 5794 17620 5894 17658
rect 5794 17586 5810 17620
rect 5878 17586 5894 17620
rect 5794 17570 5894 17586
rect 5952 17620 6052 17658
rect 5952 17586 5968 17620
rect 6036 17586 6052 17620
rect 5952 17570 6052 17586
rect 6110 17620 6210 17658
rect 6110 17586 6126 17620
rect 6194 17586 6210 17620
rect 6110 17570 6210 17586
rect 7828 23730 7928 23746
rect 7828 23696 7844 23730
rect 7912 23696 7928 23730
rect 7828 23658 7928 23696
rect 7986 23730 8086 23746
rect 7986 23696 8002 23730
rect 8070 23696 8086 23730
rect 7986 23658 8086 23696
rect 8144 23730 8244 23746
rect 8144 23696 8160 23730
rect 8228 23696 8244 23730
rect 8144 23658 8244 23696
rect 8302 23730 8402 23746
rect 8302 23696 8318 23730
rect 8386 23696 8402 23730
rect 8302 23658 8402 23696
rect 8460 23730 8560 23746
rect 8460 23696 8476 23730
rect 8544 23696 8560 23730
rect 8460 23658 8560 23696
rect 8618 23730 8718 23746
rect 8618 23696 8634 23730
rect 8702 23696 8718 23730
rect 8618 23658 8718 23696
rect 8776 23730 8876 23746
rect 8776 23696 8792 23730
rect 8860 23696 8876 23730
rect 8776 23658 8876 23696
rect 8934 23730 9034 23746
rect 8934 23696 8950 23730
rect 9018 23696 9034 23730
rect 8934 23658 9034 23696
rect 9092 23730 9192 23746
rect 9092 23696 9108 23730
rect 9176 23696 9192 23730
rect 9092 23658 9192 23696
rect 9250 23730 9350 23746
rect 9250 23696 9266 23730
rect 9334 23696 9350 23730
rect 9250 23658 9350 23696
rect 9408 23730 9508 23746
rect 9408 23696 9424 23730
rect 9492 23696 9508 23730
rect 9408 23658 9508 23696
rect 9566 23730 9666 23746
rect 9566 23696 9582 23730
rect 9650 23696 9666 23730
rect 9566 23658 9666 23696
rect 9724 23730 9824 23746
rect 9724 23696 9740 23730
rect 9808 23696 9824 23730
rect 9724 23658 9824 23696
rect 9882 23730 9982 23746
rect 9882 23696 9898 23730
rect 9966 23696 9982 23730
rect 9882 23658 9982 23696
rect 10040 23730 10140 23746
rect 10040 23696 10056 23730
rect 10124 23696 10140 23730
rect 10040 23658 10140 23696
rect 10198 23730 10298 23746
rect 10198 23696 10214 23730
rect 10282 23696 10298 23730
rect 10198 23658 10298 23696
rect 10356 23730 10456 23746
rect 10356 23696 10372 23730
rect 10440 23696 10456 23730
rect 10356 23658 10456 23696
rect 10514 23730 10614 23746
rect 10514 23696 10530 23730
rect 10598 23696 10614 23730
rect 10514 23658 10614 23696
rect 10672 23730 10772 23746
rect 10672 23696 10688 23730
rect 10756 23696 10772 23730
rect 10672 23658 10772 23696
rect 10830 23730 10930 23746
rect 10830 23696 10846 23730
rect 10914 23696 10930 23730
rect 10830 23658 10930 23696
rect 10988 23730 11088 23746
rect 10988 23696 11004 23730
rect 11072 23696 11088 23730
rect 10988 23658 11088 23696
rect 11146 23730 11246 23746
rect 11146 23696 11162 23730
rect 11230 23696 11246 23730
rect 11146 23658 11246 23696
rect 11304 23730 11404 23746
rect 11304 23696 11320 23730
rect 11388 23696 11404 23730
rect 11304 23658 11404 23696
rect 11462 23730 11562 23746
rect 11462 23696 11478 23730
rect 11546 23696 11562 23730
rect 11462 23658 11562 23696
rect 11620 23730 11720 23746
rect 11620 23696 11636 23730
rect 11704 23696 11720 23730
rect 11620 23658 11720 23696
rect 11778 23730 11878 23746
rect 11778 23696 11794 23730
rect 11862 23696 11878 23730
rect 11778 23658 11878 23696
rect 11936 23730 12036 23746
rect 11936 23696 11952 23730
rect 12020 23696 12036 23730
rect 11936 23658 12036 23696
rect 12094 23730 12194 23746
rect 12094 23696 12110 23730
rect 12178 23696 12194 23730
rect 12094 23658 12194 23696
rect 12252 23730 12352 23746
rect 12252 23696 12268 23730
rect 12336 23696 12352 23730
rect 12252 23658 12352 23696
rect 12410 23730 12510 23746
rect 12410 23696 12426 23730
rect 12494 23696 12510 23730
rect 12410 23658 12510 23696
rect 7828 17620 7928 17658
rect 7828 17586 7844 17620
rect 7912 17586 7928 17620
rect 7828 17570 7928 17586
rect 7986 17620 8086 17658
rect 7986 17586 8002 17620
rect 8070 17586 8086 17620
rect 7986 17570 8086 17586
rect 8144 17620 8244 17658
rect 8144 17586 8160 17620
rect 8228 17586 8244 17620
rect 8144 17570 8244 17586
rect 8302 17620 8402 17658
rect 8302 17586 8318 17620
rect 8386 17586 8402 17620
rect 8302 17570 8402 17586
rect 8460 17620 8560 17658
rect 8460 17586 8476 17620
rect 8544 17586 8560 17620
rect 8460 17570 8560 17586
rect 8618 17620 8718 17658
rect 8618 17586 8634 17620
rect 8702 17586 8718 17620
rect 8618 17570 8718 17586
rect 8776 17620 8876 17658
rect 8776 17586 8792 17620
rect 8860 17586 8876 17620
rect 8776 17570 8876 17586
rect 8934 17620 9034 17658
rect 8934 17586 8950 17620
rect 9018 17586 9034 17620
rect 8934 17570 9034 17586
rect 9092 17620 9192 17658
rect 9092 17586 9108 17620
rect 9176 17586 9192 17620
rect 9092 17570 9192 17586
rect 9250 17620 9350 17658
rect 9250 17586 9266 17620
rect 9334 17586 9350 17620
rect 9250 17570 9350 17586
rect 9408 17620 9508 17658
rect 9408 17586 9424 17620
rect 9492 17586 9508 17620
rect 9408 17570 9508 17586
rect 9566 17620 9666 17658
rect 9566 17586 9582 17620
rect 9650 17586 9666 17620
rect 9566 17570 9666 17586
rect 9724 17620 9824 17658
rect 9724 17586 9740 17620
rect 9808 17586 9824 17620
rect 9724 17570 9824 17586
rect 9882 17620 9982 17658
rect 9882 17586 9898 17620
rect 9966 17586 9982 17620
rect 9882 17570 9982 17586
rect 10040 17620 10140 17658
rect 10040 17586 10056 17620
rect 10124 17586 10140 17620
rect 10040 17570 10140 17586
rect 10198 17620 10298 17658
rect 10198 17586 10214 17620
rect 10282 17586 10298 17620
rect 10198 17570 10298 17586
rect 10356 17620 10456 17658
rect 10356 17586 10372 17620
rect 10440 17586 10456 17620
rect 10356 17570 10456 17586
rect 10514 17620 10614 17658
rect 10514 17586 10530 17620
rect 10598 17586 10614 17620
rect 10514 17570 10614 17586
rect 10672 17620 10772 17658
rect 10672 17586 10688 17620
rect 10756 17586 10772 17620
rect 10672 17570 10772 17586
rect 10830 17620 10930 17658
rect 10830 17586 10846 17620
rect 10914 17586 10930 17620
rect 10830 17570 10930 17586
rect 10988 17620 11088 17658
rect 10988 17586 11004 17620
rect 11072 17586 11088 17620
rect 10988 17570 11088 17586
rect 11146 17620 11246 17658
rect 11146 17586 11162 17620
rect 11230 17586 11246 17620
rect 11146 17570 11246 17586
rect 11304 17620 11404 17658
rect 11304 17586 11320 17620
rect 11388 17586 11404 17620
rect 11304 17570 11404 17586
rect 11462 17620 11562 17658
rect 11462 17586 11478 17620
rect 11546 17586 11562 17620
rect 11462 17570 11562 17586
rect 11620 17620 11720 17658
rect 11620 17586 11636 17620
rect 11704 17586 11720 17620
rect 11620 17570 11720 17586
rect 11778 17620 11878 17658
rect 11778 17586 11794 17620
rect 11862 17586 11878 17620
rect 11778 17570 11878 17586
rect 11936 17620 12036 17658
rect 11936 17586 11952 17620
rect 12020 17586 12036 17620
rect 11936 17570 12036 17586
rect 12094 17620 12194 17658
rect 12094 17586 12110 17620
rect 12178 17586 12194 17620
rect 12094 17570 12194 17586
rect 12252 17620 12352 17658
rect 12252 17586 12268 17620
rect 12336 17586 12352 17620
rect 12252 17570 12352 17586
rect 12410 17620 12510 17658
rect 12410 17586 12426 17620
rect 12494 17586 12510 17620
rect 12410 17570 12510 17586
rect 14128 23730 14228 23746
rect 14128 23696 14144 23730
rect 14212 23696 14228 23730
rect 14128 23658 14228 23696
rect 14286 23730 14386 23746
rect 14286 23696 14302 23730
rect 14370 23696 14386 23730
rect 14286 23658 14386 23696
rect 14444 23730 14544 23746
rect 14444 23696 14460 23730
rect 14528 23696 14544 23730
rect 14444 23658 14544 23696
rect 14602 23730 14702 23746
rect 14602 23696 14618 23730
rect 14686 23696 14702 23730
rect 14602 23658 14702 23696
rect 14760 23730 14860 23746
rect 14760 23696 14776 23730
rect 14844 23696 14860 23730
rect 14760 23658 14860 23696
rect 14918 23730 15018 23746
rect 14918 23696 14934 23730
rect 15002 23696 15018 23730
rect 14918 23658 15018 23696
rect 15076 23730 15176 23746
rect 15076 23696 15092 23730
rect 15160 23696 15176 23730
rect 15076 23658 15176 23696
rect 15234 23730 15334 23746
rect 15234 23696 15250 23730
rect 15318 23696 15334 23730
rect 15234 23658 15334 23696
rect 15392 23730 15492 23746
rect 15392 23696 15408 23730
rect 15476 23696 15492 23730
rect 15392 23658 15492 23696
rect 15550 23730 15650 23746
rect 15550 23696 15566 23730
rect 15634 23696 15650 23730
rect 15550 23658 15650 23696
rect 15708 23730 15808 23746
rect 15708 23696 15724 23730
rect 15792 23696 15808 23730
rect 15708 23658 15808 23696
rect 15866 23730 15966 23746
rect 15866 23696 15882 23730
rect 15950 23696 15966 23730
rect 15866 23658 15966 23696
rect 16024 23730 16124 23746
rect 16024 23696 16040 23730
rect 16108 23696 16124 23730
rect 16024 23658 16124 23696
rect 16182 23730 16282 23746
rect 16182 23696 16198 23730
rect 16266 23696 16282 23730
rect 16182 23658 16282 23696
rect 16340 23730 16440 23746
rect 16340 23696 16356 23730
rect 16424 23696 16440 23730
rect 16340 23658 16440 23696
rect 16498 23730 16598 23746
rect 16498 23696 16514 23730
rect 16582 23696 16598 23730
rect 16498 23658 16598 23696
rect 16656 23730 16756 23746
rect 16656 23696 16672 23730
rect 16740 23696 16756 23730
rect 16656 23658 16756 23696
rect 16814 23730 16914 23746
rect 16814 23696 16830 23730
rect 16898 23696 16914 23730
rect 16814 23658 16914 23696
rect 16972 23730 17072 23746
rect 16972 23696 16988 23730
rect 17056 23696 17072 23730
rect 16972 23658 17072 23696
rect 17130 23730 17230 23746
rect 17130 23696 17146 23730
rect 17214 23696 17230 23730
rect 17130 23658 17230 23696
rect 17288 23730 17388 23746
rect 17288 23696 17304 23730
rect 17372 23696 17388 23730
rect 17288 23658 17388 23696
rect 17446 23730 17546 23746
rect 17446 23696 17462 23730
rect 17530 23696 17546 23730
rect 17446 23658 17546 23696
rect 17604 23730 17704 23746
rect 17604 23696 17620 23730
rect 17688 23696 17704 23730
rect 17604 23658 17704 23696
rect 17762 23730 17862 23746
rect 17762 23696 17778 23730
rect 17846 23696 17862 23730
rect 17762 23658 17862 23696
rect 17920 23730 18020 23746
rect 17920 23696 17936 23730
rect 18004 23696 18020 23730
rect 17920 23658 18020 23696
rect 18078 23730 18178 23746
rect 18078 23696 18094 23730
rect 18162 23696 18178 23730
rect 18078 23658 18178 23696
rect 18236 23730 18336 23746
rect 18236 23696 18252 23730
rect 18320 23696 18336 23730
rect 18236 23658 18336 23696
rect 18394 23730 18494 23746
rect 18394 23696 18410 23730
rect 18478 23696 18494 23730
rect 18394 23658 18494 23696
rect 18552 23730 18652 23746
rect 18552 23696 18568 23730
rect 18636 23696 18652 23730
rect 18552 23658 18652 23696
rect 18710 23730 18810 23746
rect 18710 23696 18726 23730
rect 18794 23696 18810 23730
rect 18710 23658 18810 23696
rect 14128 17620 14228 17658
rect 14128 17586 14144 17620
rect 14212 17586 14228 17620
rect 14128 17570 14228 17586
rect 14286 17620 14386 17658
rect 14286 17586 14302 17620
rect 14370 17586 14386 17620
rect 14286 17570 14386 17586
rect 14444 17620 14544 17658
rect 14444 17586 14460 17620
rect 14528 17586 14544 17620
rect 14444 17570 14544 17586
rect 14602 17620 14702 17658
rect 14602 17586 14618 17620
rect 14686 17586 14702 17620
rect 14602 17570 14702 17586
rect 14760 17620 14860 17658
rect 14760 17586 14776 17620
rect 14844 17586 14860 17620
rect 14760 17570 14860 17586
rect 14918 17620 15018 17658
rect 14918 17586 14934 17620
rect 15002 17586 15018 17620
rect 14918 17570 15018 17586
rect 15076 17620 15176 17658
rect 15076 17586 15092 17620
rect 15160 17586 15176 17620
rect 15076 17570 15176 17586
rect 15234 17620 15334 17658
rect 15234 17586 15250 17620
rect 15318 17586 15334 17620
rect 15234 17570 15334 17586
rect 15392 17620 15492 17658
rect 15392 17586 15408 17620
rect 15476 17586 15492 17620
rect 15392 17570 15492 17586
rect 15550 17620 15650 17658
rect 15550 17586 15566 17620
rect 15634 17586 15650 17620
rect 15550 17570 15650 17586
rect 15708 17620 15808 17658
rect 15708 17586 15724 17620
rect 15792 17586 15808 17620
rect 15708 17570 15808 17586
rect 15866 17620 15966 17658
rect 15866 17586 15882 17620
rect 15950 17586 15966 17620
rect 15866 17570 15966 17586
rect 16024 17620 16124 17658
rect 16024 17586 16040 17620
rect 16108 17586 16124 17620
rect 16024 17570 16124 17586
rect 16182 17620 16282 17658
rect 16182 17586 16198 17620
rect 16266 17586 16282 17620
rect 16182 17570 16282 17586
rect 16340 17620 16440 17658
rect 16340 17586 16356 17620
rect 16424 17586 16440 17620
rect 16340 17570 16440 17586
rect 16498 17620 16598 17658
rect 16498 17586 16514 17620
rect 16582 17586 16598 17620
rect 16498 17570 16598 17586
rect 16656 17620 16756 17658
rect 16656 17586 16672 17620
rect 16740 17586 16756 17620
rect 16656 17570 16756 17586
rect 16814 17620 16914 17658
rect 16814 17586 16830 17620
rect 16898 17586 16914 17620
rect 16814 17570 16914 17586
rect 16972 17620 17072 17658
rect 16972 17586 16988 17620
rect 17056 17586 17072 17620
rect 16972 17570 17072 17586
rect 17130 17620 17230 17658
rect 17130 17586 17146 17620
rect 17214 17586 17230 17620
rect 17130 17570 17230 17586
rect 17288 17620 17388 17658
rect 17288 17586 17304 17620
rect 17372 17586 17388 17620
rect 17288 17570 17388 17586
rect 17446 17620 17546 17658
rect 17446 17586 17462 17620
rect 17530 17586 17546 17620
rect 17446 17570 17546 17586
rect 17604 17620 17704 17658
rect 17604 17586 17620 17620
rect 17688 17586 17704 17620
rect 17604 17570 17704 17586
rect 17762 17620 17862 17658
rect 17762 17586 17778 17620
rect 17846 17586 17862 17620
rect 17762 17570 17862 17586
rect 17920 17620 18020 17658
rect 17920 17586 17936 17620
rect 18004 17586 18020 17620
rect 17920 17570 18020 17586
rect 18078 17620 18178 17658
rect 18078 17586 18094 17620
rect 18162 17586 18178 17620
rect 18078 17570 18178 17586
rect 18236 17620 18336 17658
rect 18236 17586 18252 17620
rect 18320 17586 18336 17620
rect 18236 17570 18336 17586
rect 18394 17620 18494 17658
rect 18394 17586 18410 17620
rect 18478 17586 18494 17620
rect 18394 17570 18494 17586
rect 18552 17620 18652 17658
rect 18552 17586 18568 17620
rect 18636 17586 18652 17620
rect 18552 17570 18652 17586
rect 18710 17620 18810 17658
rect 18710 17586 18726 17620
rect 18794 17586 18810 17620
rect 18710 17570 18810 17586
rect 20428 23730 20528 23746
rect 20428 23696 20444 23730
rect 20512 23696 20528 23730
rect 20428 23658 20528 23696
rect 20586 23730 20686 23746
rect 20586 23696 20602 23730
rect 20670 23696 20686 23730
rect 20586 23658 20686 23696
rect 20744 23730 20844 23746
rect 20744 23696 20760 23730
rect 20828 23696 20844 23730
rect 20744 23658 20844 23696
rect 20902 23730 21002 23746
rect 20902 23696 20918 23730
rect 20986 23696 21002 23730
rect 20902 23658 21002 23696
rect 21060 23730 21160 23746
rect 21060 23696 21076 23730
rect 21144 23696 21160 23730
rect 21060 23658 21160 23696
rect 21218 23730 21318 23746
rect 21218 23696 21234 23730
rect 21302 23696 21318 23730
rect 21218 23658 21318 23696
rect 21376 23730 21476 23746
rect 21376 23696 21392 23730
rect 21460 23696 21476 23730
rect 21376 23658 21476 23696
rect 21534 23730 21634 23746
rect 21534 23696 21550 23730
rect 21618 23696 21634 23730
rect 21534 23658 21634 23696
rect 21692 23730 21792 23746
rect 21692 23696 21708 23730
rect 21776 23696 21792 23730
rect 21692 23658 21792 23696
rect 21850 23730 21950 23746
rect 21850 23696 21866 23730
rect 21934 23696 21950 23730
rect 21850 23658 21950 23696
rect 22008 23730 22108 23746
rect 22008 23696 22024 23730
rect 22092 23696 22108 23730
rect 22008 23658 22108 23696
rect 22166 23730 22266 23746
rect 22166 23696 22182 23730
rect 22250 23696 22266 23730
rect 22166 23658 22266 23696
rect 22324 23730 22424 23746
rect 22324 23696 22340 23730
rect 22408 23696 22424 23730
rect 22324 23658 22424 23696
rect 22482 23730 22582 23746
rect 22482 23696 22498 23730
rect 22566 23696 22582 23730
rect 22482 23658 22582 23696
rect 22640 23730 22740 23746
rect 22640 23696 22656 23730
rect 22724 23696 22740 23730
rect 22640 23658 22740 23696
rect 22798 23730 22898 23746
rect 22798 23696 22814 23730
rect 22882 23696 22898 23730
rect 22798 23658 22898 23696
rect 22956 23730 23056 23746
rect 22956 23696 22972 23730
rect 23040 23696 23056 23730
rect 22956 23658 23056 23696
rect 23114 23730 23214 23746
rect 23114 23696 23130 23730
rect 23198 23696 23214 23730
rect 23114 23658 23214 23696
rect 23272 23730 23372 23746
rect 23272 23696 23288 23730
rect 23356 23696 23372 23730
rect 23272 23658 23372 23696
rect 23430 23730 23530 23746
rect 23430 23696 23446 23730
rect 23514 23696 23530 23730
rect 23430 23658 23530 23696
rect 23588 23730 23688 23746
rect 23588 23696 23604 23730
rect 23672 23696 23688 23730
rect 23588 23658 23688 23696
rect 23746 23730 23846 23746
rect 23746 23696 23762 23730
rect 23830 23696 23846 23730
rect 23746 23658 23846 23696
rect 23904 23730 24004 23746
rect 23904 23696 23920 23730
rect 23988 23696 24004 23730
rect 23904 23658 24004 23696
rect 24062 23730 24162 23746
rect 24062 23696 24078 23730
rect 24146 23696 24162 23730
rect 24062 23658 24162 23696
rect 24220 23730 24320 23746
rect 24220 23696 24236 23730
rect 24304 23696 24320 23730
rect 24220 23658 24320 23696
rect 24378 23730 24478 23746
rect 24378 23696 24394 23730
rect 24462 23696 24478 23730
rect 24378 23658 24478 23696
rect 24536 23730 24636 23746
rect 24536 23696 24552 23730
rect 24620 23696 24636 23730
rect 24536 23658 24636 23696
rect 24694 23730 24794 23746
rect 24694 23696 24710 23730
rect 24778 23696 24794 23730
rect 24694 23658 24794 23696
rect 24852 23730 24952 23746
rect 24852 23696 24868 23730
rect 24936 23696 24952 23730
rect 24852 23658 24952 23696
rect 25010 23730 25110 23746
rect 25010 23696 25026 23730
rect 25094 23696 25110 23730
rect 25010 23658 25110 23696
rect 20428 17620 20528 17658
rect 20428 17586 20444 17620
rect 20512 17586 20528 17620
rect 20428 17570 20528 17586
rect 20586 17620 20686 17658
rect 20586 17586 20602 17620
rect 20670 17586 20686 17620
rect 20586 17570 20686 17586
rect 20744 17620 20844 17658
rect 20744 17586 20760 17620
rect 20828 17586 20844 17620
rect 20744 17570 20844 17586
rect 20902 17620 21002 17658
rect 20902 17586 20918 17620
rect 20986 17586 21002 17620
rect 20902 17570 21002 17586
rect 21060 17620 21160 17658
rect 21060 17586 21076 17620
rect 21144 17586 21160 17620
rect 21060 17570 21160 17586
rect 21218 17620 21318 17658
rect 21218 17586 21234 17620
rect 21302 17586 21318 17620
rect 21218 17570 21318 17586
rect 21376 17620 21476 17658
rect 21376 17586 21392 17620
rect 21460 17586 21476 17620
rect 21376 17570 21476 17586
rect 21534 17620 21634 17658
rect 21534 17586 21550 17620
rect 21618 17586 21634 17620
rect 21534 17570 21634 17586
rect 21692 17620 21792 17658
rect 21692 17586 21708 17620
rect 21776 17586 21792 17620
rect 21692 17570 21792 17586
rect 21850 17620 21950 17658
rect 21850 17586 21866 17620
rect 21934 17586 21950 17620
rect 21850 17570 21950 17586
rect 22008 17620 22108 17658
rect 22008 17586 22024 17620
rect 22092 17586 22108 17620
rect 22008 17570 22108 17586
rect 22166 17620 22266 17658
rect 22166 17586 22182 17620
rect 22250 17586 22266 17620
rect 22166 17570 22266 17586
rect 22324 17620 22424 17658
rect 22324 17586 22340 17620
rect 22408 17586 22424 17620
rect 22324 17570 22424 17586
rect 22482 17620 22582 17658
rect 22482 17586 22498 17620
rect 22566 17586 22582 17620
rect 22482 17570 22582 17586
rect 22640 17620 22740 17658
rect 22640 17586 22656 17620
rect 22724 17586 22740 17620
rect 22640 17570 22740 17586
rect 22798 17620 22898 17658
rect 22798 17586 22814 17620
rect 22882 17586 22898 17620
rect 22798 17570 22898 17586
rect 22956 17620 23056 17658
rect 22956 17586 22972 17620
rect 23040 17586 23056 17620
rect 22956 17570 23056 17586
rect 23114 17620 23214 17658
rect 23114 17586 23130 17620
rect 23198 17586 23214 17620
rect 23114 17570 23214 17586
rect 23272 17620 23372 17658
rect 23272 17586 23288 17620
rect 23356 17586 23372 17620
rect 23272 17570 23372 17586
rect 23430 17620 23530 17658
rect 23430 17586 23446 17620
rect 23514 17586 23530 17620
rect 23430 17570 23530 17586
rect 23588 17620 23688 17658
rect 23588 17586 23604 17620
rect 23672 17586 23688 17620
rect 23588 17570 23688 17586
rect 23746 17620 23846 17658
rect 23746 17586 23762 17620
rect 23830 17586 23846 17620
rect 23746 17570 23846 17586
rect 23904 17620 24004 17658
rect 23904 17586 23920 17620
rect 23988 17586 24004 17620
rect 23904 17570 24004 17586
rect 24062 17620 24162 17658
rect 24062 17586 24078 17620
rect 24146 17586 24162 17620
rect 24062 17570 24162 17586
rect 24220 17620 24320 17658
rect 24220 17586 24236 17620
rect 24304 17586 24320 17620
rect 24220 17570 24320 17586
rect 24378 17620 24478 17658
rect 24378 17586 24394 17620
rect 24462 17586 24478 17620
rect 24378 17570 24478 17586
rect 24536 17620 24636 17658
rect 24536 17586 24552 17620
rect 24620 17586 24636 17620
rect 24536 17570 24636 17586
rect 24694 17620 24794 17658
rect 24694 17586 24710 17620
rect 24778 17586 24794 17620
rect 24694 17570 24794 17586
rect 24852 17620 24952 17658
rect 24852 17586 24868 17620
rect 24936 17586 24952 17620
rect 24852 17570 24952 17586
rect 25010 17620 25110 17658
rect 25010 17586 25026 17620
rect 25094 17586 25110 17620
rect 25010 17570 25110 17586
rect 1528 15430 1628 15446
rect 1528 15396 1544 15430
rect 1612 15396 1628 15430
rect 1528 15358 1628 15396
rect 1686 15430 1786 15446
rect 1686 15396 1702 15430
rect 1770 15396 1786 15430
rect 1686 15358 1786 15396
rect 1844 15430 1944 15446
rect 1844 15396 1860 15430
rect 1928 15396 1944 15430
rect 1844 15358 1944 15396
rect 2002 15430 2102 15446
rect 2002 15396 2018 15430
rect 2086 15396 2102 15430
rect 2002 15358 2102 15396
rect 2160 15430 2260 15446
rect 2160 15396 2176 15430
rect 2244 15396 2260 15430
rect 2160 15358 2260 15396
rect 2318 15430 2418 15446
rect 2318 15396 2334 15430
rect 2402 15396 2418 15430
rect 2318 15358 2418 15396
rect 2476 15430 2576 15446
rect 2476 15396 2492 15430
rect 2560 15396 2576 15430
rect 2476 15358 2576 15396
rect 2634 15430 2734 15446
rect 2634 15396 2650 15430
rect 2718 15396 2734 15430
rect 2634 15358 2734 15396
rect 2792 15430 2892 15446
rect 2792 15396 2808 15430
rect 2876 15396 2892 15430
rect 2792 15358 2892 15396
rect 2950 15430 3050 15446
rect 2950 15396 2966 15430
rect 3034 15396 3050 15430
rect 2950 15358 3050 15396
rect 3108 15430 3208 15446
rect 3108 15396 3124 15430
rect 3192 15396 3208 15430
rect 3108 15358 3208 15396
rect 3266 15430 3366 15446
rect 3266 15396 3282 15430
rect 3350 15396 3366 15430
rect 3266 15358 3366 15396
rect 3424 15430 3524 15446
rect 3424 15396 3440 15430
rect 3508 15396 3524 15430
rect 3424 15358 3524 15396
rect 3582 15430 3682 15446
rect 3582 15396 3598 15430
rect 3666 15396 3682 15430
rect 3582 15358 3682 15396
rect 3740 15430 3840 15446
rect 3740 15396 3756 15430
rect 3824 15396 3840 15430
rect 3740 15358 3840 15396
rect 3898 15430 3998 15446
rect 3898 15396 3914 15430
rect 3982 15396 3998 15430
rect 3898 15358 3998 15396
rect 4056 15430 4156 15446
rect 4056 15396 4072 15430
rect 4140 15396 4156 15430
rect 4056 15358 4156 15396
rect 4214 15430 4314 15446
rect 4214 15396 4230 15430
rect 4298 15396 4314 15430
rect 4214 15358 4314 15396
rect 4372 15430 4472 15446
rect 4372 15396 4388 15430
rect 4456 15396 4472 15430
rect 4372 15358 4472 15396
rect 4530 15430 4630 15446
rect 4530 15396 4546 15430
rect 4614 15396 4630 15430
rect 4530 15358 4630 15396
rect 4688 15430 4788 15446
rect 4688 15396 4704 15430
rect 4772 15396 4788 15430
rect 4688 15358 4788 15396
rect 4846 15430 4946 15446
rect 4846 15396 4862 15430
rect 4930 15396 4946 15430
rect 4846 15358 4946 15396
rect 5004 15430 5104 15446
rect 5004 15396 5020 15430
rect 5088 15396 5104 15430
rect 5004 15358 5104 15396
rect 5162 15430 5262 15446
rect 5162 15396 5178 15430
rect 5246 15396 5262 15430
rect 5162 15358 5262 15396
rect 5320 15430 5420 15446
rect 5320 15396 5336 15430
rect 5404 15396 5420 15430
rect 5320 15358 5420 15396
rect 5478 15430 5578 15446
rect 5478 15396 5494 15430
rect 5562 15396 5578 15430
rect 5478 15358 5578 15396
rect 5636 15430 5736 15446
rect 5636 15396 5652 15430
rect 5720 15396 5736 15430
rect 5636 15358 5736 15396
rect 5794 15430 5894 15446
rect 5794 15396 5810 15430
rect 5878 15396 5894 15430
rect 5794 15358 5894 15396
rect 5952 15430 6052 15446
rect 5952 15396 5968 15430
rect 6036 15396 6052 15430
rect 5952 15358 6052 15396
rect 6110 15430 6210 15446
rect 6110 15396 6126 15430
rect 6194 15396 6210 15430
rect 6110 15358 6210 15396
rect 1528 9320 1628 9358
rect 1528 9286 1544 9320
rect 1612 9286 1628 9320
rect 1528 9270 1628 9286
rect 1686 9320 1786 9358
rect 1686 9286 1702 9320
rect 1770 9286 1786 9320
rect 1686 9270 1786 9286
rect 1844 9320 1944 9358
rect 1844 9286 1860 9320
rect 1928 9286 1944 9320
rect 1844 9270 1944 9286
rect 2002 9320 2102 9358
rect 2002 9286 2018 9320
rect 2086 9286 2102 9320
rect 2002 9270 2102 9286
rect 2160 9320 2260 9358
rect 2160 9286 2176 9320
rect 2244 9286 2260 9320
rect 2160 9270 2260 9286
rect 2318 9320 2418 9358
rect 2318 9286 2334 9320
rect 2402 9286 2418 9320
rect 2318 9270 2418 9286
rect 2476 9320 2576 9358
rect 2476 9286 2492 9320
rect 2560 9286 2576 9320
rect 2476 9270 2576 9286
rect 2634 9320 2734 9358
rect 2634 9286 2650 9320
rect 2718 9286 2734 9320
rect 2634 9270 2734 9286
rect 2792 9320 2892 9358
rect 2792 9286 2808 9320
rect 2876 9286 2892 9320
rect 2792 9270 2892 9286
rect 2950 9320 3050 9358
rect 2950 9286 2966 9320
rect 3034 9286 3050 9320
rect 2950 9270 3050 9286
rect 3108 9320 3208 9358
rect 3108 9286 3124 9320
rect 3192 9286 3208 9320
rect 3108 9270 3208 9286
rect 3266 9320 3366 9358
rect 3266 9286 3282 9320
rect 3350 9286 3366 9320
rect 3266 9270 3366 9286
rect 3424 9320 3524 9358
rect 3424 9286 3440 9320
rect 3508 9286 3524 9320
rect 3424 9270 3524 9286
rect 3582 9320 3682 9358
rect 3582 9286 3598 9320
rect 3666 9286 3682 9320
rect 3582 9270 3682 9286
rect 3740 9320 3840 9358
rect 3740 9286 3756 9320
rect 3824 9286 3840 9320
rect 3740 9270 3840 9286
rect 3898 9320 3998 9358
rect 3898 9286 3914 9320
rect 3982 9286 3998 9320
rect 3898 9270 3998 9286
rect 4056 9320 4156 9358
rect 4056 9286 4072 9320
rect 4140 9286 4156 9320
rect 4056 9270 4156 9286
rect 4214 9320 4314 9358
rect 4214 9286 4230 9320
rect 4298 9286 4314 9320
rect 4214 9270 4314 9286
rect 4372 9320 4472 9358
rect 4372 9286 4388 9320
rect 4456 9286 4472 9320
rect 4372 9270 4472 9286
rect 4530 9320 4630 9358
rect 4530 9286 4546 9320
rect 4614 9286 4630 9320
rect 4530 9270 4630 9286
rect 4688 9320 4788 9358
rect 4688 9286 4704 9320
rect 4772 9286 4788 9320
rect 4688 9270 4788 9286
rect 4846 9320 4946 9358
rect 4846 9286 4862 9320
rect 4930 9286 4946 9320
rect 4846 9270 4946 9286
rect 5004 9320 5104 9358
rect 5004 9286 5020 9320
rect 5088 9286 5104 9320
rect 5004 9270 5104 9286
rect 5162 9320 5262 9358
rect 5162 9286 5178 9320
rect 5246 9286 5262 9320
rect 5162 9270 5262 9286
rect 5320 9320 5420 9358
rect 5320 9286 5336 9320
rect 5404 9286 5420 9320
rect 5320 9270 5420 9286
rect 5478 9320 5578 9358
rect 5478 9286 5494 9320
rect 5562 9286 5578 9320
rect 5478 9270 5578 9286
rect 5636 9320 5736 9358
rect 5636 9286 5652 9320
rect 5720 9286 5736 9320
rect 5636 9270 5736 9286
rect 5794 9320 5894 9358
rect 5794 9286 5810 9320
rect 5878 9286 5894 9320
rect 5794 9270 5894 9286
rect 5952 9320 6052 9358
rect 5952 9286 5968 9320
rect 6036 9286 6052 9320
rect 5952 9270 6052 9286
rect 6110 9320 6210 9358
rect 6110 9286 6126 9320
rect 6194 9286 6210 9320
rect 6110 9270 6210 9286
rect 7828 15430 7928 15446
rect 7828 15396 7844 15430
rect 7912 15396 7928 15430
rect 7828 15358 7928 15396
rect 7986 15430 8086 15446
rect 7986 15396 8002 15430
rect 8070 15396 8086 15430
rect 7986 15358 8086 15396
rect 8144 15430 8244 15446
rect 8144 15396 8160 15430
rect 8228 15396 8244 15430
rect 8144 15358 8244 15396
rect 8302 15430 8402 15446
rect 8302 15396 8318 15430
rect 8386 15396 8402 15430
rect 8302 15358 8402 15396
rect 8460 15430 8560 15446
rect 8460 15396 8476 15430
rect 8544 15396 8560 15430
rect 8460 15358 8560 15396
rect 8618 15430 8718 15446
rect 8618 15396 8634 15430
rect 8702 15396 8718 15430
rect 8618 15358 8718 15396
rect 8776 15430 8876 15446
rect 8776 15396 8792 15430
rect 8860 15396 8876 15430
rect 8776 15358 8876 15396
rect 8934 15430 9034 15446
rect 8934 15396 8950 15430
rect 9018 15396 9034 15430
rect 8934 15358 9034 15396
rect 9092 15430 9192 15446
rect 9092 15396 9108 15430
rect 9176 15396 9192 15430
rect 9092 15358 9192 15396
rect 9250 15430 9350 15446
rect 9250 15396 9266 15430
rect 9334 15396 9350 15430
rect 9250 15358 9350 15396
rect 9408 15430 9508 15446
rect 9408 15396 9424 15430
rect 9492 15396 9508 15430
rect 9408 15358 9508 15396
rect 9566 15430 9666 15446
rect 9566 15396 9582 15430
rect 9650 15396 9666 15430
rect 9566 15358 9666 15396
rect 9724 15430 9824 15446
rect 9724 15396 9740 15430
rect 9808 15396 9824 15430
rect 9724 15358 9824 15396
rect 9882 15430 9982 15446
rect 9882 15396 9898 15430
rect 9966 15396 9982 15430
rect 9882 15358 9982 15396
rect 10040 15430 10140 15446
rect 10040 15396 10056 15430
rect 10124 15396 10140 15430
rect 10040 15358 10140 15396
rect 10198 15430 10298 15446
rect 10198 15396 10214 15430
rect 10282 15396 10298 15430
rect 10198 15358 10298 15396
rect 10356 15430 10456 15446
rect 10356 15396 10372 15430
rect 10440 15396 10456 15430
rect 10356 15358 10456 15396
rect 10514 15430 10614 15446
rect 10514 15396 10530 15430
rect 10598 15396 10614 15430
rect 10514 15358 10614 15396
rect 10672 15430 10772 15446
rect 10672 15396 10688 15430
rect 10756 15396 10772 15430
rect 10672 15358 10772 15396
rect 10830 15430 10930 15446
rect 10830 15396 10846 15430
rect 10914 15396 10930 15430
rect 10830 15358 10930 15396
rect 10988 15430 11088 15446
rect 10988 15396 11004 15430
rect 11072 15396 11088 15430
rect 10988 15358 11088 15396
rect 11146 15430 11246 15446
rect 11146 15396 11162 15430
rect 11230 15396 11246 15430
rect 11146 15358 11246 15396
rect 11304 15430 11404 15446
rect 11304 15396 11320 15430
rect 11388 15396 11404 15430
rect 11304 15358 11404 15396
rect 11462 15430 11562 15446
rect 11462 15396 11478 15430
rect 11546 15396 11562 15430
rect 11462 15358 11562 15396
rect 11620 15430 11720 15446
rect 11620 15396 11636 15430
rect 11704 15396 11720 15430
rect 11620 15358 11720 15396
rect 11778 15430 11878 15446
rect 11778 15396 11794 15430
rect 11862 15396 11878 15430
rect 11778 15358 11878 15396
rect 11936 15430 12036 15446
rect 11936 15396 11952 15430
rect 12020 15396 12036 15430
rect 11936 15358 12036 15396
rect 12094 15430 12194 15446
rect 12094 15396 12110 15430
rect 12178 15396 12194 15430
rect 12094 15358 12194 15396
rect 12252 15430 12352 15446
rect 12252 15396 12268 15430
rect 12336 15396 12352 15430
rect 12252 15358 12352 15396
rect 12410 15430 12510 15446
rect 12410 15396 12426 15430
rect 12494 15396 12510 15430
rect 12410 15358 12510 15396
rect 7828 9320 7928 9358
rect 7828 9286 7844 9320
rect 7912 9286 7928 9320
rect 7828 9270 7928 9286
rect 7986 9320 8086 9358
rect 7986 9286 8002 9320
rect 8070 9286 8086 9320
rect 7986 9270 8086 9286
rect 8144 9320 8244 9358
rect 8144 9286 8160 9320
rect 8228 9286 8244 9320
rect 8144 9270 8244 9286
rect 8302 9320 8402 9358
rect 8302 9286 8318 9320
rect 8386 9286 8402 9320
rect 8302 9270 8402 9286
rect 8460 9320 8560 9358
rect 8460 9286 8476 9320
rect 8544 9286 8560 9320
rect 8460 9270 8560 9286
rect 8618 9320 8718 9358
rect 8618 9286 8634 9320
rect 8702 9286 8718 9320
rect 8618 9270 8718 9286
rect 8776 9320 8876 9358
rect 8776 9286 8792 9320
rect 8860 9286 8876 9320
rect 8776 9270 8876 9286
rect 8934 9320 9034 9358
rect 8934 9286 8950 9320
rect 9018 9286 9034 9320
rect 8934 9270 9034 9286
rect 9092 9320 9192 9358
rect 9092 9286 9108 9320
rect 9176 9286 9192 9320
rect 9092 9270 9192 9286
rect 9250 9320 9350 9358
rect 9250 9286 9266 9320
rect 9334 9286 9350 9320
rect 9250 9270 9350 9286
rect 9408 9320 9508 9358
rect 9408 9286 9424 9320
rect 9492 9286 9508 9320
rect 9408 9270 9508 9286
rect 9566 9320 9666 9358
rect 9566 9286 9582 9320
rect 9650 9286 9666 9320
rect 9566 9270 9666 9286
rect 9724 9320 9824 9358
rect 9724 9286 9740 9320
rect 9808 9286 9824 9320
rect 9724 9270 9824 9286
rect 9882 9320 9982 9358
rect 9882 9286 9898 9320
rect 9966 9286 9982 9320
rect 9882 9270 9982 9286
rect 10040 9320 10140 9358
rect 10040 9286 10056 9320
rect 10124 9286 10140 9320
rect 10040 9270 10140 9286
rect 10198 9320 10298 9358
rect 10198 9286 10214 9320
rect 10282 9286 10298 9320
rect 10198 9270 10298 9286
rect 10356 9320 10456 9358
rect 10356 9286 10372 9320
rect 10440 9286 10456 9320
rect 10356 9270 10456 9286
rect 10514 9320 10614 9358
rect 10514 9286 10530 9320
rect 10598 9286 10614 9320
rect 10514 9270 10614 9286
rect 10672 9320 10772 9358
rect 10672 9286 10688 9320
rect 10756 9286 10772 9320
rect 10672 9270 10772 9286
rect 10830 9320 10930 9358
rect 10830 9286 10846 9320
rect 10914 9286 10930 9320
rect 10830 9270 10930 9286
rect 10988 9320 11088 9358
rect 10988 9286 11004 9320
rect 11072 9286 11088 9320
rect 10988 9270 11088 9286
rect 11146 9320 11246 9358
rect 11146 9286 11162 9320
rect 11230 9286 11246 9320
rect 11146 9270 11246 9286
rect 11304 9320 11404 9358
rect 11304 9286 11320 9320
rect 11388 9286 11404 9320
rect 11304 9270 11404 9286
rect 11462 9320 11562 9358
rect 11462 9286 11478 9320
rect 11546 9286 11562 9320
rect 11462 9270 11562 9286
rect 11620 9320 11720 9358
rect 11620 9286 11636 9320
rect 11704 9286 11720 9320
rect 11620 9270 11720 9286
rect 11778 9320 11878 9358
rect 11778 9286 11794 9320
rect 11862 9286 11878 9320
rect 11778 9270 11878 9286
rect 11936 9320 12036 9358
rect 11936 9286 11952 9320
rect 12020 9286 12036 9320
rect 11936 9270 12036 9286
rect 12094 9320 12194 9358
rect 12094 9286 12110 9320
rect 12178 9286 12194 9320
rect 12094 9270 12194 9286
rect 12252 9320 12352 9358
rect 12252 9286 12268 9320
rect 12336 9286 12352 9320
rect 12252 9270 12352 9286
rect 12410 9320 12510 9358
rect 12410 9286 12426 9320
rect 12494 9286 12510 9320
rect 12410 9270 12510 9286
rect 14128 15430 14228 15446
rect 14128 15396 14144 15430
rect 14212 15396 14228 15430
rect 14128 15358 14228 15396
rect 14286 15430 14386 15446
rect 14286 15396 14302 15430
rect 14370 15396 14386 15430
rect 14286 15358 14386 15396
rect 14444 15430 14544 15446
rect 14444 15396 14460 15430
rect 14528 15396 14544 15430
rect 14444 15358 14544 15396
rect 14602 15430 14702 15446
rect 14602 15396 14618 15430
rect 14686 15396 14702 15430
rect 14602 15358 14702 15396
rect 14760 15430 14860 15446
rect 14760 15396 14776 15430
rect 14844 15396 14860 15430
rect 14760 15358 14860 15396
rect 14918 15430 15018 15446
rect 14918 15396 14934 15430
rect 15002 15396 15018 15430
rect 14918 15358 15018 15396
rect 15076 15430 15176 15446
rect 15076 15396 15092 15430
rect 15160 15396 15176 15430
rect 15076 15358 15176 15396
rect 15234 15430 15334 15446
rect 15234 15396 15250 15430
rect 15318 15396 15334 15430
rect 15234 15358 15334 15396
rect 15392 15430 15492 15446
rect 15392 15396 15408 15430
rect 15476 15396 15492 15430
rect 15392 15358 15492 15396
rect 15550 15430 15650 15446
rect 15550 15396 15566 15430
rect 15634 15396 15650 15430
rect 15550 15358 15650 15396
rect 15708 15430 15808 15446
rect 15708 15396 15724 15430
rect 15792 15396 15808 15430
rect 15708 15358 15808 15396
rect 15866 15430 15966 15446
rect 15866 15396 15882 15430
rect 15950 15396 15966 15430
rect 15866 15358 15966 15396
rect 16024 15430 16124 15446
rect 16024 15396 16040 15430
rect 16108 15396 16124 15430
rect 16024 15358 16124 15396
rect 16182 15430 16282 15446
rect 16182 15396 16198 15430
rect 16266 15396 16282 15430
rect 16182 15358 16282 15396
rect 16340 15430 16440 15446
rect 16340 15396 16356 15430
rect 16424 15396 16440 15430
rect 16340 15358 16440 15396
rect 16498 15430 16598 15446
rect 16498 15396 16514 15430
rect 16582 15396 16598 15430
rect 16498 15358 16598 15396
rect 16656 15430 16756 15446
rect 16656 15396 16672 15430
rect 16740 15396 16756 15430
rect 16656 15358 16756 15396
rect 16814 15430 16914 15446
rect 16814 15396 16830 15430
rect 16898 15396 16914 15430
rect 16814 15358 16914 15396
rect 16972 15430 17072 15446
rect 16972 15396 16988 15430
rect 17056 15396 17072 15430
rect 16972 15358 17072 15396
rect 17130 15430 17230 15446
rect 17130 15396 17146 15430
rect 17214 15396 17230 15430
rect 17130 15358 17230 15396
rect 17288 15430 17388 15446
rect 17288 15396 17304 15430
rect 17372 15396 17388 15430
rect 17288 15358 17388 15396
rect 17446 15430 17546 15446
rect 17446 15396 17462 15430
rect 17530 15396 17546 15430
rect 17446 15358 17546 15396
rect 17604 15430 17704 15446
rect 17604 15396 17620 15430
rect 17688 15396 17704 15430
rect 17604 15358 17704 15396
rect 17762 15430 17862 15446
rect 17762 15396 17778 15430
rect 17846 15396 17862 15430
rect 17762 15358 17862 15396
rect 17920 15430 18020 15446
rect 17920 15396 17936 15430
rect 18004 15396 18020 15430
rect 17920 15358 18020 15396
rect 18078 15430 18178 15446
rect 18078 15396 18094 15430
rect 18162 15396 18178 15430
rect 18078 15358 18178 15396
rect 18236 15430 18336 15446
rect 18236 15396 18252 15430
rect 18320 15396 18336 15430
rect 18236 15358 18336 15396
rect 18394 15430 18494 15446
rect 18394 15396 18410 15430
rect 18478 15396 18494 15430
rect 18394 15358 18494 15396
rect 18552 15430 18652 15446
rect 18552 15396 18568 15430
rect 18636 15396 18652 15430
rect 18552 15358 18652 15396
rect 18710 15430 18810 15446
rect 18710 15396 18726 15430
rect 18794 15396 18810 15430
rect 18710 15358 18810 15396
rect 14128 9320 14228 9358
rect 14128 9286 14144 9320
rect 14212 9286 14228 9320
rect 14128 9270 14228 9286
rect 14286 9320 14386 9358
rect 14286 9286 14302 9320
rect 14370 9286 14386 9320
rect 14286 9270 14386 9286
rect 14444 9320 14544 9358
rect 14444 9286 14460 9320
rect 14528 9286 14544 9320
rect 14444 9270 14544 9286
rect 14602 9320 14702 9358
rect 14602 9286 14618 9320
rect 14686 9286 14702 9320
rect 14602 9270 14702 9286
rect 14760 9320 14860 9358
rect 14760 9286 14776 9320
rect 14844 9286 14860 9320
rect 14760 9270 14860 9286
rect 14918 9320 15018 9358
rect 14918 9286 14934 9320
rect 15002 9286 15018 9320
rect 14918 9270 15018 9286
rect 15076 9320 15176 9358
rect 15076 9286 15092 9320
rect 15160 9286 15176 9320
rect 15076 9270 15176 9286
rect 15234 9320 15334 9358
rect 15234 9286 15250 9320
rect 15318 9286 15334 9320
rect 15234 9270 15334 9286
rect 15392 9320 15492 9358
rect 15392 9286 15408 9320
rect 15476 9286 15492 9320
rect 15392 9270 15492 9286
rect 15550 9320 15650 9358
rect 15550 9286 15566 9320
rect 15634 9286 15650 9320
rect 15550 9270 15650 9286
rect 15708 9320 15808 9358
rect 15708 9286 15724 9320
rect 15792 9286 15808 9320
rect 15708 9270 15808 9286
rect 15866 9320 15966 9358
rect 15866 9286 15882 9320
rect 15950 9286 15966 9320
rect 15866 9270 15966 9286
rect 16024 9320 16124 9358
rect 16024 9286 16040 9320
rect 16108 9286 16124 9320
rect 16024 9270 16124 9286
rect 16182 9320 16282 9358
rect 16182 9286 16198 9320
rect 16266 9286 16282 9320
rect 16182 9270 16282 9286
rect 16340 9320 16440 9358
rect 16340 9286 16356 9320
rect 16424 9286 16440 9320
rect 16340 9270 16440 9286
rect 16498 9320 16598 9358
rect 16498 9286 16514 9320
rect 16582 9286 16598 9320
rect 16498 9270 16598 9286
rect 16656 9320 16756 9358
rect 16656 9286 16672 9320
rect 16740 9286 16756 9320
rect 16656 9270 16756 9286
rect 16814 9320 16914 9358
rect 16814 9286 16830 9320
rect 16898 9286 16914 9320
rect 16814 9270 16914 9286
rect 16972 9320 17072 9358
rect 16972 9286 16988 9320
rect 17056 9286 17072 9320
rect 16972 9270 17072 9286
rect 17130 9320 17230 9358
rect 17130 9286 17146 9320
rect 17214 9286 17230 9320
rect 17130 9270 17230 9286
rect 17288 9320 17388 9358
rect 17288 9286 17304 9320
rect 17372 9286 17388 9320
rect 17288 9270 17388 9286
rect 17446 9320 17546 9358
rect 17446 9286 17462 9320
rect 17530 9286 17546 9320
rect 17446 9270 17546 9286
rect 17604 9320 17704 9358
rect 17604 9286 17620 9320
rect 17688 9286 17704 9320
rect 17604 9270 17704 9286
rect 17762 9320 17862 9358
rect 17762 9286 17778 9320
rect 17846 9286 17862 9320
rect 17762 9270 17862 9286
rect 17920 9320 18020 9358
rect 17920 9286 17936 9320
rect 18004 9286 18020 9320
rect 17920 9270 18020 9286
rect 18078 9320 18178 9358
rect 18078 9286 18094 9320
rect 18162 9286 18178 9320
rect 18078 9270 18178 9286
rect 18236 9320 18336 9358
rect 18236 9286 18252 9320
rect 18320 9286 18336 9320
rect 18236 9270 18336 9286
rect 18394 9320 18494 9358
rect 18394 9286 18410 9320
rect 18478 9286 18494 9320
rect 18394 9270 18494 9286
rect 18552 9320 18652 9358
rect 18552 9286 18568 9320
rect 18636 9286 18652 9320
rect 18552 9270 18652 9286
rect 18710 9320 18810 9358
rect 18710 9286 18726 9320
rect 18794 9286 18810 9320
rect 18710 9270 18810 9286
rect 20428 15430 20528 15446
rect 20428 15396 20444 15430
rect 20512 15396 20528 15430
rect 20428 15358 20528 15396
rect 20586 15430 20686 15446
rect 20586 15396 20602 15430
rect 20670 15396 20686 15430
rect 20586 15358 20686 15396
rect 20744 15430 20844 15446
rect 20744 15396 20760 15430
rect 20828 15396 20844 15430
rect 20744 15358 20844 15396
rect 20902 15430 21002 15446
rect 20902 15396 20918 15430
rect 20986 15396 21002 15430
rect 20902 15358 21002 15396
rect 21060 15430 21160 15446
rect 21060 15396 21076 15430
rect 21144 15396 21160 15430
rect 21060 15358 21160 15396
rect 21218 15430 21318 15446
rect 21218 15396 21234 15430
rect 21302 15396 21318 15430
rect 21218 15358 21318 15396
rect 21376 15430 21476 15446
rect 21376 15396 21392 15430
rect 21460 15396 21476 15430
rect 21376 15358 21476 15396
rect 21534 15430 21634 15446
rect 21534 15396 21550 15430
rect 21618 15396 21634 15430
rect 21534 15358 21634 15396
rect 21692 15430 21792 15446
rect 21692 15396 21708 15430
rect 21776 15396 21792 15430
rect 21692 15358 21792 15396
rect 21850 15430 21950 15446
rect 21850 15396 21866 15430
rect 21934 15396 21950 15430
rect 21850 15358 21950 15396
rect 22008 15430 22108 15446
rect 22008 15396 22024 15430
rect 22092 15396 22108 15430
rect 22008 15358 22108 15396
rect 22166 15430 22266 15446
rect 22166 15396 22182 15430
rect 22250 15396 22266 15430
rect 22166 15358 22266 15396
rect 22324 15430 22424 15446
rect 22324 15396 22340 15430
rect 22408 15396 22424 15430
rect 22324 15358 22424 15396
rect 22482 15430 22582 15446
rect 22482 15396 22498 15430
rect 22566 15396 22582 15430
rect 22482 15358 22582 15396
rect 22640 15430 22740 15446
rect 22640 15396 22656 15430
rect 22724 15396 22740 15430
rect 22640 15358 22740 15396
rect 22798 15430 22898 15446
rect 22798 15396 22814 15430
rect 22882 15396 22898 15430
rect 22798 15358 22898 15396
rect 22956 15430 23056 15446
rect 22956 15396 22972 15430
rect 23040 15396 23056 15430
rect 22956 15358 23056 15396
rect 23114 15430 23214 15446
rect 23114 15396 23130 15430
rect 23198 15396 23214 15430
rect 23114 15358 23214 15396
rect 23272 15430 23372 15446
rect 23272 15396 23288 15430
rect 23356 15396 23372 15430
rect 23272 15358 23372 15396
rect 23430 15430 23530 15446
rect 23430 15396 23446 15430
rect 23514 15396 23530 15430
rect 23430 15358 23530 15396
rect 23588 15430 23688 15446
rect 23588 15396 23604 15430
rect 23672 15396 23688 15430
rect 23588 15358 23688 15396
rect 23746 15430 23846 15446
rect 23746 15396 23762 15430
rect 23830 15396 23846 15430
rect 23746 15358 23846 15396
rect 23904 15430 24004 15446
rect 23904 15396 23920 15430
rect 23988 15396 24004 15430
rect 23904 15358 24004 15396
rect 24062 15430 24162 15446
rect 24062 15396 24078 15430
rect 24146 15396 24162 15430
rect 24062 15358 24162 15396
rect 24220 15430 24320 15446
rect 24220 15396 24236 15430
rect 24304 15396 24320 15430
rect 24220 15358 24320 15396
rect 24378 15430 24478 15446
rect 24378 15396 24394 15430
rect 24462 15396 24478 15430
rect 24378 15358 24478 15396
rect 24536 15430 24636 15446
rect 24536 15396 24552 15430
rect 24620 15396 24636 15430
rect 24536 15358 24636 15396
rect 24694 15430 24794 15446
rect 24694 15396 24710 15430
rect 24778 15396 24794 15430
rect 24694 15358 24794 15396
rect 24852 15430 24952 15446
rect 24852 15396 24868 15430
rect 24936 15396 24952 15430
rect 24852 15358 24952 15396
rect 25010 15430 25110 15446
rect 25010 15396 25026 15430
rect 25094 15396 25110 15430
rect 25010 15358 25110 15396
rect 20428 9320 20528 9358
rect 20428 9286 20444 9320
rect 20512 9286 20528 9320
rect 20428 9270 20528 9286
rect 20586 9320 20686 9358
rect 20586 9286 20602 9320
rect 20670 9286 20686 9320
rect 20586 9270 20686 9286
rect 20744 9320 20844 9358
rect 20744 9286 20760 9320
rect 20828 9286 20844 9320
rect 20744 9270 20844 9286
rect 20902 9320 21002 9358
rect 20902 9286 20918 9320
rect 20986 9286 21002 9320
rect 20902 9270 21002 9286
rect 21060 9320 21160 9358
rect 21060 9286 21076 9320
rect 21144 9286 21160 9320
rect 21060 9270 21160 9286
rect 21218 9320 21318 9358
rect 21218 9286 21234 9320
rect 21302 9286 21318 9320
rect 21218 9270 21318 9286
rect 21376 9320 21476 9358
rect 21376 9286 21392 9320
rect 21460 9286 21476 9320
rect 21376 9270 21476 9286
rect 21534 9320 21634 9358
rect 21534 9286 21550 9320
rect 21618 9286 21634 9320
rect 21534 9270 21634 9286
rect 21692 9320 21792 9358
rect 21692 9286 21708 9320
rect 21776 9286 21792 9320
rect 21692 9270 21792 9286
rect 21850 9320 21950 9358
rect 21850 9286 21866 9320
rect 21934 9286 21950 9320
rect 21850 9270 21950 9286
rect 22008 9320 22108 9358
rect 22008 9286 22024 9320
rect 22092 9286 22108 9320
rect 22008 9270 22108 9286
rect 22166 9320 22266 9358
rect 22166 9286 22182 9320
rect 22250 9286 22266 9320
rect 22166 9270 22266 9286
rect 22324 9320 22424 9358
rect 22324 9286 22340 9320
rect 22408 9286 22424 9320
rect 22324 9270 22424 9286
rect 22482 9320 22582 9358
rect 22482 9286 22498 9320
rect 22566 9286 22582 9320
rect 22482 9270 22582 9286
rect 22640 9320 22740 9358
rect 22640 9286 22656 9320
rect 22724 9286 22740 9320
rect 22640 9270 22740 9286
rect 22798 9320 22898 9358
rect 22798 9286 22814 9320
rect 22882 9286 22898 9320
rect 22798 9270 22898 9286
rect 22956 9320 23056 9358
rect 22956 9286 22972 9320
rect 23040 9286 23056 9320
rect 22956 9270 23056 9286
rect 23114 9320 23214 9358
rect 23114 9286 23130 9320
rect 23198 9286 23214 9320
rect 23114 9270 23214 9286
rect 23272 9320 23372 9358
rect 23272 9286 23288 9320
rect 23356 9286 23372 9320
rect 23272 9270 23372 9286
rect 23430 9320 23530 9358
rect 23430 9286 23446 9320
rect 23514 9286 23530 9320
rect 23430 9270 23530 9286
rect 23588 9320 23688 9358
rect 23588 9286 23604 9320
rect 23672 9286 23688 9320
rect 23588 9270 23688 9286
rect 23746 9320 23846 9358
rect 23746 9286 23762 9320
rect 23830 9286 23846 9320
rect 23746 9270 23846 9286
rect 23904 9320 24004 9358
rect 23904 9286 23920 9320
rect 23988 9286 24004 9320
rect 23904 9270 24004 9286
rect 24062 9320 24162 9358
rect 24062 9286 24078 9320
rect 24146 9286 24162 9320
rect 24062 9270 24162 9286
rect 24220 9320 24320 9358
rect 24220 9286 24236 9320
rect 24304 9286 24320 9320
rect 24220 9270 24320 9286
rect 24378 9320 24478 9358
rect 24378 9286 24394 9320
rect 24462 9286 24478 9320
rect 24378 9270 24478 9286
rect 24536 9320 24636 9358
rect 24536 9286 24552 9320
rect 24620 9286 24636 9320
rect 24536 9270 24636 9286
rect 24694 9320 24794 9358
rect 24694 9286 24710 9320
rect 24778 9286 24794 9320
rect 24694 9270 24794 9286
rect 24852 9320 24952 9358
rect 24852 9286 24868 9320
rect 24936 9286 24952 9320
rect 24852 9270 24952 9286
rect 25010 9320 25110 9358
rect 25010 9286 25026 9320
rect 25094 9286 25110 9320
rect 25010 9270 25110 9286
rect 1528 8430 1628 8446
rect 1528 8396 1544 8430
rect 1612 8396 1628 8430
rect 1528 8358 1628 8396
rect 1686 8430 1786 8446
rect 1686 8396 1702 8430
rect 1770 8396 1786 8430
rect 1686 8358 1786 8396
rect 1844 8430 1944 8446
rect 1844 8396 1860 8430
rect 1928 8396 1944 8430
rect 1844 8358 1944 8396
rect 2002 8430 2102 8446
rect 2002 8396 2018 8430
rect 2086 8396 2102 8430
rect 2002 8358 2102 8396
rect 2160 8430 2260 8446
rect 2160 8396 2176 8430
rect 2244 8396 2260 8430
rect 2160 8358 2260 8396
rect 2318 8430 2418 8446
rect 2318 8396 2334 8430
rect 2402 8396 2418 8430
rect 2318 8358 2418 8396
rect 2476 8430 2576 8446
rect 2476 8396 2492 8430
rect 2560 8396 2576 8430
rect 2476 8358 2576 8396
rect 2634 8430 2734 8446
rect 2634 8396 2650 8430
rect 2718 8396 2734 8430
rect 2634 8358 2734 8396
rect 2792 8430 2892 8446
rect 2792 8396 2808 8430
rect 2876 8396 2892 8430
rect 2792 8358 2892 8396
rect 2950 8430 3050 8446
rect 2950 8396 2966 8430
rect 3034 8396 3050 8430
rect 2950 8358 3050 8396
rect 3108 8430 3208 8446
rect 3108 8396 3124 8430
rect 3192 8396 3208 8430
rect 3108 8358 3208 8396
rect 3266 8430 3366 8446
rect 3266 8396 3282 8430
rect 3350 8396 3366 8430
rect 3266 8358 3366 8396
rect 3424 8430 3524 8446
rect 3424 8396 3440 8430
rect 3508 8396 3524 8430
rect 3424 8358 3524 8396
rect 3582 8430 3682 8446
rect 3582 8396 3598 8430
rect 3666 8396 3682 8430
rect 3582 8358 3682 8396
rect 3740 8430 3840 8446
rect 3740 8396 3756 8430
rect 3824 8396 3840 8430
rect 3740 8358 3840 8396
rect 3898 8430 3998 8446
rect 3898 8396 3914 8430
rect 3982 8396 3998 8430
rect 3898 8358 3998 8396
rect 4056 8430 4156 8446
rect 4056 8396 4072 8430
rect 4140 8396 4156 8430
rect 4056 8358 4156 8396
rect 4214 8430 4314 8446
rect 4214 8396 4230 8430
rect 4298 8396 4314 8430
rect 4214 8358 4314 8396
rect 4372 8430 4472 8446
rect 4372 8396 4388 8430
rect 4456 8396 4472 8430
rect 4372 8358 4472 8396
rect 4530 8430 4630 8446
rect 4530 8396 4546 8430
rect 4614 8396 4630 8430
rect 4530 8358 4630 8396
rect 4688 8430 4788 8446
rect 4688 8396 4704 8430
rect 4772 8396 4788 8430
rect 4688 8358 4788 8396
rect 4846 8430 4946 8446
rect 4846 8396 4862 8430
rect 4930 8396 4946 8430
rect 4846 8358 4946 8396
rect 5004 8430 5104 8446
rect 5004 8396 5020 8430
rect 5088 8396 5104 8430
rect 5004 8358 5104 8396
rect 5162 8430 5262 8446
rect 5162 8396 5178 8430
rect 5246 8396 5262 8430
rect 5162 8358 5262 8396
rect 5320 8430 5420 8446
rect 5320 8396 5336 8430
rect 5404 8396 5420 8430
rect 5320 8358 5420 8396
rect 5478 8430 5578 8446
rect 5478 8396 5494 8430
rect 5562 8396 5578 8430
rect 5478 8358 5578 8396
rect 5636 8430 5736 8446
rect 5636 8396 5652 8430
rect 5720 8396 5736 8430
rect 5636 8358 5736 8396
rect 5794 8430 5894 8446
rect 5794 8396 5810 8430
rect 5878 8396 5894 8430
rect 5794 8358 5894 8396
rect 5952 8430 6052 8446
rect 5952 8396 5968 8430
rect 6036 8396 6052 8430
rect 5952 8358 6052 8396
rect 6110 8430 6210 8446
rect 6110 8396 6126 8430
rect 6194 8396 6210 8430
rect 6110 8358 6210 8396
rect 1528 2320 1628 2358
rect 1528 2286 1544 2320
rect 1612 2286 1628 2320
rect 1528 2270 1628 2286
rect 1686 2320 1786 2358
rect 1686 2286 1702 2320
rect 1770 2286 1786 2320
rect 1686 2270 1786 2286
rect 1844 2320 1944 2358
rect 1844 2286 1860 2320
rect 1928 2286 1944 2320
rect 1844 2270 1944 2286
rect 2002 2320 2102 2358
rect 2002 2286 2018 2320
rect 2086 2286 2102 2320
rect 2002 2270 2102 2286
rect 2160 2320 2260 2358
rect 2160 2286 2176 2320
rect 2244 2286 2260 2320
rect 2160 2270 2260 2286
rect 2318 2320 2418 2358
rect 2318 2286 2334 2320
rect 2402 2286 2418 2320
rect 2318 2270 2418 2286
rect 2476 2320 2576 2358
rect 2476 2286 2492 2320
rect 2560 2286 2576 2320
rect 2476 2270 2576 2286
rect 2634 2320 2734 2358
rect 2634 2286 2650 2320
rect 2718 2286 2734 2320
rect 2634 2270 2734 2286
rect 2792 2320 2892 2358
rect 2792 2286 2808 2320
rect 2876 2286 2892 2320
rect 2792 2270 2892 2286
rect 2950 2320 3050 2358
rect 2950 2286 2966 2320
rect 3034 2286 3050 2320
rect 2950 2270 3050 2286
rect 3108 2320 3208 2358
rect 3108 2286 3124 2320
rect 3192 2286 3208 2320
rect 3108 2270 3208 2286
rect 3266 2320 3366 2358
rect 3266 2286 3282 2320
rect 3350 2286 3366 2320
rect 3266 2270 3366 2286
rect 3424 2320 3524 2358
rect 3424 2286 3440 2320
rect 3508 2286 3524 2320
rect 3424 2270 3524 2286
rect 3582 2320 3682 2358
rect 3582 2286 3598 2320
rect 3666 2286 3682 2320
rect 3582 2270 3682 2286
rect 3740 2320 3840 2358
rect 3740 2286 3756 2320
rect 3824 2286 3840 2320
rect 3740 2270 3840 2286
rect 3898 2320 3998 2358
rect 3898 2286 3914 2320
rect 3982 2286 3998 2320
rect 3898 2270 3998 2286
rect 4056 2320 4156 2358
rect 4056 2286 4072 2320
rect 4140 2286 4156 2320
rect 4056 2270 4156 2286
rect 4214 2320 4314 2358
rect 4214 2286 4230 2320
rect 4298 2286 4314 2320
rect 4214 2270 4314 2286
rect 4372 2320 4472 2358
rect 4372 2286 4388 2320
rect 4456 2286 4472 2320
rect 4372 2270 4472 2286
rect 4530 2320 4630 2358
rect 4530 2286 4546 2320
rect 4614 2286 4630 2320
rect 4530 2270 4630 2286
rect 4688 2320 4788 2358
rect 4688 2286 4704 2320
rect 4772 2286 4788 2320
rect 4688 2270 4788 2286
rect 4846 2320 4946 2358
rect 4846 2286 4862 2320
rect 4930 2286 4946 2320
rect 4846 2270 4946 2286
rect 5004 2320 5104 2358
rect 5004 2286 5020 2320
rect 5088 2286 5104 2320
rect 5004 2270 5104 2286
rect 5162 2320 5262 2358
rect 5162 2286 5178 2320
rect 5246 2286 5262 2320
rect 5162 2270 5262 2286
rect 5320 2320 5420 2358
rect 5320 2286 5336 2320
rect 5404 2286 5420 2320
rect 5320 2270 5420 2286
rect 5478 2320 5578 2358
rect 5478 2286 5494 2320
rect 5562 2286 5578 2320
rect 5478 2270 5578 2286
rect 5636 2320 5736 2358
rect 5636 2286 5652 2320
rect 5720 2286 5736 2320
rect 5636 2270 5736 2286
rect 5794 2320 5894 2358
rect 5794 2286 5810 2320
rect 5878 2286 5894 2320
rect 5794 2270 5894 2286
rect 5952 2320 6052 2358
rect 5952 2286 5968 2320
rect 6036 2286 6052 2320
rect 5952 2270 6052 2286
rect 6110 2320 6210 2358
rect 6110 2286 6126 2320
rect 6194 2286 6210 2320
rect 6110 2270 6210 2286
rect 7828 8430 7928 8446
rect 7828 8396 7844 8430
rect 7912 8396 7928 8430
rect 7828 8358 7928 8396
rect 7986 8430 8086 8446
rect 7986 8396 8002 8430
rect 8070 8396 8086 8430
rect 7986 8358 8086 8396
rect 8144 8430 8244 8446
rect 8144 8396 8160 8430
rect 8228 8396 8244 8430
rect 8144 8358 8244 8396
rect 8302 8430 8402 8446
rect 8302 8396 8318 8430
rect 8386 8396 8402 8430
rect 8302 8358 8402 8396
rect 8460 8430 8560 8446
rect 8460 8396 8476 8430
rect 8544 8396 8560 8430
rect 8460 8358 8560 8396
rect 8618 8430 8718 8446
rect 8618 8396 8634 8430
rect 8702 8396 8718 8430
rect 8618 8358 8718 8396
rect 8776 8430 8876 8446
rect 8776 8396 8792 8430
rect 8860 8396 8876 8430
rect 8776 8358 8876 8396
rect 8934 8430 9034 8446
rect 8934 8396 8950 8430
rect 9018 8396 9034 8430
rect 8934 8358 9034 8396
rect 9092 8430 9192 8446
rect 9092 8396 9108 8430
rect 9176 8396 9192 8430
rect 9092 8358 9192 8396
rect 9250 8430 9350 8446
rect 9250 8396 9266 8430
rect 9334 8396 9350 8430
rect 9250 8358 9350 8396
rect 9408 8430 9508 8446
rect 9408 8396 9424 8430
rect 9492 8396 9508 8430
rect 9408 8358 9508 8396
rect 9566 8430 9666 8446
rect 9566 8396 9582 8430
rect 9650 8396 9666 8430
rect 9566 8358 9666 8396
rect 9724 8430 9824 8446
rect 9724 8396 9740 8430
rect 9808 8396 9824 8430
rect 9724 8358 9824 8396
rect 9882 8430 9982 8446
rect 9882 8396 9898 8430
rect 9966 8396 9982 8430
rect 9882 8358 9982 8396
rect 10040 8430 10140 8446
rect 10040 8396 10056 8430
rect 10124 8396 10140 8430
rect 10040 8358 10140 8396
rect 10198 8430 10298 8446
rect 10198 8396 10214 8430
rect 10282 8396 10298 8430
rect 10198 8358 10298 8396
rect 10356 8430 10456 8446
rect 10356 8396 10372 8430
rect 10440 8396 10456 8430
rect 10356 8358 10456 8396
rect 10514 8430 10614 8446
rect 10514 8396 10530 8430
rect 10598 8396 10614 8430
rect 10514 8358 10614 8396
rect 10672 8430 10772 8446
rect 10672 8396 10688 8430
rect 10756 8396 10772 8430
rect 10672 8358 10772 8396
rect 10830 8430 10930 8446
rect 10830 8396 10846 8430
rect 10914 8396 10930 8430
rect 10830 8358 10930 8396
rect 10988 8430 11088 8446
rect 10988 8396 11004 8430
rect 11072 8396 11088 8430
rect 10988 8358 11088 8396
rect 11146 8430 11246 8446
rect 11146 8396 11162 8430
rect 11230 8396 11246 8430
rect 11146 8358 11246 8396
rect 11304 8430 11404 8446
rect 11304 8396 11320 8430
rect 11388 8396 11404 8430
rect 11304 8358 11404 8396
rect 11462 8430 11562 8446
rect 11462 8396 11478 8430
rect 11546 8396 11562 8430
rect 11462 8358 11562 8396
rect 11620 8430 11720 8446
rect 11620 8396 11636 8430
rect 11704 8396 11720 8430
rect 11620 8358 11720 8396
rect 11778 8430 11878 8446
rect 11778 8396 11794 8430
rect 11862 8396 11878 8430
rect 11778 8358 11878 8396
rect 11936 8430 12036 8446
rect 11936 8396 11952 8430
rect 12020 8396 12036 8430
rect 11936 8358 12036 8396
rect 12094 8430 12194 8446
rect 12094 8396 12110 8430
rect 12178 8396 12194 8430
rect 12094 8358 12194 8396
rect 12252 8430 12352 8446
rect 12252 8396 12268 8430
rect 12336 8396 12352 8430
rect 12252 8358 12352 8396
rect 12410 8430 12510 8446
rect 12410 8396 12426 8430
rect 12494 8396 12510 8430
rect 12410 8358 12510 8396
rect 7828 2320 7928 2358
rect 7828 2286 7844 2320
rect 7912 2286 7928 2320
rect 7828 2270 7928 2286
rect 7986 2320 8086 2358
rect 7986 2286 8002 2320
rect 8070 2286 8086 2320
rect 7986 2270 8086 2286
rect 8144 2320 8244 2358
rect 8144 2286 8160 2320
rect 8228 2286 8244 2320
rect 8144 2270 8244 2286
rect 8302 2320 8402 2358
rect 8302 2286 8318 2320
rect 8386 2286 8402 2320
rect 8302 2270 8402 2286
rect 8460 2320 8560 2358
rect 8460 2286 8476 2320
rect 8544 2286 8560 2320
rect 8460 2270 8560 2286
rect 8618 2320 8718 2358
rect 8618 2286 8634 2320
rect 8702 2286 8718 2320
rect 8618 2270 8718 2286
rect 8776 2320 8876 2358
rect 8776 2286 8792 2320
rect 8860 2286 8876 2320
rect 8776 2270 8876 2286
rect 8934 2320 9034 2358
rect 8934 2286 8950 2320
rect 9018 2286 9034 2320
rect 8934 2270 9034 2286
rect 9092 2320 9192 2358
rect 9092 2286 9108 2320
rect 9176 2286 9192 2320
rect 9092 2270 9192 2286
rect 9250 2320 9350 2358
rect 9250 2286 9266 2320
rect 9334 2286 9350 2320
rect 9250 2270 9350 2286
rect 9408 2320 9508 2358
rect 9408 2286 9424 2320
rect 9492 2286 9508 2320
rect 9408 2270 9508 2286
rect 9566 2320 9666 2358
rect 9566 2286 9582 2320
rect 9650 2286 9666 2320
rect 9566 2270 9666 2286
rect 9724 2320 9824 2358
rect 9724 2286 9740 2320
rect 9808 2286 9824 2320
rect 9724 2270 9824 2286
rect 9882 2320 9982 2358
rect 9882 2286 9898 2320
rect 9966 2286 9982 2320
rect 9882 2270 9982 2286
rect 10040 2320 10140 2358
rect 10040 2286 10056 2320
rect 10124 2286 10140 2320
rect 10040 2270 10140 2286
rect 10198 2320 10298 2358
rect 10198 2286 10214 2320
rect 10282 2286 10298 2320
rect 10198 2270 10298 2286
rect 10356 2320 10456 2358
rect 10356 2286 10372 2320
rect 10440 2286 10456 2320
rect 10356 2270 10456 2286
rect 10514 2320 10614 2358
rect 10514 2286 10530 2320
rect 10598 2286 10614 2320
rect 10514 2270 10614 2286
rect 10672 2320 10772 2358
rect 10672 2286 10688 2320
rect 10756 2286 10772 2320
rect 10672 2270 10772 2286
rect 10830 2320 10930 2358
rect 10830 2286 10846 2320
rect 10914 2286 10930 2320
rect 10830 2270 10930 2286
rect 10988 2320 11088 2358
rect 10988 2286 11004 2320
rect 11072 2286 11088 2320
rect 10988 2270 11088 2286
rect 11146 2320 11246 2358
rect 11146 2286 11162 2320
rect 11230 2286 11246 2320
rect 11146 2270 11246 2286
rect 11304 2320 11404 2358
rect 11304 2286 11320 2320
rect 11388 2286 11404 2320
rect 11304 2270 11404 2286
rect 11462 2320 11562 2358
rect 11462 2286 11478 2320
rect 11546 2286 11562 2320
rect 11462 2270 11562 2286
rect 11620 2320 11720 2358
rect 11620 2286 11636 2320
rect 11704 2286 11720 2320
rect 11620 2270 11720 2286
rect 11778 2320 11878 2358
rect 11778 2286 11794 2320
rect 11862 2286 11878 2320
rect 11778 2270 11878 2286
rect 11936 2320 12036 2358
rect 11936 2286 11952 2320
rect 12020 2286 12036 2320
rect 11936 2270 12036 2286
rect 12094 2320 12194 2358
rect 12094 2286 12110 2320
rect 12178 2286 12194 2320
rect 12094 2270 12194 2286
rect 12252 2320 12352 2358
rect 12252 2286 12268 2320
rect 12336 2286 12352 2320
rect 12252 2270 12352 2286
rect 12410 2320 12510 2358
rect 12410 2286 12426 2320
rect 12494 2286 12510 2320
rect 12410 2270 12510 2286
rect 14128 8430 14228 8446
rect 14128 8396 14144 8430
rect 14212 8396 14228 8430
rect 14128 8358 14228 8396
rect 14286 8430 14386 8446
rect 14286 8396 14302 8430
rect 14370 8396 14386 8430
rect 14286 8358 14386 8396
rect 14444 8430 14544 8446
rect 14444 8396 14460 8430
rect 14528 8396 14544 8430
rect 14444 8358 14544 8396
rect 14602 8430 14702 8446
rect 14602 8396 14618 8430
rect 14686 8396 14702 8430
rect 14602 8358 14702 8396
rect 14760 8430 14860 8446
rect 14760 8396 14776 8430
rect 14844 8396 14860 8430
rect 14760 8358 14860 8396
rect 14918 8430 15018 8446
rect 14918 8396 14934 8430
rect 15002 8396 15018 8430
rect 14918 8358 15018 8396
rect 15076 8430 15176 8446
rect 15076 8396 15092 8430
rect 15160 8396 15176 8430
rect 15076 8358 15176 8396
rect 15234 8430 15334 8446
rect 15234 8396 15250 8430
rect 15318 8396 15334 8430
rect 15234 8358 15334 8396
rect 15392 8430 15492 8446
rect 15392 8396 15408 8430
rect 15476 8396 15492 8430
rect 15392 8358 15492 8396
rect 15550 8430 15650 8446
rect 15550 8396 15566 8430
rect 15634 8396 15650 8430
rect 15550 8358 15650 8396
rect 15708 8430 15808 8446
rect 15708 8396 15724 8430
rect 15792 8396 15808 8430
rect 15708 8358 15808 8396
rect 15866 8430 15966 8446
rect 15866 8396 15882 8430
rect 15950 8396 15966 8430
rect 15866 8358 15966 8396
rect 16024 8430 16124 8446
rect 16024 8396 16040 8430
rect 16108 8396 16124 8430
rect 16024 8358 16124 8396
rect 16182 8430 16282 8446
rect 16182 8396 16198 8430
rect 16266 8396 16282 8430
rect 16182 8358 16282 8396
rect 16340 8430 16440 8446
rect 16340 8396 16356 8430
rect 16424 8396 16440 8430
rect 16340 8358 16440 8396
rect 16498 8430 16598 8446
rect 16498 8396 16514 8430
rect 16582 8396 16598 8430
rect 16498 8358 16598 8396
rect 16656 8430 16756 8446
rect 16656 8396 16672 8430
rect 16740 8396 16756 8430
rect 16656 8358 16756 8396
rect 16814 8430 16914 8446
rect 16814 8396 16830 8430
rect 16898 8396 16914 8430
rect 16814 8358 16914 8396
rect 16972 8430 17072 8446
rect 16972 8396 16988 8430
rect 17056 8396 17072 8430
rect 16972 8358 17072 8396
rect 17130 8430 17230 8446
rect 17130 8396 17146 8430
rect 17214 8396 17230 8430
rect 17130 8358 17230 8396
rect 17288 8430 17388 8446
rect 17288 8396 17304 8430
rect 17372 8396 17388 8430
rect 17288 8358 17388 8396
rect 17446 8430 17546 8446
rect 17446 8396 17462 8430
rect 17530 8396 17546 8430
rect 17446 8358 17546 8396
rect 17604 8430 17704 8446
rect 17604 8396 17620 8430
rect 17688 8396 17704 8430
rect 17604 8358 17704 8396
rect 17762 8430 17862 8446
rect 17762 8396 17778 8430
rect 17846 8396 17862 8430
rect 17762 8358 17862 8396
rect 17920 8430 18020 8446
rect 17920 8396 17936 8430
rect 18004 8396 18020 8430
rect 17920 8358 18020 8396
rect 18078 8430 18178 8446
rect 18078 8396 18094 8430
rect 18162 8396 18178 8430
rect 18078 8358 18178 8396
rect 18236 8430 18336 8446
rect 18236 8396 18252 8430
rect 18320 8396 18336 8430
rect 18236 8358 18336 8396
rect 18394 8430 18494 8446
rect 18394 8396 18410 8430
rect 18478 8396 18494 8430
rect 18394 8358 18494 8396
rect 18552 8430 18652 8446
rect 18552 8396 18568 8430
rect 18636 8396 18652 8430
rect 18552 8358 18652 8396
rect 18710 8430 18810 8446
rect 18710 8396 18726 8430
rect 18794 8396 18810 8430
rect 18710 8358 18810 8396
rect 14128 2320 14228 2358
rect 14128 2286 14144 2320
rect 14212 2286 14228 2320
rect 14128 2270 14228 2286
rect 14286 2320 14386 2358
rect 14286 2286 14302 2320
rect 14370 2286 14386 2320
rect 14286 2270 14386 2286
rect 14444 2320 14544 2358
rect 14444 2286 14460 2320
rect 14528 2286 14544 2320
rect 14444 2270 14544 2286
rect 14602 2320 14702 2358
rect 14602 2286 14618 2320
rect 14686 2286 14702 2320
rect 14602 2270 14702 2286
rect 14760 2320 14860 2358
rect 14760 2286 14776 2320
rect 14844 2286 14860 2320
rect 14760 2270 14860 2286
rect 14918 2320 15018 2358
rect 14918 2286 14934 2320
rect 15002 2286 15018 2320
rect 14918 2270 15018 2286
rect 15076 2320 15176 2358
rect 15076 2286 15092 2320
rect 15160 2286 15176 2320
rect 15076 2270 15176 2286
rect 15234 2320 15334 2358
rect 15234 2286 15250 2320
rect 15318 2286 15334 2320
rect 15234 2270 15334 2286
rect 15392 2320 15492 2358
rect 15392 2286 15408 2320
rect 15476 2286 15492 2320
rect 15392 2270 15492 2286
rect 15550 2320 15650 2358
rect 15550 2286 15566 2320
rect 15634 2286 15650 2320
rect 15550 2270 15650 2286
rect 15708 2320 15808 2358
rect 15708 2286 15724 2320
rect 15792 2286 15808 2320
rect 15708 2270 15808 2286
rect 15866 2320 15966 2358
rect 15866 2286 15882 2320
rect 15950 2286 15966 2320
rect 15866 2270 15966 2286
rect 16024 2320 16124 2358
rect 16024 2286 16040 2320
rect 16108 2286 16124 2320
rect 16024 2270 16124 2286
rect 16182 2320 16282 2358
rect 16182 2286 16198 2320
rect 16266 2286 16282 2320
rect 16182 2270 16282 2286
rect 16340 2320 16440 2358
rect 16340 2286 16356 2320
rect 16424 2286 16440 2320
rect 16340 2270 16440 2286
rect 16498 2320 16598 2358
rect 16498 2286 16514 2320
rect 16582 2286 16598 2320
rect 16498 2270 16598 2286
rect 16656 2320 16756 2358
rect 16656 2286 16672 2320
rect 16740 2286 16756 2320
rect 16656 2270 16756 2286
rect 16814 2320 16914 2358
rect 16814 2286 16830 2320
rect 16898 2286 16914 2320
rect 16814 2270 16914 2286
rect 16972 2320 17072 2358
rect 16972 2286 16988 2320
rect 17056 2286 17072 2320
rect 16972 2270 17072 2286
rect 17130 2320 17230 2358
rect 17130 2286 17146 2320
rect 17214 2286 17230 2320
rect 17130 2270 17230 2286
rect 17288 2320 17388 2358
rect 17288 2286 17304 2320
rect 17372 2286 17388 2320
rect 17288 2270 17388 2286
rect 17446 2320 17546 2358
rect 17446 2286 17462 2320
rect 17530 2286 17546 2320
rect 17446 2270 17546 2286
rect 17604 2320 17704 2358
rect 17604 2286 17620 2320
rect 17688 2286 17704 2320
rect 17604 2270 17704 2286
rect 17762 2320 17862 2358
rect 17762 2286 17778 2320
rect 17846 2286 17862 2320
rect 17762 2270 17862 2286
rect 17920 2320 18020 2358
rect 17920 2286 17936 2320
rect 18004 2286 18020 2320
rect 17920 2270 18020 2286
rect 18078 2320 18178 2358
rect 18078 2286 18094 2320
rect 18162 2286 18178 2320
rect 18078 2270 18178 2286
rect 18236 2320 18336 2358
rect 18236 2286 18252 2320
rect 18320 2286 18336 2320
rect 18236 2270 18336 2286
rect 18394 2320 18494 2358
rect 18394 2286 18410 2320
rect 18478 2286 18494 2320
rect 18394 2270 18494 2286
rect 18552 2320 18652 2358
rect 18552 2286 18568 2320
rect 18636 2286 18652 2320
rect 18552 2270 18652 2286
rect 18710 2320 18810 2358
rect 18710 2286 18726 2320
rect 18794 2286 18810 2320
rect 18710 2270 18810 2286
rect 20428 8430 20528 8446
rect 20428 8396 20444 8430
rect 20512 8396 20528 8430
rect 20428 8358 20528 8396
rect 20586 8430 20686 8446
rect 20586 8396 20602 8430
rect 20670 8396 20686 8430
rect 20586 8358 20686 8396
rect 20744 8430 20844 8446
rect 20744 8396 20760 8430
rect 20828 8396 20844 8430
rect 20744 8358 20844 8396
rect 20902 8430 21002 8446
rect 20902 8396 20918 8430
rect 20986 8396 21002 8430
rect 20902 8358 21002 8396
rect 21060 8430 21160 8446
rect 21060 8396 21076 8430
rect 21144 8396 21160 8430
rect 21060 8358 21160 8396
rect 21218 8430 21318 8446
rect 21218 8396 21234 8430
rect 21302 8396 21318 8430
rect 21218 8358 21318 8396
rect 21376 8430 21476 8446
rect 21376 8396 21392 8430
rect 21460 8396 21476 8430
rect 21376 8358 21476 8396
rect 21534 8430 21634 8446
rect 21534 8396 21550 8430
rect 21618 8396 21634 8430
rect 21534 8358 21634 8396
rect 21692 8430 21792 8446
rect 21692 8396 21708 8430
rect 21776 8396 21792 8430
rect 21692 8358 21792 8396
rect 21850 8430 21950 8446
rect 21850 8396 21866 8430
rect 21934 8396 21950 8430
rect 21850 8358 21950 8396
rect 22008 8430 22108 8446
rect 22008 8396 22024 8430
rect 22092 8396 22108 8430
rect 22008 8358 22108 8396
rect 22166 8430 22266 8446
rect 22166 8396 22182 8430
rect 22250 8396 22266 8430
rect 22166 8358 22266 8396
rect 22324 8430 22424 8446
rect 22324 8396 22340 8430
rect 22408 8396 22424 8430
rect 22324 8358 22424 8396
rect 22482 8430 22582 8446
rect 22482 8396 22498 8430
rect 22566 8396 22582 8430
rect 22482 8358 22582 8396
rect 22640 8430 22740 8446
rect 22640 8396 22656 8430
rect 22724 8396 22740 8430
rect 22640 8358 22740 8396
rect 22798 8430 22898 8446
rect 22798 8396 22814 8430
rect 22882 8396 22898 8430
rect 22798 8358 22898 8396
rect 22956 8430 23056 8446
rect 22956 8396 22972 8430
rect 23040 8396 23056 8430
rect 22956 8358 23056 8396
rect 23114 8430 23214 8446
rect 23114 8396 23130 8430
rect 23198 8396 23214 8430
rect 23114 8358 23214 8396
rect 23272 8430 23372 8446
rect 23272 8396 23288 8430
rect 23356 8396 23372 8430
rect 23272 8358 23372 8396
rect 23430 8430 23530 8446
rect 23430 8396 23446 8430
rect 23514 8396 23530 8430
rect 23430 8358 23530 8396
rect 23588 8430 23688 8446
rect 23588 8396 23604 8430
rect 23672 8396 23688 8430
rect 23588 8358 23688 8396
rect 23746 8430 23846 8446
rect 23746 8396 23762 8430
rect 23830 8396 23846 8430
rect 23746 8358 23846 8396
rect 23904 8430 24004 8446
rect 23904 8396 23920 8430
rect 23988 8396 24004 8430
rect 23904 8358 24004 8396
rect 24062 8430 24162 8446
rect 24062 8396 24078 8430
rect 24146 8396 24162 8430
rect 24062 8358 24162 8396
rect 24220 8430 24320 8446
rect 24220 8396 24236 8430
rect 24304 8396 24320 8430
rect 24220 8358 24320 8396
rect 24378 8430 24478 8446
rect 24378 8396 24394 8430
rect 24462 8396 24478 8430
rect 24378 8358 24478 8396
rect 24536 8430 24636 8446
rect 24536 8396 24552 8430
rect 24620 8396 24636 8430
rect 24536 8358 24636 8396
rect 24694 8430 24794 8446
rect 24694 8396 24710 8430
rect 24778 8396 24794 8430
rect 24694 8358 24794 8396
rect 24852 8430 24952 8446
rect 24852 8396 24868 8430
rect 24936 8396 24952 8430
rect 24852 8358 24952 8396
rect 25010 8430 25110 8446
rect 25010 8396 25026 8430
rect 25094 8396 25110 8430
rect 25010 8358 25110 8396
rect 20428 2320 20528 2358
rect 20428 2286 20444 2320
rect 20512 2286 20528 2320
rect 20428 2270 20528 2286
rect 20586 2320 20686 2358
rect 20586 2286 20602 2320
rect 20670 2286 20686 2320
rect 20586 2270 20686 2286
rect 20744 2320 20844 2358
rect 20744 2286 20760 2320
rect 20828 2286 20844 2320
rect 20744 2270 20844 2286
rect 20902 2320 21002 2358
rect 20902 2286 20918 2320
rect 20986 2286 21002 2320
rect 20902 2270 21002 2286
rect 21060 2320 21160 2358
rect 21060 2286 21076 2320
rect 21144 2286 21160 2320
rect 21060 2270 21160 2286
rect 21218 2320 21318 2358
rect 21218 2286 21234 2320
rect 21302 2286 21318 2320
rect 21218 2270 21318 2286
rect 21376 2320 21476 2358
rect 21376 2286 21392 2320
rect 21460 2286 21476 2320
rect 21376 2270 21476 2286
rect 21534 2320 21634 2358
rect 21534 2286 21550 2320
rect 21618 2286 21634 2320
rect 21534 2270 21634 2286
rect 21692 2320 21792 2358
rect 21692 2286 21708 2320
rect 21776 2286 21792 2320
rect 21692 2270 21792 2286
rect 21850 2320 21950 2358
rect 21850 2286 21866 2320
rect 21934 2286 21950 2320
rect 21850 2270 21950 2286
rect 22008 2320 22108 2358
rect 22008 2286 22024 2320
rect 22092 2286 22108 2320
rect 22008 2270 22108 2286
rect 22166 2320 22266 2358
rect 22166 2286 22182 2320
rect 22250 2286 22266 2320
rect 22166 2270 22266 2286
rect 22324 2320 22424 2358
rect 22324 2286 22340 2320
rect 22408 2286 22424 2320
rect 22324 2270 22424 2286
rect 22482 2320 22582 2358
rect 22482 2286 22498 2320
rect 22566 2286 22582 2320
rect 22482 2270 22582 2286
rect 22640 2320 22740 2358
rect 22640 2286 22656 2320
rect 22724 2286 22740 2320
rect 22640 2270 22740 2286
rect 22798 2320 22898 2358
rect 22798 2286 22814 2320
rect 22882 2286 22898 2320
rect 22798 2270 22898 2286
rect 22956 2320 23056 2358
rect 22956 2286 22972 2320
rect 23040 2286 23056 2320
rect 22956 2270 23056 2286
rect 23114 2320 23214 2358
rect 23114 2286 23130 2320
rect 23198 2286 23214 2320
rect 23114 2270 23214 2286
rect 23272 2320 23372 2358
rect 23272 2286 23288 2320
rect 23356 2286 23372 2320
rect 23272 2270 23372 2286
rect 23430 2320 23530 2358
rect 23430 2286 23446 2320
rect 23514 2286 23530 2320
rect 23430 2270 23530 2286
rect 23588 2320 23688 2358
rect 23588 2286 23604 2320
rect 23672 2286 23688 2320
rect 23588 2270 23688 2286
rect 23746 2320 23846 2358
rect 23746 2286 23762 2320
rect 23830 2286 23846 2320
rect 23746 2270 23846 2286
rect 23904 2320 24004 2358
rect 23904 2286 23920 2320
rect 23988 2286 24004 2320
rect 23904 2270 24004 2286
rect 24062 2320 24162 2358
rect 24062 2286 24078 2320
rect 24146 2286 24162 2320
rect 24062 2270 24162 2286
rect 24220 2320 24320 2358
rect 24220 2286 24236 2320
rect 24304 2286 24320 2320
rect 24220 2270 24320 2286
rect 24378 2320 24478 2358
rect 24378 2286 24394 2320
rect 24462 2286 24478 2320
rect 24378 2270 24478 2286
rect 24536 2320 24636 2358
rect 24536 2286 24552 2320
rect 24620 2286 24636 2320
rect 24536 2270 24636 2286
rect 24694 2320 24794 2358
rect 24694 2286 24710 2320
rect 24778 2286 24794 2320
rect 24694 2270 24794 2286
rect 24852 2320 24952 2358
rect 24852 2286 24868 2320
rect 24936 2286 24952 2320
rect 24852 2270 24952 2286
rect 25010 2320 25110 2358
rect 25010 2286 25026 2320
rect 25094 2286 25110 2320
rect 25010 2270 25110 2286
<< polycont >>
rect -3218 40242 -3184 40276
rect -3218 38862 -3184 38896
rect 1544 45996 1612 46030
rect 1702 45996 1770 46030
rect 1860 45996 1928 46030
rect 2018 45996 2086 46030
rect 2176 45996 2244 46030
rect 2334 45996 2402 46030
rect 2492 45996 2560 46030
rect 2650 45996 2718 46030
rect 2808 45996 2876 46030
rect 2966 45996 3034 46030
rect 3124 45996 3192 46030
rect 3282 45996 3350 46030
rect 3440 45996 3508 46030
rect 3598 45996 3666 46030
rect 3756 45996 3824 46030
rect 3914 45996 3982 46030
rect 4072 45996 4140 46030
rect 4230 45996 4298 46030
rect 4388 45996 4456 46030
rect 4546 45996 4614 46030
rect 4704 45996 4772 46030
rect 4862 45996 4930 46030
rect 5020 45996 5088 46030
rect 5178 45996 5246 46030
rect 5336 45996 5404 46030
rect 5494 45996 5562 46030
rect 5652 45996 5720 46030
rect 5810 45996 5878 46030
rect 5968 45996 6036 46030
rect 6126 45996 6194 46030
rect 1544 39886 1612 39920
rect 1702 39886 1770 39920
rect 1860 39886 1928 39920
rect 2018 39886 2086 39920
rect 2176 39886 2244 39920
rect 2334 39886 2402 39920
rect 2492 39886 2560 39920
rect 2650 39886 2718 39920
rect 2808 39886 2876 39920
rect 2966 39886 3034 39920
rect 3124 39886 3192 39920
rect 3282 39886 3350 39920
rect 3440 39886 3508 39920
rect 3598 39886 3666 39920
rect 3756 39886 3824 39920
rect 3914 39886 3982 39920
rect 4072 39886 4140 39920
rect 4230 39886 4298 39920
rect 4388 39886 4456 39920
rect 4546 39886 4614 39920
rect 4704 39886 4772 39920
rect 4862 39886 4930 39920
rect 5020 39886 5088 39920
rect 5178 39886 5246 39920
rect 5336 39886 5404 39920
rect 5494 39886 5562 39920
rect 5652 39886 5720 39920
rect 5810 39886 5878 39920
rect 5968 39886 6036 39920
rect 6126 39886 6194 39920
rect 7844 45996 7912 46030
rect 8002 45996 8070 46030
rect 8160 45996 8228 46030
rect 8318 45996 8386 46030
rect 8476 45996 8544 46030
rect 8634 45996 8702 46030
rect 8792 45996 8860 46030
rect 8950 45996 9018 46030
rect 9108 45996 9176 46030
rect 9266 45996 9334 46030
rect 9424 45996 9492 46030
rect 9582 45996 9650 46030
rect 9740 45996 9808 46030
rect 9898 45996 9966 46030
rect 10056 45996 10124 46030
rect 10214 45996 10282 46030
rect 10372 45996 10440 46030
rect 10530 45996 10598 46030
rect 10688 45996 10756 46030
rect 10846 45996 10914 46030
rect 11004 45996 11072 46030
rect 11162 45996 11230 46030
rect 11320 45996 11388 46030
rect 11478 45996 11546 46030
rect 11636 45996 11704 46030
rect 11794 45996 11862 46030
rect 11952 45996 12020 46030
rect 12110 45996 12178 46030
rect 12268 45996 12336 46030
rect 12426 45996 12494 46030
rect 7844 39886 7912 39920
rect 8002 39886 8070 39920
rect 8160 39886 8228 39920
rect 8318 39886 8386 39920
rect 8476 39886 8544 39920
rect 8634 39886 8702 39920
rect 8792 39886 8860 39920
rect 8950 39886 9018 39920
rect 9108 39886 9176 39920
rect 9266 39886 9334 39920
rect 9424 39886 9492 39920
rect 9582 39886 9650 39920
rect 9740 39886 9808 39920
rect 9898 39886 9966 39920
rect 10056 39886 10124 39920
rect 10214 39886 10282 39920
rect 10372 39886 10440 39920
rect 10530 39886 10598 39920
rect 10688 39886 10756 39920
rect 10846 39886 10914 39920
rect 11004 39886 11072 39920
rect 11162 39886 11230 39920
rect 11320 39886 11388 39920
rect 11478 39886 11546 39920
rect 11636 39886 11704 39920
rect 11794 39886 11862 39920
rect 11952 39886 12020 39920
rect 12110 39886 12178 39920
rect 12268 39886 12336 39920
rect 12426 39886 12494 39920
rect 14144 45996 14212 46030
rect 14302 45996 14370 46030
rect 14460 45996 14528 46030
rect 14618 45996 14686 46030
rect 14776 45996 14844 46030
rect 14934 45996 15002 46030
rect 15092 45996 15160 46030
rect 15250 45996 15318 46030
rect 15408 45996 15476 46030
rect 15566 45996 15634 46030
rect 15724 45996 15792 46030
rect 15882 45996 15950 46030
rect 16040 45996 16108 46030
rect 16198 45996 16266 46030
rect 16356 45996 16424 46030
rect 16514 45996 16582 46030
rect 16672 45996 16740 46030
rect 16830 45996 16898 46030
rect 16988 45996 17056 46030
rect 17146 45996 17214 46030
rect 17304 45996 17372 46030
rect 17462 45996 17530 46030
rect 17620 45996 17688 46030
rect 17778 45996 17846 46030
rect 17936 45996 18004 46030
rect 18094 45996 18162 46030
rect 18252 45996 18320 46030
rect 18410 45996 18478 46030
rect 18568 45996 18636 46030
rect 18726 45996 18794 46030
rect 14144 39886 14212 39920
rect 14302 39886 14370 39920
rect 14460 39886 14528 39920
rect 14618 39886 14686 39920
rect 14776 39886 14844 39920
rect 14934 39886 15002 39920
rect 15092 39886 15160 39920
rect 15250 39886 15318 39920
rect 15408 39886 15476 39920
rect 15566 39886 15634 39920
rect 15724 39886 15792 39920
rect 15882 39886 15950 39920
rect 16040 39886 16108 39920
rect 16198 39886 16266 39920
rect 16356 39886 16424 39920
rect 16514 39886 16582 39920
rect 16672 39886 16740 39920
rect 16830 39886 16898 39920
rect 16988 39886 17056 39920
rect 17146 39886 17214 39920
rect 17304 39886 17372 39920
rect 17462 39886 17530 39920
rect 17620 39886 17688 39920
rect 17778 39886 17846 39920
rect 17936 39886 18004 39920
rect 18094 39886 18162 39920
rect 18252 39886 18320 39920
rect 18410 39886 18478 39920
rect 18568 39886 18636 39920
rect 18726 39886 18794 39920
rect 20444 45996 20512 46030
rect 20602 45996 20670 46030
rect 20760 45996 20828 46030
rect 20918 45996 20986 46030
rect 21076 45996 21144 46030
rect 21234 45996 21302 46030
rect 21392 45996 21460 46030
rect 21550 45996 21618 46030
rect 21708 45996 21776 46030
rect 21866 45996 21934 46030
rect 22024 45996 22092 46030
rect 22182 45996 22250 46030
rect 22340 45996 22408 46030
rect 22498 45996 22566 46030
rect 22656 45996 22724 46030
rect 22814 45996 22882 46030
rect 22972 45996 23040 46030
rect 23130 45996 23198 46030
rect 23288 45996 23356 46030
rect 23446 45996 23514 46030
rect 23604 45996 23672 46030
rect 23762 45996 23830 46030
rect 23920 45996 23988 46030
rect 24078 45996 24146 46030
rect 24236 45996 24304 46030
rect 24394 45996 24462 46030
rect 24552 45996 24620 46030
rect 24710 45996 24778 46030
rect 24868 45996 24936 46030
rect 25026 45996 25094 46030
rect 20444 39886 20512 39920
rect 20602 39886 20670 39920
rect 20760 39886 20828 39920
rect 20918 39886 20986 39920
rect 21076 39886 21144 39920
rect 21234 39886 21302 39920
rect 21392 39886 21460 39920
rect 21550 39886 21618 39920
rect 21708 39886 21776 39920
rect 21866 39886 21934 39920
rect 22024 39886 22092 39920
rect 22182 39886 22250 39920
rect 22340 39886 22408 39920
rect 22498 39886 22566 39920
rect 22656 39886 22724 39920
rect 22814 39886 22882 39920
rect 22972 39886 23040 39920
rect 23130 39886 23198 39920
rect 23288 39886 23356 39920
rect 23446 39886 23514 39920
rect 23604 39886 23672 39920
rect 23762 39886 23830 39920
rect 23920 39886 23988 39920
rect 24078 39886 24146 39920
rect 24236 39886 24304 39920
rect 24394 39886 24462 39920
rect 24552 39886 24620 39920
rect 24710 39886 24778 39920
rect 24868 39886 24936 39920
rect 25026 39886 25094 39920
rect 1544 38996 1612 39030
rect 1702 38996 1770 39030
rect 1860 38996 1928 39030
rect 2018 38996 2086 39030
rect 2176 38996 2244 39030
rect 2334 38996 2402 39030
rect 2492 38996 2560 39030
rect 2650 38996 2718 39030
rect 2808 38996 2876 39030
rect 2966 38996 3034 39030
rect 3124 38996 3192 39030
rect 3282 38996 3350 39030
rect 3440 38996 3508 39030
rect 3598 38996 3666 39030
rect 3756 38996 3824 39030
rect 3914 38996 3982 39030
rect 4072 38996 4140 39030
rect 4230 38996 4298 39030
rect 4388 38996 4456 39030
rect 4546 38996 4614 39030
rect 4704 38996 4772 39030
rect 4862 38996 4930 39030
rect 5020 38996 5088 39030
rect 5178 38996 5246 39030
rect 5336 38996 5404 39030
rect 5494 38996 5562 39030
rect 5652 38996 5720 39030
rect 5810 38996 5878 39030
rect 5968 38996 6036 39030
rect 6126 38996 6194 39030
rect 1544 32886 1612 32920
rect 1702 32886 1770 32920
rect 1860 32886 1928 32920
rect 2018 32886 2086 32920
rect 2176 32886 2244 32920
rect 2334 32886 2402 32920
rect 2492 32886 2560 32920
rect 2650 32886 2718 32920
rect 2808 32886 2876 32920
rect 2966 32886 3034 32920
rect 3124 32886 3192 32920
rect 3282 32886 3350 32920
rect 3440 32886 3508 32920
rect 3598 32886 3666 32920
rect 3756 32886 3824 32920
rect 3914 32886 3982 32920
rect 4072 32886 4140 32920
rect 4230 32886 4298 32920
rect 4388 32886 4456 32920
rect 4546 32886 4614 32920
rect 4704 32886 4772 32920
rect 4862 32886 4930 32920
rect 5020 32886 5088 32920
rect 5178 32886 5246 32920
rect 5336 32886 5404 32920
rect 5494 32886 5562 32920
rect 5652 32886 5720 32920
rect 5810 32886 5878 32920
rect 5968 32886 6036 32920
rect 6126 32886 6194 32920
rect 7844 38996 7912 39030
rect 8002 38996 8070 39030
rect 8160 38996 8228 39030
rect 8318 38996 8386 39030
rect 8476 38996 8544 39030
rect 8634 38996 8702 39030
rect 8792 38996 8860 39030
rect 8950 38996 9018 39030
rect 9108 38996 9176 39030
rect 9266 38996 9334 39030
rect 9424 38996 9492 39030
rect 9582 38996 9650 39030
rect 9740 38996 9808 39030
rect 9898 38996 9966 39030
rect 10056 38996 10124 39030
rect 10214 38996 10282 39030
rect 10372 38996 10440 39030
rect 10530 38996 10598 39030
rect 10688 38996 10756 39030
rect 10846 38996 10914 39030
rect 11004 38996 11072 39030
rect 11162 38996 11230 39030
rect 11320 38996 11388 39030
rect 11478 38996 11546 39030
rect 11636 38996 11704 39030
rect 11794 38996 11862 39030
rect 11952 38996 12020 39030
rect 12110 38996 12178 39030
rect 12268 38996 12336 39030
rect 12426 38996 12494 39030
rect 7844 32886 7912 32920
rect 8002 32886 8070 32920
rect 8160 32886 8228 32920
rect 8318 32886 8386 32920
rect 8476 32886 8544 32920
rect 8634 32886 8702 32920
rect 8792 32886 8860 32920
rect 8950 32886 9018 32920
rect 9108 32886 9176 32920
rect 9266 32886 9334 32920
rect 9424 32886 9492 32920
rect 9582 32886 9650 32920
rect 9740 32886 9808 32920
rect 9898 32886 9966 32920
rect 10056 32886 10124 32920
rect 10214 32886 10282 32920
rect 10372 32886 10440 32920
rect 10530 32886 10598 32920
rect 10688 32886 10756 32920
rect 10846 32886 10914 32920
rect 11004 32886 11072 32920
rect 11162 32886 11230 32920
rect 11320 32886 11388 32920
rect 11478 32886 11546 32920
rect 11636 32886 11704 32920
rect 11794 32886 11862 32920
rect 11952 32886 12020 32920
rect 12110 32886 12178 32920
rect 12268 32886 12336 32920
rect 12426 32886 12494 32920
rect 14144 38996 14212 39030
rect 14302 38996 14370 39030
rect 14460 38996 14528 39030
rect 14618 38996 14686 39030
rect 14776 38996 14844 39030
rect 14934 38996 15002 39030
rect 15092 38996 15160 39030
rect 15250 38996 15318 39030
rect 15408 38996 15476 39030
rect 15566 38996 15634 39030
rect 15724 38996 15792 39030
rect 15882 38996 15950 39030
rect 16040 38996 16108 39030
rect 16198 38996 16266 39030
rect 16356 38996 16424 39030
rect 16514 38996 16582 39030
rect 16672 38996 16740 39030
rect 16830 38996 16898 39030
rect 16988 38996 17056 39030
rect 17146 38996 17214 39030
rect 17304 38996 17372 39030
rect 17462 38996 17530 39030
rect 17620 38996 17688 39030
rect 17778 38996 17846 39030
rect 17936 38996 18004 39030
rect 18094 38996 18162 39030
rect 18252 38996 18320 39030
rect 18410 38996 18478 39030
rect 18568 38996 18636 39030
rect 18726 38996 18794 39030
rect 14144 32886 14212 32920
rect 14302 32886 14370 32920
rect 14460 32886 14528 32920
rect 14618 32886 14686 32920
rect 14776 32886 14844 32920
rect 14934 32886 15002 32920
rect 15092 32886 15160 32920
rect 15250 32886 15318 32920
rect 15408 32886 15476 32920
rect 15566 32886 15634 32920
rect 15724 32886 15792 32920
rect 15882 32886 15950 32920
rect 16040 32886 16108 32920
rect 16198 32886 16266 32920
rect 16356 32886 16424 32920
rect 16514 32886 16582 32920
rect 16672 32886 16740 32920
rect 16830 32886 16898 32920
rect 16988 32886 17056 32920
rect 17146 32886 17214 32920
rect 17304 32886 17372 32920
rect 17462 32886 17530 32920
rect 17620 32886 17688 32920
rect 17778 32886 17846 32920
rect 17936 32886 18004 32920
rect 18094 32886 18162 32920
rect 18252 32886 18320 32920
rect 18410 32886 18478 32920
rect 18568 32886 18636 32920
rect 18726 32886 18794 32920
rect 20444 38996 20512 39030
rect 20602 38996 20670 39030
rect 20760 38996 20828 39030
rect 20918 38996 20986 39030
rect 21076 38996 21144 39030
rect 21234 38996 21302 39030
rect 21392 38996 21460 39030
rect 21550 38996 21618 39030
rect 21708 38996 21776 39030
rect 21866 38996 21934 39030
rect 22024 38996 22092 39030
rect 22182 38996 22250 39030
rect 22340 38996 22408 39030
rect 22498 38996 22566 39030
rect 22656 38996 22724 39030
rect 22814 38996 22882 39030
rect 22972 38996 23040 39030
rect 23130 38996 23198 39030
rect 23288 38996 23356 39030
rect 23446 38996 23514 39030
rect 23604 38996 23672 39030
rect 23762 38996 23830 39030
rect 23920 38996 23988 39030
rect 24078 38996 24146 39030
rect 24236 38996 24304 39030
rect 24394 38996 24462 39030
rect 24552 38996 24620 39030
rect 24710 38996 24778 39030
rect 24868 38996 24936 39030
rect 25026 38996 25094 39030
rect 20444 32886 20512 32920
rect 20602 32886 20670 32920
rect 20760 32886 20828 32920
rect 20918 32886 20986 32920
rect 21076 32886 21144 32920
rect 21234 32886 21302 32920
rect 21392 32886 21460 32920
rect 21550 32886 21618 32920
rect 21708 32886 21776 32920
rect 21866 32886 21934 32920
rect 22024 32886 22092 32920
rect 22182 32886 22250 32920
rect 22340 32886 22408 32920
rect 22498 32886 22566 32920
rect 22656 32886 22724 32920
rect 22814 32886 22882 32920
rect 22972 32886 23040 32920
rect 23130 32886 23198 32920
rect 23288 32886 23356 32920
rect 23446 32886 23514 32920
rect 23604 32886 23672 32920
rect 23762 32886 23830 32920
rect 23920 32886 23988 32920
rect 24078 32886 24146 32920
rect 24236 32886 24304 32920
rect 24394 32886 24462 32920
rect 24552 32886 24620 32920
rect 24710 32886 24778 32920
rect 24868 32886 24936 32920
rect 25026 32886 25094 32920
rect 29984 40242 30018 40276
rect 29984 38862 30018 38896
rect -4218 27042 -4184 27076
rect -4218 25662 -4184 25696
rect 1544 30696 1612 30730
rect 1702 30696 1770 30730
rect 1860 30696 1928 30730
rect 2018 30696 2086 30730
rect 2176 30696 2244 30730
rect 2334 30696 2402 30730
rect 2492 30696 2560 30730
rect 2650 30696 2718 30730
rect 2808 30696 2876 30730
rect 2966 30696 3034 30730
rect 3124 30696 3192 30730
rect 3282 30696 3350 30730
rect 3440 30696 3508 30730
rect 3598 30696 3666 30730
rect 3756 30696 3824 30730
rect 3914 30696 3982 30730
rect 4072 30696 4140 30730
rect 4230 30696 4298 30730
rect 4388 30696 4456 30730
rect 4546 30696 4614 30730
rect 4704 30696 4772 30730
rect 4862 30696 4930 30730
rect 5020 30696 5088 30730
rect 5178 30696 5246 30730
rect 5336 30696 5404 30730
rect 5494 30696 5562 30730
rect 5652 30696 5720 30730
rect 5810 30696 5878 30730
rect 5968 30696 6036 30730
rect 6126 30696 6194 30730
rect 1544 24586 1612 24620
rect 1702 24586 1770 24620
rect 1860 24586 1928 24620
rect 2018 24586 2086 24620
rect 2176 24586 2244 24620
rect 2334 24586 2402 24620
rect 2492 24586 2560 24620
rect 2650 24586 2718 24620
rect 2808 24586 2876 24620
rect 2966 24586 3034 24620
rect 3124 24586 3192 24620
rect 3282 24586 3350 24620
rect 3440 24586 3508 24620
rect 3598 24586 3666 24620
rect 3756 24586 3824 24620
rect 3914 24586 3982 24620
rect 4072 24586 4140 24620
rect 4230 24586 4298 24620
rect 4388 24586 4456 24620
rect 4546 24586 4614 24620
rect 4704 24586 4772 24620
rect 4862 24586 4930 24620
rect 5020 24586 5088 24620
rect 5178 24586 5246 24620
rect 5336 24586 5404 24620
rect 5494 24586 5562 24620
rect 5652 24586 5720 24620
rect 5810 24586 5878 24620
rect 5968 24586 6036 24620
rect 6126 24586 6194 24620
rect 7844 30696 7912 30730
rect 8002 30696 8070 30730
rect 8160 30696 8228 30730
rect 8318 30696 8386 30730
rect 8476 30696 8544 30730
rect 8634 30696 8702 30730
rect 8792 30696 8860 30730
rect 8950 30696 9018 30730
rect 9108 30696 9176 30730
rect 9266 30696 9334 30730
rect 9424 30696 9492 30730
rect 9582 30696 9650 30730
rect 9740 30696 9808 30730
rect 9898 30696 9966 30730
rect 10056 30696 10124 30730
rect 10214 30696 10282 30730
rect 10372 30696 10440 30730
rect 10530 30696 10598 30730
rect 10688 30696 10756 30730
rect 10846 30696 10914 30730
rect 11004 30696 11072 30730
rect 11162 30696 11230 30730
rect 11320 30696 11388 30730
rect 11478 30696 11546 30730
rect 11636 30696 11704 30730
rect 11794 30696 11862 30730
rect 11952 30696 12020 30730
rect 12110 30696 12178 30730
rect 12268 30696 12336 30730
rect 12426 30696 12494 30730
rect 7844 24586 7912 24620
rect 8002 24586 8070 24620
rect 8160 24586 8228 24620
rect 8318 24586 8386 24620
rect 8476 24586 8544 24620
rect 8634 24586 8702 24620
rect 8792 24586 8860 24620
rect 8950 24586 9018 24620
rect 9108 24586 9176 24620
rect 9266 24586 9334 24620
rect 9424 24586 9492 24620
rect 9582 24586 9650 24620
rect 9740 24586 9808 24620
rect 9898 24586 9966 24620
rect 10056 24586 10124 24620
rect 10214 24586 10282 24620
rect 10372 24586 10440 24620
rect 10530 24586 10598 24620
rect 10688 24586 10756 24620
rect 10846 24586 10914 24620
rect 11004 24586 11072 24620
rect 11162 24586 11230 24620
rect 11320 24586 11388 24620
rect 11478 24586 11546 24620
rect 11636 24586 11704 24620
rect 11794 24586 11862 24620
rect 11952 24586 12020 24620
rect 12110 24586 12178 24620
rect 12268 24586 12336 24620
rect 12426 24586 12494 24620
rect 14144 30696 14212 30730
rect 14302 30696 14370 30730
rect 14460 30696 14528 30730
rect 14618 30696 14686 30730
rect 14776 30696 14844 30730
rect 14934 30696 15002 30730
rect 15092 30696 15160 30730
rect 15250 30696 15318 30730
rect 15408 30696 15476 30730
rect 15566 30696 15634 30730
rect 15724 30696 15792 30730
rect 15882 30696 15950 30730
rect 16040 30696 16108 30730
rect 16198 30696 16266 30730
rect 16356 30696 16424 30730
rect 16514 30696 16582 30730
rect 16672 30696 16740 30730
rect 16830 30696 16898 30730
rect 16988 30696 17056 30730
rect 17146 30696 17214 30730
rect 17304 30696 17372 30730
rect 17462 30696 17530 30730
rect 17620 30696 17688 30730
rect 17778 30696 17846 30730
rect 17936 30696 18004 30730
rect 18094 30696 18162 30730
rect 18252 30696 18320 30730
rect 18410 30696 18478 30730
rect 18568 30696 18636 30730
rect 18726 30696 18794 30730
rect 14144 24586 14212 24620
rect 14302 24586 14370 24620
rect 14460 24586 14528 24620
rect 14618 24586 14686 24620
rect 14776 24586 14844 24620
rect 14934 24586 15002 24620
rect 15092 24586 15160 24620
rect 15250 24586 15318 24620
rect 15408 24586 15476 24620
rect 15566 24586 15634 24620
rect 15724 24586 15792 24620
rect 15882 24586 15950 24620
rect 16040 24586 16108 24620
rect 16198 24586 16266 24620
rect 16356 24586 16424 24620
rect 16514 24586 16582 24620
rect 16672 24586 16740 24620
rect 16830 24586 16898 24620
rect 16988 24586 17056 24620
rect 17146 24586 17214 24620
rect 17304 24586 17372 24620
rect 17462 24586 17530 24620
rect 17620 24586 17688 24620
rect 17778 24586 17846 24620
rect 17936 24586 18004 24620
rect 18094 24586 18162 24620
rect 18252 24586 18320 24620
rect 18410 24586 18478 24620
rect 18568 24586 18636 24620
rect 18726 24586 18794 24620
rect 20444 30696 20512 30730
rect 20602 30696 20670 30730
rect 20760 30696 20828 30730
rect 20918 30696 20986 30730
rect 21076 30696 21144 30730
rect 21234 30696 21302 30730
rect 21392 30696 21460 30730
rect 21550 30696 21618 30730
rect 21708 30696 21776 30730
rect 21866 30696 21934 30730
rect 22024 30696 22092 30730
rect 22182 30696 22250 30730
rect 22340 30696 22408 30730
rect 22498 30696 22566 30730
rect 22656 30696 22724 30730
rect 22814 30696 22882 30730
rect 22972 30696 23040 30730
rect 23130 30696 23198 30730
rect 23288 30696 23356 30730
rect 23446 30696 23514 30730
rect 23604 30696 23672 30730
rect 23762 30696 23830 30730
rect 23920 30696 23988 30730
rect 24078 30696 24146 30730
rect 24236 30696 24304 30730
rect 24394 30696 24462 30730
rect 24552 30696 24620 30730
rect 24710 30696 24778 30730
rect 24868 30696 24936 30730
rect 25026 30696 25094 30730
rect 20444 24586 20512 24620
rect 20602 24586 20670 24620
rect 20760 24586 20828 24620
rect 20918 24586 20986 24620
rect 21076 24586 21144 24620
rect 21234 24586 21302 24620
rect 21392 24586 21460 24620
rect 21550 24586 21618 24620
rect 21708 24586 21776 24620
rect 21866 24586 21934 24620
rect 22024 24586 22092 24620
rect 22182 24586 22250 24620
rect 22340 24586 22408 24620
rect 22498 24586 22566 24620
rect 22656 24586 22724 24620
rect 22814 24586 22882 24620
rect 22972 24586 23040 24620
rect 23130 24586 23198 24620
rect 23288 24586 23356 24620
rect 23446 24586 23514 24620
rect 23604 24586 23672 24620
rect 23762 24586 23830 24620
rect 23920 24586 23988 24620
rect 24078 24586 24146 24620
rect 24236 24586 24304 24620
rect 24394 24586 24462 24620
rect 24552 24586 24620 24620
rect 24710 24586 24778 24620
rect 24868 24586 24936 24620
rect 25026 24586 25094 24620
rect 30984 27042 31018 27076
rect 30984 25662 31018 25696
rect 1544 23696 1612 23730
rect 1702 23696 1770 23730
rect 1860 23696 1928 23730
rect 2018 23696 2086 23730
rect 2176 23696 2244 23730
rect 2334 23696 2402 23730
rect 2492 23696 2560 23730
rect 2650 23696 2718 23730
rect 2808 23696 2876 23730
rect 2966 23696 3034 23730
rect 3124 23696 3192 23730
rect 3282 23696 3350 23730
rect 3440 23696 3508 23730
rect 3598 23696 3666 23730
rect 3756 23696 3824 23730
rect 3914 23696 3982 23730
rect 4072 23696 4140 23730
rect 4230 23696 4298 23730
rect 4388 23696 4456 23730
rect 4546 23696 4614 23730
rect 4704 23696 4772 23730
rect 4862 23696 4930 23730
rect 5020 23696 5088 23730
rect 5178 23696 5246 23730
rect 5336 23696 5404 23730
rect 5494 23696 5562 23730
rect 5652 23696 5720 23730
rect 5810 23696 5878 23730
rect 5968 23696 6036 23730
rect 6126 23696 6194 23730
rect 1544 17586 1612 17620
rect 1702 17586 1770 17620
rect 1860 17586 1928 17620
rect 2018 17586 2086 17620
rect 2176 17586 2244 17620
rect 2334 17586 2402 17620
rect 2492 17586 2560 17620
rect 2650 17586 2718 17620
rect 2808 17586 2876 17620
rect 2966 17586 3034 17620
rect 3124 17586 3192 17620
rect 3282 17586 3350 17620
rect 3440 17586 3508 17620
rect 3598 17586 3666 17620
rect 3756 17586 3824 17620
rect 3914 17586 3982 17620
rect 4072 17586 4140 17620
rect 4230 17586 4298 17620
rect 4388 17586 4456 17620
rect 4546 17586 4614 17620
rect 4704 17586 4772 17620
rect 4862 17586 4930 17620
rect 5020 17586 5088 17620
rect 5178 17586 5246 17620
rect 5336 17586 5404 17620
rect 5494 17586 5562 17620
rect 5652 17586 5720 17620
rect 5810 17586 5878 17620
rect 5968 17586 6036 17620
rect 6126 17586 6194 17620
rect 7844 23696 7912 23730
rect 8002 23696 8070 23730
rect 8160 23696 8228 23730
rect 8318 23696 8386 23730
rect 8476 23696 8544 23730
rect 8634 23696 8702 23730
rect 8792 23696 8860 23730
rect 8950 23696 9018 23730
rect 9108 23696 9176 23730
rect 9266 23696 9334 23730
rect 9424 23696 9492 23730
rect 9582 23696 9650 23730
rect 9740 23696 9808 23730
rect 9898 23696 9966 23730
rect 10056 23696 10124 23730
rect 10214 23696 10282 23730
rect 10372 23696 10440 23730
rect 10530 23696 10598 23730
rect 10688 23696 10756 23730
rect 10846 23696 10914 23730
rect 11004 23696 11072 23730
rect 11162 23696 11230 23730
rect 11320 23696 11388 23730
rect 11478 23696 11546 23730
rect 11636 23696 11704 23730
rect 11794 23696 11862 23730
rect 11952 23696 12020 23730
rect 12110 23696 12178 23730
rect 12268 23696 12336 23730
rect 12426 23696 12494 23730
rect 7844 17586 7912 17620
rect 8002 17586 8070 17620
rect 8160 17586 8228 17620
rect 8318 17586 8386 17620
rect 8476 17586 8544 17620
rect 8634 17586 8702 17620
rect 8792 17586 8860 17620
rect 8950 17586 9018 17620
rect 9108 17586 9176 17620
rect 9266 17586 9334 17620
rect 9424 17586 9492 17620
rect 9582 17586 9650 17620
rect 9740 17586 9808 17620
rect 9898 17586 9966 17620
rect 10056 17586 10124 17620
rect 10214 17586 10282 17620
rect 10372 17586 10440 17620
rect 10530 17586 10598 17620
rect 10688 17586 10756 17620
rect 10846 17586 10914 17620
rect 11004 17586 11072 17620
rect 11162 17586 11230 17620
rect 11320 17586 11388 17620
rect 11478 17586 11546 17620
rect 11636 17586 11704 17620
rect 11794 17586 11862 17620
rect 11952 17586 12020 17620
rect 12110 17586 12178 17620
rect 12268 17586 12336 17620
rect 12426 17586 12494 17620
rect 14144 23696 14212 23730
rect 14302 23696 14370 23730
rect 14460 23696 14528 23730
rect 14618 23696 14686 23730
rect 14776 23696 14844 23730
rect 14934 23696 15002 23730
rect 15092 23696 15160 23730
rect 15250 23696 15318 23730
rect 15408 23696 15476 23730
rect 15566 23696 15634 23730
rect 15724 23696 15792 23730
rect 15882 23696 15950 23730
rect 16040 23696 16108 23730
rect 16198 23696 16266 23730
rect 16356 23696 16424 23730
rect 16514 23696 16582 23730
rect 16672 23696 16740 23730
rect 16830 23696 16898 23730
rect 16988 23696 17056 23730
rect 17146 23696 17214 23730
rect 17304 23696 17372 23730
rect 17462 23696 17530 23730
rect 17620 23696 17688 23730
rect 17778 23696 17846 23730
rect 17936 23696 18004 23730
rect 18094 23696 18162 23730
rect 18252 23696 18320 23730
rect 18410 23696 18478 23730
rect 18568 23696 18636 23730
rect 18726 23696 18794 23730
rect 14144 17586 14212 17620
rect 14302 17586 14370 17620
rect 14460 17586 14528 17620
rect 14618 17586 14686 17620
rect 14776 17586 14844 17620
rect 14934 17586 15002 17620
rect 15092 17586 15160 17620
rect 15250 17586 15318 17620
rect 15408 17586 15476 17620
rect 15566 17586 15634 17620
rect 15724 17586 15792 17620
rect 15882 17586 15950 17620
rect 16040 17586 16108 17620
rect 16198 17586 16266 17620
rect 16356 17586 16424 17620
rect 16514 17586 16582 17620
rect 16672 17586 16740 17620
rect 16830 17586 16898 17620
rect 16988 17586 17056 17620
rect 17146 17586 17214 17620
rect 17304 17586 17372 17620
rect 17462 17586 17530 17620
rect 17620 17586 17688 17620
rect 17778 17586 17846 17620
rect 17936 17586 18004 17620
rect 18094 17586 18162 17620
rect 18252 17586 18320 17620
rect 18410 17586 18478 17620
rect 18568 17586 18636 17620
rect 18726 17586 18794 17620
rect 20444 23696 20512 23730
rect 20602 23696 20670 23730
rect 20760 23696 20828 23730
rect 20918 23696 20986 23730
rect 21076 23696 21144 23730
rect 21234 23696 21302 23730
rect 21392 23696 21460 23730
rect 21550 23696 21618 23730
rect 21708 23696 21776 23730
rect 21866 23696 21934 23730
rect 22024 23696 22092 23730
rect 22182 23696 22250 23730
rect 22340 23696 22408 23730
rect 22498 23696 22566 23730
rect 22656 23696 22724 23730
rect 22814 23696 22882 23730
rect 22972 23696 23040 23730
rect 23130 23696 23198 23730
rect 23288 23696 23356 23730
rect 23446 23696 23514 23730
rect 23604 23696 23672 23730
rect 23762 23696 23830 23730
rect 23920 23696 23988 23730
rect 24078 23696 24146 23730
rect 24236 23696 24304 23730
rect 24394 23696 24462 23730
rect 24552 23696 24620 23730
rect 24710 23696 24778 23730
rect 24868 23696 24936 23730
rect 25026 23696 25094 23730
rect 20444 17586 20512 17620
rect 20602 17586 20670 17620
rect 20760 17586 20828 17620
rect 20918 17586 20986 17620
rect 21076 17586 21144 17620
rect 21234 17586 21302 17620
rect 21392 17586 21460 17620
rect 21550 17586 21618 17620
rect 21708 17586 21776 17620
rect 21866 17586 21934 17620
rect 22024 17586 22092 17620
rect 22182 17586 22250 17620
rect 22340 17586 22408 17620
rect 22498 17586 22566 17620
rect 22656 17586 22724 17620
rect 22814 17586 22882 17620
rect 22972 17586 23040 17620
rect 23130 17586 23198 17620
rect 23288 17586 23356 17620
rect 23446 17586 23514 17620
rect 23604 17586 23672 17620
rect 23762 17586 23830 17620
rect 23920 17586 23988 17620
rect 24078 17586 24146 17620
rect 24236 17586 24304 17620
rect 24394 17586 24462 17620
rect 24552 17586 24620 17620
rect 24710 17586 24778 17620
rect 24868 17586 24936 17620
rect 25026 17586 25094 17620
rect 1544 15396 1612 15430
rect 1702 15396 1770 15430
rect 1860 15396 1928 15430
rect 2018 15396 2086 15430
rect 2176 15396 2244 15430
rect 2334 15396 2402 15430
rect 2492 15396 2560 15430
rect 2650 15396 2718 15430
rect 2808 15396 2876 15430
rect 2966 15396 3034 15430
rect 3124 15396 3192 15430
rect 3282 15396 3350 15430
rect 3440 15396 3508 15430
rect 3598 15396 3666 15430
rect 3756 15396 3824 15430
rect 3914 15396 3982 15430
rect 4072 15396 4140 15430
rect 4230 15396 4298 15430
rect 4388 15396 4456 15430
rect 4546 15396 4614 15430
rect 4704 15396 4772 15430
rect 4862 15396 4930 15430
rect 5020 15396 5088 15430
rect 5178 15396 5246 15430
rect 5336 15396 5404 15430
rect 5494 15396 5562 15430
rect 5652 15396 5720 15430
rect 5810 15396 5878 15430
rect 5968 15396 6036 15430
rect 6126 15396 6194 15430
rect 1544 9286 1612 9320
rect 1702 9286 1770 9320
rect 1860 9286 1928 9320
rect 2018 9286 2086 9320
rect 2176 9286 2244 9320
rect 2334 9286 2402 9320
rect 2492 9286 2560 9320
rect 2650 9286 2718 9320
rect 2808 9286 2876 9320
rect 2966 9286 3034 9320
rect 3124 9286 3192 9320
rect 3282 9286 3350 9320
rect 3440 9286 3508 9320
rect 3598 9286 3666 9320
rect 3756 9286 3824 9320
rect 3914 9286 3982 9320
rect 4072 9286 4140 9320
rect 4230 9286 4298 9320
rect 4388 9286 4456 9320
rect 4546 9286 4614 9320
rect 4704 9286 4772 9320
rect 4862 9286 4930 9320
rect 5020 9286 5088 9320
rect 5178 9286 5246 9320
rect 5336 9286 5404 9320
rect 5494 9286 5562 9320
rect 5652 9286 5720 9320
rect 5810 9286 5878 9320
rect 5968 9286 6036 9320
rect 6126 9286 6194 9320
rect 7844 15396 7912 15430
rect 8002 15396 8070 15430
rect 8160 15396 8228 15430
rect 8318 15396 8386 15430
rect 8476 15396 8544 15430
rect 8634 15396 8702 15430
rect 8792 15396 8860 15430
rect 8950 15396 9018 15430
rect 9108 15396 9176 15430
rect 9266 15396 9334 15430
rect 9424 15396 9492 15430
rect 9582 15396 9650 15430
rect 9740 15396 9808 15430
rect 9898 15396 9966 15430
rect 10056 15396 10124 15430
rect 10214 15396 10282 15430
rect 10372 15396 10440 15430
rect 10530 15396 10598 15430
rect 10688 15396 10756 15430
rect 10846 15396 10914 15430
rect 11004 15396 11072 15430
rect 11162 15396 11230 15430
rect 11320 15396 11388 15430
rect 11478 15396 11546 15430
rect 11636 15396 11704 15430
rect 11794 15396 11862 15430
rect 11952 15396 12020 15430
rect 12110 15396 12178 15430
rect 12268 15396 12336 15430
rect 12426 15396 12494 15430
rect 7844 9286 7912 9320
rect 8002 9286 8070 9320
rect 8160 9286 8228 9320
rect 8318 9286 8386 9320
rect 8476 9286 8544 9320
rect 8634 9286 8702 9320
rect 8792 9286 8860 9320
rect 8950 9286 9018 9320
rect 9108 9286 9176 9320
rect 9266 9286 9334 9320
rect 9424 9286 9492 9320
rect 9582 9286 9650 9320
rect 9740 9286 9808 9320
rect 9898 9286 9966 9320
rect 10056 9286 10124 9320
rect 10214 9286 10282 9320
rect 10372 9286 10440 9320
rect 10530 9286 10598 9320
rect 10688 9286 10756 9320
rect 10846 9286 10914 9320
rect 11004 9286 11072 9320
rect 11162 9286 11230 9320
rect 11320 9286 11388 9320
rect 11478 9286 11546 9320
rect 11636 9286 11704 9320
rect 11794 9286 11862 9320
rect 11952 9286 12020 9320
rect 12110 9286 12178 9320
rect 12268 9286 12336 9320
rect 12426 9286 12494 9320
rect 14144 15396 14212 15430
rect 14302 15396 14370 15430
rect 14460 15396 14528 15430
rect 14618 15396 14686 15430
rect 14776 15396 14844 15430
rect 14934 15396 15002 15430
rect 15092 15396 15160 15430
rect 15250 15396 15318 15430
rect 15408 15396 15476 15430
rect 15566 15396 15634 15430
rect 15724 15396 15792 15430
rect 15882 15396 15950 15430
rect 16040 15396 16108 15430
rect 16198 15396 16266 15430
rect 16356 15396 16424 15430
rect 16514 15396 16582 15430
rect 16672 15396 16740 15430
rect 16830 15396 16898 15430
rect 16988 15396 17056 15430
rect 17146 15396 17214 15430
rect 17304 15396 17372 15430
rect 17462 15396 17530 15430
rect 17620 15396 17688 15430
rect 17778 15396 17846 15430
rect 17936 15396 18004 15430
rect 18094 15396 18162 15430
rect 18252 15396 18320 15430
rect 18410 15396 18478 15430
rect 18568 15396 18636 15430
rect 18726 15396 18794 15430
rect 14144 9286 14212 9320
rect 14302 9286 14370 9320
rect 14460 9286 14528 9320
rect 14618 9286 14686 9320
rect 14776 9286 14844 9320
rect 14934 9286 15002 9320
rect 15092 9286 15160 9320
rect 15250 9286 15318 9320
rect 15408 9286 15476 9320
rect 15566 9286 15634 9320
rect 15724 9286 15792 9320
rect 15882 9286 15950 9320
rect 16040 9286 16108 9320
rect 16198 9286 16266 9320
rect 16356 9286 16424 9320
rect 16514 9286 16582 9320
rect 16672 9286 16740 9320
rect 16830 9286 16898 9320
rect 16988 9286 17056 9320
rect 17146 9286 17214 9320
rect 17304 9286 17372 9320
rect 17462 9286 17530 9320
rect 17620 9286 17688 9320
rect 17778 9286 17846 9320
rect 17936 9286 18004 9320
rect 18094 9286 18162 9320
rect 18252 9286 18320 9320
rect 18410 9286 18478 9320
rect 18568 9286 18636 9320
rect 18726 9286 18794 9320
rect 20444 15396 20512 15430
rect 20602 15396 20670 15430
rect 20760 15396 20828 15430
rect 20918 15396 20986 15430
rect 21076 15396 21144 15430
rect 21234 15396 21302 15430
rect 21392 15396 21460 15430
rect 21550 15396 21618 15430
rect 21708 15396 21776 15430
rect 21866 15396 21934 15430
rect 22024 15396 22092 15430
rect 22182 15396 22250 15430
rect 22340 15396 22408 15430
rect 22498 15396 22566 15430
rect 22656 15396 22724 15430
rect 22814 15396 22882 15430
rect 22972 15396 23040 15430
rect 23130 15396 23198 15430
rect 23288 15396 23356 15430
rect 23446 15396 23514 15430
rect 23604 15396 23672 15430
rect 23762 15396 23830 15430
rect 23920 15396 23988 15430
rect 24078 15396 24146 15430
rect 24236 15396 24304 15430
rect 24394 15396 24462 15430
rect 24552 15396 24620 15430
rect 24710 15396 24778 15430
rect 24868 15396 24936 15430
rect 25026 15396 25094 15430
rect 20444 9286 20512 9320
rect 20602 9286 20670 9320
rect 20760 9286 20828 9320
rect 20918 9286 20986 9320
rect 21076 9286 21144 9320
rect 21234 9286 21302 9320
rect 21392 9286 21460 9320
rect 21550 9286 21618 9320
rect 21708 9286 21776 9320
rect 21866 9286 21934 9320
rect 22024 9286 22092 9320
rect 22182 9286 22250 9320
rect 22340 9286 22408 9320
rect 22498 9286 22566 9320
rect 22656 9286 22724 9320
rect 22814 9286 22882 9320
rect 22972 9286 23040 9320
rect 23130 9286 23198 9320
rect 23288 9286 23356 9320
rect 23446 9286 23514 9320
rect 23604 9286 23672 9320
rect 23762 9286 23830 9320
rect 23920 9286 23988 9320
rect 24078 9286 24146 9320
rect 24236 9286 24304 9320
rect 24394 9286 24462 9320
rect 24552 9286 24620 9320
rect 24710 9286 24778 9320
rect 24868 9286 24936 9320
rect 25026 9286 25094 9320
rect 1544 8396 1612 8430
rect 1702 8396 1770 8430
rect 1860 8396 1928 8430
rect 2018 8396 2086 8430
rect 2176 8396 2244 8430
rect 2334 8396 2402 8430
rect 2492 8396 2560 8430
rect 2650 8396 2718 8430
rect 2808 8396 2876 8430
rect 2966 8396 3034 8430
rect 3124 8396 3192 8430
rect 3282 8396 3350 8430
rect 3440 8396 3508 8430
rect 3598 8396 3666 8430
rect 3756 8396 3824 8430
rect 3914 8396 3982 8430
rect 4072 8396 4140 8430
rect 4230 8396 4298 8430
rect 4388 8396 4456 8430
rect 4546 8396 4614 8430
rect 4704 8396 4772 8430
rect 4862 8396 4930 8430
rect 5020 8396 5088 8430
rect 5178 8396 5246 8430
rect 5336 8396 5404 8430
rect 5494 8396 5562 8430
rect 5652 8396 5720 8430
rect 5810 8396 5878 8430
rect 5968 8396 6036 8430
rect 6126 8396 6194 8430
rect 1544 2286 1612 2320
rect 1702 2286 1770 2320
rect 1860 2286 1928 2320
rect 2018 2286 2086 2320
rect 2176 2286 2244 2320
rect 2334 2286 2402 2320
rect 2492 2286 2560 2320
rect 2650 2286 2718 2320
rect 2808 2286 2876 2320
rect 2966 2286 3034 2320
rect 3124 2286 3192 2320
rect 3282 2286 3350 2320
rect 3440 2286 3508 2320
rect 3598 2286 3666 2320
rect 3756 2286 3824 2320
rect 3914 2286 3982 2320
rect 4072 2286 4140 2320
rect 4230 2286 4298 2320
rect 4388 2286 4456 2320
rect 4546 2286 4614 2320
rect 4704 2286 4772 2320
rect 4862 2286 4930 2320
rect 5020 2286 5088 2320
rect 5178 2286 5246 2320
rect 5336 2286 5404 2320
rect 5494 2286 5562 2320
rect 5652 2286 5720 2320
rect 5810 2286 5878 2320
rect 5968 2286 6036 2320
rect 6126 2286 6194 2320
rect 7844 8396 7912 8430
rect 8002 8396 8070 8430
rect 8160 8396 8228 8430
rect 8318 8396 8386 8430
rect 8476 8396 8544 8430
rect 8634 8396 8702 8430
rect 8792 8396 8860 8430
rect 8950 8396 9018 8430
rect 9108 8396 9176 8430
rect 9266 8396 9334 8430
rect 9424 8396 9492 8430
rect 9582 8396 9650 8430
rect 9740 8396 9808 8430
rect 9898 8396 9966 8430
rect 10056 8396 10124 8430
rect 10214 8396 10282 8430
rect 10372 8396 10440 8430
rect 10530 8396 10598 8430
rect 10688 8396 10756 8430
rect 10846 8396 10914 8430
rect 11004 8396 11072 8430
rect 11162 8396 11230 8430
rect 11320 8396 11388 8430
rect 11478 8396 11546 8430
rect 11636 8396 11704 8430
rect 11794 8396 11862 8430
rect 11952 8396 12020 8430
rect 12110 8396 12178 8430
rect 12268 8396 12336 8430
rect 12426 8396 12494 8430
rect 7844 2286 7912 2320
rect 8002 2286 8070 2320
rect 8160 2286 8228 2320
rect 8318 2286 8386 2320
rect 8476 2286 8544 2320
rect 8634 2286 8702 2320
rect 8792 2286 8860 2320
rect 8950 2286 9018 2320
rect 9108 2286 9176 2320
rect 9266 2286 9334 2320
rect 9424 2286 9492 2320
rect 9582 2286 9650 2320
rect 9740 2286 9808 2320
rect 9898 2286 9966 2320
rect 10056 2286 10124 2320
rect 10214 2286 10282 2320
rect 10372 2286 10440 2320
rect 10530 2286 10598 2320
rect 10688 2286 10756 2320
rect 10846 2286 10914 2320
rect 11004 2286 11072 2320
rect 11162 2286 11230 2320
rect 11320 2286 11388 2320
rect 11478 2286 11546 2320
rect 11636 2286 11704 2320
rect 11794 2286 11862 2320
rect 11952 2286 12020 2320
rect 12110 2286 12178 2320
rect 12268 2286 12336 2320
rect 12426 2286 12494 2320
rect 14144 8396 14212 8430
rect 14302 8396 14370 8430
rect 14460 8396 14528 8430
rect 14618 8396 14686 8430
rect 14776 8396 14844 8430
rect 14934 8396 15002 8430
rect 15092 8396 15160 8430
rect 15250 8396 15318 8430
rect 15408 8396 15476 8430
rect 15566 8396 15634 8430
rect 15724 8396 15792 8430
rect 15882 8396 15950 8430
rect 16040 8396 16108 8430
rect 16198 8396 16266 8430
rect 16356 8396 16424 8430
rect 16514 8396 16582 8430
rect 16672 8396 16740 8430
rect 16830 8396 16898 8430
rect 16988 8396 17056 8430
rect 17146 8396 17214 8430
rect 17304 8396 17372 8430
rect 17462 8396 17530 8430
rect 17620 8396 17688 8430
rect 17778 8396 17846 8430
rect 17936 8396 18004 8430
rect 18094 8396 18162 8430
rect 18252 8396 18320 8430
rect 18410 8396 18478 8430
rect 18568 8396 18636 8430
rect 18726 8396 18794 8430
rect 14144 2286 14212 2320
rect 14302 2286 14370 2320
rect 14460 2286 14528 2320
rect 14618 2286 14686 2320
rect 14776 2286 14844 2320
rect 14934 2286 15002 2320
rect 15092 2286 15160 2320
rect 15250 2286 15318 2320
rect 15408 2286 15476 2320
rect 15566 2286 15634 2320
rect 15724 2286 15792 2320
rect 15882 2286 15950 2320
rect 16040 2286 16108 2320
rect 16198 2286 16266 2320
rect 16356 2286 16424 2320
rect 16514 2286 16582 2320
rect 16672 2286 16740 2320
rect 16830 2286 16898 2320
rect 16988 2286 17056 2320
rect 17146 2286 17214 2320
rect 17304 2286 17372 2320
rect 17462 2286 17530 2320
rect 17620 2286 17688 2320
rect 17778 2286 17846 2320
rect 17936 2286 18004 2320
rect 18094 2286 18162 2320
rect 18252 2286 18320 2320
rect 18410 2286 18478 2320
rect 18568 2286 18636 2320
rect 18726 2286 18794 2320
rect 20444 8396 20512 8430
rect 20602 8396 20670 8430
rect 20760 8396 20828 8430
rect 20918 8396 20986 8430
rect 21076 8396 21144 8430
rect 21234 8396 21302 8430
rect 21392 8396 21460 8430
rect 21550 8396 21618 8430
rect 21708 8396 21776 8430
rect 21866 8396 21934 8430
rect 22024 8396 22092 8430
rect 22182 8396 22250 8430
rect 22340 8396 22408 8430
rect 22498 8396 22566 8430
rect 22656 8396 22724 8430
rect 22814 8396 22882 8430
rect 22972 8396 23040 8430
rect 23130 8396 23198 8430
rect 23288 8396 23356 8430
rect 23446 8396 23514 8430
rect 23604 8396 23672 8430
rect 23762 8396 23830 8430
rect 23920 8396 23988 8430
rect 24078 8396 24146 8430
rect 24236 8396 24304 8430
rect 24394 8396 24462 8430
rect 24552 8396 24620 8430
rect 24710 8396 24778 8430
rect 24868 8396 24936 8430
rect 25026 8396 25094 8430
rect 20444 2286 20512 2320
rect 20602 2286 20670 2320
rect 20760 2286 20828 2320
rect 20918 2286 20986 2320
rect 21076 2286 21144 2320
rect 21234 2286 21302 2320
rect 21392 2286 21460 2320
rect 21550 2286 21618 2320
rect 21708 2286 21776 2320
rect 21866 2286 21934 2320
rect 22024 2286 22092 2320
rect 22182 2286 22250 2320
rect 22340 2286 22408 2320
rect 22498 2286 22566 2320
rect 22656 2286 22724 2320
rect 22814 2286 22882 2320
rect 22972 2286 23040 2320
rect 23130 2286 23198 2320
rect 23288 2286 23356 2320
rect 23446 2286 23514 2320
rect 23604 2286 23672 2320
rect 23762 2286 23830 2320
rect 23920 2286 23988 2320
rect 24078 2286 24146 2320
rect 24236 2286 24304 2320
rect 24394 2286 24462 2320
rect 24552 2286 24620 2320
rect 24710 2286 24778 2320
rect 24868 2286 24936 2320
rect 25026 2286 25094 2320
<< xpolycontact >>
rect -4234 13418 -4164 13850
rect -4234 12666 -4164 13098
rect 30964 13418 31034 13850
rect 30964 12666 31034 13098
<< npolyres >>
rect -3234 38919 -3168 40219
rect 29968 38919 30034 40219
rect -4234 25719 -4168 27019
rect 30968 25719 31034 27019
<< ppolyres >>
rect -4234 13098 -4164 13418
rect 30964 13098 31034 13418
<< locali >>
rect 1348 46134 1444 46168
rect 6294 46134 6390 46168
rect 1348 46072 1382 46134
rect 6356 46072 6390 46134
rect 1528 45996 1544 46030
rect 1612 45996 1628 46030
rect 1686 45996 1702 46030
rect 1770 45996 1786 46030
rect 1844 45996 1860 46030
rect 1928 45996 1944 46030
rect 2002 45996 2018 46030
rect 2086 45996 2102 46030
rect 2160 45996 2176 46030
rect 2244 45996 2260 46030
rect 2318 45996 2334 46030
rect 2402 45996 2418 46030
rect 2476 45996 2492 46030
rect 2560 45996 2576 46030
rect 2634 45996 2650 46030
rect 2718 45996 2734 46030
rect 2792 45996 2808 46030
rect 2876 45996 2892 46030
rect 2950 45996 2966 46030
rect 3034 45996 3050 46030
rect 3108 45996 3124 46030
rect 3192 45996 3208 46030
rect 3266 45996 3282 46030
rect 3350 45996 3366 46030
rect 3424 45996 3440 46030
rect 3508 45996 3524 46030
rect 3582 45996 3598 46030
rect 3666 45996 3682 46030
rect 3740 45996 3756 46030
rect 3824 45996 3840 46030
rect 3898 45996 3914 46030
rect 3982 45996 3998 46030
rect 4056 45996 4072 46030
rect 4140 45996 4156 46030
rect 4214 45996 4230 46030
rect 4298 45996 4314 46030
rect 4372 45996 4388 46030
rect 4456 45996 4472 46030
rect 4530 45996 4546 46030
rect 4614 45996 4630 46030
rect 4688 45996 4704 46030
rect 4772 45996 4788 46030
rect 4846 45996 4862 46030
rect 4930 45996 4946 46030
rect 5004 45996 5020 46030
rect 5088 45996 5104 46030
rect 5162 45996 5178 46030
rect 5246 45996 5262 46030
rect 5320 45996 5336 46030
rect 5404 45996 5420 46030
rect 5478 45996 5494 46030
rect 5562 45996 5578 46030
rect 5636 45996 5652 46030
rect 5720 45996 5736 46030
rect 5794 45996 5810 46030
rect 5878 45996 5894 46030
rect 5952 45996 5968 46030
rect 6036 45996 6052 46030
rect 6110 45996 6126 46030
rect 6194 45996 6210 46030
rect 7648 46134 7744 46168
rect 12594 46134 12690 46168
rect 7648 46072 7682 46134
rect 12656 46072 12690 46134
rect 7828 45996 7844 46030
rect 7912 45996 7928 46030
rect 7986 45996 8002 46030
rect 8070 45996 8086 46030
rect 8144 45996 8160 46030
rect 8228 45996 8244 46030
rect 8302 45996 8318 46030
rect 8386 45996 8402 46030
rect 8460 45996 8476 46030
rect 8544 45996 8560 46030
rect 8618 45996 8634 46030
rect 8702 45996 8718 46030
rect 8776 45996 8792 46030
rect 8860 45996 8876 46030
rect 8934 45996 8950 46030
rect 9018 45996 9034 46030
rect 9092 45996 9108 46030
rect 9176 45996 9192 46030
rect 9250 45996 9266 46030
rect 9334 45996 9350 46030
rect 9408 45996 9424 46030
rect 9492 45996 9508 46030
rect 9566 45996 9582 46030
rect 9650 45996 9666 46030
rect 9724 45996 9740 46030
rect 9808 45996 9824 46030
rect 9882 45996 9898 46030
rect 9966 45996 9982 46030
rect 10040 45996 10056 46030
rect 10124 45996 10140 46030
rect 10198 45996 10214 46030
rect 10282 45996 10298 46030
rect 10356 45996 10372 46030
rect 10440 45996 10456 46030
rect 10514 45996 10530 46030
rect 10598 45996 10614 46030
rect 10672 45996 10688 46030
rect 10756 45996 10772 46030
rect 10830 45996 10846 46030
rect 10914 45996 10930 46030
rect 10988 45996 11004 46030
rect 11072 45996 11088 46030
rect 11146 45996 11162 46030
rect 11230 45996 11246 46030
rect 11304 45996 11320 46030
rect 11388 45996 11404 46030
rect 11462 45996 11478 46030
rect 11546 45996 11562 46030
rect 11620 45996 11636 46030
rect 11704 45996 11720 46030
rect 11778 45996 11794 46030
rect 11862 45996 11878 46030
rect 11936 45996 11952 46030
rect 12020 45996 12036 46030
rect 12094 45996 12110 46030
rect 12178 45996 12194 46030
rect 12252 45996 12268 46030
rect 12336 45996 12352 46030
rect 12410 45996 12426 46030
rect 12494 45996 12510 46030
rect 13948 46134 14044 46168
rect 18894 46134 18990 46168
rect 13948 46072 13982 46134
rect 18956 46072 18990 46134
rect 14128 45996 14144 46030
rect 14212 45996 14228 46030
rect 14286 45996 14302 46030
rect 14370 45996 14386 46030
rect 14444 45996 14460 46030
rect 14528 45996 14544 46030
rect 14602 45996 14618 46030
rect 14686 45996 14702 46030
rect 14760 45996 14776 46030
rect 14844 45996 14860 46030
rect 14918 45996 14934 46030
rect 15002 45996 15018 46030
rect 15076 45996 15092 46030
rect 15160 45996 15176 46030
rect 15234 45996 15250 46030
rect 15318 45996 15334 46030
rect 15392 45996 15408 46030
rect 15476 45996 15492 46030
rect 15550 45996 15566 46030
rect 15634 45996 15650 46030
rect 15708 45996 15724 46030
rect 15792 45996 15808 46030
rect 15866 45996 15882 46030
rect 15950 45996 15966 46030
rect 16024 45996 16040 46030
rect 16108 45996 16124 46030
rect 16182 45996 16198 46030
rect 16266 45996 16282 46030
rect 16340 45996 16356 46030
rect 16424 45996 16440 46030
rect 16498 45996 16514 46030
rect 16582 45996 16598 46030
rect 16656 45996 16672 46030
rect 16740 45996 16756 46030
rect 16814 45996 16830 46030
rect 16898 45996 16914 46030
rect 16972 45996 16988 46030
rect 17056 45996 17072 46030
rect 17130 45996 17146 46030
rect 17214 45996 17230 46030
rect 17288 45996 17304 46030
rect 17372 45996 17388 46030
rect 17446 45996 17462 46030
rect 17530 45996 17546 46030
rect 17604 45996 17620 46030
rect 17688 45996 17704 46030
rect 17762 45996 17778 46030
rect 17846 45996 17862 46030
rect 17920 45996 17936 46030
rect 18004 45996 18020 46030
rect 18078 45996 18094 46030
rect 18162 45996 18178 46030
rect 18236 45996 18252 46030
rect 18320 45996 18336 46030
rect 18394 45996 18410 46030
rect 18478 45996 18494 46030
rect 18552 45996 18568 46030
rect 18636 45996 18652 46030
rect 18710 45996 18726 46030
rect 18794 45996 18810 46030
rect 20248 46134 20344 46168
rect 25194 46134 25290 46168
rect 20248 46072 20282 46134
rect 25256 46072 25290 46134
rect 20428 45996 20444 46030
rect 20512 45996 20528 46030
rect 20586 45996 20602 46030
rect 20670 45996 20686 46030
rect 20744 45996 20760 46030
rect 20828 45996 20844 46030
rect 20902 45996 20918 46030
rect 20986 45996 21002 46030
rect 21060 45996 21076 46030
rect 21144 45996 21160 46030
rect 21218 45996 21234 46030
rect 21302 45996 21318 46030
rect 21376 45996 21392 46030
rect 21460 45996 21476 46030
rect 21534 45996 21550 46030
rect 21618 45996 21634 46030
rect 21692 45996 21708 46030
rect 21776 45996 21792 46030
rect 21850 45996 21866 46030
rect 21934 45996 21950 46030
rect 22008 45996 22024 46030
rect 22092 45996 22108 46030
rect 22166 45996 22182 46030
rect 22250 45996 22266 46030
rect 22324 45996 22340 46030
rect 22408 45996 22424 46030
rect 22482 45996 22498 46030
rect 22566 45996 22582 46030
rect 22640 45996 22656 46030
rect 22724 45996 22740 46030
rect 22798 45996 22814 46030
rect 22882 45996 22898 46030
rect 22956 45996 22972 46030
rect 23040 45996 23056 46030
rect 23114 45996 23130 46030
rect 23198 45996 23214 46030
rect 23272 45996 23288 46030
rect 23356 45996 23372 46030
rect 23430 45996 23446 46030
rect 23514 45996 23530 46030
rect 23588 45996 23604 46030
rect 23672 45996 23688 46030
rect 23746 45996 23762 46030
rect 23830 45996 23846 46030
rect 23904 45996 23920 46030
rect 23988 45996 24004 46030
rect 24062 45996 24078 46030
rect 24146 45996 24162 46030
rect 24220 45996 24236 46030
rect 24304 45996 24320 46030
rect 24378 45996 24394 46030
rect 24462 45996 24478 46030
rect 24536 45996 24552 46030
rect 24620 45996 24636 46030
rect 24694 45996 24710 46030
rect 24778 45996 24794 46030
rect 24852 45996 24868 46030
rect 24936 45996 24952 46030
rect 25010 45996 25026 46030
rect 25094 45996 25110 46030
rect -3364 40388 -3268 40422
rect -3134 40420 -3038 40422
rect -3134 40400 -2980 40420
rect -3134 40388 -3040 40400
rect -3364 40326 -3330 40388
rect -3072 40326 -3040 40388
rect -3234 40242 -3218 40276
rect -3184 40242 -3168 40276
rect -3234 38862 -3218 38896
rect -3184 38862 -3168 38896
rect -3364 38750 -3330 38812
rect -3072 38750 -3040 38812
rect -3364 38716 -3268 38750
rect -3134 38740 -3040 38750
rect -3000 38740 -2980 40400
rect 1482 45946 1516 45962
rect 1482 39954 1516 39970
rect 1640 45946 1674 45962
rect 1640 39954 1674 39970
rect 1798 45946 1832 45962
rect 1798 39954 1832 39970
rect 1956 45946 1990 45962
rect 1956 39954 1990 39970
rect 2114 45946 2148 45962
rect 2114 39954 2148 39970
rect 2272 45946 2306 45962
rect 2272 39954 2306 39970
rect 2430 45946 2464 45962
rect 2430 39954 2464 39970
rect 2588 45946 2622 45962
rect 2588 39954 2622 39970
rect 2746 45946 2780 45962
rect 2746 39954 2780 39970
rect 2904 45946 2938 45962
rect 2904 39954 2938 39970
rect 3062 45946 3096 45962
rect 3062 39954 3096 39970
rect 3220 45946 3254 45962
rect 3220 39954 3254 39970
rect 3378 45946 3412 45962
rect 3378 39954 3412 39970
rect 3536 45946 3570 45962
rect 3536 39954 3570 39970
rect 3694 45946 3728 45962
rect 3694 39954 3728 39970
rect 3852 45946 3886 45962
rect 3852 39954 3886 39970
rect 4010 45946 4044 45962
rect 4010 39954 4044 39970
rect 4168 45946 4202 45962
rect 4168 39954 4202 39970
rect 4326 45946 4360 45962
rect 4326 39954 4360 39970
rect 4484 45946 4518 45962
rect 4484 39954 4518 39970
rect 4642 45946 4676 45962
rect 4642 39954 4676 39970
rect 4800 45946 4834 45962
rect 4800 39954 4834 39970
rect 4958 45946 4992 45962
rect 4958 39954 4992 39970
rect 5116 45946 5150 45962
rect 5116 39954 5150 39970
rect 5274 45946 5308 45962
rect 5274 39954 5308 39970
rect 5432 45946 5466 45962
rect 5432 39954 5466 39970
rect 5590 45946 5624 45962
rect 5590 39954 5624 39970
rect 5748 45946 5782 45962
rect 5748 39954 5782 39970
rect 5906 45946 5940 45962
rect 5906 39954 5940 39970
rect 6064 45946 6098 45962
rect 6064 39954 6098 39970
rect 6222 45946 6256 45962
rect 6222 39954 6256 39970
rect 7782 45946 7816 45962
rect 7782 39954 7816 39970
rect 7940 45946 7974 45962
rect 7940 39954 7974 39970
rect 8098 45946 8132 45962
rect 8098 39954 8132 39970
rect 8256 45946 8290 45962
rect 8256 39954 8290 39970
rect 8414 45946 8448 45962
rect 8414 39954 8448 39970
rect 8572 45946 8606 45962
rect 8572 39954 8606 39970
rect 8730 45946 8764 45962
rect 8730 39954 8764 39970
rect 8888 45946 8922 45962
rect 8888 39954 8922 39970
rect 9046 45946 9080 45962
rect 9046 39954 9080 39970
rect 9204 45946 9238 45962
rect 9204 39954 9238 39970
rect 9362 45946 9396 45962
rect 9362 39954 9396 39970
rect 9520 45946 9554 45962
rect 9520 39954 9554 39970
rect 9678 45946 9712 45962
rect 9678 39954 9712 39970
rect 9836 45946 9870 45962
rect 9836 39954 9870 39970
rect 9994 45946 10028 45962
rect 9994 39954 10028 39970
rect 10152 45946 10186 45962
rect 10152 39954 10186 39970
rect 10310 45946 10344 45962
rect 10310 39954 10344 39970
rect 10468 45946 10502 45962
rect 10468 39954 10502 39970
rect 10626 45946 10660 45962
rect 10626 39954 10660 39970
rect 10784 45946 10818 45962
rect 10784 39954 10818 39970
rect 10942 45946 10976 45962
rect 10942 39954 10976 39970
rect 11100 45946 11134 45962
rect 11100 39954 11134 39970
rect 11258 45946 11292 45962
rect 11258 39954 11292 39970
rect 11416 45946 11450 45962
rect 11416 39954 11450 39970
rect 11574 45946 11608 45962
rect 11574 39954 11608 39970
rect 11732 45946 11766 45962
rect 11732 39954 11766 39970
rect 11890 45946 11924 45962
rect 11890 39954 11924 39970
rect 12048 45946 12082 45962
rect 12048 39954 12082 39970
rect 12206 45946 12240 45962
rect 12206 39954 12240 39970
rect 12364 45946 12398 45962
rect 12364 39954 12398 39970
rect 12522 45946 12556 45962
rect 12522 39954 12556 39970
rect 14082 45946 14116 45962
rect 14082 39954 14116 39970
rect 14240 45946 14274 45962
rect 14240 39954 14274 39970
rect 14398 45946 14432 45962
rect 14398 39954 14432 39970
rect 14556 45946 14590 45962
rect 14556 39954 14590 39970
rect 14714 45946 14748 45962
rect 14714 39954 14748 39970
rect 14872 45946 14906 45962
rect 14872 39954 14906 39970
rect 15030 45946 15064 45962
rect 15030 39954 15064 39970
rect 15188 45946 15222 45962
rect 15188 39954 15222 39970
rect 15346 45946 15380 45962
rect 15346 39954 15380 39970
rect 15504 45946 15538 45962
rect 15504 39954 15538 39970
rect 15662 45946 15696 45962
rect 15662 39954 15696 39970
rect 15820 45946 15854 45962
rect 15820 39954 15854 39970
rect 15978 45946 16012 45962
rect 15978 39954 16012 39970
rect 16136 45946 16170 45962
rect 16136 39954 16170 39970
rect 16294 45946 16328 45962
rect 16294 39954 16328 39970
rect 16452 45946 16486 45962
rect 16452 39954 16486 39970
rect 16610 45946 16644 45962
rect 16610 39954 16644 39970
rect 16768 45946 16802 45962
rect 16768 39954 16802 39970
rect 16926 45946 16960 45962
rect 16926 39954 16960 39970
rect 17084 45946 17118 45962
rect 17084 39954 17118 39970
rect 17242 45946 17276 45962
rect 17242 39954 17276 39970
rect 17400 45946 17434 45962
rect 17400 39954 17434 39970
rect 17558 45946 17592 45962
rect 17558 39954 17592 39970
rect 17716 45946 17750 45962
rect 17716 39954 17750 39970
rect 17874 45946 17908 45962
rect 17874 39954 17908 39970
rect 18032 45946 18066 45962
rect 18032 39954 18066 39970
rect 18190 45946 18224 45962
rect 18190 39954 18224 39970
rect 18348 45946 18382 45962
rect 18348 39954 18382 39970
rect 18506 45946 18540 45962
rect 18506 39954 18540 39970
rect 18664 45946 18698 45962
rect 18664 39954 18698 39970
rect 18822 45946 18856 45962
rect 18822 39954 18856 39970
rect 20382 45946 20416 45962
rect 20382 39954 20416 39970
rect 20540 45946 20574 45962
rect 20540 39954 20574 39970
rect 20698 45946 20732 45962
rect 20698 39954 20732 39970
rect 20856 45946 20890 45962
rect 20856 39954 20890 39970
rect 21014 45946 21048 45962
rect 21014 39954 21048 39970
rect 21172 45946 21206 45962
rect 21172 39954 21206 39970
rect 21330 45946 21364 45962
rect 21330 39954 21364 39970
rect 21488 45946 21522 45962
rect 21488 39954 21522 39970
rect 21646 45946 21680 45962
rect 21646 39954 21680 39970
rect 21804 45946 21838 45962
rect 21804 39954 21838 39970
rect 21962 45946 21996 45962
rect 21962 39954 21996 39970
rect 22120 45946 22154 45962
rect 22120 39954 22154 39970
rect 22278 45946 22312 45962
rect 22278 39954 22312 39970
rect 22436 45946 22470 45962
rect 22436 39954 22470 39970
rect 22594 45946 22628 45962
rect 22594 39954 22628 39970
rect 22752 45946 22786 45962
rect 22752 39954 22786 39970
rect 22910 45946 22944 45962
rect 22910 39954 22944 39970
rect 23068 45946 23102 45962
rect 23068 39954 23102 39970
rect 23226 45946 23260 45962
rect 23226 39954 23260 39970
rect 23384 45946 23418 45962
rect 23384 39954 23418 39970
rect 23542 45946 23576 45962
rect 23542 39954 23576 39970
rect 23700 45946 23734 45962
rect 23700 39954 23734 39970
rect 23858 45946 23892 45962
rect 23858 39954 23892 39970
rect 24016 45946 24050 45962
rect 24016 39954 24050 39970
rect 24174 45946 24208 45962
rect 24174 39954 24208 39970
rect 24332 45946 24366 45962
rect 24332 39954 24366 39970
rect 24490 45946 24524 45962
rect 24490 39954 24524 39970
rect 24648 45946 24682 45962
rect 24648 39954 24682 39970
rect 24806 45946 24840 45962
rect 24806 39954 24840 39970
rect 24964 45946 24998 45962
rect 24964 39954 24998 39970
rect 25122 45946 25156 45962
rect 25122 39954 25156 39970
rect 29838 40420 29934 40422
rect 29780 40400 29934 40420
rect 1528 39886 1544 39920
rect 1612 39886 1628 39920
rect 1686 39886 1702 39920
rect 1770 39886 1786 39920
rect 1844 39886 1860 39920
rect 1928 39886 1944 39920
rect 2002 39886 2018 39920
rect 2086 39886 2102 39920
rect 2160 39886 2176 39920
rect 2244 39886 2260 39920
rect 2318 39886 2334 39920
rect 2402 39886 2418 39920
rect 2476 39886 2492 39920
rect 2560 39886 2576 39920
rect 2634 39886 2650 39920
rect 2718 39886 2734 39920
rect 2792 39886 2808 39920
rect 2876 39886 2892 39920
rect 2950 39886 2966 39920
rect 3034 39886 3050 39920
rect 3108 39886 3124 39920
rect 3192 39886 3208 39920
rect 3266 39886 3282 39920
rect 3350 39886 3366 39920
rect 3424 39886 3440 39920
rect 3508 39886 3524 39920
rect 3582 39886 3598 39920
rect 3666 39886 3682 39920
rect 3740 39886 3756 39920
rect 3824 39886 3840 39920
rect 3898 39886 3914 39920
rect 3982 39886 3998 39920
rect 4056 39886 4072 39920
rect 4140 39886 4156 39920
rect 4214 39886 4230 39920
rect 4298 39886 4314 39920
rect 4372 39886 4388 39920
rect 4456 39886 4472 39920
rect 4530 39886 4546 39920
rect 4614 39886 4630 39920
rect 4688 39886 4704 39920
rect 4772 39886 4788 39920
rect 4846 39886 4862 39920
rect 4930 39886 4946 39920
rect 5004 39886 5020 39920
rect 5088 39886 5104 39920
rect 5162 39886 5178 39920
rect 5246 39886 5262 39920
rect 5320 39886 5336 39920
rect 5404 39886 5420 39920
rect 5478 39886 5494 39920
rect 5562 39886 5578 39920
rect 5636 39886 5652 39920
rect 5720 39886 5736 39920
rect 5794 39886 5810 39920
rect 5878 39886 5894 39920
rect 5952 39886 5968 39920
rect 6036 39886 6052 39920
rect 6110 39886 6126 39920
rect 6194 39886 6210 39920
rect 1348 39782 1382 39844
rect 6356 39782 6390 39844
rect 1348 39748 1444 39782
rect 6294 39748 6390 39782
rect 7828 39886 7844 39920
rect 7912 39886 7928 39920
rect 7986 39886 8002 39920
rect 8070 39886 8086 39920
rect 8144 39886 8160 39920
rect 8228 39886 8244 39920
rect 8302 39886 8318 39920
rect 8386 39886 8402 39920
rect 8460 39886 8476 39920
rect 8544 39886 8560 39920
rect 8618 39886 8634 39920
rect 8702 39886 8718 39920
rect 8776 39886 8792 39920
rect 8860 39886 8876 39920
rect 8934 39886 8950 39920
rect 9018 39886 9034 39920
rect 9092 39886 9108 39920
rect 9176 39886 9192 39920
rect 9250 39886 9266 39920
rect 9334 39886 9350 39920
rect 9408 39886 9424 39920
rect 9492 39886 9508 39920
rect 9566 39886 9582 39920
rect 9650 39886 9666 39920
rect 9724 39886 9740 39920
rect 9808 39886 9824 39920
rect 9882 39886 9898 39920
rect 9966 39886 9982 39920
rect 10040 39886 10056 39920
rect 10124 39886 10140 39920
rect 10198 39886 10214 39920
rect 10282 39886 10298 39920
rect 10356 39886 10372 39920
rect 10440 39886 10456 39920
rect 10514 39886 10530 39920
rect 10598 39886 10614 39920
rect 10672 39886 10688 39920
rect 10756 39886 10772 39920
rect 10830 39886 10846 39920
rect 10914 39886 10930 39920
rect 10988 39886 11004 39920
rect 11072 39886 11088 39920
rect 11146 39886 11162 39920
rect 11230 39886 11246 39920
rect 11304 39886 11320 39920
rect 11388 39886 11404 39920
rect 11462 39886 11478 39920
rect 11546 39886 11562 39920
rect 11620 39886 11636 39920
rect 11704 39886 11720 39920
rect 11778 39886 11794 39920
rect 11862 39886 11878 39920
rect 11936 39886 11952 39920
rect 12020 39886 12036 39920
rect 12094 39886 12110 39920
rect 12178 39886 12194 39920
rect 12252 39886 12268 39920
rect 12336 39886 12352 39920
rect 12410 39886 12426 39920
rect 12494 39886 12510 39920
rect 7648 39782 7682 39844
rect 12656 39782 12690 39844
rect 7648 39748 7744 39782
rect 12594 39748 12690 39782
rect 14128 39886 14144 39920
rect 14212 39886 14228 39920
rect 14286 39886 14302 39920
rect 14370 39886 14386 39920
rect 14444 39886 14460 39920
rect 14528 39886 14544 39920
rect 14602 39886 14618 39920
rect 14686 39886 14702 39920
rect 14760 39886 14776 39920
rect 14844 39886 14860 39920
rect 14918 39886 14934 39920
rect 15002 39886 15018 39920
rect 15076 39886 15092 39920
rect 15160 39886 15176 39920
rect 15234 39886 15250 39920
rect 15318 39886 15334 39920
rect 15392 39886 15408 39920
rect 15476 39886 15492 39920
rect 15550 39886 15566 39920
rect 15634 39886 15650 39920
rect 15708 39886 15724 39920
rect 15792 39886 15808 39920
rect 15866 39886 15882 39920
rect 15950 39886 15966 39920
rect 16024 39886 16040 39920
rect 16108 39886 16124 39920
rect 16182 39886 16198 39920
rect 16266 39886 16282 39920
rect 16340 39886 16356 39920
rect 16424 39886 16440 39920
rect 16498 39886 16514 39920
rect 16582 39886 16598 39920
rect 16656 39886 16672 39920
rect 16740 39886 16756 39920
rect 16814 39886 16830 39920
rect 16898 39886 16914 39920
rect 16972 39886 16988 39920
rect 17056 39886 17072 39920
rect 17130 39886 17146 39920
rect 17214 39886 17230 39920
rect 17288 39886 17304 39920
rect 17372 39886 17388 39920
rect 17446 39886 17462 39920
rect 17530 39886 17546 39920
rect 17604 39886 17620 39920
rect 17688 39886 17704 39920
rect 17762 39886 17778 39920
rect 17846 39886 17862 39920
rect 17920 39886 17936 39920
rect 18004 39886 18020 39920
rect 18078 39886 18094 39920
rect 18162 39886 18178 39920
rect 18236 39886 18252 39920
rect 18320 39886 18336 39920
rect 18394 39886 18410 39920
rect 18478 39886 18494 39920
rect 18552 39886 18568 39920
rect 18636 39886 18652 39920
rect 18710 39886 18726 39920
rect 18794 39886 18810 39920
rect 13948 39782 13982 39844
rect 18956 39782 18990 39844
rect 13948 39748 14044 39782
rect 18894 39748 18990 39782
rect 20428 39886 20444 39920
rect 20512 39886 20528 39920
rect 20586 39886 20602 39920
rect 20670 39886 20686 39920
rect 20744 39886 20760 39920
rect 20828 39886 20844 39920
rect 20902 39886 20918 39920
rect 20986 39886 21002 39920
rect 21060 39886 21076 39920
rect 21144 39886 21160 39920
rect 21218 39886 21234 39920
rect 21302 39886 21318 39920
rect 21376 39886 21392 39920
rect 21460 39886 21476 39920
rect 21534 39886 21550 39920
rect 21618 39886 21634 39920
rect 21692 39886 21708 39920
rect 21776 39886 21792 39920
rect 21850 39886 21866 39920
rect 21934 39886 21950 39920
rect 22008 39886 22024 39920
rect 22092 39886 22108 39920
rect 22166 39886 22182 39920
rect 22250 39886 22266 39920
rect 22324 39886 22340 39920
rect 22408 39886 22424 39920
rect 22482 39886 22498 39920
rect 22566 39886 22582 39920
rect 22640 39886 22656 39920
rect 22724 39886 22740 39920
rect 22798 39886 22814 39920
rect 22882 39886 22898 39920
rect 22956 39886 22972 39920
rect 23040 39886 23056 39920
rect 23114 39886 23130 39920
rect 23198 39886 23214 39920
rect 23272 39886 23288 39920
rect 23356 39886 23372 39920
rect 23430 39886 23446 39920
rect 23514 39886 23530 39920
rect 23588 39886 23604 39920
rect 23672 39886 23688 39920
rect 23746 39886 23762 39920
rect 23830 39886 23846 39920
rect 23904 39886 23920 39920
rect 23988 39886 24004 39920
rect 24062 39886 24078 39920
rect 24146 39886 24162 39920
rect 24220 39886 24236 39920
rect 24304 39886 24320 39920
rect 24378 39886 24394 39920
rect 24462 39886 24478 39920
rect 24536 39886 24552 39920
rect 24620 39886 24636 39920
rect 24694 39886 24710 39920
rect 24778 39886 24794 39920
rect 24852 39886 24868 39920
rect 24936 39886 24952 39920
rect 25010 39886 25026 39920
rect 25094 39886 25110 39920
rect 20248 39782 20282 39844
rect 25256 39782 25290 39844
rect 20248 39748 20344 39782
rect 25194 39748 25290 39782
rect 1348 39134 1444 39168
rect 6294 39134 6390 39168
rect 1348 39072 1382 39134
rect 6356 39072 6390 39134
rect 1528 38996 1544 39030
rect 1612 38996 1628 39030
rect 1686 38996 1702 39030
rect 1770 38996 1786 39030
rect 1844 38996 1860 39030
rect 1928 38996 1944 39030
rect 2002 38996 2018 39030
rect 2086 38996 2102 39030
rect 2160 38996 2176 39030
rect 2244 38996 2260 39030
rect 2318 38996 2334 39030
rect 2402 38996 2418 39030
rect 2476 38996 2492 39030
rect 2560 38996 2576 39030
rect 2634 38996 2650 39030
rect 2718 38996 2734 39030
rect 2792 38996 2808 39030
rect 2876 38996 2892 39030
rect 2950 38996 2966 39030
rect 3034 38996 3050 39030
rect 3108 38996 3124 39030
rect 3192 38996 3208 39030
rect 3266 38996 3282 39030
rect 3350 38996 3366 39030
rect 3424 38996 3440 39030
rect 3508 38996 3524 39030
rect 3582 38996 3598 39030
rect 3666 38996 3682 39030
rect 3740 38996 3756 39030
rect 3824 38996 3840 39030
rect 3898 38996 3914 39030
rect 3982 38996 3998 39030
rect 4056 38996 4072 39030
rect 4140 38996 4156 39030
rect 4214 38996 4230 39030
rect 4298 38996 4314 39030
rect 4372 38996 4388 39030
rect 4456 38996 4472 39030
rect 4530 38996 4546 39030
rect 4614 38996 4630 39030
rect 4688 38996 4704 39030
rect 4772 38996 4788 39030
rect 4846 38996 4862 39030
rect 4930 38996 4946 39030
rect 5004 38996 5020 39030
rect 5088 38996 5104 39030
rect 5162 38996 5178 39030
rect 5246 38996 5262 39030
rect 5320 38996 5336 39030
rect 5404 38996 5420 39030
rect 5478 38996 5494 39030
rect 5562 38996 5578 39030
rect 5636 38996 5652 39030
rect 5720 38996 5736 39030
rect 5794 38996 5810 39030
rect 5878 38996 5894 39030
rect 5952 38996 5968 39030
rect 6036 38996 6052 39030
rect 6110 38996 6126 39030
rect 6194 38996 6210 39030
rect 7648 39134 7744 39168
rect 12594 39134 12690 39168
rect 7648 39072 7682 39134
rect 12656 39072 12690 39134
rect 7828 38996 7844 39030
rect 7912 38996 7928 39030
rect 7986 38996 8002 39030
rect 8070 38996 8086 39030
rect 8144 38996 8160 39030
rect 8228 38996 8244 39030
rect 8302 38996 8318 39030
rect 8386 38996 8402 39030
rect 8460 38996 8476 39030
rect 8544 38996 8560 39030
rect 8618 38996 8634 39030
rect 8702 38996 8718 39030
rect 8776 38996 8792 39030
rect 8860 38996 8876 39030
rect 8934 38996 8950 39030
rect 9018 38996 9034 39030
rect 9092 38996 9108 39030
rect 9176 38996 9192 39030
rect 9250 38996 9266 39030
rect 9334 38996 9350 39030
rect 9408 38996 9424 39030
rect 9492 38996 9508 39030
rect 9566 38996 9582 39030
rect 9650 38996 9666 39030
rect 9724 38996 9740 39030
rect 9808 38996 9824 39030
rect 9882 38996 9898 39030
rect 9966 38996 9982 39030
rect 10040 38996 10056 39030
rect 10124 38996 10140 39030
rect 10198 38996 10214 39030
rect 10282 38996 10298 39030
rect 10356 38996 10372 39030
rect 10440 38996 10456 39030
rect 10514 38996 10530 39030
rect 10598 38996 10614 39030
rect 10672 38996 10688 39030
rect 10756 38996 10772 39030
rect 10830 38996 10846 39030
rect 10914 38996 10930 39030
rect 10988 38996 11004 39030
rect 11072 38996 11088 39030
rect 11146 38996 11162 39030
rect 11230 38996 11246 39030
rect 11304 38996 11320 39030
rect 11388 38996 11404 39030
rect 11462 38996 11478 39030
rect 11546 38996 11562 39030
rect 11620 38996 11636 39030
rect 11704 38996 11720 39030
rect 11778 38996 11794 39030
rect 11862 38996 11878 39030
rect 11936 38996 11952 39030
rect 12020 38996 12036 39030
rect 12094 38996 12110 39030
rect 12178 38996 12194 39030
rect 12252 38996 12268 39030
rect 12336 38996 12352 39030
rect 12410 38996 12426 39030
rect 12494 38996 12510 39030
rect 13948 39134 14044 39168
rect 18894 39134 18990 39168
rect 13948 39072 13982 39134
rect 18956 39072 18990 39134
rect 14128 38996 14144 39030
rect 14212 38996 14228 39030
rect 14286 38996 14302 39030
rect 14370 38996 14386 39030
rect 14444 38996 14460 39030
rect 14528 38996 14544 39030
rect 14602 38996 14618 39030
rect 14686 38996 14702 39030
rect 14760 38996 14776 39030
rect 14844 38996 14860 39030
rect 14918 38996 14934 39030
rect 15002 38996 15018 39030
rect 15076 38996 15092 39030
rect 15160 38996 15176 39030
rect 15234 38996 15250 39030
rect 15318 38996 15334 39030
rect 15392 38996 15408 39030
rect 15476 38996 15492 39030
rect 15550 38996 15566 39030
rect 15634 38996 15650 39030
rect 15708 38996 15724 39030
rect 15792 38996 15808 39030
rect 15866 38996 15882 39030
rect 15950 38996 15966 39030
rect 16024 38996 16040 39030
rect 16108 38996 16124 39030
rect 16182 38996 16198 39030
rect 16266 38996 16282 39030
rect 16340 38996 16356 39030
rect 16424 38996 16440 39030
rect 16498 38996 16514 39030
rect 16582 38996 16598 39030
rect 16656 38996 16672 39030
rect 16740 38996 16756 39030
rect 16814 38996 16830 39030
rect 16898 38996 16914 39030
rect 16972 38996 16988 39030
rect 17056 38996 17072 39030
rect 17130 38996 17146 39030
rect 17214 38996 17230 39030
rect 17288 38996 17304 39030
rect 17372 38996 17388 39030
rect 17446 38996 17462 39030
rect 17530 38996 17546 39030
rect 17604 38996 17620 39030
rect 17688 38996 17704 39030
rect 17762 38996 17778 39030
rect 17846 38996 17862 39030
rect 17920 38996 17936 39030
rect 18004 38996 18020 39030
rect 18078 38996 18094 39030
rect 18162 38996 18178 39030
rect 18236 38996 18252 39030
rect 18320 38996 18336 39030
rect 18394 38996 18410 39030
rect 18478 38996 18494 39030
rect 18552 38996 18568 39030
rect 18636 38996 18652 39030
rect 18710 38996 18726 39030
rect 18794 38996 18810 39030
rect 20248 39134 20344 39168
rect 25194 39134 25290 39168
rect 20248 39072 20282 39134
rect 25256 39072 25290 39134
rect 20428 38996 20444 39030
rect 20512 38996 20528 39030
rect 20586 38996 20602 39030
rect 20670 38996 20686 39030
rect 20744 38996 20760 39030
rect 20828 38996 20844 39030
rect 20902 38996 20918 39030
rect 20986 38996 21002 39030
rect 21060 38996 21076 39030
rect 21144 38996 21160 39030
rect 21218 38996 21234 39030
rect 21302 38996 21318 39030
rect 21376 38996 21392 39030
rect 21460 38996 21476 39030
rect 21534 38996 21550 39030
rect 21618 38996 21634 39030
rect 21692 38996 21708 39030
rect 21776 38996 21792 39030
rect 21850 38996 21866 39030
rect 21934 38996 21950 39030
rect 22008 38996 22024 39030
rect 22092 38996 22108 39030
rect 22166 38996 22182 39030
rect 22250 38996 22266 39030
rect 22324 38996 22340 39030
rect 22408 38996 22424 39030
rect 22482 38996 22498 39030
rect 22566 38996 22582 39030
rect 22640 38996 22656 39030
rect 22724 38996 22740 39030
rect 22798 38996 22814 39030
rect 22882 38996 22898 39030
rect 22956 38996 22972 39030
rect 23040 38996 23056 39030
rect 23114 38996 23130 39030
rect 23198 38996 23214 39030
rect 23272 38996 23288 39030
rect 23356 38996 23372 39030
rect 23430 38996 23446 39030
rect 23514 38996 23530 39030
rect 23588 38996 23604 39030
rect 23672 38996 23688 39030
rect 23746 38996 23762 39030
rect 23830 38996 23846 39030
rect 23904 38996 23920 39030
rect 23988 38996 24004 39030
rect 24062 38996 24078 39030
rect 24146 38996 24162 39030
rect 24220 38996 24236 39030
rect 24304 38996 24320 39030
rect 24378 38996 24394 39030
rect 24462 38996 24478 39030
rect 24536 38996 24552 39030
rect 24620 38996 24636 39030
rect 24694 38996 24710 39030
rect 24778 38996 24794 39030
rect 24852 38996 24868 39030
rect 24936 38996 24952 39030
rect 25010 38996 25026 39030
rect 25094 38996 25110 39030
rect -3134 38720 -2980 38740
rect -3134 38716 -3038 38720
rect 1482 38946 1516 38962
rect 1482 32954 1516 32970
rect 1640 38946 1674 38962
rect 1640 32954 1674 32970
rect 1798 38946 1832 38962
rect 1798 32954 1832 32970
rect 1956 38946 1990 38962
rect 1956 32954 1990 32970
rect 2114 38946 2148 38962
rect 2114 32954 2148 32970
rect 2272 38946 2306 38962
rect 2272 32954 2306 32970
rect 2430 38946 2464 38962
rect 2430 32954 2464 32970
rect 2588 38946 2622 38962
rect 2588 32954 2622 32970
rect 2746 38946 2780 38962
rect 2746 32954 2780 32970
rect 2904 38946 2938 38962
rect 2904 32954 2938 32970
rect 3062 38946 3096 38962
rect 3062 32954 3096 32970
rect 3220 38946 3254 38962
rect 3220 32954 3254 32970
rect 3378 38946 3412 38962
rect 3378 32954 3412 32970
rect 3536 38946 3570 38962
rect 3536 32954 3570 32970
rect 3694 38946 3728 38962
rect 3694 32954 3728 32970
rect 3852 38946 3886 38962
rect 3852 32954 3886 32970
rect 4010 38946 4044 38962
rect 4010 32954 4044 32970
rect 4168 38946 4202 38962
rect 4168 32954 4202 32970
rect 4326 38946 4360 38962
rect 4326 32954 4360 32970
rect 4484 38946 4518 38962
rect 4484 32954 4518 32970
rect 4642 38946 4676 38962
rect 4642 32954 4676 32970
rect 4800 38946 4834 38962
rect 4800 32954 4834 32970
rect 4958 38946 4992 38962
rect 4958 32954 4992 32970
rect 5116 38946 5150 38962
rect 5116 32954 5150 32970
rect 5274 38946 5308 38962
rect 5274 32954 5308 32970
rect 5432 38946 5466 38962
rect 5432 32954 5466 32970
rect 5590 38946 5624 38962
rect 5590 32954 5624 32970
rect 5748 38946 5782 38962
rect 5748 32954 5782 32970
rect 5906 38946 5940 38962
rect 5906 32954 5940 32970
rect 6064 38946 6098 38962
rect 6064 32954 6098 32970
rect 6222 38946 6256 38962
rect 6222 32954 6256 32970
rect 7782 38946 7816 38962
rect 7782 32954 7816 32970
rect 7940 38946 7974 38962
rect 7940 32954 7974 32970
rect 8098 38946 8132 38962
rect 8098 32954 8132 32970
rect 8256 38946 8290 38962
rect 8256 32954 8290 32970
rect 8414 38946 8448 38962
rect 8414 32954 8448 32970
rect 8572 38946 8606 38962
rect 8572 32954 8606 32970
rect 8730 38946 8764 38962
rect 8730 32954 8764 32970
rect 8888 38946 8922 38962
rect 8888 32954 8922 32970
rect 9046 38946 9080 38962
rect 9046 32954 9080 32970
rect 9204 38946 9238 38962
rect 9204 32954 9238 32970
rect 9362 38946 9396 38962
rect 9362 32954 9396 32970
rect 9520 38946 9554 38962
rect 9520 32954 9554 32970
rect 9678 38946 9712 38962
rect 9678 32954 9712 32970
rect 9836 38946 9870 38962
rect 9836 32954 9870 32970
rect 9994 38946 10028 38962
rect 9994 32954 10028 32970
rect 10152 38946 10186 38962
rect 10152 32954 10186 32970
rect 10310 38946 10344 38962
rect 10310 32954 10344 32970
rect 10468 38946 10502 38962
rect 10468 32954 10502 32970
rect 10626 38946 10660 38962
rect 10626 32954 10660 32970
rect 10784 38946 10818 38962
rect 10784 32954 10818 32970
rect 10942 38946 10976 38962
rect 10942 32954 10976 32970
rect 11100 38946 11134 38962
rect 11100 32954 11134 32970
rect 11258 38946 11292 38962
rect 11258 32954 11292 32970
rect 11416 38946 11450 38962
rect 11416 32954 11450 32970
rect 11574 38946 11608 38962
rect 11574 32954 11608 32970
rect 11732 38946 11766 38962
rect 11732 32954 11766 32970
rect 11890 38946 11924 38962
rect 11890 32954 11924 32970
rect 12048 38946 12082 38962
rect 12048 32954 12082 32970
rect 12206 38946 12240 38962
rect 12206 32954 12240 32970
rect 12364 38946 12398 38962
rect 12364 32954 12398 32970
rect 12522 38946 12556 38962
rect 12522 32954 12556 32970
rect 14082 38946 14116 38962
rect 14082 32954 14116 32970
rect 14240 38946 14274 38962
rect 14240 32954 14274 32970
rect 14398 38946 14432 38962
rect 14398 32954 14432 32970
rect 14556 38946 14590 38962
rect 14556 32954 14590 32970
rect 14714 38946 14748 38962
rect 14714 32954 14748 32970
rect 14872 38946 14906 38962
rect 14872 32954 14906 32970
rect 15030 38946 15064 38962
rect 15030 32954 15064 32970
rect 15188 38946 15222 38962
rect 15188 32954 15222 32970
rect 15346 38946 15380 38962
rect 15346 32954 15380 32970
rect 15504 38946 15538 38962
rect 15504 32954 15538 32970
rect 15662 38946 15696 38962
rect 15662 32954 15696 32970
rect 15820 38946 15854 38962
rect 15820 32954 15854 32970
rect 15978 38946 16012 38962
rect 15978 32954 16012 32970
rect 16136 38946 16170 38962
rect 16136 32954 16170 32970
rect 16294 38946 16328 38962
rect 16294 32954 16328 32970
rect 16452 38946 16486 38962
rect 16452 32954 16486 32970
rect 16610 38946 16644 38962
rect 16610 32954 16644 32970
rect 16768 38946 16802 38962
rect 16768 32954 16802 32970
rect 16926 38946 16960 38962
rect 16926 32954 16960 32970
rect 17084 38946 17118 38962
rect 17084 32954 17118 32970
rect 17242 38946 17276 38962
rect 17242 32954 17276 32970
rect 17400 38946 17434 38962
rect 17400 32954 17434 32970
rect 17558 38946 17592 38962
rect 17558 32954 17592 32970
rect 17716 38946 17750 38962
rect 17716 32954 17750 32970
rect 17874 38946 17908 38962
rect 17874 32954 17908 32970
rect 18032 38946 18066 38962
rect 18032 32954 18066 32970
rect 18190 38946 18224 38962
rect 18190 32954 18224 32970
rect 18348 38946 18382 38962
rect 18348 32954 18382 32970
rect 18506 38946 18540 38962
rect 18506 32954 18540 32970
rect 18664 38946 18698 38962
rect 18664 32954 18698 32970
rect 18822 38946 18856 38962
rect 18822 32954 18856 32970
rect 20382 38946 20416 38962
rect 20382 32954 20416 32970
rect 20540 38946 20574 38962
rect 20540 32954 20574 32970
rect 20698 38946 20732 38962
rect 20698 32954 20732 32970
rect 20856 38946 20890 38962
rect 20856 32954 20890 32970
rect 21014 38946 21048 38962
rect 21014 32954 21048 32970
rect 21172 38946 21206 38962
rect 21172 32954 21206 32970
rect 21330 38946 21364 38962
rect 21330 32954 21364 32970
rect 21488 38946 21522 38962
rect 21488 32954 21522 32970
rect 21646 38946 21680 38962
rect 21646 32954 21680 32970
rect 21804 38946 21838 38962
rect 21804 32954 21838 32970
rect 21962 38946 21996 38962
rect 21962 32954 21996 32970
rect 22120 38946 22154 38962
rect 22120 32954 22154 32970
rect 22278 38946 22312 38962
rect 22278 32954 22312 32970
rect 22436 38946 22470 38962
rect 22436 32954 22470 32970
rect 22594 38946 22628 38962
rect 22594 32954 22628 32970
rect 22752 38946 22786 38962
rect 22752 32954 22786 32970
rect 22910 38946 22944 38962
rect 22910 32954 22944 32970
rect 23068 38946 23102 38962
rect 23068 32954 23102 32970
rect 23226 38946 23260 38962
rect 23226 32954 23260 32970
rect 23384 38946 23418 38962
rect 23384 32954 23418 32970
rect 23542 38946 23576 38962
rect 23542 32954 23576 32970
rect 23700 38946 23734 38962
rect 23700 32954 23734 32970
rect 23858 38946 23892 38962
rect 23858 32954 23892 32970
rect 24016 38946 24050 38962
rect 24016 32954 24050 32970
rect 24174 38946 24208 38962
rect 24174 32954 24208 32970
rect 24332 38946 24366 38962
rect 24332 32954 24366 32970
rect 24490 38946 24524 38962
rect 24490 32954 24524 32970
rect 24648 38946 24682 38962
rect 24648 32954 24682 32970
rect 24806 38946 24840 38962
rect 24806 32954 24840 32970
rect 24964 38946 24998 38962
rect 24964 32954 24998 32970
rect 25122 38946 25156 38962
rect 25122 32954 25156 32970
rect 29780 38720 29800 40400
rect 29840 40388 29934 40400
rect 30068 40388 30164 40422
rect 29840 40326 29872 40388
rect 30130 40326 30164 40388
rect 29968 40242 29984 40276
rect 30018 40242 30034 40276
rect 29968 38862 29984 38896
rect 30018 38862 30034 38896
rect 29840 38750 29872 38812
rect 30130 38750 30164 38812
rect 29840 38720 29934 38750
rect 29780 38716 29934 38720
rect 30068 38716 30164 38750
rect 29780 38700 29860 38716
rect 1528 32886 1544 32920
rect 1612 32886 1628 32920
rect 1686 32886 1702 32920
rect 1770 32886 1786 32920
rect 1844 32886 1860 32920
rect 1928 32886 1944 32920
rect 2002 32886 2018 32920
rect 2086 32886 2102 32920
rect 2160 32886 2176 32920
rect 2244 32886 2260 32920
rect 2318 32886 2334 32920
rect 2402 32886 2418 32920
rect 2476 32886 2492 32920
rect 2560 32886 2576 32920
rect 2634 32886 2650 32920
rect 2718 32886 2734 32920
rect 2792 32886 2808 32920
rect 2876 32886 2892 32920
rect 2950 32886 2966 32920
rect 3034 32886 3050 32920
rect 3108 32886 3124 32920
rect 3192 32886 3208 32920
rect 3266 32886 3282 32920
rect 3350 32886 3366 32920
rect 3424 32886 3440 32920
rect 3508 32886 3524 32920
rect 3582 32886 3598 32920
rect 3666 32886 3682 32920
rect 3740 32886 3756 32920
rect 3824 32886 3840 32920
rect 3898 32886 3914 32920
rect 3982 32886 3998 32920
rect 4056 32886 4072 32920
rect 4140 32886 4156 32920
rect 4214 32886 4230 32920
rect 4298 32886 4314 32920
rect 4372 32886 4388 32920
rect 4456 32886 4472 32920
rect 4530 32886 4546 32920
rect 4614 32886 4630 32920
rect 4688 32886 4704 32920
rect 4772 32886 4788 32920
rect 4846 32886 4862 32920
rect 4930 32886 4946 32920
rect 5004 32886 5020 32920
rect 5088 32886 5104 32920
rect 5162 32886 5178 32920
rect 5246 32886 5262 32920
rect 5320 32886 5336 32920
rect 5404 32886 5420 32920
rect 5478 32886 5494 32920
rect 5562 32886 5578 32920
rect 5636 32886 5652 32920
rect 5720 32886 5736 32920
rect 5794 32886 5810 32920
rect 5878 32886 5894 32920
rect 5952 32886 5968 32920
rect 6036 32886 6052 32920
rect 6110 32886 6126 32920
rect 6194 32886 6210 32920
rect 1348 32782 1382 32844
rect 6356 32782 6390 32844
rect 1348 32748 1444 32782
rect 6294 32748 6390 32782
rect 7828 32886 7844 32920
rect 7912 32886 7928 32920
rect 7986 32886 8002 32920
rect 8070 32886 8086 32920
rect 8144 32886 8160 32920
rect 8228 32886 8244 32920
rect 8302 32886 8318 32920
rect 8386 32886 8402 32920
rect 8460 32886 8476 32920
rect 8544 32886 8560 32920
rect 8618 32886 8634 32920
rect 8702 32886 8718 32920
rect 8776 32886 8792 32920
rect 8860 32886 8876 32920
rect 8934 32886 8950 32920
rect 9018 32886 9034 32920
rect 9092 32886 9108 32920
rect 9176 32886 9192 32920
rect 9250 32886 9266 32920
rect 9334 32886 9350 32920
rect 9408 32886 9424 32920
rect 9492 32886 9508 32920
rect 9566 32886 9582 32920
rect 9650 32886 9666 32920
rect 9724 32886 9740 32920
rect 9808 32886 9824 32920
rect 9882 32886 9898 32920
rect 9966 32886 9982 32920
rect 10040 32886 10056 32920
rect 10124 32886 10140 32920
rect 10198 32886 10214 32920
rect 10282 32886 10298 32920
rect 10356 32886 10372 32920
rect 10440 32886 10456 32920
rect 10514 32886 10530 32920
rect 10598 32886 10614 32920
rect 10672 32886 10688 32920
rect 10756 32886 10772 32920
rect 10830 32886 10846 32920
rect 10914 32886 10930 32920
rect 10988 32886 11004 32920
rect 11072 32886 11088 32920
rect 11146 32886 11162 32920
rect 11230 32886 11246 32920
rect 11304 32886 11320 32920
rect 11388 32886 11404 32920
rect 11462 32886 11478 32920
rect 11546 32886 11562 32920
rect 11620 32886 11636 32920
rect 11704 32886 11720 32920
rect 11778 32886 11794 32920
rect 11862 32886 11878 32920
rect 11936 32886 11952 32920
rect 12020 32886 12036 32920
rect 12094 32886 12110 32920
rect 12178 32886 12194 32920
rect 12252 32886 12268 32920
rect 12336 32886 12352 32920
rect 12410 32886 12426 32920
rect 12494 32886 12510 32920
rect 7648 32782 7682 32844
rect 12656 32782 12690 32844
rect 7648 32748 7744 32782
rect 12594 32748 12690 32782
rect 14128 32886 14144 32920
rect 14212 32886 14228 32920
rect 14286 32886 14302 32920
rect 14370 32886 14386 32920
rect 14444 32886 14460 32920
rect 14528 32886 14544 32920
rect 14602 32886 14618 32920
rect 14686 32886 14702 32920
rect 14760 32886 14776 32920
rect 14844 32886 14860 32920
rect 14918 32886 14934 32920
rect 15002 32886 15018 32920
rect 15076 32886 15092 32920
rect 15160 32886 15176 32920
rect 15234 32886 15250 32920
rect 15318 32886 15334 32920
rect 15392 32886 15408 32920
rect 15476 32886 15492 32920
rect 15550 32886 15566 32920
rect 15634 32886 15650 32920
rect 15708 32886 15724 32920
rect 15792 32886 15808 32920
rect 15866 32886 15882 32920
rect 15950 32886 15966 32920
rect 16024 32886 16040 32920
rect 16108 32886 16124 32920
rect 16182 32886 16198 32920
rect 16266 32886 16282 32920
rect 16340 32886 16356 32920
rect 16424 32886 16440 32920
rect 16498 32886 16514 32920
rect 16582 32886 16598 32920
rect 16656 32886 16672 32920
rect 16740 32886 16756 32920
rect 16814 32886 16830 32920
rect 16898 32886 16914 32920
rect 16972 32886 16988 32920
rect 17056 32886 17072 32920
rect 17130 32886 17146 32920
rect 17214 32886 17230 32920
rect 17288 32886 17304 32920
rect 17372 32886 17388 32920
rect 17446 32886 17462 32920
rect 17530 32886 17546 32920
rect 17604 32886 17620 32920
rect 17688 32886 17704 32920
rect 17762 32886 17778 32920
rect 17846 32886 17862 32920
rect 17920 32886 17936 32920
rect 18004 32886 18020 32920
rect 18078 32886 18094 32920
rect 18162 32886 18178 32920
rect 18236 32886 18252 32920
rect 18320 32886 18336 32920
rect 18394 32886 18410 32920
rect 18478 32886 18494 32920
rect 18552 32886 18568 32920
rect 18636 32886 18652 32920
rect 18710 32886 18726 32920
rect 18794 32886 18810 32920
rect 13948 32782 13982 32844
rect 18956 32782 18990 32844
rect 13948 32748 14044 32782
rect 18894 32748 18990 32782
rect 20428 32886 20444 32920
rect 20512 32886 20528 32920
rect 20586 32886 20602 32920
rect 20670 32886 20686 32920
rect 20744 32886 20760 32920
rect 20828 32886 20844 32920
rect 20902 32886 20918 32920
rect 20986 32886 21002 32920
rect 21060 32886 21076 32920
rect 21144 32886 21160 32920
rect 21218 32886 21234 32920
rect 21302 32886 21318 32920
rect 21376 32886 21392 32920
rect 21460 32886 21476 32920
rect 21534 32886 21550 32920
rect 21618 32886 21634 32920
rect 21692 32886 21708 32920
rect 21776 32886 21792 32920
rect 21850 32886 21866 32920
rect 21934 32886 21950 32920
rect 22008 32886 22024 32920
rect 22092 32886 22108 32920
rect 22166 32886 22182 32920
rect 22250 32886 22266 32920
rect 22324 32886 22340 32920
rect 22408 32886 22424 32920
rect 22482 32886 22498 32920
rect 22566 32886 22582 32920
rect 22640 32886 22656 32920
rect 22724 32886 22740 32920
rect 22798 32886 22814 32920
rect 22882 32886 22898 32920
rect 22956 32886 22972 32920
rect 23040 32886 23056 32920
rect 23114 32886 23130 32920
rect 23198 32886 23214 32920
rect 23272 32886 23288 32920
rect 23356 32886 23372 32920
rect 23430 32886 23446 32920
rect 23514 32886 23530 32920
rect 23588 32886 23604 32920
rect 23672 32886 23688 32920
rect 23746 32886 23762 32920
rect 23830 32886 23846 32920
rect 23904 32886 23920 32920
rect 23988 32886 24004 32920
rect 24062 32886 24078 32920
rect 24146 32886 24162 32920
rect 24220 32886 24236 32920
rect 24304 32886 24320 32920
rect 24378 32886 24394 32920
rect 24462 32886 24478 32920
rect 24536 32886 24552 32920
rect 24620 32886 24636 32920
rect 24694 32886 24710 32920
rect 24778 32886 24794 32920
rect 24852 32886 24868 32920
rect 24936 32886 24952 32920
rect 25010 32886 25026 32920
rect 25094 32886 25110 32920
rect 20248 32782 20282 32844
rect 25256 32782 25290 32844
rect 20248 32748 20344 32782
rect 25194 32748 25290 32782
rect 1348 30834 1444 30868
rect 6294 30834 6390 30868
rect 1348 30772 1382 30834
rect 6356 30772 6390 30834
rect 1528 30696 1544 30730
rect 1612 30696 1628 30730
rect 1686 30696 1702 30730
rect 1770 30696 1786 30730
rect 1844 30696 1860 30730
rect 1928 30696 1944 30730
rect 2002 30696 2018 30730
rect 2086 30696 2102 30730
rect 2160 30696 2176 30730
rect 2244 30696 2260 30730
rect 2318 30696 2334 30730
rect 2402 30696 2418 30730
rect 2476 30696 2492 30730
rect 2560 30696 2576 30730
rect 2634 30696 2650 30730
rect 2718 30696 2734 30730
rect 2792 30696 2808 30730
rect 2876 30696 2892 30730
rect 2950 30696 2966 30730
rect 3034 30696 3050 30730
rect 3108 30696 3124 30730
rect 3192 30696 3208 30730
rect 3266 30696 3282 30730
rect 3350 30696 3366 30730
rect 3424 30696 3440 30730
rect 3508 30696 3524 30730
rect 3582 30696 3598 30730
rect 3666 30696 3682 30730
rect 3740 30696 3756 30730
rect 3824 30696 3840 30730
rect 3898 30696 3914 30730
rect 3982 30696 3998 30730
rect 4056 30696 4072 30730
rect 4140 30696 4156 30730
rect 4214 30696 4230 30730
rect 4298 30696 4314 30730
rect 4372 30696 4388 30730
rect 4456 30696 4472 30730
rect 4530 30696 4546 30730
rect 4614 30696 4630 30730
rect 4688 30696 4704 30730
rect 4772 30696 4788 30730
rect 4846 30696 4862 30730
rect 4930 30696 4946 30730
rect 5004 30696 5020 30730
rect 5088 30696 5104 30730
rect 5162 30696 5178 30730
rect 5246 30696 5262 30730
rect 5320 30696 5336 30730
rect 5404 30696 5420 30730
rect 5478 30696 5494 30730
rect 5562 30696 5578 30730
rect 5636 30696 5652 30730
rect 5720 30696 5736 30730
rect 5794 30696 5810 30730
rect 5878 30696 5894 30730
rect 5952 30696 5968 30730
rect 6036 30696 6052 30730
rect 6110 30696 6126 30730
rect 6194 30696 6210 30730
rect 7648 30834 7744 30868
rect 12594 30834 12690 30868
rect 7648 30772 7682 30834
rect 12656 30772 12690 30834
rect 7828 30696 7844 30730
rect 7912 30696 7928 30730
rect 7986 30696 8002 30730
rect 8070 30696 8086 30730
rect 8144 30696 8160 30730
rect 8228 30696 8244 30730
rect 8302 30696 8318 30730
rect 8386 30696 8402 30730
rect 8460 30696 8476 30730
rect 8544 30696 8560 30730
rect 8618 30696 8634 30730
rect 8702 30696 8718 30730
rect 8776 30696 8792 30730
rect 8860 30696 8876 30730
rect 8934 30696 8950 30730
rect 9018 30696 9034 30730
rect 9092 30696 9108 30730
rect 9176 30696 9192 30730
rect 9250 30696 9266 30730
rect 9334 30696 9350 30730
rect 9408 30696 9424 30730
rect 9492 30696 9508 30730
rect 9566 30696 9582 30730
rect 9650 30696 9666 30730
rect 9724 30696 9740 30730
rect 9808 30696 9824 30730
rect 9882 30696 9898 30730
rect 9966 30696 9982 30730
rect 10040 30696 10056 30730
rect 10124 30696 10140 30730
rect 10198 30696 10214 30730
rect 10282 30696 10298 30730
rect 10356 30696 10372 30730
rect 10440 30696 10456 30730
rect 10514 30696 10530 30730
rect 10598 30696 10614 30730
rect 10672 30696 10688 30730
rect 10756 30696 10772 30730
rect 10830 30696 10846 30730
rect 10914 30696 10930 30730
rect 10988 30696 11004 30730
rect 11072 30696 11088 30730
rect 11146 30696 11162 30730
rect 11230 30696 11246 30730
rect 11304 30696 11320 30730
rect 11388 30696 11404 30730
rect 11462 30696 11478 30730
rect 11546 30696 11562 30730
rect 11620 30696 11636 30730
rect 11704 30696 11720 30730
rect 11778 30696 11794 30730
rect 11862 30696 11878 30730
rect 11936 30696 11952 30730
rect 12020 30696 12036 30730
rect 12094 30696 12110 30730
rect 12178 30696 12194 30730
rect 12252 30696 12268 30730
rect 12336 30696 12352 30730
rect 12410 30696 12426 30730
rect 12494 30696 12510 30730
rect 13948 30834 14044 30868
rect 18894 30834 18990 30868
rect 13948 30772 13982 30834
rect 18956 30772 18990 30834
rect 14128 30696 14144 30730
rect 14212 30696 14228 30730
rect 14286 30696 14302 30730
rect 14370 30696 14386 30730
rect 14444 30696 14460 30730
rect 14528 30696 14544 30730
rect 14602 30696 14618 30730
rect 14686 30696 14702 30730
rect 14760 30696 14776 30730
rect 14844 30696 14860 30730
rect 14918 30696 14934 30730
rect 15002 30696 15018 30730
rect 15076 30696 15092 30730
rect 15160 30696 15176 30730
rect 15234 30696 15250 30730
rect 15318 30696 15334 30730
rect 15392 30696 15408 30730
rect 15476 30696 15492 30730
rect 15550 30696 15566 30730
rect 15634 30696 15650 30730
rect 15708 30696 15724 30730
rect 15792 30696 15808 30730
rect 15866 30696 15882 30730
rect 15950 30696 15966 30730
rect 16024 30696 16040 30730
rect 16108 30696 16124 30730
rect 16182 30696 16198 30730
rect 16266 30696 16282 30730
rect 16340 30696 16356 30730
rect 16424 30696 16440 30730
rect 16498 30696 16514 30730
rect 16582 30696 16598 30730
rect 16656 30696 16672 30730
rect 16740 30696 16756 30730
rect 16814 30696 16830 30730
rect 16898 30696 16914 30730
rect 16972 30696 16988 30730
rect 17056 30696 17072 30730
rect 17130 30696 17146 30730
rect 17214 30696 17230 30730
rect 17288 30696 17304 30730
rect 17372 30696 17388 30730
rect 17446 30696 17462 30730
rect 17530 30696 17546 30730
rect 17604 30696 17620 30730
rect 17688 30696 17704 30730
rect 17762 30696 17778 30730
rect 17846 30696 17862 30730
rect 17920 30696 17936 30730
rect 18004 30696 18020 30730
rect 18078 30696 18094 30730
rect 18162 30696 18178 30730
rect 18236 30696 18252 30730
rect 18320 30696 18336 30730
rect 18394 30696 18410 30730
rect 18478 30696 18494 30730
rect 18552 30696 18568 30730
rect 18636 30696 18652 30730
rect 18710 30696 18726 30730
rect 18794 30696 18810 30730
rect 20248 30834 20344 30868
rect 25194 30834 25290 30868
rect 20248 30772 20282 30834
rect 25256 30772 25290 30834
rect 20428 30696 20444 30730
rect 20512 30696 20528 30730
rect 20586 30696 20602 30730
rect 20670 30696 20686 30730
rect 20744 30696 20760 30730
rect 20828 30696 20844 30730
rect 20902 30696 20918 30730
rect 20986 30696 21002 30730
rect 21060 30696 21076 30730
rect 21144 30696 21160 30730
rect 21218 30696 21234 30730
rect 21302 30696 21318 30730
rect 21376 30696 21392 30730
rect 21460 30696 21476 30730
rect 21534 30696 21550 30730
rect 21618 30696 21634 30730
rect 21692 30696 21708 30730
rect 21776 30696 21792 30730
rect 21850 30696 21866 30730
rect 21934 30696 21950 30730
rect 22008 30696 22024 30730
rect 22092 30696 22108 30730
rect 22166 30696 22182 30730
rect 22250 30696 22266 30730
rect 22324 30696 22340 30730
rect 22408 30696 22424 30730
rect 22482 30696 22498 30730
rect 22566 30696 22582 30730
rect 22640 30696 22656 30730
rect 22724 30696 22740 30730
rect 22798 30696 22814 30730
rect 22882 30696 22898 30730
rect 22956 30696 22972 30730
rect 23040 30696 23056 30730
rect 23114 30696 23130 30730
rect 23198 30696 23214 30730
rect 23272 30696 23288 30730
rect 23356 30696 23372 30730
rect 23430 30696 23446 30730
rect 23514 30696 23530 30730
rect 23588 30696 23604 30730
rect 23672 30696 23688 30730
rect 23746 30696 23762 30730
rect 23830 30696 23846 30730
rect 23904 30696 23920 30730
rect 23988 30696 24004 30730
rect 24062 30696 24078 30730
rect 24146 30696 24162 30730
rect 24220 30696 24236 30730
rect 24304 30696 24320 30730
rect 24378 30696 24394 30730
rect 24462 30696 24478 30730
rect 24536 30696 24552 30730
rect 24620 30696 24636 30730
rect 24694 30696 24710 30730
rect 24778 30696 24794 30730
rect 24852 30696 24868 30730
rect 24936 30696 24952 30730
rect 25010 30696 25026 30730
rect 25094 30696 25110 30730
rect -4364 27188 -4268 27222
rect -4134 27220 -4038 27222
rect -4134 27200 -3980 27220
rect -4134 27188 -4040 27200
rect -4364 27126 -4330 27188
rect -4072 27126 -4040 27188
rect -4234 27042 -4218 27076
rect -4184 27042 -4168 27076
rect -4234 25662 -4218 25696
rect -4184 25662 -4168 25696
rect -4364 25550 -4330 25612
rect -4072 25550 -4040 25612
rect -4364 25516 -4268 25550
rect -4134 25540 -4040 25550
rect -4000 25540 -3980 27200
rect -4134 25520 -3980 25540
rect -4134 25516 -4038 25520
rect 1482 30646 1516 30662
rect 1482 24654 1516 24670
rect 1640 30646 1674 30662
rect 1640 24654 1674 24670
rect 1798 30646 1832 30662
rect 1798 24654 1832 24670
rect 1956 30646 1990 30662
rect 1956 24654 1990 24670
rect 2114 30646 2148 30662
rect 2114 24654 2148 24670
rect 2272 30646 2306 30662
rect 2272 24654 2306 24670
rect 2430 30646 2464 30662
rect 2430 24654 2464 24670
rect 2588 30646 2622 30662
rect 2588 24654 2622 24670
rect 2746 30646 2780 30662
rect 2746 24654 2780 24670
rect 2904 30646 2938 30662
rect 2904 24654 2938 24670
rect 3062 30646 3096 30662
rect 3062 24654 3096 24670
rect 3220 30646 3254 30662
rect 3220 24654 3254 24670
rect 3378 30646 3412 30662
rect 3378 24654 3412 24670
rect 3536 30646 3570 30662
rect 3536 24654 3570 24670
rect 3694 30646 3728 30662
rect 3694 24654 3728 24670
rect 3852 30646 3886 30662
rect 3852 24654 3886 24670
rect 4010 30646 4044 30662
rect 4010 24654 4044 24670
rect 4168 30646 4202 30662
rect 4168 24654 4202 24670
rect 4326 30646 4360 30662
rect 4326 24654 4360 24670
rect 4484 30646 4518 30662
rect 4484 24654 4518 24670
rect 4642 30646 4676 30662
rect 4642 24654 4676 24670
rect 4800 30646 4834 30662
rect 4800 24654 4834 24670
rect 4958 30646 4992 30662
rect 4958 24654 4992 24670
rect 5116 30646 5150 30662
rect 5116 24654 5150 24670
rect 5274 30646 5308 30662
rect 5274 24654 5308 24670
rect 5432 30646 5466 30662
rect 5432 24654 5466 24670
rect 5590 30646 5624 30662
rect 5590 24654 5624 24670
rect 5748 30646 5782 30662
rect 5748 24654 5782 24670
rect 5906 30646 5940 30662
rect 5906 24654 5940 24670
rect 6064 30646 6098 30662
rect 6064 24654 6098 24670
rect 6222 30646 6256 30662
rect 6222 24654 6256 24670
rect 7782 30646 7816 30662
rect 7782 24654 7816 24670
rect 7940 30646 7974 30662
rect 7940 24654 7974 24670
rect 8098 30646 8132 30662
rect 8098 24654 8132 24670
rect 8256 30646 8290 30662
rect 8256 24654 8290 24670
rect 8414 30646 8448 30662
rect 8414 24654 8448 24670
rect 8572 30646 8606 30662
rect 8572 24654 8606 24670
rect 8730 30646 8764 30662
rect 8730 24654 8764 24670
rect 8888 30646 8922 30662
rect 8888 24654 8922 24670
rect 9046 30646 9080 30662
rect 9046 24654 9080 24670
rect 9204 30646 9238 30662
rect 9204 24654 9238 24670
rect 9362 30646 9396 30662
rect 9362 24654 9396 24670
rect 9520 30646 9554 30662
rect 9520 24654 9554 24670
rect 9678 30646 9712 30662
rect 9678 24654 9712 24670
rect 9836 30646 9870 30662
rect 9836 24654 9870 24670
rect 9994 30646 10028 30662
rect 9994 24654 10028 24670
rect 10152 30646 10186 30662
rect 10152 24654 10186 24670
rect 10310 30646 10344 30662
rect 10310 24654 10344 24670
rect 10468 30646 10502 30662
rect 10468 24654 10502 24670
rect 10626 30646 10660 30662
rect 10626 24654 10660 24670
rect 10784 30646 10818 30662
rect 10784 24654 10818 24670
rect 10942 30646 10976 30662
rect 10942 24654 10976 24670
rect 11100 30646 11134 30662
rect 11100 24654 11134 24670
rect 11258 30646 11292 30662
rect 11258 24654 11292 24670
rect 11416 30646 11450 30662
rect 11416 24654 11450 24670
rect 11574 30646 11608 30662
rect 11574 24654 11608 24670
rect 11732 30646 11766 30662
rect 11732 24654 11766 24670
rect 11890 30646 11924 30662
rect 11890 24654 11924 24670
rect 12048 30646 12082 30662
rect 12048 24654 12082 24670
rect 12206 30646 12240 30662
rect 12206 24654 12240 24670
rect 12364 30646 12398 30662
rect 12364 24654 12398 24670
rect 12522 30646 12556 30662
rect 12522 24654 12556 24670
rect 14082 30646 14116 30662
rect 14082 24654 14116 24670
rect 14240 30646 14274 30662
rect 14240 24654 14274 24670
rect 14398 30646 14432 30662
rect 14398 24654 14432 24670
rect 14556 30646 14590 30662
rect 14556 24654 14590 24670
rect 14714 30646 14748 30662
rect 14714 24654 14748 24670
rect 14872 30646 14906 30662
rect 14872 24654 14906 24670
rect 15030 30646 15064 30662
rect 15030 24654 15064 24670
rect 15188 30646 15222 30662
rect 15188 24654 15222 24670
rect 15346 30646 15380 30662
rect 15346 24654 15380 24670
rect 15504 30646 15538 30662
rect 15504 24654 15538 24670
rect 15662 30646 15696 30662
rect 15662 24654 15696 24670
rect 15820 30646 15854 30662
rect 15820 24654 15854 24670
rect 15978 30646 16012 30662
rect 15978 24654 16012 24670
rect 16136 30646 16170 30662
rect 16136 24654 16170 24670
rect 16294 30646 16328 30662
rect 16294 24654 16328 24670
rect 16452 30646 16486 30662
rect 16452 24654 16486 24670
rect 16610 30646 16644 30662
rect 16610 24654 16644 24670
rect 16768 30646 16802 30662
rect 16768 24654 16802 24670
rect 16926 30646 16960 30662
rect 16926 24654 16960 24670
rect 17084 30646 17118 30662
rect 17084 24654 17118 24670
rect 17242 30646 17276 30662
rect 17242 24654 17276 24670
rect 17400 30646 17434 30662
rect 17400 24654 17434 24670
rect 17558 30646 17592 30662
rect 17558 24654 17592 24670
rect 17716 30646 17750 30662
rect 17716 24654 17750 24670
rect 17874 30646 17908 30662
rect 17874 24654 17908 24670
rect 18032 30646 18066 30662
rect 18032 24654 18066 24670
rect 18190 30646 18224 30662
rect 18190 24654 18224 24670
rect 18348 30646 18382 30662
rect 18348 24654 18382 24670
rect 18506 30646 18540 30662
rect 18506 24654 18540 24670
rect 18664 30646 18698 30662
rect 18664 24654 18698 24670
rect 18822 30646 18856 30662
rect 18822 24654 18856 24670
rect 20382 30646 20416 30662
rect 20382 24654 20416 24670
rect 20540 30646 20574 30662
rect 20540 24654 20574 24670
rect 20698 30646 20732 30662
rect 20698 24654 20732 24670
rect 20856 30646 20890 30662
rect 20856 24654 20890 24670
rect 21014 30646 21048 30662
rect 21014 24654 21048 24670
rect 21172 30646 21206 30662
rect 21172 24654 21206 24670
rect 21330 30646 21364 30662
rect 21330 24654 21364 24670
rect 21488 30646 21522 30662
rect 21488 24654 21522 24670
rect 21646 30646 21680 30662
rect 21646 24654 21680 24670
rect 21804 30646 21838 30662
rect 21804 24654 21838 24670
rect 21962 30646 21996 30662
rect 21962 24654 21996 24670
rect 22120 30646 22154 30662
rect 22120 24654 22154 24670
rect 22278 30646 22312 30662
rect 22278 24654 22312 24670
rect 22436 30646 22470 30662
rect 22436 24654 22470 24670
rect 22594 30646 22628 30662
rect 22594 24654 22628 24670
rect 22752 30646 22786 30662
rect 22752 24654 22786 24670
rect 22910 30646 22944 30662
rect 22910 24654 22944 24670
rect 23068 30646 23102 30662
rect 23068 24654 23102 24670
rect 23226 30646 23260 30662
rect 23226 24654 23260 24670
rect 23384 30646 23418 30662
rect 23384 24654 23418 24670
rect 23542 30646 23576 30662
rect 23542 24654 23576 24670
rect 23700 30646 23734 30662
rect 23700 24654 23734 24670
rect 23858 30646 23892 30662
rect 23858 24654 23892 24670
rect 24016 30646 24050 30662
rect 24016 24654 24050 24670
rect 24174 30646 24208 30662
rect 24174 24654 24208 24670
rect 24332 30646 24366 30662
rect 24332 24654 24366 24670
rect 24490 30646 24524 30662
rect 24490 24654 24524 24670
rect 24648 30646 24682 30662
rect 24648 24654 24682 24670
rect 24806 30646 24840 30662
rect 24806 24654 24840 24670
rect 24964 30646 24998 30662
rect 24964 24654 24998 24670
rect 25122 30646 25156 30662
rect 25122 24654 25156 24670
rect 30838 27188 30934 27222
rect 31068 27188 31164 27222
rect 30838 27126 30872 27188
rect 30780 26980 30838 27000
rect 31130 27126 31164 27188
rect 30968 27042 30984 27076
rect 31018 27042 31034 27076
rect 30780 26020 30800 26980
rect 30780 26000 30838 26020
rect 30968 25662 30984 25696
rect 31018 25662 31034 25696
rect 30838 25550 30872 25612
rect 31130 25550 31164 25612
rect 30838 25516 30934 25550
rect 31068 25516 31164 25550
rect 1528 24586 1544 24620
rect 1612 24586 1628 24620
rect 1686 24586 1702 24620
rect 1770 24586 1786 24620
rect 1844 24586 1860 24620
rect 1928 24586 1944 24620
rect 2002 24586 2018 24620
rect 2086 24586 2102 24620
rect 2160 24586 2176 24620
rect 2244 24586 2260 24620
rect 2318 24586 2334 24620
rect 2402 24586 2418 24620
rect 2476 24586 2492 24620
rect 2560 24586 2576 24620
rect 2634 24586 2650 24620
rect 2718 24586 2734 24620
rect 2792 24586 2808 24620
rect 2876 24586 2892 24620
rect 2950 24586 2966 24620
rect 3034 24586 3050 24620
rect 3108 24586 3124 24620
rect 3192 24586 3208 24620
rect 3266 24586 3282 24620
rect 3350 24586 3366 24620
rect 3424 24586 3440 24620
rect 3508 24586 3524 24620
rect 3582 24586 3598 24620
rect 3666 24586 3682 24620
rect 3740 24586 3756 24620
rect 3824 24586 3840 24620
rect 3898 24586 3914 24620
rect 3982 24586 3998 24620
rect 4056 24586 4072 24620
rect 4140 24586 4156 24620
rect 4214 24586 4230 24620
rect 4298 24586 4314 24620
rect 4372 24586 4388 24620
rect 4456 24586 4472 24620
rect 4530 24586 4546 24620
rect 4614 24586 4630 24620
rect 4688 24586 4704 24620
rect 4772 24586 4788 24620
rect 4846 24586 4862 24620
rect 4930 24586 4946 24620
rect 5004 24586 5020 24620
rect 5088 24586 5104 24620
rect 5162 24586 5178 24620
rect 5246 24586 5262 24620
rect 5320 24586 5336 24620
rect 5404 24586 5420 24620
rect 5478 24586 5494 24620
rect 5562 24586 5578 24620
rect 5636 24586 5652 24620
rect 5720 24586 5736 24620
rect 5794 24586 5810 24620
rect 5878 24586 5894 24620
rect 5952 24586 5968 24620
rect 6036 24586 6052 24620
rect 6110 24586 6126 24620
rect 6194 24586 6210 24620
rect 1348 24482 1382 24544
rect 6356 24482 6390 24544
rect 1348 24448 1444 24482
rect 6294 24448 6390 24482
rect 7828 24586 7844 24620
rect 7912 24586 7928 24620
rect 7986 24586 8002 24620
rect 8070 24586 8086 24620
rect 8144 24586 8160 24620
rect 8228 24586 8244 24620
rect 8302 24586 8318 24620
rect 8386 24586 8402 24620
rect 8460 24586 8476 24620
rect 8544 24586 8560 24620
rect 8618 24586 8634 24620
rect 8702 24586 8718 24620
rect 8776 24586 8792 24620
rect 8860 24586 8876 24620
rect 8934 24586 8950 24620
rect 9018 24586 9034 24620
rect 9092 24586 9108 24620
rect 9176 24586 9192 24620
rect 9250 24586 9266 24620
rect 9334 24586 9350 24620
rect 9408 24586 9424 24620
rect 9492 24586 9508 24620
rect 9566 24586 9582 24620
rect 9650 24586 9666 24620
rect 9724 24586 9740 24620
rect 9808 24586 9824 24620
rect 9882 24586 9898 24620
rect 9966 24586 9982 24620
rect 10040 24586 10056 24620
rect 10124 24586 10140 24620
rect 10198 24586 10214 24620
rect 10282 24586 10298 24620
rect 10356 24586 10372 24620
rect 10440 24586 10456 24620
rect 10514 24586 10530 24620
rect 10598 24586 10614 24620
rect 10672 24586 10688 24620
rect 10756 24586 10772 24620
rect 10830 24586 10846 24620
rect 10914 24586 10930 24620
rect 10988 24586 11004 24620
rect 11072 24586 11088 24620
rect 11146 24586 11162 24620
rect 11230 24586 11246 24620
rect 11304 24586 11320 24620
rect 11388 24586 11404 24620
rect 11462 24586 11478 24620
rect 11546 24586 11562 24620
rect 11620 24586 11636 24620
rect 11704 24586 11720 24620
rect 11778 24586 11794 24620
rect 11862 24586 11878 24620
rect 11936 24586 11952 24620
rect 12020 24586 12036 24620
rect 12094 24586 12110 24620
rect 12178 24586 12194 24620
rect 12252 24586 12268 24620
rect 12336 24586 12352 24620
rect 12410 24586 12426 24620
rect 12494 24586 12510 24620
rect 7648 24482 7682 24544
rect 12656 24482 12690 24544
rect 7648 24448 7744 24482
rect 12594 24448 12690 24482
rect 14128 24586 14144 24620
rect 14212 24586 14228 24620
rect 14286 24586 14302 24620
rect 14370 24586 14386 24620
rect 14444 24586 14460 24620
rect 14528 24586 14544 24620
rect 14602 24586 14618 24620
rect 14686 24586 14702 24620
rect 14760 24586 14776 24620
rect 14844 24586 14860 24620
rect 14918 24586 14934 24620
rect 15002 24586 15018 24620
rect 15076 24586 15092 24620
rect 15160 24586 15176 24620
rect 15234 24586 15250 24620
rect 15318 24586 15334 24620
rect 15392 24586 15408 24620
rect 15476 24586 15492 24620
rect 15550 24586 15566 24620
rect 15634 24586 15650 24620
rect 15708 24586 15724 24620
rect 15792 24586 15808 24620
rect 15866 24586 15882 24620
rect 15950 24586 15966 24620
rect 16024 24586 16040 24620
rect 16108 24586 16124 24620
rect 16182 24586 16198 24620
rect 16266 24586 16282 24620
rect 16340 24586 16356 24620
rect 16424 24586 16440 24620
rect 16498 24586 16514 24620
rect 16582 24586 16598 24620
rect 16656 24586 16672 24620
rect 16740 24586 16756 24620
rect 16814 24586 16830 24620
rect 16898 24586 16914 24620
rect 16972 24586 16988 24620
rect 17056 24586 17072 24620
rect 17130 24586 17146 24620
rect 17214 24586 17230 24620
rect 17288 24586 17304 24620
rect 17372 24586 17388 24620
rect 17446 24586 17462 24620
rect 17530 24586 17546 24620
rect 17604 24586 17620 24620
rect 17688 24586 17704 24620
rect 17762 24586 17778 24620
rect 17846 24586 17862 24620
rect 17920 24586 17936 24620
rect 18004 24586 18020 24620
rect 18078 24586 18094 24620
rect 18162 24586 18178 24620
rect 18236 24586 18252 24620
rect 18320 24586 18336 24620
rect 18394 24586 18410 24620
rect 18478 24586 18494 24620
rect 18552 24586 18568 24620
rect 18636 24586 18652 24620
rect 18710 24586 18726 24620
rect 18794 24586 18810 24620
rect 13948 24482 13982 24544
rect 18956 24482 18990 24544
rect 13948 24448 14044 24482
rect 18894 24448 18990 24482
rect 20428 24586 20444 24620
rect 20512 24586 20528 24620
rect 20586 24586 20602 24620
rect 20670 24586 20686 24620
rect 20744 24586 20760 24620
rect 20828 24586 20844 24620
rect 20902 24586 20918 24620
rect 20986 24586 21002 24620
rect 21060 24586 21076 24620
rect 21144 24586 21160 24620
rect 21218 24586 21234 24620
rect 21302 24586 21318 24620
rect 21376 24586 21392 24620
rect 21460 24586 21476 24620
rect 21534 24586 21550 24620
rect 21618 24586 21634 24620
rect 21692 24586 21708 24620
rect 21776 24586 21792 24620
rect 21850 24586 21866 24620
rect 21934 24586 21950 24620
rect 22008 24586 22024 24620
rect 22092 24586 22108 24620
rect 22166 24586 22182 24620
rect 22250 24586 22266 24620
rect 22324 24586 22340 24620
rect 22408 24586 22424 24620
rect 22482 24586 22498 24620
rect 22566 24586 22582 24620
rect 22640 24586 22656 24620
rect 22724 24586 22740 24620
rect 22798 24586 22814 24620
rect 22882 24586 22898 24620
rect 22956 24586 22972 24620
rect 23040 24586 23056 24620
rect 23114 24586 23130 24620
rect 23198 24586 23214 24620
rect 23272 24586 23288 24620
rect 23356 24586 23372 24620
rect 23430 24586 23446 24620
rect 23514 24586 23530 24620
rect 23588 24586 23604 24620
rect 23672 24586 23688 24620
rect 23746 24586 23762 24620
rect 23830 24586 23846 24620
rect 23904 24586 23920 24620
rect 23988 24586 24004 24620
rect 24062 24586 24078 24620
rect 24146 24586 24162 24620
rect 24220 24586 24236 24620
rect 24304 24586 24320 24620
rect 24378 24586 24394 24620
rect 24462 24586 24478 24620
rect 24536 24586 24552 24620
rect 24620 24586 24636 24620
rect 24694 24586 24710 24620
rect 24778 24586 24794 24620
rect 24852 24586 24868 24620
rect 24936 24586 24952 24620
rect 25010 24586 25026 24620
rect 25094 24586 25110 24620
rect 20248 24482 20282 24544
rect 25256 24482 25290 24544
rect 20248 24448 20344 24482
rect 25194 24448 25290 24482
rect 1348 23834 1444 23868
rect 6294 23834 6390 23868
rect 1348 23772 1382 23834
rect 6356 23772 6390 23834
rect 1528 23696 1544 23730
rect 1612 23696 1628 23730
rect 1686 23696 1702 23730
rect 1770 23696 1786 23730
rect 1844 23696 1860 23730
rect 1928 23696 1944 23730
rect 2002 23696 2018 23730
rect 2086 23696 2102 23730
rect 2160 23696 2176 23730
rect 2244 23696 2260 23730
rect 2318 23696 2334 23730
rect 2402 23696 2418 23730
rect 2476 23696 2492 23730
rect 2560 23696 2576 23730
rect 2634 23696 2650 23730
rect 2718 23696 2734 23730
rect 2792 23696 2808 23730
rect 2876 23696 2892 23730
rect 2950 23696 2966 23730
rect 3034 23696 3050 23730
rect 3108 23696 3124 23730
rect 3192 23696 3208 23730
rect 3266 23696 3282 23730
rect 3350 23696 3366 23730
rect 3424 23696 3440 23730
rect 3508 23696 3524 23730
rect 3582 23696 3598 23730
rect 3666 23696 3682 23730
rect 3740 23696 3756 23730
rect 3824 23696 3840 23730
rect 3898 23696 3914 23730
rect 3982 23696 3998 23730
rect 4056 23696 4072 23730
rect 4140 23696 4156 23730
rect 4214 23696 4230 23730
rect 4298 23696 4314 23730
rect 4372 23696 4388 23730
rect 4456 23696 4472 23730
rect 4530 23696 4546 23730
rect 4614 23696 4630 23730
rect 4688 23696 4704 23730
rect 4772 23696 4788 23730
rect 4846 23696 4862 23730
rect 4930 23696 4946 23730
rect 5004 23696 5020 23730
rect 5088 23696 5104 23730
rect 5162 23696 5178 23730
rect 5246 23696 5262 23730
rect 5320 23696 5336 23730
rect 5404 23696 5420 23730
rect 5478 23696 5494 23730
rect 5562 23696 5578 23730
rect 5636 23696 5652 23730
rect 5720 23696 5736 23730
rect 5794 23696 5810 23730
rect 5878 23696 5894 23730
rect 5952 23696 5968 23730
rect 6036 23696 6052 23730
rect 6110 23696 6126 23730
rect 6194 23696 6210 23730
rect 7648 23834 7744 23868
rect 12594 23834 12690 23868
rect 7648 23772 7682 23834
rect 12656 23772 12690 23834
rect 7828 23696 7844 23730
rect 7912 23696 7928 23730
rect 7986 23696 8002 23730
rect 8070 23696 8086 23730
rect 8144 23696 8160 23730
rect 8228 23696 8244 23730
rect 8302 23696 8318 23730
rect 8386 23696 8402 23730
rect 8460 23696 8476 23730
rect 8544 23696 8560 23730
rect 8618 23696 8634 23730
rect 8702 23696 8718 23730
rect 8776 23696 8792 23730
rect 8860 23696 8876 23730
rect 8934 23696 8950 23730
rect 9018 23696 9034 23730
rect 9092 23696 9108 23730
rect 9176 23696 9192 23730
rect 9250 23696 9266 23730
rect 9334 23696 9350 23730
rect 9408 23696 9424 23730
rect 9492 23696 9508 23730
rect 9566 23696 9582 23730
rect 9650 23696 9666 23730
rect 9724 23696 9740 23730
rect 9808 23696 9824 23730
rect 9882 23696 9898 23730
rect 9966 23696 9982 23730
rect 10040 23696 10056 23730
rect 10124 23696 10140 23730
rect 10198 23696 10214 23730
rect 10282 23696 10298 23730
rect 10356 23696 10372 23730
rect 10440 23696 10456 23730
rect 10514 23696 10530 23730
rect 10598 23696 10614 23730
rect 10672 23696 10688 23730
rect 10756 23696 10772 23730
rect 10830 23696 10846 23730
rect 10914 23696 10930 23730
rect 10988 23696 11004 23730
rect 11072 23696 11088 23730
rect 11146 23696 11162 23730
rect 11230 23696 11246 23730
rect 11304 23696 11320 23730
rect 11388 23696 11404 23730
rect 11462 23696 11478 23730
rect 11546 23696 11562 23730
rect 11620 23696 11636 23730
rect 11704 23696 11720 23730
rect 11778 23696 11794 23730
rect 11862 23696 11878 23730
rect 11936 23696 11952 23730
rect 12020 23696 12036 23730
rect 12094 23696 12110 23730
rect 12178 23696 12194 23730
rect 12252 23696 12268 23730
rect 12336 23696 12352 23730
rect 12410 23696 12426 23730
rect 12494 23696 12510 23730
rect 13948 23834 14044 23868
rect 18894 23834 18990 23868
rect 13948 23772 13982 23834
rect 18956 23772 18990 23834
rect 14128 23696 14144 23730
rect 14212 23696 14228 23730
rect 14286 23696 14302 23730
rect 14370 23696 14386 23730
rect 14444 23696 14460 23730
rect 14528 23696 14544 23730
rect 14602 23696 14618 23730
rect 14686 23696 14702 23730
rect 14760 23696 14776 23730
rect 14844 23696 14860 23730
rect 14918 23696 14934 23730
rect 15002 23696 15018 23730
rect 15076 23696 15092 23730
rect 15160 23696 15176 23730
rect 15234 23696 15250 23730
rect 15318 23696 15334 23730
rect 15392 23696 15408 23730
rect 15476 23696 15492 23730
rect 15550 23696 15566 23730
rect 15634 23696 15650 23730
rect 15708 23696 15724 23730
rect 15792 23696 15808 23730
rect 15866 23696 15882 23730
rect 15950 23696 15966 23730
rect 16024 23696 16040 23730
rect 16108 23696 16124 23730
rect 16182 23696 16198 23730
rect 16266 23696 16282 23730
rect 16340 23696 16356 23730
rect 16424 23696 16440 23730
rect 16498 23696 16514 23730
rect 16582 23696 16598 23730
rect 16656 23696 16672 23730
rect 16740 23696 16756 23730
rect 16814 23696 16830 23730
rect 16898 23696 16914 23730
rect 16972 23696 16988 23730
rect 17056 23696 17072 23730
rect 17130 23696 17146 23730
rect 17214 23696 17230 23730
rect 17288 23696 17304 23730
rect 17372 23696 17388 23730
rect 17446 23696 17462 23730
rect 17530 23696 17546 23730
rect 17604 23696 17620 23730
rect 17688 23696 17704 23730
rect 17762 23696 17778 23730
rect 17846 23696 17862 23730
rect 17920 23696 17936 23730
rect 18004 23696 18020 23730
rect 18078 23696 18094 23730
rect 18162 23696 18178 23730
rect 18236 23696 18252 23730
rect 18320 23696 18336 23730
rect 18394 23696 18410 23730
rect 18478 23696 18494 23730
rect 18552 23696 18568 23730
rect 18636 23696 18652 23730
rect 18710 23696 18726 23730
rect 18794 23696 18810 23730
rect 20248 23834 20344 23868
rect 25194 23834 25290 23868
rect 20248 23772 20282 23834
rect 25256 23772 25290 23834
rect 20428 23696 20444 23730
rect 20512 23696 20528 23730
rect 20586 23696 20602 23730
rect 20670 23696 20686 23730
rect 20744 23696 20760 23730
rect 20828 23696 20844 23730
rect 20902 23696 20918 23730
rect 20986 23696 21002 23730
rect 21060 23696 21076 23730
rect 21144 23696 21160 23730
rect 21218 23696 21234 23730
rect 21302 23696 21318 23730
rect 21376 23696 21392 23730
rect 21460 23696 21476 23730
rect 21534 23696 21550 23730
rect 21618 23696 21634 23730
rect 21692 23696 21708 23730
rect 21776 23696 21792 23730
rect 21850 23696 21866 23730
rect 21934 23696 21950 23730
rect 22008 23696 22024 23730
rect 22092 23696 22108 23730
rect 22166 23696 22182 23730
rect 22250 23696 22266 23730
rect 22324 23696 22340 23730
rect 22408 23696 22424 23730
rect 22482 23696 22498 23730
rect 22566 23696 22582 23730
rect 22640 23696 22656 23730
rect 22724 23696 22740 23730
rect 22798 23696 22814 23730
rect 22882 23696 22898 23730
rect 22956 23696 22972 23730
rect 23040 23696 23056 23730
rect 23114 23696 23130 23730
rect 23198 23696 23214 23730
rect 23272 23696 23288 23730
rect 23356 23696 23372 23730
rect 23430 23696 23446 23730
rect 23514 23696 23530 23730
rect 23588 23696 23604 23730
rect 23672 23696 23688 23730
rect 23746 23696 23762 23730
rect 23830 23696 23846 23730
rect 23904 23696 23920 23730
rect 23988 23696 24004 23730
rect 24062 23696 24078 23730
rect 24146 23696 24162 23730
rect 24220 23696 24236 23730
rect 24304 23696 24320 23730
rect 24378 23696 24394 23730
rect 24462 23696 24478 23730
rect 24536 23696 24552 23730
rect 24620 23696 24636 23730
rect 24694 23696 24710 23730
rect 24778 23696 24794 23730
rect 24852 23696 24868 23730
rect 24936 23696 24952 23730
rect 25010 23696 25026 23730
rect 25094 23696 25110 23730
rect 1482 23646 1516 23662
rect 1482 17654 1516 17670
rect 1640 23646 1674 23662
rect 1640 17654 1674 17670
rect 1798 23646 1832 23662
rect 1798 17654 1832 17670
rect 1956 23646 1990 23662
rect 1956 17654 1990 17670
rect 2114 23646 2148 23662
rect 2114 17654 2148 17670
rect 2272 23646 2306 23662
rect 2272 17654 2306 17670
rect 2430 23646 2464 23662
rect 2430 17654 2464 17670
rect 2588 23646 2622 23662
rect 2588 17654 2622 17670
rect 2746 23646 2780 23662
rect 2746 17654 2780 17670
rect 2904 23646 2938 23662
rect 2904 17654 2938 17670
rect 3062 23646 3096 23662
rect 3062 17654 3096 17670
rect 3220 23646 3254 23662
rect 3220 17654 3254 17670
rect 3378 23646 3412 23662
rect 3378 17654 3412 17670
rect 3536 23646 3570 23662
rect 3536 17654 3570 17670
rect 3694 23646 3728 23662
rect 3694 17654 3728 17670
rect 3852 23646 3886 23662
rect 3852 17654 3886 17670
rect 4010 23646 4044 23662
rect 4010 17654 4044 17670
rect 4168 23646 4202 23662
rect 4168 17654 4202 17670
rect 4326 23646 4360 23662
rect 4326 17654 4360 17670
rect 4484 23646 4518 23662
rect 4484 17654 4518 17670
rect 4642 23646 4676 23662
rect 4642 17654 4676 17670
rect 4800 23646 4834 23662
rect 4800 17654 4834 17670
rect 4958 23646 4992 23662
rect 4958 17654 4992 17670
rect 5116 23646 5150 23662
rect 5116 17654 5150 17670
rect 5274 23646 5308 23662
rect 5274 17654 5308 17670
rect 5432 23646 5466 23662
rect 5432 17654 5466 17670
rect 5590 23646 5624 23662
rect 5590 17654 5624 17670
rect 5748 23646 5782 23662
rect 5748 17654 5782 17670
rect 5906 23646 5940 23662
rect 5906 17654 5940 17670
rect 6064 23646 6098 23662
rect 6064 17654 6098 17670
rect 6222 23646 6256 23662
rect 6222 17654 6256 17670
rect 7782 23646 7816 23662
rect 7782 17654 7816 17670
rect 7940 23646 7974 23662
rect 7940 17654 7974 17670
rect 8098 23646 8132 23662
rect 8098 17654 8132 17670
rect 8256 23646 8290 23662
rect 8256 17654 8290 17670
rect 8414 23646 8448 23662
rect 8414 17654 8448 17670
rect 8572 23646 8606 23662
rect 8572 17654 8606 17670
rect 8730 23646 8764 23662
rect 8730 17654 8764 17670
rect 8888 23646 8922 23662
rect 8888 17654 8922 17670
rect 9046 23646 9080 23662
rect 9046 17654 9080 17670
rect 9204 23646 9238 23662
rect 9204 17654 9238 17670
rect 9362 23646 9396 23662
rect 9362 17654 9396 17670
rect 9520 23646 9554 23662
rect 9520 17654 9554 17670
rect 9678 23646 9712 23662
rect 9678 17654 9712 17670
rect 9836 23646 9870 23662
rect 9836 17654 9870 17670
rect 9994 23646 10028 23662
rect 9994 17654 10028 17670
rect 10152 23646 10186 23662
rect 10152 17654 10186 17670
rect 10310 23646 10344 23662
rect 10310 17654 10344 17670
rect 10468 23646 10502 23662
rect 10468 17654 10502 17670
rect 10626 23646 10660 23662
rect 10626 17654 10660 17670
rect 10784 23646 10818 23662
rect 10784 17654 10818 17670
rect 10942 23646 10976 23662
rect 10942 17654 10976 17670
rect 11100 23646 11134 23662
rect 11100 17654 11134 17670
rect 11258 23646 11292 23662
rect 11258 17654 11292 17670
rect 11416 23646 11450 23662
rect 11416 17654 11450 17670
rect 11574 23646 11608 23662
rect 11574 17654 11608 17670
rect 11732 23646 11766 23662
rect 11732 17654 11766 17670
rect 11890 23646 11924 23662
rect 11890 17654 11924 17670
rect 12048 23646 12082 23662
rect 12048 17654 12082 17670
rect 12206 23646 12240 23662
rect 12206 17654 12240 17670
rect 12364 23646 12398 23662
rect 12364 17654 12398 17670
rect 12522 23646 12556 23662
rect 12522 17654 12556 17670
rect 14082 23646 14116 23662
rect 14082 17654 14116 17670
rect 14240 23646 14274 23662
rect 14240 17654 14274 17670
rect 14398 23646 14432 23662
rect 14398 17654 14432 17670
rect 14556 23646 14590 23662
rect 14556 17654 14590 17670
rect 14714 23646 14748 23662
rect 14714 17654 14748 17670
rect 14872 23646 14906 23662
rect 14872 17654 14906 17670
rect 15030 23646 15064 23662
rect 15030 17654 15064 17670
rect 15188 23646 15222 23662
rect 15188 17654 15222 17670
rect 15346 23646 15380 23662
rect 15346 17654 15380 17670
rect 15504 23646 15538 23662
rect 15504 17654 15538 17670
rect 15662 23646 15696 23662
rect 15662 17654 15696 17670
rect 15820 23646 15854 23662
rect 15820 17654 15854 17670
rect 15978 23646 16012 23662
rect 15978 17654 16012 17670
rect 16136 23646 16170 23662
rect 16136 17654 16170 17670
rect 16294 23646 16328 23662
rect 16294 17654 16328 17670
rect 16452 23646 16486 23662
rect 16452 17654 16486 17670
rect 16610 23646 16644 23662
rect 16610 17654 16644 17670
rect 16768 23646 16802 23662
rect 16768 17654 16802 17670
rect 16926 23646 16960 23662
rect 16926 17654 16960 17670
rect 17084 23646 17118 23662
rect 17084 17654 17118 17670
rect 17242 23646 17276 23662
rect 17242 17654 17276 17670
rect 17400 23646 17434 23662
rect 17400 17654 17434 17670
rect 17558 23646 17592 23662
rect 17558 17654 17592 17670
rect 17716 23646 17750 23662
rect 17716 17654 17750 17670
rect 17874 23646 17908 23662
rect 17874 17654 17908 17670
rect 18032 23646 18066 23662
rect 18032 17654 18066 17670
rect 18190 23646 18224 23662
rect 18190 17654 18224 17670
rect 18348 23646 18382 23662
rect 18348 17654 18382 17670
rect 18506 23646 18540 23662
rect 18506 17654 18540 17670
rect 18664 23646 18698 23662
rect 18664 17654 18698 17670
rect 18822 23646 18856 23662
rect 18822 17654 18856 17670
rect 20382 23646 20416 23662
rect 20382 17654 20416 17670
rect 20540 23646 20574 23662
rect 20540 17654 20574 17670
rect 20698 23646 20732 23662
rect 20698 17654 20732 17670
rect 20856 23646 20890 23662
rect 20856 17654 20890 17670
rect 21014 23646 21048 23662
rect 21014 17654 21048 17670
rect 21172 23646 21206 23662
rect 21172 17654 21206 17670
rect 21330 23646 21364 23662
rect 21330 17654 21364 17670
rect 21488 23646 21522 23662
rect 21488 17654 21522 17670
rect 21646 23646 21680 23662
rect 21646 17654 21680 17670
rect 21804 23646 21838 23662
rect 21804 17654 21838 17670
rect 21962 23646 21996 23662
rect 21962 17654 21996 17670
rect 22120 23646 22154 23662
rect 22120 17654 22154 17670
rect 22278 23646 22312 23662
rect 22278 17654 22312 17670
rect 22436 23646 22470 23662
rect 22436 17654 22470 17670
rect 22594 23646 22628 23662
rect 22594 17654 22628 17670
rect 22752 23646 22786 23662
rect 22752 17654 22786 17670
rect 22910 23646 22944 23662
rect 22910 17654 22944 17670
rect 23068 23646 23102 23662
rect 23068 17654 23102 17670
rect 23226 23646 23260 23662
rect 23226 17654 23260 17670
rect 23384 23646 23418 23662
rect 23384 17654 23418 17670
rect 23542 23646 23576 23662
rect 23542 17654 23576 17670
rect 23700 23646 23734 23662
rect 23700 17654 23734 17670
rect 23858 23646 23892 23662
rect 23858 17654 23892 17670
rect 24016 23646 24050 23662
rect 24016 17654 24050 17670
rect 24174 23646 24208 23662
rect 24174 17654 24208 17670
rect 24332 23646 24366 23662
rect 24332 17654 24366 17670
rect 24490 23646 24524 23662
rect 24490 17654 24524 17670
rect 24648 23646 24682 23662
rect 24648 17654 24682 17670
rect 24806 23646 24840 23662
rect 24806 17654 24840 17670
rect 24964 23646 24998 23662
rect 24964 17654 24998 17670
rect 25122 23646 25156 23662
rect 25122 17654 25156 17670
rect 1528 17586 1544 17620
rect 1612 17586 1628 17620
rect 1686 17586 1702 17620
rect 1770 17586 1786 17620
rect 1844 17586 1860 17620
rect 1928 17586 1944 17620
rect 2002 17586 2018 17620
rect 2086 17586 2102 17620
rect 2160 17586 2176 17620
rect 2244 17586 2260 17620
rect 2318 17586 2334 17620
rect 2402 17586 2418 17620
rect 2476 17586 2492 17620
rect 2560 17586 2576 17620
rect 2634 17586 2650 17620
rect 2718 17586 2734 17620
rect 2792 17586 2808 17620
rect 2876 17586 2892 17620
rect 2950 17586 2966 17620
rect 3034 17586 3050 17620
rect 3108 17586 3124 17620
rect 3192 17586 3208 17620
rect 3266 17586 3282 17620
rect 3350 17586 3366 17620
rect 3424 17586 3440 17620
rect 3508 17586 3524 17620
rect 3582 17586 3598 17620
rect 3666 17586 3682 17620
rect 3740 17586 3756 17620
rect 3824 17586 3840 17620
rect 3898 17586 3914 17620
rect 3982 17586 3998 17620
rect 4056 17586 4072 17620
rect 4140 17586 4156 17620
rect 4214 17586 4230 17620
rect 4298 17586 4314 17620
rect 4372 17586 4388 17620
rect 4456 17586 4472 17620
rect 4530 17586 4546 17620
rect 4614 17586 4630 17620
rect 4688 17586 4704 17620
rect 4772 17586 4788 17620
rect 4846 17586 4862 17620
rect 4930 17586 4946 17620
rect 5004 17586 5020 17620
rect 5088 17586 5104 17620
rect 5162 17586 5178 17620
rect 5246 17586 5262 17620
rect 5320 17586 5336 17620
rect 5404 17586 5420 17620
rect 5478 17586 5494 17620
rect 5562 17586 5578 17620
rect 5636 17586 5652 17620
rect 5720 17586 5736 17620
rect 5794 17586 5810 17620
rect 5878 17586 5894 17620
rect 5952 17586 5968 17620
rect 6036 17586 6052 17620
rect 6110 17586 6126 17620
rect 6194 17586 6210 17620
rect 1348 17482 1382 17544
rect 6356 17482 6390 17544
rect 1348 17448 1444 17482
rect 6294 17448 6390 17482
rect 7828 17586 7844 17620
rect 7912 17586 7928 17620
rect 7986 17586 8002 17620
rect 8070 17586 8086 17620
rect 8144 17586 8160 17620
rect 8228 17586 8244 17620
rect 8302 17586 8318 17620
rect 8386 17586 8402 17620
rect 8460 17586 8476 17620
rect 8544 17586 8560 17620
rect 8618 17586 8634 17620
rect 8702 17586 8718 17620
rect 8776 17586 8792 17620
rect 8860 17586 8876 17620
rect 8934 17586 8950 17620
rect 9018 17586 9034 17620
rect 9092 17586 9108 17620
rect 9176 17586 9192 17620
rect 9250 17586 9266 17620
rect 9334 17586 9350 17620
rect 9408 17586 9424 17620
rect 9492 17586 9508 17620
rect 9566 17586 9582 17620
rect 9650 17586 9666 17620
rect 9724 17586 9740 17620
rect 9808 17586 9824 17620
rect 9882 17586 9898 17620
rect 9966 17586 9982 17620
rect 10040 17586 10056 17620
rect 10124 17586 10140 17620
rect 10198 17586 10214 17620
rect 10282 17586 10298 17620
rect 10356 17586 10372 17620
rect 10440 17586 10456 17620
rect 10514 17586 10530 17620
rect 10598 17586 10614 17620
rect 10672 17586 10688 17620
rect 10756 17586 10772 17620
rect 10830 17586 10846 17620
rect 10914 17586 10930 17620
rect 10988 17586 11004 17620
rect 11072 17586 11088 17620
rect 11146 17586 11162 17620
rect 11230 17586 11246 17620
rect 11304 17586 11320 17620
rect 11388 17586 11404 17620
rect 11462 17586 11478 17620
rect 11546 17586 11562 17620
rect 11620 17586 11636 17620
rect 11704 17586 11720 17620
rect 11778 17586 11794 17620
rect 11862 17586 11878 17620
rect 11936 17586 11952 17620
rect 12020 17586 12036 17620
rect 12094 17586 12110 17620
rect 12178 17586 12194 17620
rect 12252 17586 12268 17620
rect 12336 17586 12352 17620
rect 12410 17586 12426 17620
rect 12494 17586 12510 17620
rect 7648 17482 7682 17544
rect 12656 17482 12690 17544
rect 7648 17448 7744 17482
rect 12594 17448 12690 17482
rect 14128 17586 14144 17620
rect 14212 17586 14228 17620
rect 14286 17586 14302 17620
rect 14370 17586 14386 17620
rect 14444 17586 14460 17620
rect 14528 17586 14544 17620
rect 14602 17586 14618 17620
rect 14686 17586 14702 17620
rect 14760 17586 14776 17620
rect 14844 17586 14860 17620
rect 14918 17586 14934 17620
rect 15002 17586 15018 17620
rect 15076 17586 15092 17620
rect 15160 17586 15176 17620
rect 15234 17586 15250 17620
rect 15318 17586 15334 17620
rect 15392 17586 15408 17620
rect 15476 17586 15492 17620
rect 15550 17586 15566 17620
rect 15634 17586 15650 17620
rect 15708 17586 15724 17620
rect 15792 17586 15808 17620
rect 15866 17586 15882 17620
rect 15950 17586 15966 17620
rect 16024 17586 16040 17620
rect 16108 17586 16124 17620
rect 16182 17586 16198 17620
rect 16266 17586 16282 17620
rect 16340 17586 16356 17620
rect 16424 17586 16440 17620
rect 16498 17586 16514 17620
rect 16582 17586 16598 17620
rect 16656 17586 16672 17620
rect 16740 17586 16756 17620
rect 16814 17586 16830 17620
rect 16898 17586 16914 17620
rect 16972 17586 16988 17620
rect 17056 17586 17072 17620
rect 17130 17586 17146 17620
rect 17214 17586 17230 17620
rect 17288 17586 17304 17620
rect 17372 17586 17388 17620
rect 17446 17586 17462 17620
rect 17530 17586 17546 17620
rect 17604 17586 17620 17620
rect 17688 17586 17704 17620
rect 17762 17586 17778 17620
rect 17846 17586 17862 17620
rect 17920 17586 17936 17620
rect 18004 17586 18020 17620
rect 18078 17586 18094 17620
rect 18162 17586 18178 17620
rect 18236 17586 18252 17620
rect 18320 17586 18336 17620
rect 18394 17586 18410 17620
rect 18478 17586 18494 17620
rect 18552 17586 18568 17620
rect 18636 17586 18652 17620
rect 18710 17586 18726 17620
rect 18794 17586 18810 17620
rect 13948 17482 13982 17544
rect 18956 17482 18990 17544
rect 13948 17448 14044 17482
rect 18894 17448 18990 17482
rect 20428 17586 20444 17620
rect 20512 17586 20528 17620
rect 20586 17586 20602 17620
rect 20670 17586 20686 17620
rect 20744 17586 20760 17620
rect 20828 17586 20844 17620
rect 20902 17586 20918 17620
rect 20986 17586 21002 17620
rect 21060 17586 21076 17620
rect 21144 17586 21160 17620
rect 21218 17586 21234 17620
rect 21302 17586 21318 17620
rect 21376 17586 21392 17620
rect 21460 17586 21476 17620
rect 21534 17586 21550 17620
rect 21618 17586 21634 17620
rect 21692 17586 21708 17620
rect 21776 17586 21792 17620
rect 21850 17586 21866 17620
rect 21934 17586 21950 17620
rect 22008 17586 22024 17620
rect 22092 17586 22108 17620
rect 22166 17586 22182 17620
rect 22250 17586 22266 17620
rect 22324 17586 22340 17620
rect 22408 17586 22424 17620
rect 22482 17586 22498 17620
rect 22566 17586 22582 17620
rect 22640 17586 22656 17620
rect 22724 17586 22740 17620
rect 22798 17586 22814 17620
rect 22882 17586 22898 17620
rect 22956 17586 22972 17620
rect 23040 17586 23056 17620
rect 23114 17586 23130 17620
rect 23198 17586 23214 17620
rect 23272 17586 23288 17620
rect 23356 17586 23372 17620
rect 23430 17586 23446 17620
rect 23514 17586 23530 17620
rect 23588 17586 23604 17620
rect 23672 17586 23688 17620
rect 23746 17586 23762 17620
rect 23830 17586 23846 17620
rect 23904 17586 23920 17620
rect 23988 17586 24004 17620
rect 24062 17586 24078 17620
rect 24146 17586 24162 17620
rect 24220 17586 24236 17620
rect 24304 17586 24320 17620
rect 24378 17586 24394 17620
rect 24462 17586 24478 17620
rect 24536 17586 24552 17620
rect 24620 17586 24636 17620
rect 24694 17586 24710 17620
rect 24778 17586 24794 17620
rect 24852 17586 24868 17620
rect 24936 17586 24952 17620
rect 25010 17586 25026 17620
rect 25094 17586 25110 17620
rect 20248 17482 20282 17544
rect 25256 17482 25290 17544
rect 20248 17448 20344 17482
rect 25194 17448 25290 17482
rect 1348 15534 1444 15568
rect 6294 15534 6390 15568
rect 1348 15472 1382 15534
rect 6356 15472 6390 15534
rect 1528 15396 1544 15430
rect 1612 15396 1628 15430
rect 1686 15396 1702 15430
rect 1770 15396 1786 15430
rect 1844 15396 1860 15430
rect 1928 15396 1944 15430
rect 2002 15396 2018 15430
rect 2086 15396 2102 15430
rect 2160 15396 2176 15430
rect 2244 15396 2260 15430
rect 2318 15396 2334 15430
rect 2402 15396 2418 15430
rect 2476 15396 2492 15430
rect 2560 15396 2576 15430
rect 2634 15396 2650 15430
rect 2718 15396 2734 15430
rect 2792 15396 2808 15430
rect 2876 15396 2892 15430
rect 2950 15396 2966 15430
rect 3034 15396 3050 15430
rect 3108 15396 3124 15430
rect 3192 15396 3208 15430
rect 3266 15396 3282 15430
rect 3350 15396 3366 15430
rect 3424 15396 3440 15430
rect 3508 15396 3524 15430
rect 3582 15396 3598 15430
rect 3666 15396 3682 15430
rect 3740 15396 3756 15430
rect 3824 15396 3840 15430
rect 3898 15396 3914 15430
rect 3982 15396 3998 15430
rect 4056 15396 4072 15430
rect 4140 15396 4156 15430
rect 4214 15396 4230 15430
rect 4298 15396 4314 15430
rect 4372 15396 4388 15430
rect 4456 15396 4472 15430
rect 4530 15396 4546 15430
rect 4614 15396 4630 15430
rect 4688 15396 4704 15430
rect 4772 15396 4788 15430
rect 4846 15396 4862 15430
rect 4930 15396 4946 15430
rect 5004 15396 5020 15430
rect 5088 15396 5104 15430
rect 5162 15396 5178 15430
rect 5246 15396 5262 15430
rect 5320 15396 5336 15430
rect 5404 15396 5420 15430
rect 5478 15396 5494 15430
rect 5562 15396 5578 15430
rect 5636 15396 5652 15430
rect 5720 15396 5736 15430
rect 5794 15396 5810 15430
rect 5878 15396 5894 15430
rect 5952 15396 5968 15430
rect 6036 15396 6052 15430
rect 6110 15396 6126 15430
rect 6194 15396 6210 15430
rect 7648 15534 7744 15568
rect 12594 15534 12690 15568
rect 7648 15472 7682 15534
rect 12656 15472 12690 15534
rect 7828 15396 7844 15430
rect 7912 15396 7928 15430
rect 7986 15396 8002 15430
rect 8070 15396 8086 15430
rect 8144 15396 8160 15430
rect 8228 15396 8244 15430
rect 8302 15396 8318 15430
rect 8386 15396 8402 15430
rect 8460 15396 8476 15430
rect 8544 15396 8560 15430
rect 8618 15396 8634 15430
rect 8702 15396 8718 15430
rect 8776 15396 8792 15430
rect 8860 15396 8876 15430
rect 8934 15396 8950 15430
rect 9018 15396 9034 15430
rect 9092 15396 9108 15430
rect 9176 15396 9192 15430
rect 9250 15396 9266 15430
rect 9334 15396 9350 15430
rect 9408 15396 9424 15430
rect 9492 15396 9508 15430
rect 9566 15396 9582 15430
rect 9650 15396 9666 15430
rect 9724 15396 9740 15430
rect 9808 15396 9824 15430
rect 9882 15396 9898 15430
rect 9966 15396 9982 15430
rect 10040 15396 10056 15430
rect 10124 15396 10140 15430
rect 10198 15396 10214 15430
rect 10282 15396 10298 15430
rect 10356 15396 10372 15430
rect 10440 15396 10456 15430
rect 10514 15396 10530 15430
rect 10598 15396 10614 15430
rect 10672 15396 10688 15430
rect 10756 15396 10772 15430
rect 10830 15396 10846 15430
rect 10914 15396 10930 15430
rect 10988 15396 11004 15430
rect 11072 15396 11088 15430
rect 11146 15396 11162 15430
rect 11230 15396 11246 15430
rect 11304 15396 11320 15430
rect 11388 15396 11404 15430
rect 11462 15396 11478 15430
rect 11546 15396 11562 15430
rect 11620 15396 11636 15430
rect 11704 15396 11720 15430
rect 11778 15396 11794 15430
rect 11862 15396 11878 15430
rect 11936 15396 11952 15430
rect 12020 15396 12036 15430
rect 12094 15396 12110 15430
rect 12178 15396 12194 15430
rect 12252 15396 12268 15430
rect 12336 15396 12352 15430
rect 12410 15396 12426 15430
rect 12494 15396 12510 15430
rect 13948 15534 14044 15568
rect 18894 15534 18990 15568
rect 13948 15472 13982 15534
rect 18956 15472 18990 15534
rect 14128 15396 14144 15430
rect 14212 15396 14228 15430
rect 14286 15396 14302 15430
rect 14370 15396 14386 15430
rect 14444 15396 14460 15430
rect 14528 15396 14544 15430
rect 14602 15396 14618 15430
rect 14686 15396 14702 15430
rect 14760 15396 14776 15430
rect 14844 15396 14860 15430
rect 14918 15396 14934 15430
rect 15002 15396 15018 15430
rect 15076 15396 15092 15430
rect 15160 15396 15176 15430
rect 15234 15396 15250 15430
rect 15318 15396 15334 15430
rect 15392 15396 15408 15430
rect 15476 15396 15492 15430
rect 15550 15396 15566 15430
rect 15634 15396 15650 15430
rect 15708 15396 15724 15430
rect 15792 15396 15808 15430
rect 15866 15396 15882 15430
rect 15950 15396 15966 15430
rect 16024 15396 16040 15430
rect 16108 15396 16124 15430
rect 16182 15396 16198 15430
rect 16266 15396 16282 15430
rect 16340 15396 16356 15430
rect 16424 15396 16440 15430
rect 16498 15396 16514 15430
rect 16582 15396 16598 15430
rect 16656 15396 16672 15430
rect 16740 15396 16756 15430
rect 16814 15396 16830 15430
rect 16898 15396 16914 15430
rect 16972 15396 16988 15430
rect 17056 15396 17072 15430
rect 17130 15396 17146 15430
rect 17214 15396 17230 15430
rect 17288 15396 17304 15430
rect 17372 15396 17388 15430
rect 17446 15396 17462 15430
rect 17530 15396 17546 15430
rect 17604 15396 17620 15430
rect 17688 15396 17704 15430
rect 17762 15396 17778 15430
rect 17846 15396 17862 15430
rect 17920 15396 17936 15430
rect 18004 15396 18020 15430
rect 18078 15396 18094 15430
rect 18162 15396 18178 15430
rect 18236 15396 18252 15430
rect 18320 15396 18336 15430
rect 18394 15396 18410 15430
rect 18478 15396 18494 15430
rect 18552 15396 18568 15430
rect 18636 15396 18652 15430
rect 18710 15396 18726 15430
rect 18794 15396 18810 15430
rect 20248 15534 20344 15568
rect 25194 15534 25290 15568
rect 20248 15472 20282 15534
rect 25256 15472 25290 15534
rect 20428 15396 20444 15430
rect 20512 15396 20528 15430
rect 20586 15396 20602 15430
rect 20670 15396 20686 15430
rect 20744 15396 20760 15430
rect 20828 15396 20844 15430
rect 20902 15396 20918 15430
rect 20986 15396 21002 15430
rect 21060 15396 21076 15430
rect 21144 15396 21160 15430
rect 21218 15396 21234 15430
rect 21302 15396 21318 15430
rect 21376 15396 21392 15430
rect 21460 15396 21476 15430
rect 21534 15396 21550 15430
rect 21618 15396 21634 15430
rect 21692 15396 21708 15430
rect 21776 15396 21792 15430
rect 21850 15396 21866 15430
rect 21934 15396 21950 15430
rect 22008 15396 22024 15430
rect 22092 15396 22108 15430
rect 22166 15396 22182 15430
rect 22250 15396 22266 15430
rect 22324 15396 22340 15430
rect 22408 15396 22424 15430
rect 22482 15396 22498 15430
rect 22566 15396 22582 15430
rect 22640 15396 22656 15430
rect 22724 15396 22740 15430
rect 22798 15396 22814 15430
rect 22882 15396 22898 15430
rect 22956 15396 22972 15430
rect 23040 15396 23056 15430
rect 23114 15396 23130 15430
rect 23198 15396 23214 15430
rect 23272 15396 23288 15430
rect 23356 15396 23372 15430
rect 23430 15396 23446 15430
rect 23514 15396 23530 15430
rect 23588 15396 23604 15430
rect 23672 15396 23688 15430
rect 23746 15396 23762 15430
rect 23830 15396 23846 15430
rect 23904 15396 23920 15430
rect 23988 15396 24004 15430
rect 24062 15396 24078 15430
rect 24146 15396 24162 15430
rect 24220 15396 24236 15430
rect 24304 15396 24320 15430
rect 24378 15396 24394 15430
rect 24462 15396 24478 15430
rect 24536 15396 24552 15430
rect 24620 15396 24636 15430
rect 24694 15396 24710 15430
rect 24778 15396 24794 15430
rect 24852 15396 24868 15430
rect 24936 15396 24952 15430
rect 25010 15396 25026 15430
rect 25094 15396 25110 15430
rect -4364 13946 -4268 13980
rect -4130 13960 -4034 13980
rect -4130 13946 -3980 13960
rect -4364 13884 -4330 13946
rect -4068 13940 -3980 13946
rect -4068 13884 -4040 13940
rect -4364 12570 -4330 12632
rect -4068 12570 -4040 12632
rect -4364 12536 -4268 12570
rect -4130 12560 -4040 12570
rect -4000 12560 -3980 13940
rect -4130 12540 -3980 12560
rect -4130 12536 -4034 12540
rect 1482 15346 1516 15362
rect 1482 9354 1516 9370
rect 1640 15346 1674 15362
rect 1640 9354 1674 9370
rect 1798 15346 1832 15362
rect 1798 9354 1832 9370
rect 1956 15346 1990 15362
rect 1956 9354 1990 9370
rect 2114 15346 2148 15362
rect 2114 9354 2148 9370
rect 2272 15346 2306 15362
rect 2272 9354 2306 9370
rect 2430 15346 2464 15362
rect 2430 9354 2464 9370
rect 2588 15346 2622 15362
rect 2588 9354 2622 9370
rect 2746 15346 2780 15362
rect 2746 9354 2780 9370
rect 2904 15346 2938 15362
rect 2904 9354 2938 9370
rect 3062 15346 3096 15362
rect 3062 9354 3096 9370
rect 3220 15346 3254 15362
rect 3220 9354 3254 9370
rect 3378 15346 3412 15362
rect 3378 9354 3412 9370
rect 3536 15346 3570 15362
rect 3536 9354 3570 9370
rect 3694 15346 3728 15362
rect 3694 9354 3728 9370
rect 3852 15346 3886 15362
rect 3852 9354 3886 9370
rect 4010 15346 4044 15362
rect 4010 9354 4044 9370
rect 4168 15346 4202 15362
rect 4168 9354 4202 9370
rect 4326 15346 4360 15362
rect 4326 9354 4360 9370
rect 4484 15346 4518 15362
rect 4484 9354 4518 9370
rect 4642 15346 4676 15362
rect 4642 9354 4676 9370
rect 4800 15346 4834 15362
rect 4800 9354 4834 9370
rect 4958 15346 4992 15362
rect 4958 9354 4992 9370
rect 5116 15346 5150 15362
rect 5116 9354 5150 9370
rect 5274 15346 5308 15362
rect 5274 9354 5308 9370
rect 5432 15346 5466 15362
rect 5432 9354 5466 9370
rect 5590 15346 5624 15362
rect 5590 9354 5624 9370
rect 5748 15346 5782 15362
rect 5748 9354 5782 9370
rect 5906 15346 5940 15362
rect 5906 9354 5940 9370
rect 6064 15346 6098 15362
rect 6064 9354 6098 9370
rect 6222 15346 6256 15362
rect 6222 9354 6256 9370
rect 7782 15346 7816 15362
rect 7782 9354 7816 9370
rect 7940 15346 7974 15362
rect 7940 9354 7974 9370
rect 8098 15346 8132 15362
rect 8098 9354 8132 9370
rect 8256 15346 8290 15362
rect 8256 9354 8290 9370
rect 8414 15346 8448 15362
rect 8414 9354 8448 9370
rect 8572 15346 8606 15362
rect 8572 9354 8606 9370
rect 8730 15346 8764 15362
rect 8730 9354 8764 9370
rect 8888 15346 8922 15362
rect 8888 9354 8922 9370
rect 9046 15346 9080 15362
rect 9046 9354 9080 9370
rect 9204 15346 9238 15362
rect 9204 9354 9238 9370
rect 9362 15346 9396 15362
rect 9362 9354 9396 9370
rect 9520 15346 9554 15362
rect 9520 9354 9554 9370
rect 9678 15346 9712 15362
rect 9678 9354 9712 9370
rect 9836 15346 9870 15362
rect 9836 9354 9870 9370
rect 9994 15346 10028 15362
rect 9994 9354 10028 9370
rect 10152 15346 10186 15362
rect 10152 9354 10186 9370
rect 10310 15346 10344 15362
rect 10310 9354 10344 9370
rect 10468 15346 10502 15362
rect 10468 9354 10502 9370
rect 10626 15346 10660 15362
rect 10626 9354 10660 9370
rect 10784 15346 10818 15362
rect 10784 9354 10818 9370
rect 10942 15346 10976 15362
rect 10942 9354 10976 9370
rect 11100 15346 11134 15362
rect 11100 9354 11134 9370
rect 11258 15346 11292 15362
rect 11258 9354 11292 9370
rect 11416 15346 11450 15362
rect 11416 9354 11450 9370
rect 11574 15346 11608 15362
rect 11574 9354 11608 9370
rect 11732 15346 11766 15362
rect 11732 9354 11766 9370
rect 11890 15346 11924 15362
rect 11890 9354 11924 9370
rect 12048 15346 12082 15362
rect 12048 9354 12082 9370
rect 12206 15346 12240 15362
rect 12206 9354 12240 9370
rect 12364 15346 12398 15362
rect 12364 9354 12398 9370
rect 12522 15346 12556 15362
rect 12522 9354 12556 9370
rect 14082 15346 14116 15362
rect 14082 9354 14116 9370
rect 14240 15346 14274 15362
rect 14240 9354 14274 9370
rect 14398 15346 14432 15362
rect 14398 9354 14432 9370
rect 14556 15346 14590 15362
rect 14556 9354 14590 9370
rect 14714 15346 14748 15362
rect 14714 9354 14748 9370
rect 14872 15346 14906 15362
rect 14872 9354 14906 9370
rect 15030 15346 15064 15362
rect 15030 9354 15064 9370
rect 15188 15346 15222 15362
rect 15188 9354 15222 9370
rect 15346 15346 15380 15362
rect 15346 9354 15380 9370
rect 15504 15346 15538 15362
rect 15504 9354 15538 9370
rect 15662 15346 15696 15362
rect 15662 9354 15696 9370
rect 15820 15346 15854 15362
rect 15820 9354 15854 9370
rect 15978 15346 16012 15362
rect 15978 9354 16012 9370
rect 16136 15346 16170 15362
rect 16136 9354 16170 9370
rect 16294 15346 16328 15362
rect 16294 9354 16328 9370
rect 16452 15346 16486 15362
rect 16452 9354 16486 9370
rect 16610 15346 16644 15362
rect 16610 9354 16644 9370
rect 16768 15346 16802 15362
rect 16768 9354 16802 9370
rect 16926 15346 16960 15362
rect 16926 9354 16960 9370
rect 17084 15346 17118 15362
rect 17084 9354 17118 9370
rect 17242 15346 17276 15362
rect 17242 9354 17276 9370
rect 17400 15346 17434 15362
rect 17400 9354 17434 9370
rect 17558 15346 17592 15362
rect 17558 9354 17592 9370
rect 17716 15346 17750 15362
rect 17716 9354 17750 9370
rect 17874 15346 17908 15362
rect 17874 9354 17908 9370
rect 18032 15346 18066 15362
rect 18032 9354 18066 9370
rect 18190 15346 18224 15362
rect 18190 9354 18224 9370
rect 18348 15346 18382 15362
rect 18348 9354 18382 9370
rect 18506 15346 18540 15362
rect 18506 9354 18540 9370
rect 18664 15346 18698 15362
rect 18664 9354 18698 9370
rect 18822 15346 18856 15362
rect 18822 9354 18856 9370
rect 20382 15346 20416 15362
rect 20382 9354 20416 9370
rect 20540 15346 20574 15362
rect 20540 9354 20574 9370
rect 20698 15346 20732 15362
rect 20698 9354 20732 9370
rect 20856 15346 20890 15362
rect 20856 9354 20890 9370
rect 21014 15346 21048 15362
rect 21014 9354 21048 9370
rect 21172 15346 21206 15362
rect 21172 9354 21206 9370
rect 21330 15346 21364 15362
rect 21330 9354 21364 9370
rect 21488 15346 21522 15362
rect 21488 9354 21522 9370
rect 21646 15346 21680 15362
rect 21646 9354 21680 9370
rect 21804 15346 21838 15362
rect 21804 9354 21838 9370
rect 21962 15346 21996 15362
rect 21962 9354 21996 9370
rect 22120 15346 22154 15362
rect 22120 9354 22154 9370
rect 22278 15346 22312 15362
rect 22278 9354 22312 9370
rect 22436 15346 22470 15362
rect 22436 9354 22470 9370
rect 22594 15346 22628 15362
rect 22594 9354 22628 9370
rect 22752 15346 22786 15362
rect 22752 9354 22786 9370
rect 22910 15346 22944 15362
rect 22910 9354 22944 9370
rect 23068 15346 23102 15362
rect 23068 9354 23102 9370
rect 23226 15346 23260 15362
rect 23226 9354 23260 9370
rect 23384 15346 23418 15362
rect 23384 9354 23418 9370
rect 23542 15346 23576 15362
rect 23542 9354 23576 9370
rect 23700 15346 23734 15362
rect 23700 9354 23734 9370
rect 23858 15346 23892 15362
rect 23858 9354 23892 9370
rect 24016 15346 24050 15362
rect 24016 9354 24050 9370
rect 24174 15346 24208 15362
rect 24174 9354 24208 9370
rect 24332 15346 24366 15362
rect 24332 9354 24366 9370
rect 24490 15346 24524 15362
rect 24490 9354 24524 9370
rect 24648 15346 24682 15362
rect 24648 9354 24682 9370
rect 24806 15346 24840 15362
rect 24806 9354 24840 9370
rect 24964 15346 24998 15362
rect 24964 9354 24998 9370
rect 25122 15346 25156 15362
rect 25122 9354 25156 9370
rect 30780 13980 30860 14000
rect 30780 12520 30800 13980
rect 30840 13946 30930 13980
rect 31068 13946 31164 13980
rect 30840 13884 30868 13946
rect 31130 13884 31164 13946
rect 30840 12570 30868 12632
rect 31130 12570 31164 12632
rect 30840 12536 30930 12570
rect 31068 12536 31164 12570
rect 30840 12520 30860 12536
rect 30780 12500 30860 12520
rect 1528 9286 1544 9320
rect 1612 9286 1628 9320
rect 1686 9286 1702 9320
rect 1770 9286 1786 9320
rect 1844 9286 1860 9320
rect 1928 9286 1944 9320
rect 2002 9286 2018 9320
rect 2086 9286 2102 9320
rect 2160 9286 2176 9320
rect 2244 9286 2260 9320
rect 2318 9286 2334 9320
rect 2402 9286 2418 9320
rect 2476 9286 2492 9320
rect 2560 9286 2576 9320
rect 2634 9286 2650 9320
rect 2718 9286 2734 9320
rect 2792 9286 2808 9320
rect 2876 9286 2892 9320
rect 2950 9286 2966 9320
rect 3034 9286 3050 9320
rect 3108 9286 3124 9320
rect 3192 9286 3208 9320
rect 3266 9286 3282 9320
rect 3350 9286 3366 9320
rect 3424 9286 3440 9320
rect 3508 9286 3524 9320
rect 3582 9286 3598 9320
rect 3666 9286 3682 9320
rect 3740 9286 3756 9320
rect 3824 9286 3840 9320
rect 3898 9286 3914 9320
rect 3982 9286 3998 9320
rect 4056 9286 4072 9320
rect 4140 9286 4156 9320
rect 4214 9286 4230 9320
rect 4298 9286 4314 9320
rect 4372 9286 4388 9320
rect 4456 9286 4472 9320
rect 4530 9286 4546 9320
rect 4614 9286 4630 9320
rect 4688 9286 4704 9320
rect 4772 9286 4788 9320
rect 4846 9286 4862 9320
rect 4930 9286 4946 9320
rect 5004 9286 5020 9320
rect 5088 9286 5104 9320
rect 5162 9286 5178 9320
rect 5246 9286 5262 9320
rect 5320 9286 5336 9320
rect 5404 9286 5420 9320
rect 5478 9286 5494 9320
rect 5562 9286 5578 9320
rect 5636 9286 5652 9320
rect 5720 9286 5736 9320
rect 5794 9286 5810 9320
rect 5878 9286 5894 9320
rect 5952 9286 5968 9320
rect 6036 9286 6052 9320
rect 6110 9286 6126 9320
rect 6194 9286 6210 9320
rect 1348 9182 1382 9244
rect 6356 9182 6390 9244
rect 1348 9148 1444 9182
rect 6294 9148 6390 9182
rect 7828 9286 7844 9320
rect 7912 9286 7928 9320
rect 7986 9286 8002 9320
rect 8070 9286 8086 9320
rect 8144 9286 8160 9320
rect 8228 9286 8244 9320
rect 8302 9286 8318 9320
rect 8386 9286 8402 9320
rect 8460 9286 8476 9320
rect 8544 9286 8560 9320
rect 8618 9286 8634 9320
rect 8702 9286 8718 9320
rect 8776 9286 8792 9320
rect 8860 9286 8876 9320
rect 8934 9286 8950 9320
rect 9018 9286 9034 9320
rect 9092 9286 9108 9320
rect 9176 9286 9192 9320
rect 9250 9286 9266 9320
rect 9334 9286 9350 9320
rect 9408 9286 9424 9320
rect 9492 9286 9508 9320
rect 9566 9286 9582 9320
rect 9650 9286 9666 9320
rect 9724 9286 9740 9320
rect 9808 9286 9824 9320
rect 9882 9286 9898 9320
rect 9966 9286 9982 9320
rect 10040 9286 10056 9320
rect 10124 9286 10140 9320
rect 10198 9286 10214 9320
rect 10282 9286 10298 9320
rect 10356 9286 10372 9320
rect 10440 9286 10456 9320
rect 10514 9286 10530 9320
rect 10598 9286 10614 9320
rect 10672 9286 10688 9320
rect 10756 9286 10772 9320
rect 10830 9286 10846 9320
rect 10914 9286 10930 9320
rect 10988 9286 11004 9320
rect 11072 9286 11088 9320
rect 11146 9286 11162 9320
rect 11230 9286 11246 9320
rect 11304 9286 11320 9320
rect 11388 9286 11404 9320
rect 11462 9286 11478 9320
rect 11546 9286 11562 9320
rect 11620 9286 11636 9320
rect 11704 9286 11720 9320
rect 11778 9286 11794 9320
rect 11862 9286 11878 9320
rect 11936 9286 11952 9320
rect 12020 9286 12036 9320
rect 12094 9286 12110 9320
rect 12178 9286 12194 9320
rect 12252 9286 12268 9320
rect 12336 9286 12352 9320
rect 12410 9286 12426 9320
rect 12494 9286 12510 9320
rect 7648 9182 7682 9244
rect 12656 9182 12690 9244
rect 7648 9148 7744 9182
rect 12594 9148 12690 9182
rect 14128 9286 14144 9320
rect 14212 9286 14228 9320
rect 14286 9286 14302 9320
rect 14370 9286 14386 9320
rect 14444 9286 14460 9320
rect 14528 9286 14544 9320
rect 14602 9286 14618 9320
rect 14686 9286 14702 9320
rect 14760 9286 14776 9320
rect 14844 9286 14860 9320
rect 14918 9286 14934 9320
rect 15002 9286 15018 9320
rect 15076 9286 15092 9320
rect 15160 9286 15176 9320
rect 15234 9286 15250 9320
rect 15318 9286 15334 9320
rect 15392 9286 15408 9320
rect 15476 9286 15492 9320
rect 15550 9286 15566 9320
rect 15634 9286 15650 9320
rect 15708 9286 15724 9320
rect 15792 9286 15808 9320
rect 15866 9286 15882 9320
rect 15950 9286 15966 9320
rect 16024 9286 16040 9320
rect 16108 9286 16124 9320
rect 16182 9286 16198 9320
rect 16266 9286 16282 9320
rect 16340 9286 16356 9320
rect 16424 9286 16440 9320
rect 16498 9286 16514 9320
rect 16582 9286 16598 9320
rect 16656 9286 16672 9320
rect 16740 9286 16756 9320
rect 16814 9286 16830 9320
rect 16898 9286 16914 9320
rect 16972 9286 16988 9320
rect 17056 9286 17072 9320
rect 17130 9286 17146 9320
rect 17214 9286 17230 9320
rect 17288 9286 17304 9320
rect 17372 9286 17388 9320
rect 17446 9286 17462 9320
rect 17530 9286 17546 9320
rect 17604 9286 17620 9320
rect 17688 9286 17704 9320
rect 17762 9286 17778 9320
rect 17846 9286 17862 9320
rect 17920 9286 17936 9320
rect 18004 9286 18020 9320
rect 18078 9286 18094 9320
rect 18162 9286 18178 9320
rect 18236 9286 18252 9320
rect 18320 9286 18336 9320
rect 18394 9286 18410 9320
rect 18478 9286 18494 9320
rect 18552 9286 18568 9320
rect 18636 9286 18652 9320
rect 18710 9286 18726 9320
rect 18794 9286 18810 9320
rect 13948 9182 13982 9244
rect 18956 9182 18990 9244
rect 13948 9148 14044 9182
rect 18894 9148 18990 9182
rect 20428 9286 20444 9320
rect 20512 9286 20528 9320
rect 20586 9286 20602 9320
rect 20670 9286 20686 9320
rect 20744 9286 20760 9320
rect 20828 9286 20844 9320
rect 20902 9286 20918 9320
rect 20986 9286 21002 9320
rect 21060 9286 21076 9320
rect 21144 9286 21160 9320
rect 21218 9286 21234 9320
rect 21302 9286 21318 9320
rect 21376 9286 21392 9320
rect 21460 9286 21476 9320
rect 21534 9286 21550 9320
rect 21618 9286 21634 9320
rect 21692 9286 21708 9320
rect 21776 9286 21792 9320
rect 21850 9286 21866 9320
rect 21934 9286 21950 9320
rect 22008 9286 22024 9320
rect 22092 9286 22108 9320
rect 22166 9286 22182 9320
rect 22250 9286 22266 9320
rect 22324 9286 22340 9320
rect 22408 9286 22424 9320
rect 22482 9286 22498 9320
rect 22566 9286 22582 9320
rect 22640 9286 22656 9320
rect 22724 9286 22740 9320
rect 22798 9286 22814 9320
rect 22882 9286 22898 9320
rect 22956 9286 22972 9320
rect 23040 9286 23056 9320
rect 23114 9286 23130 9320
rect 23198 9286 23214 9320
rect 23272 9286 23288 9320
rect 23356 9286 23372 9320
rect 23430 9286 23446 9320
rect 23514 9286 23530 9320
rect 23588 9286 23604 9320
rect 23672 9286 23688 9320
rect 23746 9286 23762 9320
rect 23830 9286 23846 9320
rect 23904 9286 23920 9320
rect 23988 9286 24004 9320
rect 24062 9286 24078 9320
rect 24146 9286 24162 9320
rect 24220 9286 24236 9320
rect 24304 9286 24320 9320
rect 24378 9286 24394 9320
rect 24462 9286 24478 9320
rect 24536 9286 24552 9320
rect 24620 9286 24636 9320
rect 24694 9286 24710 9320
rect 24778 9286 24794 9320
rect 24852 9286 24868 9320
rect 24936 9286 24952 9320
rect 25010 9286 25026 9320
rect 25094 9286 25110 9320
rect 20248 9182 20282 9244
rect 25256 9182 25290 9244
rect 20248 9148 20344 9182
rect 25194 9148 25290 9182
rect 1348 8534 1444 8568
rect 6294 8534 6390 8568
rect 1348 8472 1382 8534
rect 6356 8472 6390 8534
rect 1528 8396 1544 8430
rect 1612 8396 1628 8430
rect 1686 8396 1702 8430
rect 1770 8396 1786 8430
rect 1844 8396 1860 8430
rect 1928 8396 1944 8430
rect 2002 8396 2018 8430
rect 2086 8396 2102 8430
rect 2160 8396 2176 8430
rect 2244 8396 2260 8430
rect 2318 8396 2334 8430
rect 2402 8396 2418 8430
rect 2476 8396 2492 8430
rect 2560 8396 2576 8430
rect 2634 8396 2650 8430
rect 2718 8396 2734 8430
rect 2792 8396 2808 8430
rect 2876 8396 2892 8430
rect 2950 8396 2966 8430
rect 3034 8396 3050 8430
rect 3108 8396 3124 8430
rect 3192 8396 3208 8430
rect 3266 8396 3282 8430
rect 3350 8396 3366 8430
rect 3424 8396 3440 8430
rect 3508 8396 3524 8430
rect 3582 8396 3598 8430
rect 3666 8396 3682 8430
rect 3740 8396 3756 8430
rect 3824 8396 3840 8430
rect 3898 8396 3914 8430
rect 3982 8396 3998 8430
rect 4056 8396 4072 8430
rect 4140 8396 4156 8430
rect 4214 8396 4230 8430
rect 4298 8396 4314 8430
rect 4372 8396 4388 8430
rect 4456 8396 4472 8430
rect 4530 8396 4546 8430
rect 4614 8396 4630 8430
rect 4688 8396 4704 8430
rect 4772 8396 4788 8430
rect 4846 8396 4862 8430
rect 4930 8396 4946 8430
rect 5004 8396 5020 8430
rect 5088 8396 5104 8430
rect 5162 8396 5178 8430
rect 5246 8396 5262 8430
rect 5320 8396 5336 8430
rect 5404 8396 5420 8430
rect 5478 8396 5494 8430
rect 5562 8396 5578 8430
rect 5636 8396 5652 8430
rect 5720 8396 5736 8430
rect 5794 8396 5810 8430
rect 5878 8396 5894 8430
rect 5952 8396 5968 8430
rect 6036 8396 6052 8430
rect 6110 8396 6126 8430
rect 6194 8396 6210 8430
rect 7648 8534 7744 8568
rect 12594 8534 12690 8568
rect 7648 8472 7682 8534
rect 12656 8472 12690 8534
rect 7828 8396 7844 8430
rect 7912 8396 7928 8430
rect 7986 8396 8002 8430
rect 8070 8396 8086 8430
rect 8144 8396 8160 8430
rect 8228 8396 8244 8430
rect 8302 8396 8318 8430
rect 8386 8396 8402 8430
rect 8460 8396 8476 8430
rect 8544 8396 8560 8430
rect 8618 8396 8634 8430
rect 8702 8396 8718 8430
rect 8776 8396 8792 8430
rect 8860 8396 8876 8430
rect 8934 8396 8950 8430
rect 9018 8396 9034 8430
rect 9092 8396 9108 8430
rect 9176 8396 9192 8430
rect 9250 8396 9266 8430
rect 9334 8396 9350 8430
rect 9408 8396 9424 8430
rect 9492 8396 9508 8430
rect 9566 8396 9582 8430
rect 9650 8396 9666 8430
rect 9724 8396 9740 8430
rect 9808 8396 9824 8430
rect 9882 8396 9898 8430
rect 9966 8396 9982 8430
rect 10040 8396 10056 8430
rect 10124 8396 10140 8430
rect 10198 8396 10214 8430
rect 10282 8396 10298 8430
rect 10356 8396 10372 8430
rect 10440 8396 10456 8430
rect 10514 8396 10530 8430
rect 10598 8396 10614 8430
rect 10672 8396 10688 8430
rect 10756 8396 10772 8430
rect 10830 8396 10846 8430
rect 10914 8396 10930 8430
rect 10988 8396 11004 8430
rect 11072 8396 11088 8430
rect 11146 8396 11162 8430
rect 11230 8396 11246 8430
rect 11304 8396 11320 8430
rect 11388 8396 11404 8430
rect 11462 8396 11478 8430
rect 11546 8396 11562 8430
rect 11620 8396 11636 8430
rect 11704 8396 11720 8430
rect 11778 8396 11794 8430
rect 11862 8396 11878 8430
rect 11936 8396 11952 8430
rect 12020 8396 12036 8430
rect 12094 8396 12110 8430
rect 12178 8396 12194 8430
rect 12252 8396 12268 8430
rect 12336 8396 12352 8430
rect 12410 8396 12426 8430
rect 12494 8396 12510 8430
rect 13948 8534 14044 8568
rect 18894 8534 18990 8568
rect 13948 8472 13982 8534
rect 18956 8472 18990 8534
rect 14128 8396 14144 8430
rect 14212 8396 14228 8430
rect 14286 8396 14302 8430
rect 14370 8396 14386 8430
rect 14444 8396 14460 8430
rect 14528 8396 14544 8430
rect 14602 8396 14618 8430
rect 14686 8396 14702 8430
rect 14760 8396 14776 8430
rect 14844 8396 14860 8430
rect 14918 8396 14934 8430
rect 15002 8396 15018 8430
rect 15076 8396 15092 8430
rect 15160 8396 15176 8430
rect 15234 8396 15250 8430
rect 15318 8396 15334 8430
rect 15392 8396 15408 8430
rect 15476 8396 15492 8430
rect 15550 8396 15566 8430
rect 15634 8396 15650 8430
rect 15708 8396 15724 8430
rect 15792 8396 15808 8430
rect 15866 8396 15882 8430
rect 15950 8396 15966 8430
rect 16024 8396 16040 8430
rect 16108 8396 16124 8430
rect 16182 8396 16198 8430
rect 16266 8396 16282 8430
rect 16340 8396 16356 8430
rect 16424 8396 16440 8430
rect 16498 8396 16514 8430
rect 16582 8396 16598 8430
rect 16656 8396 16672 8430
rect 16740 8396 16756 8430
rect 16814 8396 16830 8430
rect 16898 8396 16914 8430
rect 16972 8396 16988 8430
rect 17056 8396 17072 8430
rect 17130 8396 17146 8430
rect 17214 8396 17230 8430
rect 17288 8396 17304 8430
rect 17372 8396 17388 8430
rect 17446 8396 17462 8430
rect 17530 8396 17546 8430
rect 17604 8396 17620 8430
rect 17688 8396 17704 8430
rect 17762 8396 17778 8430
rect 17846 8396 17862 8430
rect 17920 8396 17936 8430
rect 18004 8396 18020 8430
rect 18078 8396 18094 8430
rect 18162 8396 18178 8430
rect 18236 8396 18252 8430
rect 18320 8396 18336 8430
rect 18394 8396 18410 8430
rect 18478 8396 18494 8430
rect 18552 8396 18568 8430
rect 18636 8396 18652 8430
rect 18710 8396 18726 8430
rect 18794 8396 18810 8430
rect 20248 8534 20344 8568
rect 25194 8534 25290 8568
rect 20248 8472 20282 8534
rect 25256 8472 25290 8534
rect 20428 8396 20444 8430
rect 20512 8396 20528 8430
rect 20586 8396 20602 8430
rect 20670 8396 20686 8430
rect 20744 8396 20760 8430
rect 20828 8396 20844 8430
rect 20902 8396 20918 8430
rect 20986 8396 21002 8430
rect 21060 8396 21076 8430
rect 21144 8396 21160 8430
rect 21218 8396 21234 8430
rect 21302 8396 21318 8430
rect 21376 8396 21392 8430
rect 21460 8396 21476 8430
rect 21534 8396 21550 8430
rect 21618 8396 21634 8430
rect 21692 8396 21708 8430
rect 21776 8396 21792 8430
rect 21850 8396 21866 8430
rect 21934 8396 21950 8430
rect 22008 8396 22024 8430
rect 22092 8396 22108 8430
rect 22166 8396 22182 8430
rect 22250 8396 22266 8430
rect 22324 8396 22340 8430
rect 22408 8396 22424 8430
rect 22482 8396 22498 8430
rect 22566 8396 22582 8430
rect 22640 8396 22656 8430
rect 22724 8396 22740 8430
rect 22798 8396 22814 8430
rect 22882 8396 22898 8430
rect 22956 8396 22972 8430
rect 23040 8396 23056 8430
rect 23114 8396 23130 8430
rect 23198 8396 23214 8430
rect 23272 8396 23288 8430
rect 23356 8396 23372 8430
rect 23430 8396 23446 8430
rect 23514 8396 23530 8430
rect 23588 8396 23604 8430
rect 23672 8396 23688 8430
rect 23746 8396 23762 8430
rect 23830 8396 23846 8430
rect 23904 8396 23920 8430
rect 23988 8396 24004 8430
rect 24062 8396 24078 8430
rect 24146 8396 24162 8430
rect 24220 8396 24236 8430
rect 24304 8396 24320 8430
rect 24378 8396 24394 8430
rect 24462 8396 24478 8430
rect 24536 8396 24552 8430
rect 24620 8396 24636 8430
rect 24694 8396 24710 8430
rect 24778 8396 24794 8430
rect 24852 8396 24868 8430
rect 24936 8396 24952 8430
rect 25010 8396 25026 8430
rect 25094 8396 25110 8430
rect 1482 8346 1516 8362
rect 1482 2354 1516 2370
rect 1640 8346 1674 8362
rect 1640 2354 1674 2370
rect 1798 8346 1832 8362
rect 1798 2354 1832 2370
rect 1956 8346 1990 8362
rect 1956 2354 1990 2370
rect 2114 8346 2148 8362
rect 2114 2354 2148 2370
rect 2272 8346 2306 8362
rect 2272 2354 2306 2370
rect 2430 8346 2464 8362
rect 2430 2354 2464 2370
rect 2588 8346 2622 8362
rect 2588 2354 2622 2370
rect 2746 8346 2780 8362
rect 2746 2354 2780 2370
rect 2904 8346 2938 8362
rect 2904 2354 2938 2370
rect 3062 8346 3096 8362
rect 3062 2354 3096 2370
rect 3220 8346 3254 8362
rect 3220 2354 3254 2370
rect 3378 8346 3412 8362
rect 3378 2354 3412 2370
rect 3536 8346 3570 8362
rect 3536 2354 3570 2370
rect 3694 8346 3728 8362
rect 3694 2354 3728 2370
rect 3852 8346 3886 8362
rect 3852 2354 3886 2370
rect 4010 8346 4044 8362
rect 4010 2354 4044 2370
rect 4168 8346 4202 8362
rect 4168 2354 4202 2370
rect 4326 8346 4360 8362
rect 4326 2354 4360 2370
rect 4484 8346 4518 8362
rect 4484 2354 4518 2370
rect 4642 8346 4676 8362
rect 4642 2354 4676 2370
rect 4800 8346 4834 8362
rect 4800 2354 4834 2370
rect 4958 8346 4992 8362
rect 4958 2354 4992 2370
rect 5116 8346 5150 8362
rect 5116 2354 5150 2370
rect 5274 8346 5308 8362
rect 5274 2354 5308 2370
rect 5432 8346 5466 8362
rect 5432 2354 5466 2370
rect 5590 8346 5624 8362
rect 5590 2354 5624 2370
rect 5748 8346 5782 8362
rect 5748 2354 5782 2370
rect 5906 8346 5940 8362
rect 5906 2354 5940 2370
rect 6064 8346 6098 8362
rect 6064 2354 6098 2370
rect 6222 8346 6256 8362
rect 6222 2354 6256 2370
rect 7782 8346 7816 8362
rect 7782 2354 7816 2370
rect 7940 8346 7974 8362
rect 7940 2354 7974 2370
rect 8098 8346 8132 8362
rect 8098 2354 8132 2370
rect 8256 8346 8290 8362
rect 8256 2354 8290 2370
rect 8414 8346 8448 8362
rect 8414 2354 8448 2370
rect 8572 8346 8606 8362
rect 8572 2354 8606 2370
rect 8730 8346 8764 8362
rect 8730 2354 8764 2370
rect 8888 8346 8922 8362
rect 8888 2354 8922 2370
rect 9046 8346 9080 8362
rect 9046 2354 9080 2370
rect 9204 8346 9238 8362
rect 9204 2354 9238 2370
rect 9362 8346 9396 8362
rect 9362 2354 9396 2370
rect 9520 8346 9554 8362
rect 9520 2354 9554 2370
rect 9678 8346 9712 8362
rect 9678 2354 9712 2370
rect 9836 8346 9870 8362
rect 9836 2354 9870 2370
rect 9994 8346 10028 8362
rect 9994 2354 10028 2370
rect 10152 8346 10186 8362
rect 10152 2354 10186 2370
rect 10310 8346 10344 8362
rect 10310 2354 10344 2370
rect 10468 8346 10502 8362
rect 10468 2354 10502 2370
rect 10626 8346 10660 8362
rect 10626 2354 10660 2370
rect 10784 8346 10818 8362
rect 10784 2354 10818 2370
rect 10942 8346 10976 8362
rect 10942 2354 10976 2370
rect 11100 8346 11134 8362
rect 11100 2354 11134 2370
rect 11258 8346 11292 8362
rect 11258 2354 11292 2370
rect 11416 8346 11450 8362
rect 11416 2354 11450 2370
rect 11574 8346 11608 8362
rect 11574 2354 11608 2370
rect 11732 8346 11766 8362
rect 11732 2354 11766 2370
rect 11890 8346 11924 8362
rect 11890 2354 11924 2370
rect 12048 8346 12082 8362
rect 12048 2354 12082 2370
rect 12206 8346 12240 8362
rect 12206 2354 12240 2370
rect 12364 8346 12398 8362
rect 12364 2354 12398 2370
rect 12522 8346 12556 8362
rect 12522 2354 12556 2370
rect 14082 8346 14116 8362
rect 14082 2354 14116 2370
rect 14240 8346 14274 8362
rect 14240 2354 14274 2370
rect 14398 8346 14432 8362
rect 14398 2354 14432 2370
rect 14556 8346 14590 8362
rect 14556 2354 14590 2370
rect 14714 8346 14748 8362
rect 14714 2354 14748 2370
rect 14872 8346 14906 8362
rect 14872 2354 14906 2370
rect 15030 8346 15064 8362
rect 15030 2354 15064 2370
rect 15188 8346 15222 8362
rect 15188 2354 15222 2370
rect 15346 8346 15380 8362
rect 15346 2354 15380 2370
rect 15504 8346 15538 8362
rect 15504 2354 15538 2370
rect 15662 8346 15696 8362
rect 15662 2354 15696 2370
rect 15820 8346 15854 8362
rect 15820 2354 15854 2370
rect 15978 8346 16012 8362
rect 15978 2354 16012 2370
rect 16136 8346 16170 8362
rect 16136 2354 16170 2370
rect 16294 8346 16328 8362
rect 16294 2354 16328 2370
rect 16452 8346 16486 8362
rect 16452 2354 16486 2370
rect 16610 8346 16644 8362
rect 16610 2354 16644 2370
rect 16768 8346 16802 8362
rect 16768 2354 16802 2370
rect 16926 8346 16960 8362
rect 16926 2354 16960 2370
rect 17084 8346 17118 8362
rect 17084 2354 17118 2370
rect 17242 8346 17276 8362
rect 17242 2354 17276 2370
rect 17400 8346 17434 8362
rect 17400 2354 17434 2370
rect 17558 8346 17592 8362
rect 17558 2354 17592 2370
rect 17716 8346 17750 8362
rect 17716 2354 17750 2370
rect 17874 8346 17908 8362
rect 17874 2354 17908 2370
rect 18032 8346 18066 8362
rect 18032 2354 18066 2370
rect 18190 8346 18224 8362
rect 18190 2354 18224 2370
rect 18348 8346 18382 8362
rect 18348 2354 18382 2370
rect 18506 8346 18540 8362
rect 18506 2354 18540 2370
rect 18664 8346 18698 8362
rect 18664 2354 18698 2370
rect 18822 8346 18856 8362
rect 18822 2354 18856 2370
rect 20382 8346 20416 8362
rect 20382 2354 20416 2370
rect 20540 8346 20574 8362
rect 20540 2354 20574 2370
rect 20698 8346 20732 8362
rect 20698 2354 20732 2370
rect 20856 8346 20890 8362
rect 20856 2354 20890 2370
rect 21014 8346 21048 8362
rect 21014 2354 21048 2370
rect 21172 8346 21206 8362
rect 21172 2354 21206 2370
rect 21330 8346 21364 8362
rect 21330 2354 21364 2370
rect 21488 8346 21522 8362
rect 21488 2354 21522 2370
rect 21646 8346 21680 8362
rect 21646 2354 21680 2370
rect 21804 8346 21838 8362
rect 21804 2354 21838 2370
rect 21962 8346 21996 8362
rect 21962 2354 21996 2370
rect 22120 8346 22154 8362
rect 22120 2354 22154 2370
rect 22278 8346 22312 8362
rect 22278 2354 22312 2370
rect 22436 8346 22470 8362
rect 22436 2354 22470 2370
rect 22594 8346 22628 8362
rect 22594 2354 22628 2370
rect 22752 8346 22786 8362
rect 22752 2354 22786 2370
rect 22910 8346 22944 8362
rect 22910 2354 22944 2370
rect 23068 8346 23102 8362
rect 23068 2354 23102 2370
rect 23226 8346 23260 8362
rect 23226 2354 23260 2370
rect 23384 8346 23418 8362
rect 23384 2354 23418 2370
rect 23542 8346 23576 8362
rect 23542 2354 23576 2370
rect 23700 8346 23734 8362
rect 23700 2354 23734 2370
rect 23858 8346 23892 8362
rect 23858 2354 23892 2370
rect 24016 8346 24050 8362
rect 24016 2354 24050 2370
rect 24174 8346 24208 8362
rect 24174 2354 24208 2370
rect 24332 8346 24366 8362
rect 24332 2354 24366 2370
rect 24490 8346 24524 8362
rect 24490 2354 24524 2370
rect 24648 8346 24682 8362
rect 24648 2354 24682 2370
rect 24806 8346 24840 8362
rect 24806 2354 24840 2370
rect 24964 8346 24998 8362
rect 24964 2354 24998 2370
rect 25122 8346 25156 8362
rect 25122 2354 25156 2370
rect 1528 2286 1544 2320
rect 1612 2286 1628 2320
rect 1686 2286 1702 2320
rect 1770 2286 1786 2320
rect 1844 2286 1860 2320
rect 1928 2286 1944 2320
rect 2002 2286 2018 2320
rect 2086 2286 2102 2320
rect 2160 2286 2176 2320
rect 2244 2286 2260 2320
rect 2318 2286 2334 2320
rect 2402 2286 2418 2320
rect 2476 2286 2492 2320
rect 2560 2286 2576 2320
rect 2634 2286 2650 2320
rect 2718 2286 2734 2320
rect 2792 2286 2808 2320
rect 2876 2286 2892 2320
rect 2950 2286 2966 2320
rect 3034 2286 3050 2320
rect 3108 2286 3124 2320
rect 3192 2286 3208 2320
rect 3266 2286 3282 2320
rect 3350 2286 3366 2320
rect 3424 2286 3440 2320
rect 3508 2286 3524 2320
rect 3582 2286 3598 2320
rect 3666 2286 3682 2320
rect 3740 2286 3756 2320
rect 3824 2286 3840 2320
rect 3898 2286 3914 2320
rect 3982 2286 3998 2320
rect 4056 2286 4072 2320
rect 4140 2286 4156 2320
rect 4214 2286 4230 2320
rect 4298 2286 4314 2320
rect 4372 2286 4388 2320
rect 4456 2286 4472 2320
rect 4530 2286 4546 2320
rect 4614 2286 4630 2320
rect 4688 2286 4704 2320
rect 4772 2286 4788 2320
rect 4846 2286 4862 2320
rect 4930 2286 4946 2320
rect 5004 2286 5020 2320
rect 5088 2286 5104 2320
rect 5162 2286 5178 2320
rect 5246 2286 5262 2320
rect 5320 2286 5336 2320
rect 5404 2286 5420 2320
rect 5478 2286 5494 2320
rect 5562 2286 5578 2320
rect 5636 2286 5652 2320
rect 5720 2286 5736 2320
rect 5794 2286 5810 2320
rect 5878 2286 5894 2320
rect 5952 2286 5968 2320
rect 6036 2286 6052 2320
rect 6110 2286 6126 2320
rect 6194 2286 6210 2320
rect 1348 2182 1382 2244
rect 6356 2182 6390 2244
rect 1348 2148 1444 2182
rect 6294 2148 6390 2182
rect 7828 2286 7844 2320
rect 7912 2286 7928 2320
rect 7986 2286 8002 2320
rect 8070 2286 8086 2320
rect 8144 2286 8160 2320
rect 8228 2286 8244 2320
rect 8302 2286 8318 2320
rect 8386 2286 8402 2320
rect 8460 2286 8476 2320
rect 8544 2286 8560 2320
rect 8618 2286 8634 2320
rect 8702 2286 8718 2320
rect 8776 2286 8792 2320
rect 8860 2286 8876 2320
rect 8934 2286 8950 2320
rect 9018 2286 9034 2320
rect 9092 2286 9108 2320
rect 9176 2286 9192 2320
rect 9250 2286 9266 2320
rect 9334 2286 9350 2320
rect 9408 2286 9424 2320
rect 9492 2286 9508 2320
rect 9566 2286 9582 2320
rect 9650 2286 9666 2320
rect 9724 2286 9740 2320
rect 9808 2286 9824 2320
rect 9882 2286 9898 2320
rect 9966 2286 9982 2320
rect 10040 2286 10056 2320
rect 10124 2286 10140 2320
rect 10198 2286 10214 2320
rect 10282 2286 10298 2320
rect 10356 2286 10372 2320
rect 10440 2286 10456 2320
rect 10514 2286 10530 2320
rect 10598 2286 10614 2320
rect 10672 2286 10688 2320
rect 10756 2286 10772 2320
rect 10830 2286 10846 2320
rect 10914 2286 10930 2320
rect 10988 2286 11004 2320
rect 11072 2286 11088 2320
rect 11146 2286 11162 2320
rect 11230 2286 11246 2320
rect 11304 2286 11320 2320
rect 11388 2286 11404 2320
rect 11462 2286 11478 2320
rect 11546 2286 11562 2320
rect 11620 2286 11636 2320
rect 11704 2286 11720 2320
rect 11778 2286 11794 2320
rect 11862 2286 11878 2320
rect 11936 2286 11952 2320
rect 12020 2286 12036 2320
rect 12094 2286 12110 2320
rect 12178 2286 12194 2320
rect 12252 2286 12268 2320
rect 12336 2286 12352 2320
rect 12410 2286 12426 2320
rect 12494 2286 12510 2320
rect 7648 2182 7682 2244
rect 12656 2182 12690 2244
rect 7648 2148 7744 2182
rect 12594 2148 12690 2182
rect 14128 2286 14144 2320
rect 14212 2286 14228 2320
rect 14286 2286 14302 2320
rect 14370 2286 14386 2320
rect 14444 2286 14460 2320
rect 14528 2286 14544 2320
rect 14602 2286 14618 2320
rect 14686 2286 14702 2320
rect 14760 2286 14776 2320
rect 14844 2286 14860 2320
rect 14918 2286 14934 2320
rect 15002 2286 15018 2320
rect 15076 2286 15092 2320
rect 15160 2286 15176 2320
rect 15234 2286 15250 2320
rect 15318 2286 15334 2320
rect 15392 2286 15408 2320
rect 15476 2286 15492 2320
rect 15550 2286 15566 2320
rect 15634 2286 15650 2320
rect 15708 2286 15724 2320
rect 15792 2286 15808 2320
rect 15866 2286 15882 2320
rect 15950 2286 15966 2320
rect 16024 2286 16040 2320
rect 16108 2286 16124 2320
rect 16182 2286 16198 2320
rect 16266 2286 16282 2320
rect 16340 2286 16356 2320
rect 16424 2286 16440 2320
rect 16498 2286 16514 2320
rect 16582 2286 16598 2320
rect 16656 2286 16672 2320
rect 16740 2286 16756 2320
rect 16814 2286 16830 2320
rect 16898 2286 16914 2320
rect 16972 2286 16988 2320
rect 17056 2286 17072 2320
rect 17130 2286 17146 2320
rect 17214 2286 17230 2320
rect 17288 2286 17304 2320
rect 17372 2286 17388 2320
rect 17446 2286 17462 2320
rect 17530 2286 17546 2320
rect 17604 2286 17620 2320
rect 17688 2286 17704 2320
rect 17762 2286 17778 2320
rect 17846 2286 17862 2320
rect 17920 2286 17936 2320
rect 18004 2286 18020 2320
rect 18078 2286 18094 2320
rect 18162 2286 18178 2320
rect 18236 2286 18252 2320
rect 18320 2286 18336 2320
rect 18394 2286 18410 2320
rect 18478 2286 18494 2320
rect 18552 2286 18568 2320
rect 18636 2286 18652 2320
rect 18710 2286 18726 2320
rect 18794 2286 18810 2320
rect 13948 2182 13982 2244
rect 18956 2182 18990 2244
rect 13948 2148 14044 2182
rect 18894 2148 18990 2182
rect 20428 2286 20444 2320
rect 20512 2286 20528 2320
rect 20586 2286 20602 2320
rect 20670 2286 20686 2320
rect 20744 2286 20760 2320
rect 20828 2286 20844 2320
rect 20902 2286 20918 2320
rect 20986 2286 21002 2320
rect 21060 2286 21076 2320
rect 21144 2286 21160 2320
rect 21218 2286 21234 2320
rect 21302 2286 21318 2320
rect 21376 2286 21392 2320
rect 21460 2286 21476 2320
rect 21534 2286 21550 2320
rect 21618 2286 21634 2320
rect 21692 2286 21708 2320
rect 21776 2286 21792 2320
rect 21850 2286 21866 2320
rect 21934 2286 21950 2320
rect 22008 2286 22024 2320
rect 22092 2286 22108 2320
rect 22166 2286 22182 2320
rect 22250 2286 22266 2320
rect 22324 2286 22340 2320
rect 22408 2286 22424 2320
rect 22482 2286 22498 2320
rect 22566 2286 22582 2320
rect 22640 2286 22656 2320
rect 22724 2286 22740 2320
rect 22798 2286 22814 2320
rect 22882 2286 22898 2320
rect 22956 2286 22972 2320
rect 23040 2286 23056 2320
rect 23114 2286 23130 2320
rect 23198 2286 23214 2320
rect 23272 2286 23288 2320
rect 23356 2286 23372 2320
rect 23430 2286 23446 2320
rect 23514 2286 23530 2320
rect 23588 2286 23604 2320
rect 23672 2286 23688 2320
rect 23746 2286 23762 2320
rect 23830 2286 23846 2320
rect 23904 2286 23920 2320
rect 23988 2286 24004 2320
rect 24062 2286 24078 2320
rect 24146 2286 24162 2320
rect 24220 2286 24236 2320
rect 24304 2286 24320 2320
rect 24378 2286 24394 2320
rect 24462 2286 24478 2320
rect 24536 2286 24552 2320
rect 24620 2286 24636 2320
rect 24694 2286 24710 2320
rect 24778 2286 24794 2320
rect 24852 2286 24868 2320
rect 24936 2286 24952 2320
rect 25010 2286 25026 2320
rect 25094 2286 25110 2320
rect 20248 2182 20282 2244
rect 25256 2182 25290 2244
rect 20248 2148 20344 2182
rect 25194 2148 25290 2182
<< viali >>
rect 1536 46168 6259 46170
rect 7836 46168 12559 46170
rect 14136 46168 18859 46170
rect 20436 46168 25159 46170
rect 1536 46134 6259 46168
rect 1536 46132 6259 46134
rect 1544 45996 1612 46030
rect 1702 45996 1770 46030
rect 1860 45996 1928 46030
rect 2018 45996 2086 46030
rect 2176 45996 2244 46030
rect 2334 45996 2402 46030
rect 2492 45996 2560 46030
rect 2650 45996 2718 46030
rect 2808 45996 2876 46030
rect 2966 45996 3034 46030
rect 3124 45996 3192 46030
rect 3282 45996 3350 46030
rect 3440 45996 3508 46030
rect 3598 45996 3666 46030
rect 3756 45996 3824 46030
rect 3914 45996 3982 46030
rect 4072 45996 4140 46030
rect 4230 45996 4298 46030
rect 4388 45996 4456 46030
rect 4546 45996 4614 46030
rect 4704 45996 4772 46030
rect 4862 45996 4930 46030
rect 5020 45996 5088 46030
rect 5178 45996 5246 46030
rect 5336 45996 5404 46030
rect 5494 45996 5562 46030
rect 5652 45996 5720 46030
rect 5810 45996 5878 46030
rect 5968 45996 6036 46030
rect 6126 45996 6194 46030
rect 7836 46134 12559 46168
rect 7836 46132 12559 46134
rect 7844 45996 7912 46030
rect 8002 45996 8070 46030
rect 8160 45996 8228 46030
rect 8318 45996 8386 46030
rect 8476 45996 8544 46030
rect 8634 45996 8702 46030
rect 8792 45996 8860 46030
rect 8950 45996 9018 46030
rect 9108 45996 9176 46030
rect 9266 45996 9334 46030
rect 9424 45996 9492 46030
rect 9582 45996 9650 46030
rect 9740 45996 9808 46030
rect 9898 45996 9966 46030
rect 10056 45996 10124 46030
rect 10214 45996 10282 46030
rect 10372 45996 10440 46030
rect 10530 45996 10598 46030
rect 10688 45996 10756 46030
rect 10846 45996 10914 46030
rect 11004 45996 11072 46030
rect 11162 45996 11230 46030
rect 11320 45996 11388 46030
rect 11478 45996 11546 46030
rect 11636 45996 11704 46030
rect 11794 45996 11862 46030
rect 11952 45996 12020 46030
rect 12110 45996 12178 46030
rect 12268 45996 12336 46030
rect 12426 45996 12494 46030
rect 14136 46134 18859 46168
rect 14136 46132 18859 46134
rect 14144 45996 14212 46030
rect 14302 45996 14370 46030
rect 14460 45996 14528 46030
rect 14618 45996 14686 46030
rect 14776 45996 14844 46030
rect 14934 45996 15002 46030
rect 15092 45996 15160 46030
rect 15250 45996 15318 46030
rect 15408 45996 15476 46030
rect 15566 45996 15634 46030
rect 15724 45996 15792 46030
rect 15882 45996 15950 46030
rect 16040 45996 16108 46030
rect 16198 45996 16266 46030
rect 16356 45996 16424 46030
rect 16514 45996 16582 46030
rect 16672 45996 16740 46030
rect 16830 45996 16898 46030
rect 16988 45996 17056 46030
rect 17146 45996 17214 46030
rect 17304 45996 17372 46030
rect 17462 45996 17530 46030
rect 17620 45996 17688 46030
rect 17778 45996 17846 46030
rect 17936 45996 18004 46030
rect 18094 45996 18162 46030
rect 18252 45996 18320 46030
rect 18410 45996 18478 46030
rect 18568 45996 18636 46030
rect 18726 45996 18794 46030
rect 20436 46134 25159 46168
rect 20436 46132 25159 46134
rect 20444 45996 20512 46030
rect 20602 45996 20670 46030
rect 20760 45996 20828 46030
rect 20918 45996 20986 46030
rect 21076 45996 21144 46030
rect 21234 45996 21302 46030
rect 21392 45996 21460 46030
rect 21550 45996 21618 46030
rect 21708 45996 21776 46030
rect 21866 45996 21934 46030
rect 22024 45996 22092 46030
rect 22182 45996 22250 46030
rect 22340 45996 22408 46030
rect 22498 45996 22566 46030
rect 22656 45996 22724 46030
rect 22814 45996 22882 46030
rect 22972 45996 23040 46030
rect 23130 45996 23198 46030
rect 23288 45996 23356 46030
rect 23446 45996 23514 46030
rect 23604 45996 23672 46030
rect 23762 45996 23830 46030
rect 23920 45996 23988 46030
rect 24078 45996 24146 46030
rect 24236 45996 24304 46030
rect 24394 45996 24462 46030
rect 24552 45996 24620 46030
rect 24710 45996 24778 46030
rect 24868 45996 24936 46030
rect 25026 45996 25094 46030
rect -3040 40326 -3000 40400
rect -3218 40242 -3184 40276
rect -3218 40236 -3184 40242
rect -3218 38896 -3184 38902
rect -3218 38862 -3184 38896
rect -3040 38812 -3038 40326
rect -3038 38812 -3000 40326
rect -3040 38740 -3000 38812
rect 1346 39936 1348 45980
rect 1348 39936 1382 45980
rect 1382 39936 1384 45980
rect 1482 39970 1516 45946
rect 1640 39970 1674 45946
rect 1798 39970 1832 45946
rect 1956 39970 1990 45946
rect 2114 39970 2148 45946
rect 2272 39970 2306 45946
rect 2430 39970 2464 45946
rect 2588 39970 2622 45946
rect 2746 39970 2780 45946
rect 2904 39970 2938 45946
rect 3062 39970 3096 45946
rect 3220 39970 3254 45946
rect 3378 39970 3412 45946
rect 3536 39970 3570 45946
rect 3694 39970 3728 45946
rect 3852 39970 3886 45946
rect 4010 39970 4044 45946
rect 4168 39970 4202 45946
rect 4326 39970 4360 45946
rect 4484 39970 4518 45946
rect 4642 39970 4676 45946
rect 4800 39970 4834 45946
rect 4958 39970 4992 45946
rect 5116 39970 5150 45946
rect 5274 39970 5308 45946
rect 5432 39970 5466 45946
rect 5590 39970 5624 45946
rect 5748 39970 5782 45946
rect 5906 39970 5940 45946
rect 6064 39970 6098 45946
rect 6222 39970 6256 45946
rect 6354 39936 6356 45980
rect 6356 39936 6390 45980
rect 6390 39936 6392 45980
rect 7646 39936 7648 45980
rect 7648 39936 7682 45980
rect 7682 39936 7684 45980
rect 7782 39970 7816 45946
rect 7940 39970 7974 45946
rect 8098 39970 8132 45946
rect 8256 39970 8290 45946
rect 8414 39970 8448 45946
rect 8572 39970 8606 45946
rect 8730 39970 8764 45946
rect 8888 39970 8922 45946
rect 9046 39970 9080 45946
rect 9204 39970 9238 45946
rect 9362 39970 9396 45946
rect 9520 39970 9554 45946
rect 9678 39970 9712 45946
rect 9836 39970 9870 45946
rect 9994 39970 10028 45946
rect 10152 39970 10186 45946
rect 10310 39970 10344 45946
rect 10468 39970 10502 45946
rect 10626 39970 10660 45946
rect 10784 39970 10818 45946
rect 10942 39970 10976 45946
rect 11100 39970 11134 45946
rect 11258 39970 11292 45946
rect 11416 39970 11450 45946
rect 11574 39970 11608 45946
rect 11732 39970 11766 45946
rect 11890 39970 11924 45946
rect 12048 39970 12082 45946
rect 12206 39970 12240 45946
rect 12364 39970 12398 45946
rect 12522 39970 12556 45946
rect 12654 39936 12656 45980
rect 12656 39936 12690 45980
rect 12690 39936 12692 45980
rect 13946 39936 13948 45980
rect 13948 39936 13982 45980
rect 13982 39936 13984 45980
rect 14082 39970 14116 45946
rect 14240 39970 14274 45946
rect 14398 39970 14432 45946
rect 14556 39970 14590 45946
rect 14714 39970 14748 45946
rect 14872 39970 14906 45946
rect 15030 39970 15064 45946
rect 15188 39970 15222 45946
rect 15346 39970 15380 45946
rect 15504 39970 15538 45946
rect 15662 39970 15696 45946
rect 15820 39970 15854 45946
rect 15978 39970 16012 45946
rect 16136 39970 16170 45946
rect 16294 39970 16328 45946
rect 16452 39970 16486 45946
rect 16610 39970 16644 45946
rect 16768 39970 16802 45946
rect 16926 39970 16960 45946
rect 17084 39970 17118 45946
rect 17242 39970 17276 45946
rect 17400 39970 17434 45946
rect 17558 39970 17592 45946
rect 17716 39970 17750 45946
rect 17874 39970 17908 45946
rect 18032 39970 18066 45946
rect 18190 39970 18224 45946
rect 18348 39970 18382 45946
rect 18506 39970 18540 45946
rect 18664 39970 18698 45946
rect 18822 39970 18856 45946
rect 18954 39936 18956 45980
rect 18956 39936 18990 45980
rect 18990 39936 18992 45980
rect 20246 39936 20248 45980
rect 20248 39936 20282 45980
rect 20282 39936 20284 45980
rect 20382 39970 20416 45946
rect 20540 39970 20574 45946
rect 20698 39970 20732 45946
rect 20856 39970 20890 45946
rect 21014 39970 21048 45946
rect 21172 39970 21206 45946
rect 21330 39970 21364 45946
rect 21488 39970 21522 45946
rect 21646 39970 21680 45946
rect 21804 39970 21838 45946
rect 21962 39970 21996 45946
rect 22120 39970 22154 45946
rect 22278 39970 22312 45946
rect 22436 39970 22470 45946
rect 22594 39970 22628 45946
rect 22752 39970 22786 45946
rect 22910 39970 22944 45946
rect 23068 39970 23102 45946
rect 23226 39970 23260 45946
rect 23384 39970 23418 45946
rect 23542 39970 23576 45946
rect 23700 39970 23734 45946
rect 23858 39970 23892 45946
rect 24016 39970 24050 45946
rect 24174 39970 24208 45946
rect 24332 39970 24366 45946
rect 24490 39970 24524 45946
rect 24648 39970 24682 45946
rect 24806 39970 24840 45946
rect 24964 39970 24998 45946
rect 25122 39970 25156 45946
rect 25254 39936 25256 45980
rect 25256 39936 25290 45980
rect 25290 39936 25292 45980
rect 1544 39886 1612 39920
rect 1702 39886 1770 39920
rect 1860 39886 1928 39920
rect 2018 39886 2086 39920
rect 2176 39886 2244 39920
rect 2334 39886 2402 39920
rect 2492 39886 2560 39920
rect 2650 39886 2718 39920
rect 2808 39886 2876 39920
rect 2966 39886 3034 39920
rect 3124 39886 3192 39920
rect 3282 39886 3350 39920
rect 3440 39886 3508 39920
rect 3598 39886 3666 39920
rect 3756 39886 3824 39920
rect 3914 39886 3982 39920
rect 4072 39886 4140 39920
rect 4230 39886 4298 39920
rect 4388 39886 4456 39920
rect 4546 39886 4614 39920
rect 4704 39886 4772 39920
rect 4862 39886 4930 39920
rect 5020 39886 5088 39920
rect 5178 39886 5246 39920
rect 5336 39886 5404 39920
rect 5494 39886 5562 39920
rect 5652 39886 5720 39920
rect 5810 39886 5878 39920
rect 5968 39886 6036 39920
rect 6126 39886 6194 39920
rect 1536 39782 6202 39784
rect 1536 39748 6202 39782
rect 7844 39886 7912 39920
rect 8002 39886 8070 39920
rect 8160 39886 8228 39920
rect 8318 39886 8386 39920
rect 8476 39886 8544 39920
rect 8634 39886 8702 39920
rect 8792 39886 8860 39920
rect 8950 39886 9018 39920
rect 9108 39886 9176 39920
rect 9266 39886 9334 39920
rect 9424 39886 9492 39920
rect 9582 39886 9650 39920
rect 9740 39886 9808 39920
rect 9898 39886 9966 39920
rect 10056 39886 10124 39920
rect 10214 39886 10282 39920
rect 10372 39886 10440 39920
rect 10530 39886 10598 39920
rect 10688 39886 10756 39920
rect 10846 39886 10914 39920
rect 11004 39886 11072 39920
rect 11162 39886 11230 39920
rect 11320 39886 11388 39920
rect 11478 39886 11546 39920
rect 11636 39886 11704 39920
rect 11794 39886 11862 39920
rect 11952 39886 12020 39920
rect 12110 39886 12178 39920
rect 12268 39886 12336 39920
rect 12426 39886 12494 39920
rect 7836 39782 12502 39784
rect 7836 39748 12502 39782
rect 14144 39886 14212 39920
rect 14302 39886 14370 39920
rect 14460 39886 14528 39920
rect 14618 39886 14686 39920
rect 14776 39886 14844 39920
rect 14934 39886 15002 39920
rect 15092 39886 15160 39920
rect 15250 39886 15318 39920
rect 15408 39886 15476 39920
rect 15566 39886 15634 39920
rect 15724 39886 15792 39920
rect 15882 39886 15950 39920
rect 16040 39886 16108 39920
rect 16198 39886 16266 39920
rect 16356 39886 16424 39920
rect 16514 39886 16582 39920
rect 16672 39886 16740 39920
rect 16830 39886 16898 39920
rect 16988 39886 17056 39920
rect 17146 39886 17214 39920
rect 17304 39886 17372 39920
rect 17462 39886 17530 39920
rect 17620 39886 17688 39920
rect 17778 39886 17846 39920
rect 17936 39886 18004 39920
rect 18094 39886 18162 39920
rect 18252 39886 18320 39920
rect 18410 39886 18478 39920
rect 18568 39886 18636 39920
rect 18726 39886 18794 39920
rect 14136 39782 18802 39784
rect 14136 39748 18802 39782
rect 20444 39886 20512 39920
rect 20602 39886 20670 39920
rect 20760 39886 20828 39920
rect 20918 39886 20986 39920
rect 21076 39886 21144 39920
rect 21234 39886 21302 39920
rect 21392 39886 21460 39920
rect 21550 39886 21618 39920
rect 21708 39886 21776 39920
rect 21866 39886 21934 39920
rect 22024 39886 22092 39920
rect 22182 39886 22250 39920
rect 22340 39886 22408 39920
rect 22498 39886 22566 39920
rect 22656 39886 22724 39920
rect 22814 39886 22882 39920
rect 22972 39886 23040 39920
rect 23130 39886 23198 39920
rect 23288 39886 23356 39920
rect 23446 39886 23514 39920
rect 23604 39886 23672 39920
rect 23762 39886 23830 39920
rect 23920 39886 23988 39920
rect 24078 39886 24146 39920
rect 24236 39886 24304 39920
rect 24394 39886 24462 39920
rect 24552 39886 24620 39920
rect 24710 39886 24778 39920
rect 24868 39886 24936 39920
rect 25026 39886 25094 39920
rect 20436 39782 25102 39784
rect 20436 39748 25102 39782
rect 1536 39746 6202 39748
rect 7836 39746 12502 39748
rect 14136 39746 18802 39748
rect 20436 39746 25102 39748
rect 1536 39168 6259 39170
rect 7836 39168 12559 39170
rect 14136 39168 18859 39170
rect 20436 39168 25159 39170
rect 1536 39134 6259 39168
rect 1536 39132 6259 39134
rect 1544 38996 1612 39030
rect 1702 38996 1770 39030
rect 1860 38996 1928 39030
rect 2018 38996 2086 39030
rect 2176 38996 2244 39030
rect 2334 38996 2402 39030
rect 2492 38996 2560 39030
rect 2650 38996 2718 39030
rect 2808 38996 2876 39030
rect 2966 38996 3034 39030
rect 3124 38996 3192 39030
rect 3282 38996 3350 39030
rect 3440 38996 3508 39030
rect 3598 38996 3666 39030
rect 3756 38996 3824 39030
rect 3914 38996 3982 39030
rect 4072 38996 4140 39030
rect 4230 38996 4298 39030
rect 4388 38996 4456 39030
rect 4546 38996 4614 39030
rect 4704 38996 4772 39030
rect 4862 38996 4930 39030
rect 5020 38996 5088 39030
rect 5178 38996 5246 39030
rect 5336 38996 5404 39030
rect 5494 38996 5562 39030
rect 5652 38996 5720 39030
rect 5810 38996 5878 39030
rect 5968 38996 6036 39030
rect 6126 38996 6194 39030
rect 7836 39134 12559 39168
rect 7836 39132 12559 39134
rect 7844 38996 7912 39030
rect 8002 38996 8070 39030
rect 8160 38996 8228 39030
rect 8318 38996 8386 39030
rect 8476 38996 8544 39030
rect 8634 38996 8702 39030
rect 8792 38996 8860 39030
rect 8950 38996 9018 39030
rect 9108 38996 9176 39030
rect 9266 38996 9334 39030
rect 9424 38996 9492 39030
rect 9582 38996 9650 39030
rect 9740 38996 9808 39030
rect 9898 38996 9966 39030
rect 10056 38996 10124 39030
rect 10214 38996 10282 39030
rect 10372 38996 10440 39030
rect 10530 38996 10598 39030
rect 10688 38996 10756 39030
rect 10846 38996 10914 39030
rect 11004 38996 11072 39030
rect 11162 38996 11230 39030
rect 11320 38996 11388 39030
rect 11478 38996 11546 39030
rect 11636 38996 11704 39030
rect 11794 38996 11862 39030
rect 11952 38996 12020 39030
rect 12110 38996 12178 39030
rect 12268 38996 12336 39030
rect 12426 38996 12494 39030
rect 14136 39134 18859 39168
rect 14136 39132 18859 39134
rect 14144 38996 14212 39030
rect 14302 38996 14370 39030
rect 14460 38996 14528 39030
rect 14618 38996 14686 39030
rect 14776 38996 14844 39030
rect 14934 38996 15002 39030
rect 15092 38996 15160 39030
rect 15250 38996 15318 39030
rect 15408 38996 15476 39030
rect 15566 38996 15634 39030
rect 15724 38996 15792 39030
rect 15882 38996 15950 39030
rect 16040 38996 16108 39030
rect 16198 38996 16266 39030
rect 16356 38996 16424 39030
rect 16514 38996 16582 39030
rect 16672 38996 16740 39030
rect 16830 38996 16898 39030
rect 16988 38996 17056 39030
rect 17146 38996 17214 39030
rect 17304 38996 17372 39030
rect 17462 38996 17530 39030
rect 17620 38996 17688 39030
rect 17778 38996 17846 39030
rect 17936 38996 18004 39030
rect 18094 38996 18162 39030
rect 18252 38996 18320 39030
rect 18410 38996 18478 39030
rect 18568 38996 18636 39030
rect 18726 38996 18794 39030
rect 20436 39134 25159 39168
rect 20436 39132 25159 39134
rect 20444 38996 20512 39030
rect 20602 38996 20670 39030
rect 20760 38996 20828 39030
rect 20918 38996 20986 39030
rect 21076 38996 21144 39030
rect 21234 38996 21302 39030
rect 21392 38996 21460 39030
rect 21550 38996 21618 39030
rect 21708 38996 21776 39030
rect 21866 38996 21934 39030
rect 22024 38996 22092 39030
rect 22182 38996 22250 39030
rect 22340 38996 22408 39030
rect 22498 38996 22566 39030
rect 22656 38996 22724 39030
rect 22814 38996 22882 39030
rect 22972 38996 23040 39030
rect 23130 38996 23198 39030
rect 23288 38996 23356 39030
rect 23446 38996 23514 39030
rect 23604 38996 23672 39030
rect 23762 38996 23830 39030
rect 23920 38996 23988 39030
rect 24078 38996 24146 39030
rect 24236 38996 24304 39030
rect 24394 38996 24462 39030
rect 24552 38996 24620 39030
rect 24710 38996 24778 39030
rect 24868 38996 24936 39030
rect 25026 38996 25094 39030
rect 1346 32936 1348 38980
rect 1348 32936 1382 38980
rect 1382 32936 1384 38980
rect 1482 32970 1516 38946
rect 1640 32970 1674 38946
rect 1798 32970 1832 38946
rect 1956 32970 1990 38946
rect 2114 32970 2148 38946
rect 2272 32970 2306 38946
rect 2430 32970 2464 38946
rect 2588 32970 2622 38946
rect 2746 32970 2780 38946
rect 2904 32970 2938 38946
rect 3062 32970 3096 38946
rect 3220 32970 3254 38946
rect 3378 32970 3412 38946
rect 3536 32970 3570 38946
rect 3694 32970 3728 38946
rect 3852 32970 3886 38946
rect 4010 32970 4044 38946
rect 4168 32970 4202 38946
rect 4326 32970 4360 38946
rect 4484 32970 4518 38946
rect 4642 32970 4676 38946
rect 4800 32970 4834 38946
rect 4958 32970 4992 38946
rect 5116 32970 5150 38946
rect 5274 32970 5308 38946
rect 5432 32970 5466 38946
rect 5590 32970 5624 38946
rect 5748 32970 5782 38946
rect 5906 32970 5940 38946
rect 6064 32970 6098 38946
rect 6222 32970 6256 38946
rect 6354 32936 6356 38980
rect 6356 32936 6390 38980
rect 6390 32936 6392 38980
rect 7646 32936 7648 38980
rect 7648 32936 7682 38980
rect 7682 32936 7684 38980
rect 7782 32970 7816 38946
rect 7940 32970 7974 38946
rect 8098 32970 8132 38946
rect 8256 32970 8290 38946
rect 8414 32970 8448 38946
rect 8572 32970 8606 38946
rect 8730 32970 8764 38946
rect 8888 32970 8922 38946
rect 9046 32970 9080 38946
rect 9204 32970 9238 38946
rect 9362 32970 9396 38946
rect 9520 32970 9554 38946
rect 9678 32970 9712 38946
rect 9836 32970 9870 38946
rect 9994 32970 10028 38946
rect 10152 32970 10186 38946
rect 10310 32970 10344 38946
rect 10468 32970 10502 38946
rect 10626 32970 10660 38946
rect 10784 32970 10818 38946
rect 10942 32970 10976 38946
rect 11100 32970 11134 38946
rect 11258 32970 11292 38946
rect 11416 32970 11450 38946
rect 11574 32970 11608 38946
rect 11732 32970 11766 38946
rect 11890 32970 11924 38946
rect 12048 32970 12082 38946
rect 12206 32970 12240 38946
rect 12364 32970 12398 38946
rect 12522 32970 12556 38946
rect 12654 32936 12656 38980
rect 12656 32936 12690 38980
rect 12690 32936 12692 38980
rect 13946 32936 13948 38980
rect 13948 32936 13982 38980
rect 13982 32936 13984 38980
rect 14082 32970 14116 38946
rect 14240 32970 14274 38946
rect 14398 32970 14432 38946
rect 14556 32970 14590 38946
rect 14714 32970 14748 38946
rect 14872 32970 14906 38946
rect 15030 32970 15064 38946
rect 15188 32970 15222 38946
rect 15346 32970 15380 38946
rect 15504 32970 15538 38946
rect 15662 32970 15696 38946
rect 15820 32970 15854 38946
rect 15978 32970 16012 38946
rect 16136 32970 16170 38946
rect 16294 32970 16328 38946
rect 16452 32970 16486 38946
rect 16610 32970 16644 38946
rect 16768 32970 16802 38946
rect 16926 32970 16960 38946
rect 17084 32970 17118 38946
rect 17242 32970 17276 38946
rect 17400 32970 17434 38946
rect 17558 32970 17592 38946
rect 17716 32970 17750 38946
rect 17874 32970 17908 38946
rect 18032 32970 18066 38946
rect 18190 32970 18224 38946
rect 18348 32970 18382 38946
rect 18506 32970 18540 38946
rect 18664 32970 18698 38946
rect 18822 32970 18856 38946
rect 18954 32936 18956 38980
rect 18956 32936 18990 38980
rect 18990 32936 18992 38980
rect 20246 32936 20248 38980
rect 20248 32936 20282 38980
rect 20282 32936 20284 38980
rect 20382 32970 20416 38946
rect 20540 32970 20574 38946
rect 20698 32970 20732 38946
rect 20856 32970 20890 38946
rect 21014 32970 21048 38946
rect 21172 32970 21206 38946
rect 21330 32970 21364 38946
rect 21488 32970 21522 38946
rect 21646 32970 21680 38946
rect 21804 32970 21838 38946
rect 21962 32970 21996 38946
rect 22120 32970 22154 38946
rect 22278 32970 22312 38946
rect 22436 32970 22470 38946
rect 22594 32970 22628 38946
rect 22752 32970 22786 38946
rect 22910 32970 22944 38946
rect 23068 32970 23102 38946
rect 23226 32970 23260 38946
rect 23384 32970 23418 38946
rect 23542 32970 23576 38946
rect 23700 32970 23734 38946
rect 23858 32970 23892 38946
rect 24016 32970 24050 38946
rect 24174 32970 24208 38946
rect 24332 32970 24366 38946
rect 24490 32970 24524 38946
rect 24648 32970 24682 38946
rect 24806 32970 24840 38946
rect 24964 32970 24998 38946
rect 25122 32970 25156 38946
rect 25254 32936 25256 38980
rect 25256 32936 25290 38980
rect 25290 32936 25292 38980
rect 29800 40326 29840 40400
rect 29800 38812 29838 40326
rect 29838 38812 29840 40326
rect 29984 40242 30018 40276
rect 29984 40236 30018 40242
rect 29984 38896 30018 38902
rect 29984 38862 30018 38896
rect 29800 38720 29840 38812
rect 1544 32886 1612 32920
rect 1702 32886 1770 32920
rect 1860 32886 1928 32920
rect 2018 32886 2086 32920
rect 2176 32886 2244 32920
rect 2334 32886 2402 32920
rect 2492 32886 2560 32920
rect 2650 32886 2718 32920
rect 2808 32886 2876 32920
rect 2966 32886 3034 32920
rect 3124 32886 3192 32920
rect 3282 32886 3350 32920
rect 3440 32886 3508 32920
rect 3598 32886 3666 32920
rect 3756 32886 3824 32920
rect 3914 32886 3982 32920
rect 4072 32886 4140 32920
rect 4230 32886 4298 32920
rect 4388 32886 4456 32920
rect 4546 32886 4614 32920
rect 4704 32886 4772 32920
rect 4862 32886 4930 32920
rect 5020 32886 5088 32920
rect 5178 32886 5246 32920
rect 5336 32886 5404 32920
rect 5494 32886 5562 32920
rect 5652 32886 5720 32920
rect 5810 32886 5878 32920
rect 5968 32886 6036 32920
rect 6126 32886 6194 32920
rect 1536 32782 6202 32784
rect 1536 32748 6202 32782
rect 7844 32886 7912 32920
rect 8002 32886 8070 32920
rect 8160 32886 8228 32920
rect 8318 32886 8386 32920
rect 8476 32886 8544 32920
rect 8634 32886 8702 32920
rect 8792 32886 8860 32920
rect 8950 32886 9018 32920
rect 9108 32886 9176 32920
rect 9266 32886 9334 32920
rect 9424 32886 9492 32920
rect 9582 32886 9650 32920
rect 9740 32886 9808 32920
rect 9898 32886 9966 32920
rect 10056 32886 10124 32920
rect 10214 32886 10282 32920
rect 10372 32886 10440 32920
rect 10530 32886 10598 32920
rect 10688 32886 10756 32920
rect 10846 32886 10914 32920
rect 11004 32886 11072 32920
rect 11162 32886 11230 32920
rect 11320 32886 11388 32920
rect 11478 32886 11546 32920
rect 11636 32886 11704 32920
rect 11794 32886 11862 32920
rect 11952 32886 12020 32920
rect 12110 32886 12178 32920
rect 12268 32886 12336 32920
rect 12426 32886 12494 32920
rect 7836 32782 12502 32784
rect 7836 32748 12502 32782
rect 14144 32886 14212 32920
rect 14302 32886 14370 32920
rect 14460 32886 14528 32920
rect 14618 32886 14686 32920
rect 14776 32886 14844 32920
rect 14934 32886 15002 32920
rect 15092 32886 15160 32920
rect 15250 32886 15318 32920
rect 15408 32886 15476 32920
rect 15566 32886 15634 32920
rect 15724 32886 15792 32920
rect 15882 32886 15950 32920
rect 16040 32886 16108 32920
rect 16198 32886 16266 32920
rect 16356 32886 16424 32920
rect 16514 32886 16582 32920
rect 16672 32886 16740 32920
rect 16830 32886 16898 32920
rect 16988 32886 17056 32920
rect 17146 32886 17214 32920
rect 17304 32886 17372 32920
rect 17462 32886 17530 32920
rect 17620 32886 17688 32920
rect 17778 32886 17846 32920
rect 17936 32886 18004 32920
rect 18094 32886 18162 32920
rect 18252 32886 18320 32920
rect 18410 32886 18478 32920
rect 18568 32886 18636 32920
rect 18726 32886 18794 32920
rect 14136 32782 18802 32784
rect 14136 32748 18802 32782
rect 20444 32886 20512 32920
rect 20602 32886 20670 32920
rect 20760 32886 20828 32920
rect 20918 32886 20986 32920
rect 21076 32886 21144 32920
rect 21234 32886 21302 32920
rect 21392 32886 21460 32920
rect 21550 32886 21618 32920
rect 21708 32886 21776 32920
rect 21866 32886 21934 32920
rect 22024 32886 22092 32920
rect 22182 32886 22250 32920
rect 22340 32886 22408 32920
rect 22498 32886 22566 32920
rect 22656 32886 22724 32920
rect 22814 32886 22882 32920
rect 22972 32886 23040 32920
rect 23130 32886 23198 32920
rect 23288 32886 23356 32920
rect 23446 32886 23514 32920
rect 23604 32886 23672 32920
rect 23762 32886 23830 32920
rect 23920 32886 23988 32920
rect 24078 32886 24146 32920
rect 24236 32886 24304 32920
rect 24394 32886 24462 32920
rect 24552 32886 24620 32920
rect 24710 32886 24778 32920
rect 24868 32886 24936 32920
rect 25026 32886 25094 32920
rect 20436 32782 25102 32784
rect 20436 32748 25102 32782
rect 1536 32746 6202 32748
rect 7836 32746 12502 32748
rect 14136 32746 18802 32748
rect 20436 32746 25102 32748
rect 1536 30868 6259 30870
rect 7836 30868 12559 30870
rect 14136 30868 18859 30870
rect 20436 30868 25159 30870
rect 1536 30834 6259 30868
rect 1536 30832 6259 30834
rect 1544 30696 1612 30730
rect 1702 30696 1770 30730
rect 1860 30696 1928 30730
rect 2018 30696 2086 30730
rect 2176 30696 2244 30730
rect 2334 30696 2402 30730
rect 2492 30696 2560 30730
rect 2650 30696 2718 30730
rect 2808 30696 2876 30730
rect 2966 30696 3034 30730
rect 3124 30696 3192 30730
rect 3282 30696 3350 30730
rect 3440 30696 3508 30730
rect 3598 30696 3666 30730
rect 3756 30696 3824 30730
rect 3914 30696 3982 30730
rect 4072 30696 4140 30730
rect 4230 30696 4298 30730
rect 4388 30696 4456 30730
rect 4546 30696 4614 30730
rect 4704 30696 4772 30730
rect 4862 30696 4930 30730
rect 5020 30696 5088 30730
rect 5178 30696 5246 30730
rect 5336 30696 5404 30730
rect 5494 30696 5562 30730
rect 5652 30696 5720 30730
rect 5810 30696 5878 30730
rect 5968 30696 6036 30730
rect 6126 30696 6194 30730
rect 7836 30834 12559 30868
rect 7836 30832 12559 30834
rect 7844 30696 7912 30730
rect 8002 30696 8070 30730
rect 8160 30696 8228 30730
rect 8318 30696 8386 30730
rect 8476 30696 8544 30730
rect 8634 30696 8702 30730
rect 8792 30696 8860 30730
rect 8950 30696 9018 30730
rect 9108 30696 9176 30730
rect 9266 30696 9334 30730
rect 9424 30696 9492 30730
rect 9582 30696 9650 30730
rect 9740 30696 9808 30730
rect 9898 30696 9966 30730
rect 10056 30696 10124 30730
rect 10214 30696 10282 30730
rect 10372 30696 10440 30730
rect 10530 30696 10598 30730
rect 10688 30696 10756 30730
rect 10846 30696 10914 30730
rect 11004 30696 11072 30730
rect 11162 30696 11230 30730
rect 11320 30696 11388 30730
rect 11478 30696 11546 30730
rect 11636 30696 11704 30730
rect 11794 30696 11862 30730
rect 11952 30696 12020 30730
rect 12110 30696 12178 30730
rect 12268 30696 12336 30730
rect 12426 30696 12494 30730
rect 14136 30834 18859 30868
rect 14136 30832 18859 30834
rect 14144 30696 14212 30730
rect 14302 30696 14370 30730
rect 14460 30696 14528 30730
rect 14618 30696 14686 30730
rect 14776 30696 14844 30730
rect 14934 30696 15002 30730
rect 15092 30696 15160 30730
rect 15250 30696 15318 30730
rect 15408 30696 15476 30730
rect 15566 30696 15634 30730
rect 15724 30696 15792 30730
rect 15882 30696 15950 30730
rect 16040 30696 16108 30730
rect 16198 30696 16266 30730
rect 16356 30696 16424 30730
rect 16514 30696 16582 30730
rect 16672 30696 16740 30730
rect 16830 30696 16898 30730
rect 16988 30696 17056 30730
rect 17146 30696 17214 30730
rect 17304 30696 17372 30730
rect 17462 30696 17530 30730
rect 17620 30696 17688 30730
rect 17778 30696 17846 30730
rect 17936 30696 18004 30730
rect 18094 30696 18162 30730
rect 18252 30696 18320 30730
rect 18410 30696 18478 30730
rect 18568 30696 18636 30730
rect 18726 30696 18794 30730
rect 20436 30834 25159 30868
rect 20436 30832 25159 30834
rect 20444 30696 20512 30730
rect 20602 30696 20670 30730
rect 20760 30696 20828 30730
rect 20918 30696 20986 30730
rect 21076 30696 21144 30730
rect 21234 30696 21302 30730
rect 21392 30696 21460 30730
rect 21550 30696 21618 30730
rect 21708 30696 21776 30730
rect 21866 30696 21934 30730
rect 22024 30696 22092 30730
rect 22182 30696 22250 30730
rect 22340 30696 22408 30730
rect 22498 30696 22566 30730
rect 22656 30696 22724 30730
rect 22814 30696 22882 30730
rect 22972 30696 23040 30730
rect 23130 30696 23198 30730
rect 23288 30696 23356 30730
rect 23446 30696 23514 30730
rect 23604 30696 23672 30730
rect 23762 30696 23830 30730
rect 23920 30696 23988 30730
rect 24078 30696 24146 30730
rect 24236 30696 24304 30730
rect 24394 30696 24462 30730
rect 24552 30696 24620 30730
rect 24710 30696 24778 30730
rect 24868 30696 24936 30730
rect 25026 30696 25094 30730
rect -4040 27126 -4000 27200
rect -4218 27042 -4184 27076
rect -4218 27036 -4184 27042
rect -4218 25696 -4184 25702
rect -4218 25662 -4184 25696
rect -4040 25612 -4038 27126
rect -4038 25612 -4000 27126
rect -4040 25540 -4000 25612
rect 1346 24636 1348 30680
rect 1348 24636 1382 30680
rect 1382 24636 1384 30680
rect 1482 24670 1516 30646
rect 1640 24670 1674 30646
rect 1798 24670 1832 30646
rect 1956 24670 1990 30646
rect 2114 24670 2148 30646
rect 2272 24670 2306 30646
rect 2430 24670 2464 30646
rect 2588 24670 2622 30646
rect 2746 24670 2780 30646
rect 2904 24670 2938 30646
rect 3062 24670 3096 30646
rect 3220 24670 3254 30646
rect 3378 24670 3412 30646
rect 3536 24670 3570 30646
rect 3694 24670 3728 30646
rect 3852 24670 3886 30646
rect 4010 24670 4044 30646
rect 4168 24670 4202 30646
rect 4326 24670 4360 30646
rect 4484 24670 4518 30646
rect 4642 24670 4676 30646
rect 4800 24670 4834 30646
rect 4958 24670 4992 30646
rect 5116 24670 5150 30646
rect 5274 24670 5308 30646
rect 5432 24670 5466 30646
rect 5590 24670 5624 30646
rect 5748 24670 5782 30646
rect 5906 24670 5940 30646
rect 6064 24670 6098 30646
rect 6222 24670 6256 30646
rect 6354 24636 6356 30680
rect 6356 24636 6390 30680
rect 6390 24636 6392 30680
rect 7646 24636 7648 30680
rect 7648 24636 7682 30680
rect 7682 24636 7684 30680
rect 7782 24670 7816 30646
rect 7940 24670 7974 30646
rect 8098 24670 8132 30646
rect 8256 24670 8290 30646
rect 8414 24670 8448 30646
rect 8572 24670 8606 30646
rect 8730 24670 8764 30646
rect 8888 24670 8922 30646
rect 9046 24670 9080 30646
rect 9204 24670 9238 30646
rect 9362 24670 9396 30646
rect 9520 24670 9554 30646
rect 9678 24670 9712 30646
rect 9836 24670 9870 30646
rect 9994 24670 10028 30646
rect 10152 24670 10186 30646
rect 10310 24670 10344 30646
rect 10468 24670 10502 30646
rect 10626 24670 10660 30646
rect 10784 24670 10818 30646
rect 10942 24670 10976 30646
rect 11100 24670 11134 30646
rect 11258 24670 11292 30646
rect 11416 24670 11450 30646
rect 11574 24670 11608 30646
rect 11732 24670 11766 30646
rect 11890 24670 11924 30646
rect 12048 24670 12082 30646
rect 12206 24670 12240 30646
rect 12364 24670 12398 30646
rect 12522 24670 12556 30646
rect 12654 24636 12656 30680
rect 12656 24636 12690 30680
rect 12690 24636 12692 30680
rect 13946 24636 13948 30680
rect 13948 24636 13982 30680
rect 13982 24636 13984 30680
rect 14082 24670 14116 30646
rect 14240 24670 14274 30646
rect 14398 24670 14432 30646
rect 14556 24670 14590 30646
rect 14714 24670 14748 30646
rect 14872 24670 14906 30646
rect 15030 24670 15064 30646
rect 15188 24670 15222 30646
rect 15346 24670 15380 30646
rect 15504 24670 15538 30646
rect 15662 24670 15696 30646
rect 15820 24670 15854 30646
rect 15978 24670 16012 30646
rect 16136 24670 16170 30646
rect 16294 24670 16328 30646
rect 16452 24670 16486 30646
rect 16610 24670 16644 30646
rect 16768 24670 16802 30646
rect 16926 24670 16960 30646
rect 17084 24670 17118 30646
rect 17242 24670 17276 30646
rect 17400 24670 17434 30646
rect 17558 24670 17592 30646
rect 17716 24670 17750 30646
rect 17874 24670 17908 30646
rect 18032 24670 18066 30646
rect 18190 24670 18224 30646
rect 18348 24670 18382 30646
rect 18506 24670 18540 30646
rect 18664 24670 18698 30646
rect 18822 24670 18856 30646
rect 18954 24636 18956 30680
rect 18956 24636 18990 30680
rect 18990 24636 18992 30680
rect 20246 24636 20248 30680
rect 20248 24636 20282 30680
rect 20282 24636 20284 30680
rect 20382 24670 20416 30646
rect 20540 24670 20574 30646
rect 20698 24670 20732 30646
rect 20856 24670 20890 30646
rect 21014 24670 21048 30646
rect 21172 24670 21206 30646
rect 21330 24670 21364 30646
rect 21488 24670 21522 30646
rect 21646 24670 21680 30646
rect 21804 24670 21838 30646
rect 21962 24670 21996 30646
rect 22120 24670 22154 30646
rect 22278 24670 22312 30646
rect 22436 24670 22470 30646
rect 22594 24670 22628 30646
rect 22752 24670 22786 30646
rect 22910 24670 22944 30646
rect 23068 24670 23102 30646
rect 23226 24670 23260 30646
rect 23384 24670 23418 30646
rect 23542 24670 23576 30646
rect 23700 24670 23734 30646
rect 23858 24670 23892 30646
rect 24016 24670 24050 30646
rect 24174 24670 24208 30646
rect 24332 24670 24366 30646
rect 24490 24670 24524 30646
rect 24648 24670 24682 30646
rect 24806 24670 24840 30646
rect 24964 24670 24998 30646
rect 25122 24670 25156 30646
rect 25254 24636 25256 30680
rect 25256 24636 25290 30680
rect 25290 24636 25292 30680
rect 30984 27042 31018 27076
rect 30984 27036 31018 27042
rect 30800 26020 30838 26980
rect 30838 26020 30840 26980
rect 30984 25696 31018 25702
rect 30984 25662 31018 25696
rect 1544 24586 1612 24620
rect 1702 24586 1770 24620
rect 1860 24586 1928 24620
rect 2018 24586 2086 24620
rect 2176 24586 2244 24620
rect 2334 24586 2402 24620
rect 2492 24586 2560 24620
rect 2650 24586 2718 24620
rect 2808 24586 2876 24620
rect 2966 24586 3034 24620
rect 3124 24586 3192 24620
rect 3282 24586 3350 24620
rect 3440 24586 3508 24620
rect 3598 24586 3666 24620
rect 3756 24586 3824 24620
rect 3914 24586 3982 24620
rect 4072 24586 4140 24620
rect 4230 24586 4298 24620
rect 4388 24586 4456 24620
rect 4546 24586 4614 24620
rect 4704 24586 4772 24620
rect 4862 24586 4930 24620
rect 5020 24586 5088 24620
rect 5178 24586 5246 24620
rect 5336 24586 5404 24620
rect 5494 24586 5562 24620
rect 5652 24586 5720 24620
rect 5810 24586 5878 24620
rect 5968 24586 6036 24620
rect 6126 24586 6194 24620
rect 1536 24482 6202 24484
rect 1536 24448 6202 24482
rect 7844 24586 7912 24620
rect 8002 24586 8070 24620
rect 8160 24586 8228 24620
rect 8318 24586 8386 24620
rect 8476 24586 8544 24620
rect 8634 24586 8702 24620
rect 8792 24586 8860 24620
rect 8950 24586 9018 24620
rect 9108 24586 9176 24620
rect 9266 24586 9334 24620
rect 9424 24586 9492 24620
rect 9582 24586 9650 24620
rect 9740 24586 9808 24620
rect 9898 24586 9966 24620
rect 10056 24586 10124 24620
rect 10214 24586 10282 24620
rect 10372 24586 10440 24620
rect 10530 24586 10598 24620
rect 10688 24586 10756 24620
rect 10846 24586 10914 24620
rect 11004 24586 11072 24620
rect 11162 24586 11230 24620
rect 11320 24586 11388 24620
rect 11478 24586 11546 24620
rect 11636 24586 11704 24620
rect 11794 24586 11862 24620
rect 11952 24586 12020 24620
rect 12110 24586 12178 24620
rect 12268 24586 12336 24620
rect 12426 24586 12494 24620
rect 7836 24482 12502 24484
rect 7836 24448 12502 24482
rect 14144 24586 14212 24620
rect 14302 24586 14370 24620
rect 14460 24586 14528 24620
rect 14618 24586 14686 24620
rect 14776 24586 14844 24620
rect 14934 24586 15002 24620
rect 15092 24586 15160 24620
rect 15250 24586 15318 24620
rect 15408 24586 15476 24620
rect 15566 24586 15634 24620
rect 15724 24586 15792 24620
rect 15882 24586 15950 24620
rect 16040 24586 16108 24620
rect 16198 24586 16266 24620
rect 16356 24586 16424 24620
rect 16514 24586 16582 24620
rect 16672 24586 16740 24620
rect 16830 24586 16898 24620
rect 16988 24586 17056 24620
rect 17146 24586 17214 24620
rect 17304 24586 17372 24620
rect 17462 24586 17530 24620
rect 17620 24586 17688 24620
rect 17778 24586 17846 24620
rect 17936 24586 18004 24620
rect 18094 24586 18162 24620
rect 18252 24586 18320 24620
rect 18410 24586 18478 24620
rect 18568 24586 18636 24620
rect 18726 24586 18794 24620
rect 14136 24482 18802 24484
rect 14136 24448 18802 24482
rect 20444 24586 20512 24620
rect 20602 24586 20670 24620
rect 20760 24586 20828 24620
rect 20918 24586 20986 24620
rect 21076 24586 21144 24620
rect 21234 24586 21302 24620
rect 21392 24586 21460 24620
rect 21550 24586 21618 24620
rect 21708 24586 21776 24620
rect 21866 24586 21934 24620
rect 22024 24586 22092 24620
rect 22182 24586 22250 24620
rect 22340 24586 22408 24620
rect 22498 24586 22566 24620
rect 22656 24586 22724 24620
rect 22814 24586 22882 24620
rect 22972 24586 23040 24620
rect 23130 24586 23198 24620
rect 23288 24586 23356 24620
rect 23446 24586 23514 24620
rect 23604 24586 23672 24620
rect 23762 24586 23830 24620
rect 23920 24586 23988 24620
rect 24078 24586 24146 24620
rect 24236 24586 24304 24620
rect 24394 24586 24462 24620
rect 24552 24586 24620 24620
rect 24710 24586 24778 24620
rect 24868 24586 24936 24620
rect 25026 24586 25094 24620
rect 20436 24482 25102 24484
rect 20436 24448 25102 24482
rect 1536 24446 6202 24448
rect 7836 24446 12502 24448
rect 14136 24446 18802 24448
rect 20436 24446 25102 24448
rect 1536 23868 6259 23870
rect 7836 23868 12559 23870
rect 14136 23868 18859 23870
rect 20436 23868 25159 23870
rect 1536 23834 6259 23868
rect 1536 23832 6259 23834
rect 1544 23696 1612 23730
rect 1702 23696 1770 23730
rect 1860 23696 1928 23730
rect 2018 23696 2086 23730
rect 2176 23696 2244 23730
rect 2334 23696 2402 23730
rect 2492 23696 2560 23730
rect 2650 23696 2718 23730
rect 2808 23696 2876 23730
rect 2966 23696 3034 23730
rect 3124 23696 3192 23730
rect 3282 23696 3350 23730
rect 3440 23696 3508 23730
rect 3598 23696 3666 23730
rect 3756 23696 3824 23730
rect 3914 23696 3982 23730
rect 4072 23696 4140 23730
rect 4230 23696 4298 23730
rect 4388 23696 4456 23730
rect 4546 23696 4614 23730
rect 4704 23696 4772 23730
rect 4862 23696 4930 23730
rect 5020 23696 5088 23730
rect 5178 23696 5246 23730
rect 5336 23696 5404 23730
rect 5494 23696 5562 23730
rect 5652 23696 5720 23730
rect 5810 23696 5878 23730
rect 5968 23696 6036 23730
rect 6126 23696 6194 23730
rect 7836 23834 12559 23868
rect 7836 23832 12559 23834
rect 7844 23696 7912 23730
rect 8002 23696 8070 23730
rect 8160 23696 8228 23730
rect 8318 23696 8386 23730
rect 8476 23696 8544 23730
rect 8634 23696 8702 23730
rect 8792 23696 8860 23730
rect 8950 23696 9018 23730
rect 9108 23696 9176 23730
rect 9266 23696 9334 23730
rect 9424 23696 9492 23730
rect 9582 23696 9650 23730
rect 9740 23696 9808 23730
rect 9898 23696 9966 23730
rect 10056 23696 10124 23730
rect 10214 23696 10282 23730
rect 10372 23696 10440 23730
rect 10530 23696 10598 23730
rect 10688 23696 10756 23730
rect 10846 23696 10914 23730
rect 11004 23696 11072 23730
rect 11162 23696 11230 23730
rect 11320 23696 11388 23730
rect 11478 23696 11546 23730
rect 11636 23696 11704 23730
rect 11794 23696 11862 23730
rect 11952 23696 12020 23730
rect 12110 23696 12178 23730
rect 12268 23696 12336 23730
rect 12426 23696 12494 23730
rect 14136 23834 18859 23868
rect 14136 23832 18859 23834
rect 14144 23696 14212 23730
rect 14302 23696 14370 23730
rect 14460 23696 14528 23730
rect 14618 23696 14686 23730
rect 14776 23696 14844 23730
rect 14934 23696 15002 23730
rect 15092 23696 15160 23730
rect 15250 23696 15318 23730
rect 15408 23696 15476 23730
rect 15566 23696 15634 23730
rect 15724 23696 15792 23730
rect 15882 23696 15950 23730
rect 16040 23696 16108 23730
rect 16198 23696 16266 23730
rect 16356 23696 16424 23730
rect 16514 23696 16582 23730
rect 16672 23696 16740 23730
rect 16830 23696 16898 23730
rect 16988 23696 17056 23730
rect 17146 23696 17214 23730
rect 17304 23696 17372 23730
rect 17462 23696 17530 23730
rect 17620 23696 17688 23730
rect 17778 23696 17846 23730
rect 17936 23696 18004 23730
rect 18094 23696 18162 23730
rect 18252 23696 18320 23730
rect 18410 23696 18478 23730
rect 18568 23696 18636 23730
rect 18726 23696 18794 23730
rect 20436 23834 25159 23868
rect 20436 23832 25159 23834
rect 20444 23696 20512 23730
rect 20602 23696 20670 23730
rect 20760 23696 20828 23730
rect 20918 23696 20986 23730
rect 21076 23696 21144 23730
rect 21234 23696 21302 23730
rect 21392 23696 21460 23730
rect 21550 23696 21618 23730
rect 21708 23696 21776 23730
rect 21866 23696 21934 23730
rect 22024 23696 22092 23730
rect 22182 23696 22250 23730
rect 22340 23696 22408 23730
rect 22498 23696 22566 23730
rect 22656 23696 22724 23730
rect 22814 23696 22882 23730
rect 22972 23696 23040 23730
rect 23130 23696 23198 23730
rect 23288 23696 23356 23730
rect 23446 23696 23514 23730
rect 23604 23696 23672 23730
rect 23762 23696 23830 23730
rect 23920 23696 23988 23730
rect 24078 23696 24146 23730
rect 24236 23696 24304 23730
rect 24394 23696 24462 23730
rect 24552 23696 24620 23730
rect 24710 23696 24778 23730
rect 24868 23696 24936 23730
rect 25026 23696 25094 23730
rect 1346 17636 1348 23680
rect 1348 17636 1382 23680
rect 1382 17636 1384 23680
rect 1482 17670 1516 23646
rect 1640 17670 1674 23646
rect 1798 17670 1832 23646
rect 1956 17670 1990 23646
rect 2114 17670 2148 23646
rect 2272 17670 2306 23646
rect 2430 17670 2464 23646
rect 2588 17670 2622 23646
rect 2746 17670 2780 23646
rect 2904 17670 2938 23646
rect 3062 17670 3096 23646
rect 3220 17670 3254 23646
rect 3378 17670 3412 23646
rect 3536 17670 3570 23646
rect 3694 17670 3728 23646
rect 3852 17670 3886 23646
rect 4010 17670 4044 23646
rect 4168 17670 4202 23646
rect 4326 17670 4360 23646
rect 4484 17670 4518 23646
rect 4642 17670 4676 23646
rect 4800 17670 4834 23646
rect 4958 17670 4992 23646
rect 5116 17670 5150 23646
rect 5274 17670 5308 23646
rect 5432 17670 5466 23646
rect 5590 17670 5624 23646
rect 5748 17670 5782 23646
rect 5906 17670 5940 23646
rect 6064 17670 6098 23646
rect 6222 17670 6256 23646
rect 6354 17636 6356 23680
rect 6356 17636 6390 23680
rect 6390 17636 6392 23680
rect 7646 17636 7648 23680
rect 7648 17636 7682 23680
rect 7682 17636 7684 23680
rect 7782 17670 7816 23646
rect 7940 17670 7974 23646
rect 8098 17670 8132 23646
rect 8256 17670 8290 23646
rect 8414 17670 8448 23646
rect 8572 17670 8606 23646
rect 8730 17670 8764 23646
rect 8888 17670 8922 23646
rect 9046 17670 9080 23646
rect 9204 17670 9238 23646
rect 9362 17670 9396 23646
rect 9520 17670 9554 23646
rect 9678 17670 9712 23646
rect 9836 17670 9870 23646
rect 9994 17670 10028 23646
rect 10152 17670 10186 23646
rect 10310 17670 10344 23646
rect 10468 17670 10502 23646
rect 10626 17670 10660 23646
rect 10784 17670 10818 23646
rect 10942 17670 10976 23646
rect 11100 17670 11134 23646
rect 11258 17670 11292 23646
rect 11416 17670 11450 23646
rect 11574 17670 11608 23646
rect 11732 17670 11766 23646
rect 11890 17670 11924 23646
rect 12048 17670 12082 23646
rect 12206 17670 12240 23646
rect 12364 17670 12398 23646
rect 12522 17670 12556 23646
rect 12654 17636 12656 23680
rect 12656 17636 12690 23680
rect 12690 17636 12692 23680
rect 13946 17636 13948 23680
rect 13948 17636 13982 23680
rect 13982 17636 13984 23680
rect 14082 17670 14116 23646
rect 14240 17670 14274 23646
rect 14398 17670 14432 23646
rect 14556 17670 14590 23646
rect 14714 17670 14748 23646
rect 14872 17670 14906 23646
rect 15030 17670 15064 23646
rect 15188 17670 15222 23646
rect 15346 17670 15380 23646
rect 15504 17670 15538 23646
rect 15662 17670 15696 23646
rect 15820 17670 15854 23646
rect 15978 17670 16012 23646
rect 16136 17670 16170 23646
rect 16294 17670 16328 23646
rect 16452 17670 16486 23646
rect 16610 17670 16644 23646
rect 16768 17670 16802 23646
rect 16926 17670 16960 23646
rect 17084 17670 17118 23646
rect 17242 17670 17276 23646
rect 17400 17670 17434 23646
rect 17558 17670 17592 23646
rect 17716 17670 17750 23646
rect 17874 17670 17908 23646
rect 18032 17670 18066 23646
rect 18190 17670 18224 23646
rect 18348 17670 18382 23646
rect 18506 17670 18540 23646
rect 18664 17670 18698 23646
rect 18822 17670 18856 23646
rect 18954 17636 18956 23680
rect 18956 17636 18990 23680
rect 18990 17636 18992 23680
rect 20246 17636 20248 23680
rect 20248 17636 20282 23680
rect 20282 17636 20284 23680
rect 20382 17670 20416 23646
rect 20540 17670 20574 23646
rect 20698 17670 20732 23646
rect 20856 17670 20890 23646
rect 21014 17670 21048 23646
rect 21172 17670 21206 23646
rect 21330 17670 21364 23646
rect 21488 17670 21522 23646
rect 21646 17670 21680 23646
rect 21804 17670 21838 23646
rect 21962 17670 21996 23646
rect 22120 17670 22154 23646
rect 22278 17670 22312 23646
rect 22436 17670 22470 23646
rect 22594 17670 22628 23646
rect 22752 17670 22786 23646
rect 22910 17670 22944 23646
rect 23068 17670 23102 23646
rect 23226 17670 23260 23646
rect 23384 17670 23418 23646
rect 23542 17670 23576 23646
rect 23700 17670 23734 23646
rect 23858 17670 23892 23646
rect 24016 17670 24050 23646
rect 24174 17670 24208 23646
rect 24332 17670 24366 23646
rect 24490 17670 24524 23646
rect 24648 17670 24682 23646
rect 24806 17670 24840 23646
rect 24964 17670 24998 23646
rect 25122 17670 25156 23646
rect 25254 17636 25256 23680
rect 25256 17636 25290 23680
rect 25290 17636 25292 23680
rect 1544 17586 1612 17620
rect 1702 17586 1770 17620
rect 1860 17586 1928 17620
rect 2018 17586 2086 17620
rect 2176 17586 2244 17620
rect 2334 17586 2402 17620
rect 2492 17586 2560 17620
rect 2650 17586 2718 17620
rect 2808 17586 2876 17620
rect 2966 17586 3034 17620
rect 3124 17586 3192 17620
rect 3282 17586 3350 17620
rect 3440 17586 3508 17620
rect 3598 17586 3666 17620
rect 3756 17586 3824 17620
rect 3914 17586 3982 17620
rect 4072 17586 4140 17620
rect 4230 17586 4298 17620
rect 4388 17586 4456 17620
rect 4546 17586 4614 17620
rect 4704 17586 4772 17620
rect 4862 17586 4930 17620
rect 5020 17586 5088 17620
rect 5178 17586 5246 17620
rect 5336 17586 5404 17620
rect 5494 17586 5562 17620
rect 5652 17586 5720 17620
rect 5810 17586 5878 17620
rect 5968 17586 6036 17620
rect 6126 17586 6194 17620
rect 1536 17482 6202 17484
rect 1536 17448 6202 17482
rect 7844 17586 7912 17620
rect 8002 17586 8070 17620
rect 8160 17586 8228 17620
rect 8318 17586 8386 17620
rect 8476 17586 8544 17620
rect 8634 17586 8702 17620
rect 8792 17586 8860 17620
rect 8950 17586 9018 17620
rect 9108 17586 9176 17620
rect 9266 17586 9334 17620
rect 9424 17586 9492 17620
rect 9582 17586 9650 17620
rect 9740 17586 9808 17620
rect 9898 17586 9966 17620
rect 10056 17586 10124 17620
rect 10214 17586 10282 17620
rect 10372 17586 10440 17620
rect 10530 17586 10598 17620
rect 10688 17586 10756 17620
rect 10846 17586 10914 17620
rect 11004 17586 11072 17620
rect 11162 17586 11230 17620
rect 11320 17586 11388 17620
rect 11478 17586 11546 17620
rect 11636 17586 11704 17620
rect 11794 17586 11862 17620
rect 11952 17586 12020 17620
rect 12110 17586 12178 17620
rect 12268 17586 12336 17620
rect 12426 17586 12494 17620
rect 7836 17482 12502 17484
rect 7836 17448 12502 17482
rect 14144 17586 14212 17620
rect 14302 17586 14370 17620
rect 14460 17586 14528 17620
rect 14618 17586 14686 17620
rect 14776 17586 14844 17620
rect 14934 17586 15002 17620
rect 15092 17586 15160 17620
rect 15250 17586 15318 17620
rect 15408 17586 15476 17620
rect 15566 17586 15634 17620
rect 15724 17586 15792 17620
rect 15882 17586 15950 17620
rect 16040 17586 16108 17620
rect 16198 17586 16266 17620
rect 16356 17586 16424 17620
rect 16514 17586 16582 17620
rect 16672 17586 16740 17620
rect 16830 17586 16898 17620
rect 16988 17586 17056 17620
rect 17146 17586 17214 17620
rect 17304 17586 17372 17620
rect 17462 17586 17530 17620
rect 17620 17586 17688 17620
rect 17778 17586 17846 17620
rect 17936 17586 18004 17620
rect 18094 17586 18162 17620
rect 18252 17586 18320 17620
rect 18410 17586 18478 17620
rect 18568 17586 18636 17620
rect 18726 17586 18794 17620
rect 14136 17482 18802 17484
rect 14136 17448 18802 17482
rect 20444 17586 20512 17620
rect 20602 17586 20670 17620
rect 20760 17586 20828 17620
rect 20918 17586 20986 17620
rect 21076 17586 21144 17620
rect 21234 17586 21302 17620
rect 21392 17586 21460 17620
rect 21550 17586 21618 17620
rect 21708 17586 21776 17620
rect 21866 17586 21934 17620
rect 22024 17586 22092 17620
rect 22182 17586 22250 17620
rect 22340 17586 22408 17620
rect 22498 17586 22566 17620
rect 22656 17586 22724 17620
rect 22814 17586 22882 17620
rect 22972 17586 23040 17620
rect 23130 17586 23198 17620
rect 23288 17586 23356 17620
rect 23446 17586 23514 17620
rect 23604 17586 23672 17620
rect 23762 17586 23830 17620
rect 23920 17586 23988 17620
rect 24078 17586 24146 17620
rect 24236 17586 24304 17620
rect 24394 17586 24462 17620
rect 24552 17586 24620 17620
rect 24710 17586 24778 17620
rect 24868 17586 24936 17620
rect 25026 17586 25094 17620
rect 20436 17482 25102 17484
rect 20436 17448 25102 17482
rect 1536 17446 6202 17448
rect 7836 17446 12502 17448
rect 14136 17446 18802 17448
rect 20436 17446 25102 17448
rect 1536 15568 6259 15570
rect 7836 15568 12559 15570
rect 14136 15568 18859 15570
rect 20436 15568 25159 15570
rect 1536 15534 6259 15568
rect 1536 15532 6259 15534
rect 1544 15396 1612 15430
rect 1702 15396 1770 15430
rect 1860 15396 1928 15430
rect 2018 15396 2086 15430
rect 2176 15396 2244 15430
rect 2334 15396 2402 15430
rect 2492 15396 2560 15430
rect 2650 15396 2718 15430
rect 2808 15396 2876 15430
rect 2966 15396 3034 15430
rect 3124 15396 3192 15430
rect 3282 15396 3350 15430
rect 3440 15396 3508 15430
rect 3598 15396 3666 15430
rect 3756 15396 3824 15430
rect 3914 15396 3982 15430
rect 4072 15396 4140 15430
rect 4230 15396 4298 15430
rect 4388 15396 4456 15430
rect 4546 15396 4614 15430
rect 4704 15396 4772 15430
rect 4862 15396 4930 15430
rect 5020 15396 5088 15430
rect 5178 15396 5246 15430
rect 5336 15396 5404 15430
rect 5494 15396 5562 15430
rect 5652 15396 5720 15430
rect 5810 15396 5878 15430
rect 5968 15396 6036 15430
rect 6126 15396 6194 15430
rect 7836 15534 12559 15568
rect 7836 15532 12559 15534
rect 7844 15396 7912 15430
rect 8002 15396 8070 15430
rect 8160 15396 8228 15430
rect 8318 15396 8386 15430
rect 8476 15396 8544 15430
rect 8634 15396 8702 15430
rect 8792 15396 8860 15430
rect 8950 15396 9018 15430
rect 9108 15396 9176 15430
rect 9266 15396 9334 15430
rect 9424 15396 9492 15430
rect 9582 15396 9650 15430
rect 9740 15396 9808 15430
rect 9898 15396 9966 15430
rect 10056 15396 10124 15430
rect 10214 15396 10282 15430
rect 10372 15396 10440 15430
rect 10530 15396 10598 15430
rect 10688 15396 10756 15430
rect 10846 15396 10914 15430
rect 11004 15396 11072 15430
rect 11162 15396 11230 15430
rect 11320 15396 11388 15430
rect 11478 15396 11546 15430
rect 11636 15396 11704 15430
rect 11794 15396 11862 15430
rect 11952 15396 12020 15430
rect 12110 15396 12178 15430
rect 12268 15396 12336 15430
rect 12426 15396 12494 15430
rect 14136 15534 18859 15568
rect 14136 15532 18859 15534
rect 14144 15396 14212 15430
rect 14302 15396 14370 15430
rect 14460 15396 14528 15430
rect 14618 15396 14686 15430
rect 14776 15396 14844 15430
rect 14934 15396 15002 15430
rect 15092 15396 15160 15430
rect 15250 15396 15318 15430
rect 15408 15396 15476 15430
rect 15566 15396 15634 15430
rect 15724 15396 15792 15430
rect 15882 15396 15950 15430
rect 16040 15396 16108 15430
rect 16198 15396 16266 15430
rect 16356 15396 16424 15430
rect 16514 15396 16582 15430
rect 16672 15396 16740 15430
rect 16830 15396 16898 15430
rect 16988 15396 17056 15430
rect 17146 15396 17214 15430
rect 17304 15396 17372 15430
rect 17462 15396 17530 15430
rect 17620 15396 17688 15430
rect 17778 15396 17846 15430
rect 17936 15396 18004 15430
rect 18094 15396 18162 15430
rect 18252 15396 18320 15430
rect 18410 15396 18478 15430
rect 18568 15396 18636 15430
rect 18726 15396 18794 15430
rect 20436 15534 25159 15568
rect 20436 15532 25159 15534
rect 20444 15396 20512 15430
rect 20602 15396 20670 15430
rect 20760 15396 20828 15430
rect 20918 15396 20986 15430
rect 21076 15396 21144 15430
rect 21234 15396 21302 15430
rect 21392 15396 21460 15430
rect 21550 15396 21618 15430
rect 21708 15396 21776 15430
rect 21866 15396 21934 15430
rect 22024 15396 22092 15430
rect 22182 15396 22250 15430
rect 22340 15396 22408 15430
rect 22498 15396 22566 15430
rect 22656 15396 22724 15430
rect 22814 15396 22882 15430
rect 22972 15396 23040 15430
rect 23130 15396 23198 15430
rect 23288 15396 23356 15430
rect 23446 15396 23514 15430
rect 23604 15396 23672 15430
rect 23762 15396 23830 15430
rect 23920 15396 23988 15430
rect 24078 15396 24146 15430
rect 24236 15396 24304 15430
rect 24394 15396 24462 15430
rect 24552 15396 24620 15430
rect 24710 15396 24778 15430
rect 24868 15396 24936 15430
rect 25026 15396 25094 15430
rect -4040 13884 -4000 13940
rect -4218 13435 -4180 13832
rect -4218 12684 -4180 13081
rect -4040 12632 -4034 13884
rect -4034 12632 -4000 13884
rect -4040 12560 -4000 12632
rect 1346 9336 1348 15380
rect 1348 9336 1382 15380
rect 1382 9336 1384 15380
rect 1482 9370 1516 15346
rect 1640 9370 1674 15346
rect 1798 9370 1832 15346
rect 1956 9370 1990 15346
rect 2114 9370 2148 15346
rect 2272 9370 2306 15346
rect 2430 9370 2464 15346
rect 2588 9370 2622 15346
rect 2746 9370 2780 15346
rect 2904 9370 2938 15346
rect 3062 9370 3096 15346
rect 3220 9370 3254 15346
rect 3378 9370 3412 15346
rect 3536 9370 3570 15346
rect 3694 9370 3728 15346
rect 3852 9370 3886 15346
rect 4010 9370 4044 15346
rect 4168 9370 4202 15346
rect 4326 9370 4360 15346
rect 4484 9370 4518 15346
rect 4642 9370 4676 15346
rect 4800 9370 4834 15346
rect 4958 9370 4992 15346
rect 5116 9370 5150 15346
rect 5274 9370 5308 15346
rect 5432 9370 5466 15346
rect 5590 9370 5624 15346
rect 5748 9370 5782 15346
rect 5906 9370 5940 15346
rect 6064 9370 6098 15346
rect 6222 9370 6256 15346
rect 6354 9336 6356 15380
rect 6356 9336 6390 15380
rect 6390 9336 6392 15380
rect 7646 9336 7648 15380
rect 7648 9336 7682 15380
rect 7682 9336 7684 15380
rect 7782 9370 7816 15346
rect 7940 9370 7974 15346
rect 8098 9370 8132 15346
rect 8256 9370 8290 15346
rect 8414 9370 8448 15346
rect 8572 9370 8606 15346
rect 8730 9370 8764 15346
rect 8888 9370 8922 15346
rect 9046 9370 9080 15346
rect 9204 9370 9238 15346
rect 9362 9370 9396 15346
rect 9520 9370 9554 15346
rect 9678 9370 9712 15346
rect 9836 9370 9870 15346
rect 9994 9370 10028 15346
rect 10152 9370 10186 15346
rect 10310 9370 10344 15346
rect 10468 9370 10502 15346
rect 10626 9370 10660 15346
rect 10784 9370 10818 15346
rect 10942 9370 10976 15346
rect 11100 9370 11134 15346
rect 11258 9370 11292 15346
rect 11416 9370 11450 15346
rect 11574 9370 11608 15346
rect 11732 9370 11766 15346
rect 11890 9370 11924 15346
rect 12048 9370 12082 15346
rect 12206 9370 12240 15346
rect 12364 9370 12398 15346
rect 12522 9370 12556 15346
rect 12654 9336 12656 15380
rect 12656 9336 12690 15380
rect 12690 9336 12692 15380
rect 13946 9336 13948 15380
rect 13948 9336 13982 15380
rect 13982 9336 13984 15380
rect 14082 9370 14116 15346
rect 14240 9370 14274 15346
rect 14398 9370 14432 15346
rect 14556 9370 14590 15346
rect 14714 9370 14748 15346
rect 14872 9370 14906 15346
rect 15030 9370 15064 15346
rect 15188 9370 15222 15346
rect 15346 9370 15380 15346
rect 15504 9370 15538 15346
rect 15662 9370 15696 15346
rect 15820 9370 15854 15346
rect 15978 9370 16012 15346
rect 16136 9370 16170 15346
rect 16294 9370 16328 15346
rect 16452 9370 16486 15346
rect 16610 9370 16644 15346
rect 16768 9370 16802 15346
rect 16926 9370 16960 15346
rect 17084 9370 17118 15346
rect 17242 9370 17276 15346
rect 17400 9370 17434 15346
rect 17558 9370 17592 15346
rect 17716 9370 17750 15346
rect 17874 9370 17908 15346
rect 18032 9370 18066 15346
rect 18190 9370 18224 15346
rect 18348 9370 18382 15346
rect 18506 9370 18540 15346
rect 18664 9370 18698 15346
rect 18822 9370 18856 15346
rect 18954 9336 18956 15380
rect 18956 9336 18990 15380
rect 18990 9336 18992 15380
rect 20246 9336 20248 15380
rect 20248 9336 20282 15380
rect 20282 9336 20284 15380
rect 20382 9370 20416 15346
rect 20540 9370 20574 15346
rect 20698 9370 20732 15346
rect 20856 9370 20890 15346
rect 21014 9370 21048 15346
rect 21172 9370 21206 15346
rect 21330 9370 21364 15346
rect 21488 9370 21522 15346
rect 21646 9370 21680 15346
rect 21804 9370 21838 15346
rect 21962 9370 21996 15346
rect 22120 9370 22154 15346
rect 22278 9370 22312 15346
rect 22436 9370 22470 15346
rect 22594 9370 22628 15346
rect 22752 9370 22786 15346
rect 22910 9370 22944 15346
rect 23068 9370 23102 15346
rect 23226 9370 23260 15346
rect 23384 9370 23418 15346
rect 23542 9370 23576 15346
rect 23700 9370 23734 15346
rect 23858 9370 23892 15346
rect 24016 9370 24050 15346
rect 24174 9370 24208 15346
rect 24332 9370 24366 15346
rect 24490 9370 24524 15346
rect 24648 9370 24682 15346
rect 24806 9370 24840 15346
rect 24964 9370 24998 15346
rect 25122 9370 25156 15346
rect 25254 9336 25256 15380
rect 25256 9336 25290 15380
rect 25290 9336 25292 15380
rect 30800 13884 30840 13980
rect 30800 12632 30834 13884
rect 30834 12632 30840 13884
rect 30980 13435 31018 13832
rect 30980 12684 31018 13081
rect 30800 12520 30840 12632
rect 1544 9286 1612 9320
rect 1702 9286 1770 9320
rect 1860 9286 1928 9320
rect 2018 9286 2086 9320
rect 2176 9286 2244 9320
rect 2334 9286 2402 9320
rect 2492 9286 2560 9320
rect 2650 9286 2718 9320
rect 2808 9286 2876 9320
rect 2966 9286 3034 9320
rect 3124 9286 3192 9320
rect 3282 9286 3350 9320
rect 3440 9286 3508 9320
rect 3598 9286 3666 9320
rect 3756 9286 3824 9320
rect 3914 9286 3982 9320
rect 4072 9286 4140 9320
rect 4230 9286 4298 9320
rect 4388 9286 4456 9320
rect 4546 9286 4614 9320
rect 4704 9286 4772 9320
rect 4862 9286 4930 9320
rect 5020 9286 5088 9320
rect 5178 9286 5246 9320
rect 5336 9286 5404 9320
rect 5494 9286 5562 9320
rect 5652 9286 5720 9320
rect 5810 9286 5878 9320
rect 5968 9286 6036 9320
rect 6126 9286 6194 9320
rect 1536 9182 6202 9184
rect 1536 9148 6202 9182
rect 7844 9286 7912 9320
rect 8002 9286 8070 9320
rect 8160 9286 8228 9320
rect 8318 9286 8386 9320
rect 8476 9286 8544 9320
rect 8634 9286 8702 9320
rect 8792 9286 8860 9320
rect 8950 9286 9018 9320
rect 9108 9286 9176 9320
rect 9266 9286 9334 9320
rect 9424 9286 9492 9320
rect 9582 9286 9650 9320
rect 9740 9286 9808 9320
rect 9898 9286 9966 9320
rect 10056 9286 10124 9320
rect 10214 9286 10282 9320
rect 10372 9286 10440 9320
rect 10530 9286 10598 9320
rect 10688 9286 10756 9320
rect 10846 9286 10914 9320
rect 11004 9286 11072 9320
rect 11162 9286 11230 9320
rect 11320 9286 11388 9320
rect 11478 9286 11546 9320
rect 11636 9286 11704 9320
rect 11794 9286 11862 9320
rect 11952 9286 12020 9320
rect 12110 9286 12178 9320
rect 12268 9286 12336 9320
rect 12426 9286 12494 9320
rect 7836 9182 12502 9184
rect 7836 9148 12502 9182
rect 14144 9286 14212 9320
rect 14302 9286 14370 9320
rect 14460 9286 14528 9320
rect 14618 9286 14686 9320
rect 14776 9286 14844 9320
rect 14934 9286 15002 9320
rect 15092 9286 15160 9320
rect 15250 9286 15318 9320
rect 15408 9286 15476 9320
rect 15566 9286 15634 9320
rect 15724 9286 15792 9320
rect 15882 9286 15950 9320
rect 16040 9286 16108 9320
rect 16198 9286 16266 9320
rect 16356 9286 16424 9320
rect 16514 9286 16582 9320
rect 16672 9286 16740 9320
rect 16830 9286 16898 9320
rect 16988 9286 17056 9320
rect 17146 9286 17214 9320
rect 17304 9286 17372 9320
rect 17462 9286 17530 9320
rect 17620 9286 17688 9320
rect 17778 9286 17846 9320
rect 17936 9286 18004 9320
rect 18094 9286 18162 9320
rect 18252 9286 18320 9320
rect 18410 9286 18478 9320
rect 18568 9286 18636 9320
rect 18726 9286 18794 9320
rect 14136 9182 18802 9184
rect 14136 9148 18802 9182
rect 20444 9286 20512 9320
rect 20602 9286 20670 9320
rect 20760 9286 20828 9320
rect 20918 9286 20986 9320
rect 21076 9286 21144 9320
rect 21234 9286 21302 9320
rect 21392 9286 21460 9320
rect 21550 9286 21618 9320
rect 21708 9286 21776 9320
rect 21866 9286 21934 9320
rect 22024 9286 22092 9320
rect 22182 9286 22250 9320
rect 22340 9286 22408 9320
rect 22498 9286 22566 9320
rect 22656 9286 22724 9320
rect 22814 9286 22882 9320
rect 22972 9286 23040 9320
rect 23130 9286 23198 9320
rect 23288 9286 23356 9320
rect 23446 9286 23514 9320
rect 23604 9286 23672 9320
rect 23762 9286 23830 9320
rect 23920 9286 23988 9320
rect 24078 9286 24146 9320
rect 24236 9286 24304 9320
rect 24394 9286 24462 9320
rect 24552 9286 24620 9320
rect 24710 9286 24778 9320
rect 24868 9286 24936 9320
rect 25026 9286 25094 9320
rect 20436 9182 25102 9184
rect 20436 9148 25102 9182
rect 1536 9146 6202 9148
rect 7836 9146 12502 9148
rect 14136 9146 18802 9148
rect 20436 9146 25102 9148
rect 1536 8568 6259 8570
rect 7836 8568 12559 8570
rect 14136 8568 18859 8570
rect 20436 8568 25159 8570
rect 1536 8534 6259 8568
rect 1536 8532 6259 8534
rect 1544 8396 1612 8430
rect 1702 8396 1770 8430
rect 1860 8396 1928 8430
rect 2018 8396 2086 8430
rect 2176 8396 2244 8430
rect 2334 8396 2402 8430
rect 2492 8396 2560 8430
rect 2650 8396 2718 8430
rect 2808 8396 2876 8430
rect 2966 8396 3034 8430
rect 3124 8396 3192 8430
rect 3282 8396 3350 8430
rect 3440 8396 3508 8430
rect 3598 8396 3666 8430
rect 3756 8396 3824 8430
rect 3914 8396 3982 8430
rect 4072 8396 4140 8430
rect 4230 8396 4298 8430
rect 4388 8396 4456 8430
rect 4546 8396 4614 8430
rect 4704 8396 4772 8430
rect 4862 8396 4930 8430
rect 5020 8396 5088 8430
rect 5178 8396 5246 8430
rect 5336 8396 5404 8430
rect 5494 8396 5562 8430
rect 5652 8396 5720 8430
rect 5810 8396 5878 8430
rect 5968 8396 6036 8430
rect 6126 8396 6194 8430
rect 7836 8534 12559 8568
rect 7836 8532 12559 8534
rect 7844 8396 7912 8430
rect 8002 8396 8070 8430
rect 8160 8396 8228 8430
rect 8318 8396 8386 8430
rect 8476 8396 8544 8430
rect 8634 8396 8702 8430
rect 8792 8396 8860 8430
rect 8950 8396 9018 8430
rect 9108 8396 9176 8430
rect 9266 8396 9334 8430
rect 9424 8396 9492 8430
rect 9582 8396 9650 8430
rect 9740 8396 9808 8430
rect 9898 8396 9966 8430
rect 10056 8396 10124 8430
rect 10214 8396 10282 8430
rect 10372 8396 10440 8430
rect 10530 8396 10598 8430
rect 10688 8396 10756 8430
rect 10846 8396 10914 8430
rect 11004 8396 11072 8430
rect 11162 8396 11230 8430
rect 11320 8396 11388 8430
rect 11478 8396 11546 8430
rect 11636 8396 11704 8430
rect 11794 8396 11862 8430
rect 11952 8396 12020 8430
rect 12110 8396 12178 8430
rect 12268 8396 12336 8430
rect 12426 8396 12494 8430
rect 14136 8534 18859 8568
rect 14136 8532 18859 8534
rect 14144 8396 14212 8430
rect 14302 8396 14370 8430
rect 14460 8396 14528 8430
rect 14618 8396 14686 8430
rect 14776 8396 14844 8430
rect 14934 8396 15002 8430
rect 15092 8396 15160 8430
rect 15250 8396 15318 8430
rect 15408 8396 15476 8430
rect 15566 8396 15634 8430
rect 15724 8396 15792 8430
rect 15882 8396 15950 8430
rect 16040 8396 16108 8430
rect 16198 8396 16266 8430
rect 16356 8396 16424 8430
rect 16514 8396 16582 8430
rect 16672 8396 16740 8430
rect 16830 8396 16898 8430
rect 16988 8396 17056 8430
rect 17146 8396 17214 8430
rect 17304 8396 17372 8430
rect 17462 8396 17530 8430
rect 17620 8396 17688 8430
rect 17778 8396 17846 8430
rect 17936 8396 18004 8430
rect 18094 8396 18162 8430
rect 18252 8396 18320 8430
rect 18410 8396 18478 8430
rect 18568 8396 18636 8430
rect 18726 8396 18794 8430
rect 20436 8534 25159 8568
rect 20436 8532 25159 8534
rect 20444 8396 20512 8430
rect 20602 8396 20670 8430
rect 20760 8396 20828 8430
rect 20918 8396 20986 8430
rect 21076 8396 21144 8430
rect 21234 8396 21302 8430
rect 21392 8396 21460 8430
rect 21550 8396 21618 8430
rect 21708 8396 21776 8430
rect 21866 8396 21934 8430
rect 22024 8396 22092 8430
rect 22182 8396 22250 8430
rect 22340 8396 22408 8430
rect 22498 8396 22566 8430
rect 22656 8396 22724 8430
rect 22814 8396 22882 8430
rect 22972 8396 23040 8430
rect 23130 8396 23198 8430
rect 23288 8396 23356 8430
rect 23446 8396 23514 8430
rect 23604 8396 23672 8430
rect 23762 8396 23830 8430
rect 23920 8396 23988 8430
rect 24078 8396 24146 8430
rect 24236 8396 24304 8430
rect 24394 8396 24462 8430
rect 24552 8396 24620 8430
rect 24710 8396 24778 8430
rect 24868 8396 24936 8430
rect 25026 8396 25094 8430
rect 1346 2336 1348 8380
rect 1348 2336 1382 8380
rect 1382 2336 1384 8380
rect 1482 2370 1516 8346
rect 1640 2370 1674 8346
rect 1798 2370 1832 8346
rect 1956 2370 1990 8346
rect 2114 2370 2148 8346
rect 2272 2370 2306 8346
rect 2430 2370 2464 8346
rect 2588 2370 2622 8346
rect 2746 2370 2780 8346
rect 2904 2370 2938 8346
rect 3062 2370 3096 8346
rect 3220 2370 3254 8346
rect 3378 2370 3412 8346
rect 3536 2370 3570 8346
rect 3694 2370 3728 8346
rect 3852 2370 3886 8346
rect 4010 2370 4044 8346
rect 4168 2370 4202 8346
rect 4326 2370 4360 8346
rect 4484 2370 4518 8346
rect 4642 2370 4676 8346
rect 4800 2370 4834 8346
rect 4958 2370 4992 8346
rect 5116 2370 5150 8346
rect 5274 2370 5308 8346
rect 5432 2370 5466 8346
rect 5590 2370 5624 8346
rect 5748 2370 5782 8346
rect 5906 2370 5940 8346
rect 6064 2370 6098 8346
rect 6222 2370 6256 8346
rect 6354 2336 6356 8380
rect 6356 2336 6390 8380
rect 6390 2336 6392 8380
rect 7646 2336 7648 8380
rect 7648 2336 7682 8380
rect 7682 2336 7684 8380
rect 7782 2370 7816 8346
rect 7940 2370 7974 8346
rect 8098 2370 8132 8346
rect 8256 2370 8290 8346
rect 8414 2370 8448 8346
rect 8572 2370 8606 8346
rect 8730 2370 8764 8346
rect 8888 2370 8922 8346
rect 9046 2370 9080 8346
rect 9204 2370 9238 8346
rect 9362 2370 9396 8346
rect 9520 2370 9554 8346
rect 9678 2370 9712 8346
rect 9836 2370 9870 8346
rect 9994 2370 10028 8346
rect 10152 2370 10186 8346
rect 10310 2370 10344 8346
rect 10468 2370 10502 8346
rect 10626 2370 10660 8346
rect 10784 2370 10818 8346
rect 10942 2370 10976 8346
rect 11100 2370 11134 8346
rect 11258 2370 11292 8346
rect 11416 2370 11450 8346
rect 11574 2370 11608 8346
rect 11732 2370 11766 8346
rect 11890 2370 11924 8346
rect 12048 2370 12082 8346
rect 12206 2370 12240 8346
rect 12364 2370 12398 8346
rect 12522 2370 12556 8346
rect 12654 2336 12656 8380
rect 12656 2336 12690 8380
rect 12690 2336 12692 8380
rect 13946 2336 13948 8380
rect 13948 2336 13982 8380
rect 13982 2336 13984 8380
rect 14082 2370 14116 8346
rect 14240 2370 14274 8346
rect 14398 2370 14432 8346
rect 14556 2370 14590 8346
rect 14714 2370 14748 8346
rect 14872 2370 14906 8346
rect 15030 2370 15064 8346
rect 15188 2370 15222 8346
rect 15346 2370 15380 8346
rect 15504 2370 15538 8346
rect 15662 2370 15696 8346
rect 15820 2370 15854 8346
rect 15978 2370 16012 8346
rect 16136 2370 16170 8346
rect 16294 2370 16328 8346
rect 16452 2370 16486 8346
rect 16610 2370 16644 8346
rect 16768 2370 16802 8346
rect 16926 2370 16960 8346
rect 17084 2370 17118 8346
rect 17242 2370 17276 8346
rect 17400 2370 17434 8346
rect 17558 2370 17592 8346
rect 17716 2370 17750 8346
rect 17874 2370 17908 8346
rect 18032 2370 18066 8346
rect 18190 2370 18224 8346
rect 18348 2370 18382 8346
rect 18506 2370 18540 8346
rect 18664 2370 18698 8346
rect 18822 2370 18856 8346
rect 18954 2336 18956 8380
rect 18956 2336 18990 8380
rect 18990 2336 18992 8380
rect 20246 2336 20248 8380
rect 20248 2336 20282 8380
rect 20282 2336 20284 8380
rect 20382 2370 20416 8346
rect 20540 2370 20574 8346
rect 20698 2370 20732 8346
rect 20856 2370 20890 8346
rect 21014 2370 21048 8346
rect 21172 2370 21206 8346
rect 21330 2370 21364 8346
rect 21488 2370 21522 8346
rect 21646 2370 21680 8346
rect 21804 2370 21838 8346
rect 21962 2370 21996 8346
rect 22120 2370 22154 8346
rect 22278 2370 22312 8346
rect 22436 2370 22470 8346
rect 22594 2370 22628 8346
rect 22752 2370 22786 8346
rect 22910 2370 22944 8346
rect 23068 2370 23102 8346
rect 23226 2370 23260 8346
rect 23384 2370 23418 8346
rect 23542 2370 23576 8346
rect 23700 2370 23734 8346
rect 23858 2370 23892 8346
rect 24016 2370 24050 8346
rect 24174 2370 24208 8346
rect 24332 2370 24366 8346
rect 24490 2370 24524 8346
rect 24648 2370 24682 8346
rect 24806 2370 24840 8346
rect 24964 2370 24998 8346
rect 25122 2370 25156 8346
rect 25254 2336 25256 8380
rect 25256 2336 25290 8380
rect 25290 2336 25292 8380
rect 1544 2286 1612 2320
rect 1702 2286 1770 2320
rect 1860 2286 1928 2320
rect 2018 2286 2086 2320
rect 2176 2286 2244 2320
rect 2334 2286 2402 2320
rect 2492 2286 2560 2320
rect 2650 2286 2718 2320
rect 2808 2286 2876 2320
rect 2966 2286 3034 2320
rect 3124 2286 3192 2320
rect 3282 2286 3350 2320
rect 3440 2286 3508 2320
rect 3598 2286 3666 2320
rect 3756 2286 3824 2320
rect 3914 2286 3982 2320
rect 4072 2286 4140 2320
rect 4230 2286 4298 2320
rect 4388 2286 4456 2320
rect 4546 2286 4614 2320
rect 4704 2286 4772 2320
rect 4862 2286 4930 2320
rect 5020 2286 5088 2320
rect 5178 2286 5246 2320
rect 5336 2286 5404 2320
rect 5494 2286 5562 2320
rect 5652 2286 5720 2320
rect 5810 2286 5878 2320
rect 5968 2286 6036 2320
rect 6126 2286 6194 2320
rect 1536 2182 6202 2184
rect 1536 2148 6202 2182
rect 7844 2286 7912 2320
rect 8002 2286 8070 2320
rect 8160 2286 8228 2320
rect 8318 2286 8386 2320
rect 8476 2286 8544 2320
rect 8634 2286 8702 2320
rect 8792 2286 8860 2320
rect 8950 2286 9018 2320
rect 9108 2286 9176 2320
rect 9266 2286 9334 2320
rect 9424 2286 9492 2320
rect 9582 2286 9650 2320
rect 9740 2286 9808 2320
rect 9898 2286 9966 2320
rect 10056 2286 10124 2320
rect 10214 2286 10282 2320
rect 10372 2286 10440 2320
rect 10530 2286 10598 2320
rect 10688 2286 10756 2320
rect 10846 2286 10914 2320
rect 11004 2286 11072 2320
rect 11162 2286 11230 2320
rect 11320 2286 11388 2320
rect 11478 2286 11546 2320
rect 11636 2286 11704 2320
rect 11794 2286 11862 2320
rect 11952 2286 12020 2320
rect 12110 2286 12178 2320
rect 12268 2286 12336 2320
rect 12426 2286 12494 2320
rect 7836 2182 12502 2184
rect 7836 2148 12502 2182
rect 14144 2286 14212 2320
rect 14302 2286 14370 2320
rect 14460 2286 14528 2320
rect 14618 2286 14686 2320
rect 14776 2286 14844 2320
rect 14934 2286 15002 2320
rect 15092 2286 15160 2320
rect 15250 2286 15318 2320
rect 15408 2286 15476 2320
rect 15566 2286 15634 2320
rect 15724 2286 15792 2320
rect 15882 2286 15950 2320
rect 16040 2286 16108 2320
rect 16198 2286 16266 2320
rect 16356 2286 16424 2320
rect 16514 2286 16582 2320
rect 16672 2286 16740 2320
rect 16830 2286 16898 2320
rect 16988 2286 17056 2320
rect 17146 2286 17214 2320
rect 17304 2286 17372 2320
rect 17462 2286 17530 2320
rect 17620 2286 17688 2320
rect 17778 2286 17846 2320
rect 17936 2286 18004 2320
rect 18094 2286 18162 2320
rect 18252 2286 18320 2320
rect 18410 2286 18478 2320
rect 18568 2286 18636 2320
rect 18726 2286 18794 2320
rect 14136 2182 18802 2184
rect 14136 2148 18802 2182
rect 20444 2286 20512 2320
rect 20602 2286 20670 2320
rect 20760 2286 20828 2320
rect 20918 2286 20986 2320
rect 21076 2286 21144 2320
rect 21234 2286 21302 2320
rect 21392 2286 21460 2320
rect 21550 2286 21618 2320
rect 21708 2286 21776 2320
rect 21866 2286 21934 2320
rect 22024 2286 22092 2320
rect 22182 2286 22250 2320
rect 22340 2286 22408 2320
rect 22498 2286 22566 2320
rect 22656 2286 22724 2320
rect 22814 2286 22882 2320
rect 22972 2286 23040 2320
rect 23130 2286 23198 2320
rect 23288 2286 23356 2320
rect 23446 2286 23514 2320
rect 23604 2286 23672 2320
rect 23762 2286 23830 2320
rect 23920 2286 23988 2320
rect 24078 2286 24146 2320
rect 24236 2286 24304 2320
rect 24394 2286 24462 2320
rect 24552 2286 24620 2320
rect 24710 2286 24778 2320
rect 24868 2286 24936 2320
rect 25026 2286 25094 2320
rect 20436 2182 25102 2184
rect 20436 2148 25102 2182
rect 1536 2146 6202 2148
rect 7836 2146 12502 2148
rect 14136 2146 18802 2148
rect 20436 2146 25102 2148
<< metal1 >>
rect 0 47480 26500 47500
rect 0 47410 150 47480
rect 350 47410 650 47480
rect 850 47410 1150 47480
rect 1350 47410 1650 47480
rect 1850 47410 2150 47480
rect 2350 47410 2650 47480
rect 2850 47410 3150 47480
rect 3350 47410 3650 47480
rect 3850 47410 4150 47480
rect 4350 47410 4650 47480
rect 4850 47410 5150 47480
rect 5350 47410 5650 47480
rect 5850 47410 6150 47480
rect 6350 47410 6650 47480
rect 6850 47410 7150 47480
rect 7350 47410 7650 47480
rect 7850 47410 8150 47480
rect 8350 47410 8650 47480
rect 8850 47410 9150 47480
rect 9350 47410 9650 47480
rect 9850 47410 10150 47480
rect 10350 47410 10650 47480
rect 10850 47410 11150 47480
rect 11350 47410 11650 47480
rect 11850 47410 12150 47480
rect 12350 47410 12650 47480
rect 12850 47410 13150 47480
rect 13350 47410 13650 47480
rect 13850 47410 14150 47480
rect 14350 47410 14650 47480
rect 14850 47410 15150 47480
rect 15350 47410 15650 47480
rect 15850 47410 16150 47480
rect 16350 47410 16650 47480
rect 16850 47410 17150 47480
rect 17350 47410 17650 47480
rect 17850 47410 18150 47480
rect 18350 47410 18650 47480
rect 18850 47410 19150 47480
rect 19350 47410 19650 47480
rect 19850 47410 20150 47480
rect 20350 47410 20650 47480
rect 20850 47410 21150 47480
rect 21350 47410 21650 47480
rect 21850 47410 22150 47480
rect 22350 47410 22650 47480
rect 22850 47410 23150 47480
rect 23350 47410 23650 47480
rect 23850 47410 24150 47480
rect 24350 47410 24650 47480
rect 24850 47410 25150 47480
rect 25350 47410 25650 47480
rect 25850 47410 26150 47480
rect 26350 47410 26500 47480
rect 0 47400 26500 47410
rect 0 47380 120 47400
rect 380 47380 620 47400
rect 880 47380 1120 47400
rect 1380 47380 1620 47400
rect 1880 47380 2120 47400
rect 2380 47380 2620 47400
rect 2880 47380 3120 47400
rect 3380 47380 3620 47400
rect 3880 47380 4120 47400
rect 4380 47380 4620 47400
rect 4880 47380 5120 47400
rect 5380 47380 5620 47400
rect 5880 47380 6120 47400
rect 6380 47380 6620 47400
rect 6880 47380 7120 47400
rect 7380 47380 7620 47400
rect 7880 47380 8120 47400
rect 8380 47380 8620 47400
rect 8880 47380 9120 47400
rect 9380 47380 9620 47400
rect 9880 47380 10120 47400
rect 10380 47380 10620 47400
rect 10880 47380 11120 47400
rect 11380 47380 11620 47400
rect 11880 47380 12120 47400
rect 12380 47380 12620 47400
rect 12880 47380 13120 47400
rect 13380 47380 13620 47400
rect 13880 47380 14120 47400
rect 14380 47380 14620 47400
rect 14880 47380 15120 47400
rect 15380 47380 15620 47400
rect 15880 47380 16120 47400
rect 16380 47380 16620 47400
rect 16880 47380 17120 47400
rect 17380 47380 17620 47400
rect 17880 47380 18120 47400
rect 18380 47380 18620 47400
rect 18880 47380 19120 47400
rect 19380 47380 19620 47400
rect 19880 47380 20120 47400
rect 20380 47380 20620 47400
rect 20880 47380 21120 47400
rect 21380 47380 21620 47400
rect 21880 47380 22120 47400
rect 22380 47380 22620 47400
rect 22880 47380 23120 47400
rect 23380 47380 23620 47400
rect 23880 47380 24120 47400
rect 24380 47380 24620 47400
rect 24880 47380 25120 47400
rect 25380 47380 25620 47400
rect 25880 47380 26120 47400
rect 26380 47380 26500 47400
rect 0 47350 100 47380
rect 0 47150 20 47350
rect 90 47150 100 47350
rect 0 47120 100 47150
rect 400 47350 600 47380
rect 400 47150 410 47350
rect 480 47150 520 47350
rect 590 47150 600 47350
rect 400 47120 600 47150
rect 900 47350 1100 47380
rect 900 47150 910 47350
rect 980 47150 1020 47350
rect 1090 47150 1100 47350
rect 900 47120 1100 47150
rect 1400 47350 1600 47380
rect 1400 47150 1410 47350
rect 1480 47150 1520 47350
rect 1590 47150 1600 47350
rect 1400 47120 1600 47150
rect 1900 47350 2100 47380
rect 1900 47150 1910 47350
rect 1980 47150 2020 47350
rect 2090 47150 2100 47350
rect 1900 47120 2100 47150
rect 2400 47350 2600 47380
rect 2400 47150 2410 47350
rect 2480 47150 2520 47350
rect 2590 47150 2600 47350
rect 2400 47120 2600 47150
rect 2900 47350 3100 47380
rect 2900 47150 2910 47350
rect 2980 47150 3020 47350
rect 3090 47150 3100 47350
rect 2900 47120 3100 47150
rect 3400 47350 3600 47380
rect 3400 47150 3410 47350
rect 3480 47150 3520 47350
rect 3590 47150 3600 47350
rect 3400 47120 3600 47150
rect 3900 47350 4100 47380
rect 3900 47150 3910 47350
rect 3980 47150 4020 47350
rect 4090 47150 4100 47350
rect 3900 47120 4100 47150
rect 4400 47350 4600 47380
rect 4400 47150 4410 47350
rect 4480 47150 4520 47350
rect 4590 47150 4600 47350
rect 4400 47120 4600 47150
rect 4900 47350 5100 47380
rect 4900 47150 4910 47350
rect 4980 47150 5020 47350
rect 5090 47150 5100 47350
rect 4900 47120 5100 47150
rect 5400 47350 5600 47380
rect 5400 47150 5410 47350
rect 5480 47150 5520 47350
rect 5590 47150 5600 47350
rect 5400 47120 5600 47150
rect 5900 47350 6100 47380
rect 5900 47150 5910 47350
rect 5980 47150 6020 47350
rect 6090 47150 6100 47350
rect 5900 47120 6100 47150
rect 6400 47350 6600 47380
rect 6400 47150 6410 47350
rect 6480 47150 6520 47350
rect 6590 47150 6600 47350
rect 6400 47120 6600 47150
rect 6900 47350 7100 47380
rect 6900 47150 6910 47350
rect 6980 47150 7020 47350
rect 7090 47150 7100 47350
rect 6900 47120 7100 47150
rect 7400 47350 7600 47380
rect 7400 47150 7410 47350
rect 7480 47150 7520 47350
rect 7590 47150 7600 47350
rect 7400 47120 7600 47150
rect 7900 47350 8100 47380
rect 7900 47150 7910 47350
rect 7980 47150 8020 47350
rect 8090 47150 8100 47350
rect 7900 47120 8100 47150
rect 8400 47350 8600 47380
rect 8400 47150 8410 47350
rect 8480 47150 8520 47350
rect 8590 47150 8600 47350
rect 8400 47120 8600 47150
rect 8900 47350 9100 47380
rect 8900 47150 8910 47350
rect 8980 47150 9020 47350
rect 9090 47150 9100 47350
rect 8900 47120 9100 47150
rect 9400 47350 9600 47380
rect 9400 47150 9410 47350
rect 9480 47150 9520 47350
rect 9590 47150 9600 47350
rect 9400 47120 9600 47150
rect 9900 47350 10100 47380
rect 9900 47150 9910 47350
rect 9980 47150 10020 47350
rect 10090 47150 10100 47350
rect 9900 47120 10100 47150
rect 10400 47350 10600 47380
rect 10400 47150 10410 47350
rect 10480 47150 10520 47350
rect 10590 47150 10600 47350
rect 10400 47120 10600 47150
rect 10900 47350 11100 47380
rect 10900 47150 10910 47350
rect 10980 47150 11020 47350
rect 11090 47150 11100 47350
rect 10900 47120 11100 47150
rect 11400 47350 11600 47380
rect 11400 47150 11410 47350
rect 11480 47150 11520 47350
rect 11590 47150 11600 47350
rect 11400 47120 11600 47150
rect 11900 47350 12100 47380
rect 11900 47150 11910 47350
rect 11980 47150 12020 47350
rect 12090 47150 12100 47350
rect 11900 47120 12100 47150
rect 12400 47350 12600 47380
rect 12400 47150 12410 47350
rect 12480 47150 12520 47350
rect 12590 47150 12600 47350
rect 12400 47120 12600 47150
rect 12900 47350 13100 47380
rect 12900 47150 12910 47350
rect 12980 47150 13020 47350
rect 13090 47150 13100 47350
rect 12900 47120 13100 47150
rect 13400 47350 13600 47380
rect 13400 47150 13410 47350
rect 13480 47150 13520 47350
rect 13590 47150 13600 47350
rect 13400 47120 13600 47150
rect 13900 47350 14100 47380
rect 13900 47150 13910 47350
rect 13980 47150 14020 47350
rect 14090 47150 14100 47350
rect 13900 47120 14100 47150
rect 14400 47350 14600 47380
rect 14400 47150 14410 47350
rect 14480 47150 14520 47350
rect 14590 47150 14600 47350
rect 14400 47120 14600 47150
rect 14900 47350 15100 47380
rect 14900 47150 14910 47350
rect 14980 47150 15020 47350
rect 15090 47150 15100 47350
rect 14900 47120 15100 47150
rect 15400 47350 15600 47380
rect 15400 47150 15410 47350
rect 15480 47150 15520 47350
rect 15590 47150 15600 47350
rect 15400 47120 15600 47150
rect 15900 47350 16100 47380
rect 15900 47150 15910 47350
rect 15980 47150 16020 47350
rect 16090 47150 16100 47350
rect 15900 47120 16100 47150
rect 16400 47350 16600 47380
rect 16400 47150 16410 47350
rect 16480 47150 16520 47350
rect 16590 47150 16600 47350
rect 16400 47120 16600 47150
rect 16900 47350 17100 47380
rect 16900 47150 16910 47350
rect 16980 47150 17020 47350
rect 17090 47150 17100 47350
rect 16900 47120 17100 47150
rect 17400 47350 17600 47380
rect 17400 47150 17410 47350
rect 17480 47150 17520 47350
rect 17590 47150 17600 47350
rect 17400 47120 17600 47150
rect 17900 47350 18100 47380
rect 17900 47150 17910 47350
rect 17980 47150 18020 47350
rect 18090 47150 18100 47350
rect 17900 47120 18100 47150
rect 18400 47350 18600 47380
rect 18400 47150 18410 47350
rect 18480 47150 18520 47350
rect 18590 47150 18600 47350
rect 18400 47120 18600 47150
rect 18900 47350 19100 47380
rect 18900 47150 18910 47350
rect 18980 47150 19020 47350
rect 19090 47150 19100 47350
rect 18900 47120 19100 47150
rect 19400 47350 19600 47380
rect 19400 47150 19410 47350
rect 19480 47150 19520 47350
rect 19590 47150 19600 47350
rect 19400 47120 19600 47150
rect 19900 47350 20100 47380
rect 19900 47150 19910 47350
rect 19980 47150 20020 47350
rect 20090 47150 20100 47350
rect 19900 47120 20100 47150
rect 20400 47350 20600 47380
rect 20400 47150 20410 47350
rect 20480 47150 20520 47350
rect 20590 47150 20600 47350
rect 20400 47120 20600 47150
rect 20900 47350 21100 47380
rect 20900 47150 20910 47350
rect 20980 47150 21020 47350
rect 21090 47150 21100 47350
rect 20900 47120 21100 47150
rect 21400 47350 21600 47380
rect 21400 47150 21410 47350
rect 21480 47150 21520 47350
rect 21590 47150 21600 47350
rect 21400 47120 21600 47150
rect 21900 47350 22100 47380
rect 21900 47150 21910 47350
rect 21980 47150 22020 47350
rect 22090 47150 22100 47350
rect 21900 47120 22100 47150
rect 22400 47350 22600 47380
rect 22400 47150 22410 47350
rect 22480 47150 22520 47350
rect 22590 47150 22600 47350
rect 22400 47120 22600 47150
rect 22900 47350 23100 47380
rect 22900 47150 22910 47350
rect 22980 47150 23020 47350
rect 23090 47150 23100 47350
rect 22900 47120 23100 47150
rect 23400 47350 23600 47380
rect 23400 47150 23410 47350
rect 23480 47150 23520 47350
rect 23590 47150 23600 47350
rect 23400 47120 23600 47150
rect 23900 47350 24100 47380
rect 23900 47150 23910 47350
rect 23980 47150 24020 47350
rect 24090 47150 24100 47350
rect 23900 47120 24100 47150
rect 24400 47350 24600 47380
rect 24400 47150 24410 47350
rect 24480 47150 24520 47350
rect 24590 47150 24600 47350
rect 24400 47120 24600 47150
rect 24900 47350 25100 47380
rect 24900 47150 24910 47350
rect 24980 47150 25020 47350
rect 25090 47150 25100 47350
rect 24900 47120 25100 47150
rect 25400 47350 25600 47380
rect 25400 47150 25410 47350
rect 25480 47150 25520 47350
rect 25590 47150 25600 47350
rect 25400 47120 25600 47150
rect 25900 47350 26100 47380
rect 25900 47150 25910 47350
rect 25980 47150 26020 47350
rect 26090 47150 26100 47350
rect 25900 47120 26100 47150
rect 26400 47350 26500 47380
rect 26400 47150 26410 47350
rect 26480 47150 26500 47350
rect 26400 47120 26500 47150
rect 0 47100 120 47120
rect 380 47100 620 47120
rect 880 47100 1120 47120
rect 1380 47100 1620 47120
rect 1880 47100 2120 47120
rect 2380 47100 2620 47120
rect 2880 47100 3120 47120
rect 3380 47100 3620 47120
rect 3880 47100 4120 47120
rect 4380 47100 4620 47120
rect 4880 47100 5120 47120
rect 5380 47100 5620 47120
rect 5880 47100 6120 47120
rect 6380 47100 6620 47120
rect 6880 47100 7120 47120
rect 7380 47100 7620 47120
rect 7880 47100 8120 47120
rect 8380 47100 8620 47120
rect 8880 47100 9120 47120
rect 9380 47100 9620 47120
rect 9880 47100 10120 47120
rect 10380 47100 10620 47120
rect 10880 47100 11120 47120
rect 11380 47100 11620 47120
rect 11880 47100 12120 47120
rect 12380 47100 12620 47120
rect 12880 47100 13120 47120
rect 13380 47100 13620 47120
rect 13880 47100 14120 47120
rect 14380 47100 14620 47120
rect 14880 47100 15120 47120
rect 15380 47100 15620 47120
rect 15880 47100 16120 47120
rect 16380 47100 16620 47120
rect 16880 47100 17120 47120
rect 17380 47100 17620 47120
rect 17880 47100 18120 47120
rect 18380 47100 18620 47120
rect 18880 47100 19120 47120
rect 19380 47100 19620 47120
rect 19880 47100 20120 47120
rect 20380 47100 20620 47120
rect 20880 47100 21120 47120
rect 21380 47100 21620 47120
rect 21880 47100 22120 47120
rect 22380 47100 22620 47120
rect 22880 47100 23120 47120
rect 23380 47100 23620 47120
rect 23880 47100 24120 47120
rect 24380 47100 24620 47120
rect 24880 47100 25120 47120
rect 25380 47100 25620 47120
rect 25880 47100 26120 47120
rect 26380 47100 26500 47120
rect 0 47090 26500 47100
rect 0 47020 150 47090
rect 350 47020 650 47090
rect 850 47020 1150 47090
rect 1350 47020 1650 47090
rect 1850 47020 2150 47090
rect 2350 47020 2650 47090
rect 2850 47020 3150 47090
rect 3350 47020 3650 47090
rect 3850 47020 4150 47090
rect 4350 47020 4650 47090
rect 4850 47020 5150 47090
rect 5350 47020 5650 47090
rect 5850 47020 6150 47090
rect 6350 47020 6650 47090
rect 6850 47020 7150 47090
rect 7350 47020 7650 47090
rect 7850 47020 8150 47090
rect 8350 47020 8650 47090
rect 8850 47020 9150 47090
rect 9350 47020 9650 47090
rect 9850 47020 10150 47090
rect 10350 47020 10650 47090
rect 10850 47020 11150 47090
rect 11350 47020 11650 47090
rect 11850 47020 12150 47090
rect 12350 47020 12650 47090
rect 12850 47020 13150 47090
rect 13350 47020 13650 47090
rect 13850 47020 14150 47090
rect 14350 47020 14650 47090
rect 14850 47020 15150 47090
rect 15350 47020 15650 47090
rect 15850 47020 16150 47090
rect 16350 47020 16650 47090
rect 16850 47020 17150 47090
rect 17350 47020 17650 47090
rect 17850 47020 18150 47090
rect 18350 47020 18650 47090
rect 18850 47020 19150 47090
rect 19350 47020 19650 47090
rect 19850 47020 20150 47090
rect 20350 47020 20650 47090
rect 20850 47020 21150 47090
rect 21350 47020 21650 47090
rect 21850 47020 22150 47090
rect 22350 47020 22650 47090
rect 22850 47020 23150 47090
rect 23350 47020 23650 47090
rect 23850 47020 24150 47090
rect 24350 47020 24650 47090
rect 24850 47020 25150 47090
rect 25350 47020 25650 47090
rect 25850 47020 26150 47090
rect 26350 47020 26500 47090
rect 0 46980 26500 47020
rect 0 46910 150 46980
rect 350 46910 650 46980
rect 850 46910 1150 46980
rect 1350 46910 1650 46980
rect 1850 46910 2150 46980
rect 2350 46910 2650 46980
rect 2850 46910 3150 46980
rect 3350 46910 3650 46980
rect 3850 46910 4150 46980
rect 4350 46910 4650 46980
rect 4850 46910 5150 46980
rect 5350 46910 5650 46980
rect 5850 46910 6150 46980
rect 6350 46910 6650 46980
rect 6850 46910 7150 46980
rect 7350 46910 7650 46980
rect 7850 46910 8150 46980
rect 8350 46910 8650 46980
rect 8850 46910 9150 46980
rect 9350 46910 9650 46980
rect 9850 46910 10150 46980
rect 10350 46910 10650 46980
rect 10850 46910 11150 46980
rect 11350 46910 11650 46980
rect 11850 46910 12150 46980
rect 12350 46910 12650 46980
rect 12850 46910 13150 46980
rect 13350 46910 13650 46980
rect 13850 46910 14150 46980
rect 14350 46910 14650 46980
rect 14850 46910 15150 46980
rect 15350 46910 15650 46980
rect 15850 46910 16150 46980
rect 16350 46910 16650 46980
rect 16850 46910 17150 46980
rect 17350 46910 17650 46980
rect 17850 46910 18150 46980
rect 18350 46910 18650 46980
rect 18850 46910 19150 46980
rect 19350 46910 19650 46980
rect 19850 46910 20150 46980
rect 20350 46910 20650 46980
rect 20850 46910 21150 46980
rect 21350 46910 21650 46980
rect 21850 46910 22150 46980
rect 22350 46910 22650 46980
rect 22850 46910 23150 46980
rect 23350 46910 23650 46980
rect 23850 46910 24150 46980
rect 24350 46910 24650 46980
rect 24850 46910 25150 46980
rect 25350 46910 25650 46980
rect 25850 46910 26150 46980
rect 26350 46910 26500 46980
rect 0 46900 26500 46910
rect 0 46880 120 46900
rect 380 46880 620 46900
rect 880 46880 1120 46900
rect 1380 46880 1620 46900
rect 1880 46880 2120 46900
rect 2380 46880 2620 46900
rect 2880 46880 3120 46900
rect 3380 46880 3620 46900
rect 3880 46880 4120 46900
rect 4380 46880 4620 46900
rect 4880 46880 5120 46900
rect 5380 46880 5620 46900
rect 5880 46880 6120 46900
rect 6380 46880 6620 46900
rect 6880 46880 7120 46900
rect 7380 46880 7620 46900
rect 7880 46880 8120 46900
rect 8380 46880 8620 46900
rect 8880 46880 9120 46900
rect 9380 46880 9620 46900
rect 9880 46880 10120 46900
rect 10380 46880 10620 46900
rect 10880 46880 11120 46900
rect 11380 46880 11620 46900
rect 11880 46880 12120 46900
rect 12380 46880 12620 46900
rect 12880 46880 13120 46900
rect 13380 46880 13620 46900
rect 13880 46880 14120 46900
rect 14380 46880 14620 46900
rect 14880 46880 15120 46900
rect 15380 46880 15620 46900
rect 15880 46880 16120 46900
rect 16380 46880 16620 46900
rect 16880 46880 17120 46900
rect 17380 46880 17620 46900
rect 17880 46880 18120 46900
rect 18380 46880 18620 46900
rect 18880 46880 19120 46900
rect 19380 46880 19620 46900
rect 19880 46880 20120 46900
rect 20380 46880 20620 46900
rect 20880 46880 21120 46900
rect 21380 46880 21620 46900
rect 21880 46880 22120 46900
rect 22380 46880 22620 46900
rect 22880 46880 23120 46900
rect 23380 46880 23620 46900
rect 23880 46880 24120 46900
rect 24380 46880 24620 46900
rect 24880 46880 25120 46900
rect 25380 46880 25620 46900
rect 25880 46880 26120 46900
rect 26380 46880 26500 46900
rect 0 46850 100 46880
rect 0 46650 20 46850
rect 90 46650 100 46850
rect 0 46620 100 46650
rect 400 46850 600 46880
rect 400 46650 410 46850
rect 480 46650 520 46850
rect 590 46650 600 46850
rect 400 46620 600 46650
rect 900 46850 1100 46880
rect 900 46650 910 46850
rect 980 46650 1020 46850
rect 1090 46650 1100 46850
rect 900 46620 1100 46650
rect 1400 46850 1600 46880
rect 1400 46650 1410 46850
rect 1480 46650 1520 46850
rect 1590 46650 1600 46850
rect 1400 46620 1600 46650
rect 1900 46850 2100 46880
rect 1900 46650 1910 46850
rect 1980 46650 2020 46850
rect 2090 46650 2100 46850
rect 1900 46620 2100 46650
rect 2400 46850 2600 46880
rect 2400 46650 2410 46850
rect 2480 46650 2520 46850
rect 2590 46650 2600 46850
rect 2400 46620 2600 46650
rect 2900 46850 3100 46880
rect 2900 46650 2910 46850
rect 2980 46650 3020 46850
rect 3090 46650 3100 46850
rect 2900 46620 3100 46650
rect 3400 46850 3600 46880
rect 3400 46650 3410 46850
rect 3480 46650 3520 46850
rect 3590 46650 3600 46850
rect 3400 46620 3600 46650
rect 3900 46850 4100 46880
rect 3900 46650 3910 46850
rect 3980 46650 4020 46850
rect 4090 46650 4100 46850
rect 3900 46620 4100 46650
rect 4400 46850 4600 46880
rect 4400 46650 4410 46850
rect 4480 46650 4520 46850
rect 4590 46650 4600 46850
rect 4400 46620 4600 46650
rect 4900 46850 5100 46880
rect 4900 46650 4910 46850
rect 4980 46650 5020 46850
rect 5090 46650 5100 46850
rect 4900 46620 5100 46650
rect 5400 46850 5600 46880
rect 5400 46650 5410 46850
rect 5480 46650 5520 46850
rect 5590 46650 5600 46850
rect 5400 46620 5600 46650
rect 5900 46850 6100 46880
rect 5900 46650 5910 46850
rect 5980 46650 6020 46850
rect 6090 46650 6100 46850
rect 5900 46620 6100 46650
rect 6400 46850 6600 46880
rect 6400 46650 6410 46850
rect 6480 46650 6520 46850
rect 6590 46650 6600 46850
rect 6400 46620 6600 46650
rect 6900 46850 7100 46880
rect 6900 46650 6910 46850
rect 6980 46650 7020 46850
rect 7090 46650 7100 46850
rect 6900 46620 7100 46650
rect 7400 46850 7600 46880
rect 7400 46650 7410 46850
rect 7480 46650 7520 46850
rect 7590 46650 7600 46850
rect 7400 46620 7600 46650
rect 7900 46850 8100 46880
rect 7900 46650 7910 46850
rect 7980 46650 8020 46850
rect 8090 46650 8100 46850
rect 7900 46620 8100 46650
rect 8400 46850 8600 46880
rect 8400 46650 8410 46850
rect 8480 46650 8520 46850
rect 8590 46650 8600 46850
rect 8400 46620 8600 46650
rect 8900 46850 9100 46880
rect 8900 46650 8910 46850
rect 8980 46650 9020 46850
rect 9090 46650 9100 46850
rect 8900 46620 9100 46650
rect 9400 46850 9600 46880
rect 9400 46650 9410 46850
rect 9480 46650 9520 46850
rect 9590 46650 9600 46850
rect 9400 46620 9600 46650
rect 9900 46850 10100 46880
rect 9900 46650 9910 46850
rect 9980 46650 10020 46850
rect 10090 46650 10100 46850
rect 9900 46620 10100 46650
rect 10400 46850 10600 46880
rect 10400 46650 10410 46850
rect 10480 46650 10520 46850
rect 10590 46650 10600 46850
rect 10400 46620 10600 46650
rect 10900 46850 11100 46880
rect 10900 46650 10910 46850
rect 10980 46650 11020 46850
rect 11090 46650 11100 46850
rect 10900 46620 11100 46650
rect 11400 46850 11600 46880
rect 11400 46650 11410 46850
rect 11480 46650 11520 46850
rect 11590 46650 11600 46850
rect 11400 46620 11600 46650
rect 11900 46850 12100 46880
rect 11900 46650 11910 46850
rect 11980 46650 12020 46850
rect 12090 46650 12100 46850
rect 11900 46620 12100 46650
rect 12400 46850 12600 46880
rect 12400 46650 12410 46850
rect 12480 46650 12520 46850
rect 12590 46650 12600 46850
rect 12400 46620 12600 46650
rect 12900 46850 13100 46880
rect 12900 46650 12910 46850
rect 12980 46650 13020 46850
rect 13090 46650 13100 46850
rect 12900 46620 13100 46650
rect 13400 46850 13600 46880
rect 13400 46650 13410 46850
rect 13480 46650 13520 46850
rect 13590 46650 13600 46850
rect 13400 46620 13600 46650
rect 13900 46850 14100 46880
rect 13900 46650 13910 46850
rect 13980 46650 14020 46850
rect 14090 46650 14100 46850
rect 13900 46620 14100 46650
rect 14400 46850 14600 46880
rect 14400 46650 14410 46850
rect 14480 46650 14520 46850
rect 14590 46650 14600 46850
rect 14400 46620 14600 46650
rect 14900 46850 15100 46880
rect 14900 46650 14910 46850
rect 14980 46650 15020 46850
rect 15090 46650 15100 46850
rect 14900 46620 15100 46650
rect 15400 46850 15600 46880
rect 15400 46650 15410 46850
rect 15480 46650 15520 46850
rect 15590 46650 15600 46850
rect 15400 46620 15600 46650
rect 15900 46850 16100 46880
rect 15900 46650 15910 46850
rect 15980 46650 16020 46850
rect 16090 46650 16100 46850
rect 15900 46620 16100 46650
rect 16400 46850 16600 46880
rect 16400 46650 16410 46850
rect 16480 46650 16520 46850
rect 16590 46650 16600 46850
rect 16400 46620 16600 46650
rect 16900 46850 17100 46880
rect 16900 46650 16910 46850
rect 16980 46650 17020 46850
rect 17090 46650 17100 46850
rect 16900 46620 17100 46650
rect 17400 46850 17600 46880
rect 17400 46650 17410 46850
rect 17480 46650 17520 46850
rect 17590 46650 17600 46850
rect 17400 46620 17600 46650
rect 17900 46850 18100 46880
rect 17900 46650 17910 46850
rect 17980 46650 18020 46850
rect 18090 46650 18100 46850
rect 17900 46620 18100 46650
rect 18400 46850 18600 46880
rect 18400 46650 18410 46850
rect 18480 46650 18520 46850
rect 18590 46650 18600 46850
rect 18400 46620 18600 46650
rect 18900 46850 19100 46880
rect 18900 46650 18910 46850
rect 18980 46650 19020 46850
rect 19090 46650 19100 46850
rect 18900 46620 19100 46650
rect 19400 46850 19600 46880
rect 19400 46650 19410 46850
rect 19480 46650 19520 46850
rect 19590 46650 19600 46850
rect 19400 46620 19600 46650
rect 19900 46850 20100 46880
rect 19900 46650 19910 46850
rect 19980 46650 20020 46850
rect 20090 46650 20100 46850
rect 19900 46620 20100 46650
rect 20400 46850 20600 46880
rect 20400 46650 20410 46850
rect 20480 46650 20520 46850
rect 20590 46650 20600 46850
rect 20400 46620 20600 46650
rect 20900 46850 21100 46880
rect 20900 46650 20910 46850
rect 20980 46650 21020 46850
rect 21090 46650 21100 46850
rect 20900 46620 21100 46650
rect 21400 46850 21600 46880
rect 21400 46650 21410 46850
rect 21480 46650 21520 46850
rect 21590 46650 21600 46850
rect 21400 46620 21600 46650
rect 21900 46850 22100 46880
rect 21900 46650 21910 46850
rect 21980 46650 22020 46850
rect 22090 46650 22100 46850
rect 21900 46620 22100 46650
rect 22400 46850 22600 46880
rect 22400 46650 22410 46850
rect 22480 46650 22520 46850
rect 22590 46650 22600 46850
rect 22400 46620 22600 46650
rect 22900 46850 23100 46880
rect 22900 46650 22910 46850
rect 22980 46650 23020 46850
rect 23090 46650 23100 46850
rect 22900 46620 23100 46650
rect 23400 46850 23600 46880
rect 23400 46650 23410 46850
rect 23480 46650 23520 46850
rect 23590 46650 23600 46850
rect 23400 46620 23600 46650
rect 23900 46850 24100 46880
rect 23900 46650 23910 46850
rect 23980 46650 24020 46850
rect 24090 46650 24100 46850
rect 23900 46620 24100 46650
rect 24400 46850 24600 46880
rect 24400 46650 24410 46850
rect 24480 46650 24520 46850
rect 24590 46650 24600 46850
rect 24400 46620 24600 46650
rect 24900 46850 25100 46880
rect 24900 46650 24910 46850
rect 24980 46650 25020 46850
rect 25090 46650 25100 46850
rect 24900 46620 25100 46650
rect 25400 46850 25600 46880
rect 25400 46650 25410 46850
rect 25480 46650 25520 46850
rect 25590 46650 25600 46850
rect 25400 46620 25600 46650
rect 25900 46850 26100 46880
rect 25900 46650 25910 46850
rect 25980 46650 26020 46850
rect 26090 46650 26100 46850
rect 25900 46620 26100 46650
rect 26400 46850 26500 46880
rect 26400 46650 26410 46850
rect 26480 46650 26500 46850
rect 26400 46620 26500 46650
rect 0 46600 120 46620
rect 380 46600 620 46620
rect 880 46600 1120 46620
rect 1380 46600 1620 46620
rect 1880 46600 2120 46620
rect 2380 46600 2620 46620
rect 2880 46600 3120 46620
rect 3380 46600 3620 46620
rect 3880 46600 4120 46620
rect 4380 46600 4620 46620
rect 4880 46600 5120 46620
rect 5380 46600 5620 46620
rect 5880 46600 6120 46620
rect 6380 46600 6620 46620
rect 6880 46600 7120 46620
rect 7380 46600 7620 46620
rect 7880 46600 8120 46620
rect 8380 46600 8620 46620
rect 8880 46600 9120 46620
rect 9380 46600 9620 46620
rect 9880 46600 10120 46620
rect 10380 46600 10620 46620
rect 10880 46600 11120 46620
rect 11380 46600 11620 46620
rect 11880 46600 12120 46620
rect 12380 46600 12620 46620
rect 12880 46600 13120 46620
rect 13380 46600 13620 46620
rect 13880 46600 14120 46620
rect 14380 46600 14620 46620
rect 14880 46600 15120 46620
rect 15380 46600 15620 46620
rect 15880 46600 16120 46620
rect 16380 46600 16620 46620
rect 16880 46600 17120 46620
rect 17380 46600 17620 46620
rect 17880 46600 18120 46620
rect 18380 46600 18620 46620
rect 18880 46600 19120 46620
rect 19380 46600 19620 46620
rect 19880 46600 20120 46620
rect 20380 46600 20620 46620
rect 20880 46600 21120 46620
rect 21380 46600 21620 46620
rect 21880 46600 22120 46620
rect 22380 46600 22620 46620
rect 22880 46600 23120 46620
rect 23380 46600 23620 46620
rect 23880 46600 24120 46620
rect 24380 46600 24620 46620
rect 24880 46600 25120 46620
rect 25380 46600 25620 46620
rect 25880 46600 26120 46620
rect 26380 46600 26500 46620
rect 0 46590 26500 46600
rect 0 46520 150 46590
rect 350 46520 650 46590
rect 850 46520 1150 46590
rect 1350 46520 1650 46590
rect 1850 46520 2150 46590
rect 2350 46520 2650 46590
rect 2850 46520 3150 46590
rect 3350 46520 3650 46590
rect 3850 46520 4150 46590
rect 4350 46520 4650 46590
rect 4850 46520 5150 46590
rect 5350 46520 5650 46590
rect 5850 46520 6150 46590
rect 6350 46520 6650 46590
rect 6850 46520 7150 46590
rect 7350 46520 7650 46590
rect 7850 46520 8150 46590
rect 8350 46520 8650 46590
rect 8850 46520 9150 46590
rect 9350 46520 9650 46590
rect 9850 46520 10150 46590
rect 10350 46520 10650 46590
rect 10850 46520 11150 46590
rect 11350 46520 11650 46590
rect 11850 46520 12150 46590
rect 12350 46520 12650 46590
rect 12850 46520 13150 46590
rect 13350 46520 13650 46590
rect 13850 46520 14150 46590
rect 14350 46520 14650 46590
rect 14850 46520 15150 46590
rect 15350 46520 15650 46590
rect 15850 46520 16150 46590
rect 16350 46520 16650 46590
rect 16850 46520 17150 46590
rect 17350 46520 17650 46590
rect 17850 46520 18150 46590
rect 18350 46520 18650 46590
rect 18850 46520 19150 46590
rect 19350 46520 19650 46590
rect 19850 46520 20150 46590
rect 20350 46520 20650 46590
rect 20850 46520 21150 46590
rect 21350 46520 21650 46590
rect 21850 46520 22150 46590
rect 22350 46520 22650 46590
rect 22850 46520 23150 46590
rect 23350 46520 23650 46590
rect 23850 46520 24150 46590
rect 24350 46520 24650 46590
rect 24850 46520 25150 46590
rect 25350 46520 25650 46590
rect 25850 46520 26150 46590
rect 26350 46520 26500 46590
rect 0 46500 26500 46520
rect 0 46480 1340 46500
rect 0 46410 150 46480
rect 350 46410 650 46480
rect 850 46410 1340 46480
rect 0 46400 1340 46410
rect 0 46380 120 46400
rect 380 46380 620 46400
rect 880 46380 1340 46400
rect 0 46350 100 46380
rect 0 46150 20 46350
rect 90 46150 100 46350
rect 0 46120 100 46150
rect 400 46350 600 46380
rect 400 46150 410 46350
rect 480 46150 520 46350
rect 590 46150 600 46350
rect 400 46120 600 46150
rect 900 46350 1340 46380
rect 900 46150 910 46350
rect 980 46180 1340 46350
rect 6500 46480 7500 46500
rect 6500 46410 6650 46480
rect 6850 46410 7150 46480
rect 7350 46410 7500 46480
rect 6500 46400 7500 46410
rect 6500 46380 6620 46400
rect 6880 46380 7120 46400
rect 7380 46380 7500 46400
rect 6500 46350 6600 46380
rect 980 46170 6410 46180
rect 980 46150 1536 46170
rect 900 46132 1536 46150
rect 6259 46132 6410 46170
rect 900 46122 6410 46132
rect 900 46120 1400 46122
rect 0 46100 120 46120
rect 380 46100 620 46120
rect 880 46100 1330 46120
rect 0 46090 1330 46100
rect 0 46020 150 46090
rect 350 46020 650 46090
rect 850 46020 1330 46090
rect 0 45980 1330 46020
rect 6340 46120 6410 46122
rect 1532 46030 1552 46090
rect 6186 46030 6206 46090
rect 1532 45996 1544 46030
rect 6194 45996 6206 46030
rect 1532 45990 1552 45996
rect 6186 45990 6206 45996
rect 0 45910 150 45980
rect 350 45910 650 45980
rect 850 45910 1330 45980
rect 0 45900 1330 45910
rect 0 45880 120 45900
rect 380 45880 620 45900
rect 880 45880 1330 45900
rect 0 45850 100 45880
rect 0 45650 20 45850
rect 90 45650 100 45850
rect 0 45620 100 45650
rect 400 45850 600 45880
rect 400 45650 410 45850
rect 480 45650 520 45850
rect 590 45650 600 45850
rect 400 45620 600 45650
rect 900 45850 1330 45880
rect 900 45650 910 45850
rect 980 45650 1330 45850
rect 900 45620 1330 45650
rect 0 45600 120 45620
rect 380 45600 620 45620
rect 880 45600 1330 45620
rect 0 45590 1330 45600
rect 0 45520 150 45590
rect 350 45520 650 45590
rect 850 45520 1330 45590
rect 0 45480 1330 45520
rect 0 45410 150 45480
rect 350 45410 650 45480
rect 850 45410 1330 45480
rect 0 45400 1330 45410
rect 0 45380 120 45400
rect 380 45380 620 45400
rect 880 45380 1330 45400
rect 0 45350 100 45380
rect 0 45150 20 45350
rect 90 45150 100 45350
rect 0 45120 100 45150
rect 400 45350 600 45380
rect 400 45150 410 45350
rect 480 45150 520 45350
rect 590 45150 600 45350
rect 400 45120 600 45150
rect 900 45350 1330 45380
rect 900 45150 910 45350
rect 980 45150 1330 45350
rect 900 45120 1330 45150
rect 0 45100 120 45120
rect 380 45100 620 45120
rect 880 45100 1330 45120
rect 0 45090 1330 45100
rect 0 45020 150 45090
rect 350 45020 650 45090
rect 850 45020 1330 45090
rect 0 44980 1330 45020
rect 0 44910 150 44980
rect 350 44910 650 44980
rect 850 44910 1330 44980
rect 0 44900 1330 44910
rect 0 44880 120 44900
rect 380 44880 620 44900
rect 880 44880 1330 44900
rect 0 44850 100 44880
rect 0 44650 20 44850
rect 90 44650 100 44850
rect 0 44620 100 44650
rect 400 44850 600 44880
rect 400 44650 410 44850
rect 480 44650 520 44850
rect 590 44650 600 44850
rect 400 44620 600 44650
rect 900 44850 1330 44880
rect 900 44650 910 44850
rect 980 44650 1330 44850
rect 900 44620 1330 44650
rect 0 44600 120 44620
rect 380 44600 620 44620
rect 880 44600 1330 44620
rect 0 44590 1330 44600
rect 0 44520 150 44590
rect 350 44520 650 44590
rect 850 44520 1330 44590
rect 0 44480 1330 44520
rect 0 44410 150 44480
rect 350 44410 650 44480
rect 850 44410 1330 44480
rect 0 44400 1330 44410
rect 0 44380 120 44400
rect 380 44380 620 44400
rect 880 44380 1330 44400
rect 0 44350 100 44380
rect 0 44150 20 44350
rect 90 44150 100 44350
rect 0 44120 100 44150
rect 400 44350 600 44380
rect 400 44150 410 44350
rect 480 44150 520 44350
rect 590 44150 600 44350
rect 400 44120 600 44150
rect 900 44350 1330 44380
rect 900 44150 910 44350
rect 980 44150 1330 44350
rect 900 44120 1330 44150
rect 0 44100 120 44120
rect 380 44100 620 44120
rect 880 44100 1330 44120
rect 0 44090 1330 44100
rect 0 44020 150 44090
rect 350 44020 650 44090
rect 850 44020 1330 44090
rect 0 43980 1330 44020
rect 0 43910 150 43980
rect 350 43910 650 43980
rect 850 43910 1330 43980
rect 0 43900 1330 43910
rect 0 43880 120 43900
rect 380 43880 620 43900
rect 880 43880 1330 43900
rect 0 43850 100 43880
rect 0 43650 20 43850
rect 90 43650 100 43850
rect 0 43620 100 43650
rect 400 43850 600 43880
rect 400 43650 410 43850
rect 480 43650 520 43850
rect 590 43650 600 43850
rect 400 43620 600 43650
rect 900 43850 1330 43880
rect 900 43650 910 43850
rect 980 43650 1330 43850
rect 900 43620 1330 43650
rect 0 43600 120 43620
rect 380 43600 620 43620
rect 880 43600 1330 43620
rect 0 43590 1330 43600
rect 0 43520 150 43590
rect 350 43520 650 43590
rect 850 43520 1330 43590
rect 0 43480 1330 43520
rect 0 43410 150 43480
rect 350 43410 650 43480
rect 850 43410 1330 43480
rect 0 43400 1330 43410
rect 0 43380 120 43400
rect 380 43380 620 43400
rect 880 43380 1330 43400
rect 0 43350 100 43380
rect 0 43150 20 43350
rect 90 43150 100 43350
rect 0 43120 100 43150
rect 400 43350 600 43380
rect 400 43150 410 43350
rect 480 43150 520 43350
rect 590 43150 600 43350
rect 400 43120 600 43150
rect 900 43350 1330 43380
rect 900 43150 910 43350
rect 980 43150 1330 43350
rect 900 43120 1330 43150
rect 0 43100 120 43120
rect 380 43100 620 43120
rect 880 43100 1330 43120
rect 0 43090 1330 43100
rect 0 43020 150 43090
rect 350 43020 650 43090
rect 850 43020 1330 43090
rect 0 42980 1330 43020
rect 0 42910 150 42980
rect 350 42910 650 42980
rect 850 42910 1330 42980
rect 0 42900 1330 42910
rect 0 42880 120 42900
rect 380 42880 620 42900
rect 880 42880 1330 42900
rect 0 42850 100 42880
rect 0 42650 20 42850
rect 90 42650 100 42850
rect 0 42620 100 42650
rect 400 42850 600 42880
rect 400 42650 410 42850
rect 480 42650 520 42850
rect 590 42650 600 42850
rect 400 42620 600 42650
rect 900 42850 1330 42880
rect 900 42650 910 42850
rect 980 42650 1330 42850
rect 900 42620 1330 42650
rect 0 42600 120 42620
rect 380 42600 620 42620
rect 880 42600 1330 42620
rect 0 42590 1330 42600
rect 0 42520 150 42590
rect 350 42520 650 42590
rect 850 42520 1330 42590
rect 0 42480 1330 42520
rect 0 42410 150 42480
rect 350 42410 650 42480
rect 850 42410 1330 42480
rect 0 42400 1330 42410
rect 0 42380 120 42400
rect 380 42380 620 42400
rect 880 42380 1330 42400
rect 0 42350 100 42380
rect 0 42150 20 42350
rect 90 42150 100 42350
rect 0 42120 100 42150
rect 400 42350 600 42380
rect 400 42150 410 42350
rect 480 42150 520 42350
rect 590 42150 600 42350
rect 400 42120 600 42150
rect 900 42350 1330 42380
rect 900 42150 910 42350
rect 980 42150 1330 42350
rect 900 42120 1330 42150
rect 0 42100 120 42120
rect 380 42100 620 42120
rect 880 42100 1330 42120
rect 0 42090 1330 42100
rect 0 42020 150 42090
rect 350 42020 650 42090
rect 850 42020 1330 42090
rect 0 41980 1330 42020
rect 0 41910 150 41980
rect 350 41910 650 41980
rect 850 41910 1330 41980
rect 0 41900 1330 41910
rect 0 41880 120 41900
rect 380 41880 620 41900
rect 880 41880 1330 41900
rect 0 41850 100 41880
rect 0 41650 20 41850
rect 90 41650 100 41850
rect 0 41620 100 41650
rect 400 41850 600 41880
rect 400 41650 410 41850
rect 480 41650 520 41850
rect 590 41650 600 41850
rect 400 41620 600 41650
rect 900 41850 1330 41880
rect 900 41650 910 41850
rect 980 41650 1330 41850
rect 900 41620 1330 41650
rect 0 41600 120 41620
rect 380 41600 620 41620
rect 880 41600 1330 41620
rect 0 41590 1330 41600
rect 0 41520 150 41590
rect 350 41520 650 41590
rect 850 41520 1330 41590
rect 0 41480 1330 41520
rect 0 41410 150 41480
rect 350 41410 650 41480
rect 850 41410 1330 41480
rect 0 41400 1330 41410
rect 0 41380 120 41400
rect 380 41380 620 41400
rect 880 41380 1330 41400
rect 0 41350 100 41380
rect 0 41150 20 41350
rect 90 41150 100 41350
rect 0 41120 100 41150
rect 400 41350 600 41380
rect 400 41150 410 41350
rect 480 41150 520 41350
rect 590 41150 600 41350
rect 400 41120 600 41150
rect 900 41350 1330 41380
rect 900 41150 910 41350
rect 980 41150 1330 41350
rect 900 41120 1330 41150
rect 0 41100 120 41120
rect 380 41100 620 41120
rect 880 41100 1330 41120
rect 0 41090 1330 41100
rect 0 41020 150 41090
rect 350 41020 650 41090
rect 850 41020 1330 41090
rect 0 40980 1330 41020
rect 0 40910 150 40980
rect 350 40910 650 40980
rect 850 40910 1330 40980
rect 0 40900 1330 40910
rect 0 40880 120 40900
rect 380 40880 620 40900
rect 880 40880 1330 40900
rect 0 40850 100 40880
rect 0 40650 20 40850
rect 90 40650 100 40850
rect 0 40620 100 40650
rect 400 40850 600 40880
rect 400 40650 410 40850
rect 480 40650 520 40850
rect 590 40650 600 40850
rect 400 40620 600 40650
rect 900 40850 1330 40880
rect 900 40650 910 40850
rect 980 40650 1330 40850
rect 900 40620 1330 40650
rect 0 40600 120 40620
rect 380 40600 620 40620
rect 880 40600 1330 40620
rect 0 40590 1330 40600
rect 0 40520 150 40590
rect 350 40520 650 40590
rect 850 40520 1330 40590
rect 0 40480 1330 40520
rect -3300 40450 -3100 40460
rect -3300 40190 -3290 40450
rect -3110 40190 -3100 40450
rect -3300 40180 -3100 40190
rect -3060 40400 -2980 40420
rect -3300 38910 -3100 38920
rect -3300 38690 -3290 38910
rect -3110 38690 -3100 38910
rect -3060 38740 -3040 40400
rect -3000 40000 -2980 40400
rect 0 40410 150 40480
rect 350 40410 650 40480
rect 850 40410 1330 40480
rect 0 40400 1330 40410
rect 0 40380 120 40400
rect 380 40380 620 40400
rect 880 40380 1330 40400
rect 0 40350 100 40380
rect 0 40150 20 40350
rect 90 40150 100 40350
rect 0 40120 100 40150
rect 400 40350 600 40380
rect 400 40150 410 40350
rect 480 40150 520 40350
rect 590 40150 600 40350
rect 400 40120 600 40150
rect 900 40350 1330 40380
rect 900 40150 910 40350
rect 980 40150 1330 40350
rect 900 40120 1330 40150
rect 0 40100 120 40120
rect 380 40100 620 40120
rect 880 40100 1330 40120
rect 0 40090 1330 40100
rect 0 40020 150 40090
rect 350 40020 650 40090
rect 850 40020 1330 40090
rect 0 40000 1330 40020
rect -3000 39980 1330 40000
rect -3000 39910 -2850 39980
rect -2650 39910 -2350 39980
rect -2150 39910 -1850 39980
rect -1650 39910 -1350 39980
rect -1150 39910 -850 39980
rect -650 39910 -350 39980
rect -150 39910 150 39980
rect 350 39910 650 39980
rect 850 39910 1330 39980
rect 6500 46150 6520 46350
rect 6590 46150 6600 46350
rect 6500 46120 6600 46150
rect 6900 46350 7100 46380
rect 6900 46150 6910 46350
rect 6980 46150 7020 46350
rect 7090 46150 7100 46350
rect 6900 46120 7100 46150
rect 7400 46350 7500 46380
rect 7400 46150 7410 46350
rect 7480 46150 7500 46350
rect 13000 46480 14000 46500
rect 13000 46410 13150 46480
rect 13350 46410 13650 46480
rect 13850 46410 14000 46480
rect 13000 46400 14000 46410
rect 13000 46380 13120 46400
rect 13380 46380 13620 46400
rect 13880 46380 14000 46400
rect 13000 46350 13100 46380
rect 7400 46120 7500 46150
rect 6500 46100 6620 46120
rect 6880 46100 7120 46120
rect 7380 46100 7500 46120
rect 6500 46090 7500 46100
rect 6500 46020 6650 46090
rect 6850 46020 7150 46090
rect 7350 46020 7500 46090
rect 6500 46000 7500 46020
rect 7630 46170 12710 46180
rect 7630 46132 7836 46170
rect 12559 46132 12710 46170
rect 7630 46122 12710 46132
rect 7630 46120 7700 46122
rect 1465 45946 1531 45958
rect 1465 45938 1482 45946
rect 1516 45938 1531 45946
rect 1465 39970 1482 39978
rect 1516 39970 1531 39978
rect 1465 39958 1531 39970
rect 1623 45946 1689 45958
rect 1623 45938 1640 45946
rect 1674 45938 1689 45946
rect 1623 39970 1640 39978
rect 1674 39970 1689 39978
rect 1623 39958 1689 39970
rect 1781 45946 1847 45958
rect 1781 45938 1798 45946
rect 1832 45938 1847 45946
rect 1781 39970 1798 39978
rect 1832 39970 1847 39978
rect 1781 39958 1847 39970
rect 1939 45946 2005 45958
rect 1939 45938 1956 45946
rect 1990 45938 2005 45946
rect 1939 39970 1956 39978
rect 1990 39970 2005 39978
rect 1939 39958 2005 39970
rect 2097 45946 2163 45958
rect 2097 45938 2114 45946
rect 2148 45938 2163 45946
rect 2097 39970 2114 39978
rect 2148 39970 2163 39978
rect 2097 39958 2163 39970
rect 2255 45946 2321 45958
rect 2255 45938 2272 45946
rect 2306 45938 2321 45946
rect 2255 39970 2272 39978
rect 2306 39970 2321 39978
rect 2255 39958 2321 39970
rect 2413 45946 2479 45958
rect 2413 45938 2430 45946
rect 2464 45938 2479 45946
rect 2413 39970 2430 39978
rect 2464 39970 2479 39978
rect 2413 39958 2479 39970
rect 2571 45946 2637 45958
rect 2571 45938 2588 45946
rect 2622 45938 2637 45946
rect 2571 39970 2588 39978
rect 2622 39970 2637 39978
rect 2571 39958 2637 39970
rect 2729 45946 2795 45958
rect 2729 45938 2746 45946
rect 2780 45938 2795 45946
rect 2729 39970 2746 39978
rect 2780 39970 2795 39978
rect 2729 39958 2795 39970
rect 2887 45946 2953 45958
rect 2887 45938 2904 45946
rect 2938 45938 2953 45946
rect 2887 39970 2904 39978
rect 2938 39970 2953 39978
rect 2887 39958 2953 39970
rect 3045 45946 3111 45958
rect 3045 45938 3062 45946
rect 3096 45938 3111 45946
rect 3045 39970 3062 39978
rect 3096 39970 3111 39978
rect 3045 39958 3111 39970
rect 3203 45946 3269 45958
rect 3203 45938 3220 45946
rect 3254 45938 3269 45946
rect 3203 39970 3220 39978
rect 3254 39970 3269 39978
rect 3203 39958 3269 39970
rect 3361 45946 3427 45958
rect 3361 45938 3378 45946
rect 3412 45938 3427 45946
rect 3361 39970 3378 39978
rect 3412 39970 3427 39978
rect 3361 39958 3427 39970
rect 3519 45946 3585 45958
rect 3519 45938 3536 45946
rect 3570 45938 3585 45946
rect 3519 39970 3536 39978
rect 3570 39970 3585 39978
rect 3519 39958 3585 39970
rect 3677 45946 3743 45958
rect 3677 45938 3694 45946
rect 3728 45938 3743 45946
rect 3677 39970 3694 39978
rect 3728 39970 3743 39978
rect 3677 39958 3743 39970
rect 3835 45946 3901 45958
rect 3835 45938 3852 45946
rect 3886 45938 3901 45946
rect 3835 39970 3852 39978
rect 3886 39970 3901 39978
rect 3835 39958 3901 39970
rect 3993 45946 4059 45958
rect 3993 45938 4010 45946
rect 4044 45938 4059 45946
rect 3993 39970 4010 39978
rect 4044 39970 4059 39978
rect 3993 39958 4059 39970
rect 4151 45946 4217 45958
rect 4151 45938 4168 45946
rect 4202 45938 4217 45946
rect 4151 39970 4168 39978
rect 4202 39970 4217 39978
rect 4151 39958 4217 39970
rect 4309 45946 4375 45958
rect 4309 45938 4326 45946
rect 4360 45938 4375 45946
rect 4309 39970 4326 39978
rect 4360 39970 4375 39978
rect 4309 39958 4375 39970
rect 4467 45946 4533 45958
rect 4467 45938 4484 45946
rect 4518 45938 4533 45946
rect 4467 39970 4484 39978
rect 4518 39970 4533 39978
rect 4467 39958 4533 39970
rect 4625 45946 4691 45958
rect 4625 45938 4642 45946
rect 4676 45938 4691 45946
rect 4625 39970 4642 39978
rect 4676 39970 4691 39978
rect 4625 39958 4691 39970
rect 4783 45946 4849 45958
rect 4783 45938 4800 45946
rect 4834 45938 4849 45946
rect 4783 39970 4800 39978
rect 4834 39970 4849 39978
rect 4783 39958 4849 39970
rect 4941 45946 5007 45958
rect 4941 45938 4958 45946
rect 4992 45938 5007 45946
rect 4941 39970 4958 39978
rect 4992 39970 5007 39978
rect 4941 39958 5007 39970
rect 5099 45946 5165 45958
rect 5099 45938 5116 45946
rect 5150 45938 5165 45946
rect 5099 39970 5116 39978
rect 5150 39970 5165 39978
rect 5099 39958 5165 39970
rect 5257 45946 5323 45958
rect 5257 45938 5274 45946
rect 5308 45938 5323 45946
rect 5257 39970 5274 39978
rect 5308 39970 5323 39978
rect 5257 39958 5323 39970
rect 5415 45946 5481 45958
rect 5415 45938 5432 45946
rect 5466 45938 5481 45946
rect 5415 39970 5432 39978
rect 5466 39970 5481 39978
rect 5415 39958 5481 39970
rect 5573 45946 5639 45958
rect 5573 45938 5590 45946
rect 5624 45938 5639 45946
rect 5573 39970 5590 39978
rect 5624 39970 5639 39978
rect 5573 39958 5639 39970
rect 5731 45946 5797 45958
rect 5731 45938 5748 45946
rect 5782 45938 5797 45946
rect 5731 39970 5748 39978
rect 5782 39970 5797 39978
rect 5731 39958 5797 39970
rect 5889 45946 5955 45958
rect 5889 45938 5906 45946
rect 5940 45938 5955 45946
rect 5889 39970 5906 39978
rect 5940 39970 5955 39978
rect 5889 39958 5955 39970
rect 6047 45946 6113 45958
rect 6047 45938 6064 45946
rect 6098 45938 6113 45946
rect 6047 39970 6064 39978
rect 6098 39970 6113 39978
rect 6047 39958 6113 39970
rect 6205 45946 6271 45958
rect 6205 45938 6222 45946
rect 6256 45938 6271 45946
rect 6205 39970 6222 39978
rect 6256 39970 6271 39978
rect 6205 39958 6271 39970
rect -3000 39900 1330 39910
rect -3000 39880 -2880 39900
rect -2620 39880 -2380 39900
rect -2120 39880 -1880 39900
rect -1620 39880 -1380 39900
rect -1120 39880 -880 39900
rect -620 39880 -380 39900
rect -120 39880 120 39900
rect 380 39880 620 39900
rect 880 39880 1330 39900
rect -3000 39850 -2900 39880
rect -3000 39650 -2980 39850
rect -2910 39650 -2900 39850
rect -3000 39620 -2900 39650
rect -2600 39850 -2400 39880
rect -2600 39650 -2590 39850
rect -2520 39650 -2480 39850
rect -2410 39650 -2400 39850
rect -2600 39620 -2400 39650
rect -2100 39850 -1900 39880
rect -2100 39650 -2090 39850
rect -2020 39650 -1980 39850
rect -1910 39650 -1900 39850
rect -2100 39620 -1900 39650
rect -1600 39850 -1400 39880
rect -1600 39650 -1590 39850
rect -1520 39650 -1480 39850
rect -1410 39650 -1400 39850
rect -1600 39620 -1400 39650
rect -1100 39850 -900 39880
rect -1100 39650 -1090 39850
rect -1020 39650 -980 39850
rect -910 39650 -900 39850
rect -1100 39620 -900 39650
rect -600 39850 -400 39880
rect -600 39650 -590 39850
rect -520 39650 -480 39850
rect -410 39650 -400 39850
rect -600 39620 -400 39650
rect -100 39850 100 39880
rect -100 39650 -90 39850
rect -20 39650 20 39850
rect 90 39650 100 39850
rect -100 39620 100 39650
rect 400 39850 600 39880
rect 400 39650 410 39850
rect 480 39650 520 39850
rect 590 39650 600 39850
rect 400 39620 600 39650
rect 900 39850 1330 39880
rect 900 39650 910 39850
rect 980 39800 1330 39850
rect 1532 39920 1552 39926
rect 6186 39920 6206 39926
rect 1532 39886 1544 39920
rect 6194 39886 6206 39920
rect 1532 39826 1552 39886
rect 6186 39826 6206 39886
rect 980 39794 1400 39800
rect 6340 39794 6410 39800
rect 980 39784 6410 39794
rect 980 39746 1536 39784
rect 6202 39746 6410 39784
rect 980 39730 6410 39746
rect 12640 46120 12710 46122
rect 7832 46030 7852 46090
rect 12486 46030 12506 46090
rect 7832 45996 7844 46030
rect 12494 45996 12506 46030
rect 7832 45990 7852 45996
rect 12486 45990 12506 45996
rect 13000 46150 13020 46350
rect 13090 46150 13100 46350
rect 13000 46120 13100 46150
rect 13400 46350 13600 46380
rect 13400 46150 13410 46350
rect 13480 46150 13520 46350
rect 13590 46150 13600 46350
rect 13400 46120 13600 46150
rect 13900 46350 14000 46380
rect 13900 46150 13910 46350
rect 13980 46180 14000 46350
rect 19000 46480 20000 46500
rect 19000 46410 19150 46480
rect 19350 46410 19650 46480
rect 19850 46410 20000 46480
rect 19000 46400 20000 46410
rect 19000 46380 19120 46400
rect 19380 46380 19620 46400
rect 19880 46380 20000 46400
rect 19000 46350 19100 46380
rect 19000 46180 19020 46350
rect 13980 46170 19020 46180
rect 13980 46150 14136 46170
rect 13900 46132 14136 46150
rect 18859 46150 19020 46170
rect 19090 46150 19100 46350
rect 18859 46132 19100 46150
rect 13900 46122 19100 46132
rect 13900 46120 14000 46122
rect 13000 46100 13120 46120
rect 13380 46100 13620 46120
rect 13880 46100 13930 46120
rect 13000 46090 13930 46100
rect 13000 46020 13150 46090
rect 13350 46020 13650 46090
rect 13850 46020 13930 46090
rect 13000 46000 13930 46020
rect 7765 45946 7831 45958
rect 7765 45938 7782 45946
rect 7816 45938 7831 45946
rect 7765 39970 7782 39978
rect 7816 39970 7831 39978
rect 7765 39958 7831 39970
rect 7923 45946 7989 45958
rect 7923 45938 7940 45946
rect 7974 45938 7989 45946
rect 7923 39970 7940 39978
rect 7974 39970 7989 39978
rect 7923 39958 7989 39970
rect 8081 45946 8147 45958
rect 8081 45938 8098 45946
rect 8132 45938 8147 45946
rect 8081 39970 8098 39978
rect 8132 39970 8147 39978
rect 8081 39958 8147 39970
rect 8239 45946 8305 45958
rect 8239 45938 8256 45946
rect 8290 45938 8305 45946
rect 8239 39970 8256 39978
rect 8290 39970 8305 39978
rect 8239 39958 8305 39970
rect 8397 45946 8463 45958
rect 8397 45938 8414 45946
rect 8448 45938 8463 45946
rect 8397 39970 8414 39978
rect 8448 39970 8463 39978
rect 8397 39958 8463 39970
rect 8555 45946 8621 45958
rect 8555 45938 8572 45946
rect 8606 45938 8621 45946
rect 8555 39970 8572 39978
rect 8606 39970 8621 39978
rect 8555 39958 8621 39970
rect 8713 45946 8779 45958
rect 8713 45938 8730 45946
rect 8764 45938 8779 45946
rect 8713 39970 8730 39978
rect 8764 39970 8779 39978
rect 8713 39958 8779 39970
rect 8871 45946 8937 45958
rect 8871 45938 8888 45946
rect 8922 45938 8937 45946
rect 8871 39970 8888 39978
rect 8922 39970 8937 39978
rect 8871 39958 8937 39970
rect 9029 45946 9095 45958
rect 9029 45938 9046 45946
rect 9080 45938 9095 45946
rect 9029 39970 9046 39978
rect 9080 39970 9095 39978
rect 9029 39958 9095 39970
rect 9187 45946 9253 45958
rect 9187 45938 9204 45946
rect 9238 45938 9253 45946
rect 9187 39970 9204 39978
rect 9238 39970 9253 39978
rect 9187 39958 9253 39970
rect 9345 45946 9411 45958
rect 9345 45938 9362 45946
rect 9396 45938 9411 45946
rect 9345 39970 9362 39978
rect 9396 39970 9411 39978
rect 9345 39958 9411 39970
rect 9503 45946 9569 45958
rect 9503 45938 9520 45946
rect 9554 45938 9569 45946
rect 9503 39970 9520 39978
rect 9554 39970 9569 39978
rect 9503 39958 9569 39970
rect 9661 45946 9727 45958
rect 9661 45938 9678 45946
rect 9712 45938 9727 45946
rect 9661 39970 9678 39978
rect 9712 39970 9727 39978
rect 9661 39958 9727 39970
rect 9819 45946 9885 45958
rect 9819 45938 9836 45946
rect 9870 45938 9885 45946
rect 9819 39970 9836 39978
rect 9870 39970 9885 39978
rect 9819 39958 9885 39970
rect 9977 45946 10043 45958
rect 9977 45938 9994 45946
rect 10028 45938 10043 45946
rect 9977 39970 9994 39978
rect 10028 39970 10043 39978
rect 9977 39958 10043 39970
rect 10135 45946 10201 45958
rect 10135 45938 10152 45946
rect 10186 45938 10201 45946
rect 10135 39970 10152 39978
rect 10186 39970 10201 39978
rect 10135 39958 10201 39970
rect 10293 45946 10359 45958
rect 10293 45938 10310 45946
rect 10344 45938 10359 45946
rect 10293 39970 10310 39978
rect 10344 39970 10359 39978
rect 10293 39958 10359 39970
rect 10451 45946 10517 45958
rect 10451 45938 10468 45946
rect 10502 45938 10517 45946
rect 10451 39970 10468 39978
rect 10502 39970 10517 39978
rect 10451 39958 10517 39970
rect 10609 45946 10675 45958
rect 10609 45938 10626 45946
rect 10660 45938 10675 45946
rect 10609 39970 10626 39978
rect 10660 39970 10675 39978
rect 10609 39958 10675 39970
rect 10767 45946 10833 45958
rect 10767 45938 10784 45946
rect 10818 45938 10833 45946
rect 10767 39970 10784 39978
rect 10818 39970 10833 39978
rect 10767 39958 10833 39970
rect 10925 45946 10991 45958
rect 10925 45938 10942 45946
rect 10976 45938 10991 45946
rect 10925 39970 10942 39978
rect 10976 39970 10991 39978
rect 10925 39958 10991 39970
rect 11083 45946 11149 45958
rect 11083 45938 11100 45946
rect 11134 45938 11149 45946
rect 11083 39970 11100 39978
rect 11134 39970 11149 39978
rect 11083 39958 11149 39970
rect 11241 45946 11307 45958
rect 11241 45938 11258 45946
rect 11292 45938 11307 45946
rect 11241 39970 11258 39978
rect 11292 39970 11307 39978
rect 11241 39958 11307 39970
rect 11399 45946 11465 45958
rect 11399 45938 11416 45946
rect 11450 45938 11465 45946
rect 11399 39970 11416 39978
rect 11450 39970 11465 39978
rect 11399 39958 11465 39970
rect 11557 45946 11623 45958
rect 11557 45938 11574 45946
rect 11608 45938 11623 45946
rect 11557 39970 11574 39978
rect 11608 39970 11623 39978
rect 11557 39958 11623 39970
rect 11715 45946 11781 45958
rect 11715 45938 11732 45946
rect 11766 45938 11781 45946
rect 11715 39970 11732 39978
rect 11766 39970 11781 39978
rect 11715 39958 11781 39970
rect 11873 45946 11939 45958
rect 11873 45938 11890 45946
rect 11924 45938 11939 45946
rect 11873 39970 11890 39978
rect 11924 39970 11939 39978
rect 11873 39958 11939 39970
rect 12031 45946 12097 45958
rect 12031 45938 12048 45946
rect 12082 45938 12097 45946
rect 12031 39970 12048 39978
rect 12082 39970 12097 39978
rect 12031 39958 12097 39970
rect 12189 45946 12255 45958
rect 12189 45938 12206 45946
rect 12240 45938 12255 45946
rect 12189 39970 12206 39978
rect 12240 39970 12255 39978
rect 12189 39958 12255 39970
rect 12347 45946 12413 45958
rect 12347 45938 12364 45946
rect 12398 45938 12413 45946
rect 12347 39970 12364 39978
rect 12398 39970 12413 39978
rect 12347 39958 12413 39970
rect 12505 45946 12571 45958
rect 12505 45938 12522 45946
rect 12556 45938 12571 45946
rect 12505 39970 12522 39978
rect 12556 39970 12571 39978
rect 12505 39958 12571 39970
rect 7832 39920 7852 39926
rect 12486 39920 12506 39926
rect 7832 39886 7844 39920
rect 12494 39886 12506 39920
rect 7832 39826 7852 39886
rect 12486 39826 12506 39886
rect 7630 39794 7700 39800
rect 12640 39794 12710 39800
rect 7630 39784 12710 39794
rect 7630 39746 7836 39784
rect 12502 39746 12710 39784
rect 7630 39730 12710 39746
rect 18940 46120 19100 46122
rect 19400 46350 19600 46380
rect 19400 46150 19410 46350
rect 19480 46150 19520 46350
rect 19590 46150 19600 46350
rect 19400 46120 19600 46150
rect 19900 46350 20000 46380
rect 19900 46150 19910 46350
rect 19980 46150 20000 46350
rect 25260 46480 26500 46500
rect 25260 46410 25650 46480
rect 25850 46410 26150 46480
rect 26350 46410 26500 46480
rect 25260 46400 26500 46410
rect 25260 46380 25620 46400
rect 25880 46380 26120 46400
rect 26380 46380 26500 46400
rect 25260 46350 25600 46380
rect 25260 46180 25520 46350
rect 19900 46120 20000 46150
rect 14132 46030 14152 46090
rect 18786 46030 18806 46090
rect 14132 45996 14144 46030
rect 18794 45996 18806 46030
rect 14132 45990 14152 45996
rect 18786 45990 18806 45996
rect 19010 46100 19120 46120
rect 19380 46100 19620 46120
rect 19880 46100 20000 46120
rect 19010 46090 20000 46100
rect 19010 46020 19150 46090
rect 19350 46020 19650 46090
rect 19850 46020 20000 46090
rect 19010 46000 20000 46020
rect 20230 46170 25520 46180
rect 20230 46132 20436 46170
rect 25159 46150 25520 46170
rect 25590 46150 25600 46350
rect 25159 46132 25600 46150
rect 20230 46122 25600 46132
rect 20230 46120 20300 46122
rect 14065 45946 14131 45958
rect 14065 45938 14082 45946
rect 14116 45938 14131 45946
rect 14065 39970 14082 39978
rect 14116 39970 14131 39978
rect 14065 39958 14131 39970
rect 14223 45946 14289 45958
rect 14223 45938 14240 45946
rect 14274 45938 14289 45946
rect 14223 39970 14240 39978
rect 14274 39970 14289 39978
rect 14223 39958 14289 39970
rect 14381 45946 14447 45958
rect 14381 45938 14398 45946
rect 14432 45938 14447 45946
rect 14381 39970 14398 39978
rect 14432 39970 14447 39978
rect 14381 39958 14447 39970
rect 14539 45946 14605 45958
rect 14539 45938 14556 45946
rect 14590 45938 14605 45946
rect 14539 39970 14556 39978
rect 14590 39970 14605 39978
rect 14539 39958 14605 39970
rect 14697 45946 14763 45958
rect 14697 45938 14714 45946
rect 14748 45938 14763 45946
rect 14697 39970 14714 39978
rect 14748 39970 14763 39978
rect 14697 39958 14763 39970
rect 14855 45946 14921 45958
rect 14855 45938 14872 45946
rect 14906 45938 14921 45946
rect 14855 39970 14872 39978
rect 14906 39970 14921 39978
rect 14855 39958 14921 39970
rect 15013 45946 15079 45958
rect 15013 45938 15030 45946
rect 15064 45938 15079 45946
rect 15013 39970 15030 39978
rect 15064 39970 15079 39978
rect 15013 39958 15079 39970
rect 15171 45946 15237 45958
rect 15171 45938 15188 45946
rect 15222 45938 15237 45946
rect 15171 39970 15188 39978
rect 15222 39970 15237 39978
rect 15171 39958 15237 39970
rect 15329 45946 15395 45958
rect 15329 45938 15346 45946
rect 15380 45938 15395 45946
rect 15329 39970 15346 39978
rect 15380 39970 15395 39978
rect 15329 39958 15395 39970
rect 15487 45946 15553 45958
rect 15487 45938 15504 45946
rect 15538 45938 15553 45946
rect 15487 39970 15504 39978
rect 15538 39970 15553 39978
rect 15487 39958 15553 39970
rect 15645 45946 15711 45958
rect 15645 45938 15662 45946
rect 15696 45938 15711 45946
rect 15645 39970 15662 39978
rect 15696 39970 15711 39978
rect 15645 39958 15711 39970
rect 15803 45946 15869 45958
rect 15803 45938 15820 45946
rect 15854 45938 15869 45946
rect 15803 39970 15820 39978
rect 15854 39970 15869 39978
rect 15803 39958 15869 39970
rect 15961 45946 16027 45958
rect 15961 45938 15978 45946
rect 16012 45938 16027 45946
rect 15961 39970 15978 39978
rect 16012 39970 16027 39978
rect 15961 39958 16027 39970
rect 16119 45946 16185 45958
rect 16119 45938 16136 45946
rect 16170 45938 16185 45946
rect 16119 39970 16136 39978
rect 16170 39970 16185 39978
rect 16119 39958 16185 39970
rect 16277 45946 16343 45958
rect 16277 45938 16294 45946
rect 16328 45938 16343 45946
rect 16277 39970 16294 39978
rect 16328 39970 16343 39978
rect 16277 39958 16343 39970
rect 16435 45946 16501 45958
rect 16435 45938 16452 45946
rect 16486 45938 16501 45946
rect 16435 39970 16452 39978
rect 16486 39970 16501 39978
rect 16435 39958 16501 39970
rect 16593 45946 16659 45958
rect 16593 45938 16610 45946
rect 16644 45938 16659 45946
rect 16593 39970 16610 39978
rect 16644 39970 16659 39978
rect 16593 39958 16659 39970
rect 16751 45946 16817 45958
rect 16751 45938 16768 45946
rect 16802 45938 16817 45946
rect 16751 39970 16768 39978
rect 16802 39970 16817 39978
rect 16751 39958 16817 39970
rect 16909 45946 16975 45958
rect 16909 45938 16926 45946
rect 16960 45938 16975 45946
rect 16909 39970 16926 39978
rect 16960 39970 16975 39978
rect 16909 39958 16975 39970
rect 17067 45946 17133 45958
rect 17067 45938 17084 45946
rect 17118 45938 17133 45946
rect 17067 39970 17084 39978
rect 17118 39970 17133 39978
rect 17067 39958 17133 39970
rect 17225 45946 17291 45958
rect 17225 45938 17242 45946
rect 17276 45938 17291 45946
rect 17225 39970 17242 39978
rect 17276 39970 17291 39978
rect 17225 39958 17291 39970
rect 17383 45946 17449 45958
rect 17383 45938 17400 45946
rect 17434 45938 17449 45946
rect 17383 39970 17400 39978
rect 17434 39970 17449 39978
rect 17383 39958 17449 39970
rect 17541 45946 17607 45958
rect 17541 45938 17558 45946
rect 17592 45938 17607 45946
rect 17541 39970 17558 39978
rect 17592 39970 17607 39978
rect 17541 39958 17607 39970
rect 17699 45946 17765 45958
rect 17699 45938 17716 45946
rect 17750 45938 17765 45946
rect 17699 39970 17716 39978
rect 17750 39970 17765 39978
rect 17699 39958 17765 39970
rect 17857 45946 17923 45958
rect 17857 45938 17874 45946
rect 17908 45938 17923 45946
rect 17857 39970 17874 39978
rect 17908 39970 17923 39978
rect 17857 39958 17923 39970
rect 18015 45946 18081 45958
rect 18015 45938 18032 45946
rect 18066 45938 18081 45946
rect 18015 39970 18032 39978
rect 18066 39970 18081 39978
rect 18015 39958 18081 39970
rect 18173 45946 18239 45958
rect 18173 45938 18190 45946
rect 18224 45938 18239 45946
rect 18173 39970 18190 39978
rect 18224 39970 18239 39978
rect 18173 39958 18239 39970
rect 18331 45946 18397 45958
rect 18331 45938 18348 45946
rect 18382 45938 18397 45946
rect 18331 39970 18348 39978
rect 18382 39970 18397 39978
rect 18331 39958 18397 39970
rect 18489 45946 18555 45958
rect 18489 45938 18506 45946
rect 18540 45938 18555 45946
rect 18489 39970 18506 39978
rect 18540 39970 18555 39978
rect 18489 39958 18555 39970
rect 18647 45946 18713 45958
rect 18647 45938 18664 45946
rect 18698 45938 18713 45946
rect 18647 39970 18664 39978
rect 18698 39970 18713 39978
rect 18647 39958 18713 39970
rect 18805 45946 18871 45958
rect 18805 45938 18822 45946
rect 18856 45938 18871 45946
rect 18805 39970 18822 39978
rect 18856 39970 18871 39978
rect 18805 39958 18871 39970
rect 14132 39920 14152 39926
rect 18786 39920 18806 39926
rect 14132 39886 14144 39920
rect 18794 39886 18806 39920
rect 14132 39826 14152 39886
rect 18786 39826 18806 39886
rect 13930 39794 14000 39800
rect 18940 39794 19010 39800
rect 13930 39784 19010 39794
rect 13930 39746 14136 39784
rect 18802 39746 19010 39784
rect 13930 39730 19010 39746
rect 25240 46120 25600 46122
rect 25900 46350 26100 46380
rect 25900 46150 25910 46350
rect 25980 46150 26020 46350
rect 26090 46150 26100 46350
rect 25900 46120 26100 46150
rect 26400 46350 26500 46380
rect 26400 46150 26410 46350
rect 26480 46150 26500 46350
rect 26400 46120 26500 46150
rect 20432 46030 20452 46090
rect 25086 46030 25106 46090
rect 20432 45996 20444 46030
rect 25094 45996 25106 46030
rect 20432 45990 20452 45996
rect 25086 45990 25106 45996
rect 25310 46100 25620 46120
rect 25880 46100 26120 46120
rect 26380 46100 26500 46120
rect 25310 46090 26500 46100
rect 25310 46020 25650 46090
rect 25850 46020 26150 46090
rect 26350 46020 26500 46090
rect 25310 45980 26500 46020
rect 20365 45946 20431 45958
rect 20365 45938 20382 45946
rect 20416 45938 20431 45946
rect 20365 39970 20382 39978
rect 20416 39970 20431 39978
rect 20365 39958 20431 39970
rect 20523 45946 20589 45958
rect 20523 45938 20540 45946
rect 20574 45938 20589 45946
rect 20523 39970 20540 39978
rect 20574 39970 20589 39978
rect 20523 39958 20589 39970
rect 20681 45946 20747 45958
rect 20681 45938 20698 45946
rect 20732 45938 20747 45946
rect 20681 39970 20698 39978
rect 20732 39970 20747 39978
rect 20681 39958 20747 39970
rect 20839 45946 20905 45958
rect 20839 45938 20856 45946
rect 20890 45938 20905 45946
rect 20839 39970 20856 39978
rect 20890 39970 20905 39978
rect 20839 39958 20905 39970
rect 20997 45946 21063 45958
rect 20997 45938 21014 45946
rect 21048 45938 21063 45946
rect 20997 39970 21014 39978
rect 21048 39970 21063 39978
rect 20997 39958 21063 39970
rect 21155 45946 21221 45958
rect 21155 45938 21172 45946
rect 21206 45938 21221 45946
rect 21155 39970 21172 39978
rect 21206 39970 21221 39978
rect 21155 39958 21221 39970
rect 21313 45946 21379 45958
rect 21313 45938 21330 45946
rect 21364 45938 21379 45946
rect 21313 39970 21330 39978
rect 21364 39970 21379 39978
rect 21313 39958 21379 39970
rect 21471 45946 21537 45958
rect 21471 45938 21488 45946
rect 21522 45938 21537 45946
rect 21471 39970 21488 39978
rect 21522 39970 21537 39978
rect 21471 39958 21537 39970
rect 21629 45946 21695 45958
rect 21629 45938 21646 45946
rect 21680 45938 21695 45946
rect 21629 39970 21646 39978
rect 21680 39970 21695 39978
rect 21629 39958 21695 39970
rect 21787 45946 21853 45958
rect 21787 45938 21804 45946
rect 21838 45938 21853 45946
rect 21787 39970 21804 39978
rect 21838 39970 21853 39978
rect 21787 39958 21853 39970
rect 21945 45946 22011 45958
rect 21945 45938 21962 45946
rect 21996 45938 22011 45946
rect 21945 39970 21962 39978
rect 21996 39970 22011 39978
rect 21945 39958 22011 39970
rect 22103 45946 22169 45958
rect 22103 45938 22120 45946
rect 22154 45938 22169 45946
rect 22103 39970 22120 39978
rect 22154 39970 22169 39978
rect 22103 39958 22169 39970
rect 22261 45946 22327 45958
rect 22261 45938 22278 45946
rect 22312 45938 22327 45946
rect 22261 39970 22278 39978
rect 22312 39970 22327 39978
rect 22261 39958 22327 39970
rect 22419 45946 22485 45958
rect 22419 45938 22436 45946
rect 22470 45938 22485 45946
rect 22419 39970 22436 39978
rect 22470 39970 22485 39978
rect 22419 39958 22485 39970
rect 22577 45946 22643 45958
rect 22577 45938 22594 45946
rect 22628 45938 22643 45946
rect 22577 39970 22594 39978
rect 22628 39970 22643 39978
rect 22577 39958 22643 39970
rect 22735 45946 22801 45958
rect 22735 45938 22752 45946
rect 22786 45938 22801 45946
rect 22735 39970 22752 39978
rect 22786 39970 22801 39978
rect 22735 39958 22801 39970
rect 22893 45946 22959 45958
rect 22893 45938 22910 45946
rect 22944 45938 22959 45946
rect 22893 39970 22910 39978
rect 22944 39970 22959 39978
rect 22893 39958 22959 39970
rect 23051 45946 23117 45958
rect 23051 45938 23068 45946
rect 23102 45938 23117 45946
rect 23051 39970 23068 39978
rect 23102 39970 23117 39978
rect 23051 39958 23117 39970
rect 23209 45946 23275 45958
rect 23209 45938 23226 45946
rect 23260 45938 23275 45946
rect 23209 39970 23226 39978
rect 23260 39970 23275 39978
rect 23209 39958 23275 39970
rect 23367 45946 23433 45958
rect 23367 45938 23384 45946
rect 23418 45938 23433 45946
rect 23367 39970 23384 39978
rect 23418 39970 23433 39978
rect 23367 39958 23433 39970
rect 23525 45946 23591 45958
rect 23525 45938 23542 45946
rect 23576 45938 23591 45946
rect 23525 39970 23542 39978
rect 23576 39970 23591 39978
rect 23525 39958 23591 39970
rect 23683 45946 23749 45958
rect 23683 45938 23700 45946
rect 23734 45938 23749 45946
rect 23683 39970 23700 39978
rect 23734 39970 23749 39978
rect 23683 39958 23749 39970
rect 23841 45946 23907 45958
rect 23841 45938 23858 45946
rect 23892 45938 23907 45946
rect 23841 39970 23858 39978
rect 23892 39970 23907 39978
rect 23841 39958 23907 39970
rect 23999 45946 24065 45958
rect 23999 45938 24016 45946
rect 24050 45938 24065 45946
rect 23999 39970 24016 39978
rect 24050 39970 24065 39978
rect 23999 39958 24065 39970
rect 24157 45946 24223 45958
rect 24157 45938 24174 45946
rect 24208 45938 24223 45946
rect 24157 39970 24174 39978
rect 24208 39970 24223 39978
rect 24157 39958 24223 39970
rect 24315 45946 24381 45958
rect 24315 45938 24332 45946
rect 24366 45938 24381 45946
rect 24315 39970 24332 39978
rect 24366 39970 24381 39978
rect 24315 39958 24381 39970
rect 24473 45946 24539 45958
rect 24473 45938 24490 45946
rect 24524 45938 24539 45946
rect 24473 39970 24490 39978
rect 24524 39970 24539 39978
rect 24473 39958 24539 39970
rect 24631 45946 24697 45958
rect 24631 45938 24648 45946
rect 24682 45938 24697 45946
rect 24631 39970 24648 39978
rect 24682 39970 24697 39978
rect 24631 39958 24697 39970
rect 24789 45946 24855 45958
rect 24789 45938 24806 45946
rect 24840 45938 24855 45946
rect 24789 39970 24806 39978
rect 24840 39970 24855 39978
rect 24789 39958 24855 39970
rect 24947 45946 25013 45958
rect 24947 45938 24964 45946
rect 24998 45938 25013 45946
rect 24947 39970 24964 39978
rect 24998 39970 25013 39978
rect 24947 39958 25013 39970
rect 25105 45946 25171 45958
rect 25105 45938 25122 45946
rect 25156 45938 25171 45946
rect 25105 39970 25122 39978
rect 25156 39970 25171 39978
rect 25105 39958 25171 39970
rect 25310 45910 25650 45980
rect 25850 45910 26150 45980
rect 26350 45910 26500 45980
rect 25310 45900 26500 45910
rect 25310 45880 25620 45900
rect 25880 45880 26120 45900
rect 26380 45880 26500 45900
rect 25310 45850 25600 45880
rect 25310 45650 25520 45850
rect 25590 45650 25600 45850
rect 25310 45620 25600 45650
rect 25900 45850 26100 45880
rect 25900 45650 25910 45850
rect 25980 45650 26020 45850
rect 26090 45650 26100 45850
rect 25900 45620 26100 45650
rect 26400 45850 26500 45880
rect 26400 45650 26410 45850
rect 26480 45650 26500 45850
rect 26400 45620 26500 45650
rect 25310 45600 25620 45620
rect 25880 45600 26120 45620
rect 26380 45600 26500 45620
rect 25310 45590 26500 45600
rect 25310 45520 25650 45590
rect 25850 45520 26150 45590
rect 26350 45520 26500 45590
rect 25310 45480 26500 45520
rect 25310 45410 25650 45480
rect 25850 45410 26150 45480
rect 26350 45410 26500 45480
rect 25310 45400 26500 45410
rect 25310 45380 25620 45400
rect 25880 45380 26120 45400
rect 26380 45380 26500 45400
rect 25310 45350 25600 45380
rect 25310 45150 25520 45350
rect 25590 45150 25600 45350
rect 25310 45120 25600 45150
rect 25900 45350 26100 45380
rect 25900 45150 25910 45350
rect 25980 45150 26020 45350
rect 26090 45150 26100 45350
rect 25900 45120 26100 45150
rect 26400 45350 26500 45380
rect 26400 45150 26410 45350
rect 26480 45150 26500 45350
rect 26400 45120 26500 45150
rect 25310 45100 25620 45120
rect 25880 45100 26120 45120
rect 26380 45100 26500 45120
rect 25310 45090 26500 45100
rect 25310 45020 25650 45090
rect 25850 45020 26150 45090
rect 26350 45020 26500 45090
rect 25310 44980 26500 45020
rect 25310 44910 25650 44980
rect 25850 44910 26150 44980
rect 26350 44910 26500 44980
rect 25310 44900 26500 44910
rect 25310 44880 25620 44900
rect 25880 44880 26120 44900
rect 26380 44880 26500 44900
rect 25310 44850 25600 44880
rect 25310 44650 25520 44850
rect 25590 44650 25600 44850
rect 25310 44620 25600 44650
rect 25900 44850 26100 44880
rect 25900 44650 25910 44850
rect 25980 44650 26020 44850
rect 26090 44650 26100 44850
rect 25900 44620 26100 44650
rect 26400 44850 26500 44880
rect 26400 44650 26410 44850
rect 26480 44650 26500 44850
rect 26400 44620 26500 44650
rect 25310 44600 25620 44620
rect 25880 44600 26120 44620
rect 26380 44600 26500 44620
rect 25310 44590 26500 44600
rect 25310 44520 25650 44590
rect 25850 44520 26150 44590
rect 26350 44520 26500 44590
rect 25310 44480 26500 44520
rect 25310 44410 25650 44480
rect 25850 44410 26150 44480
rect 26350 44410 26500 44480
rect 25310 44400 26500 44410
rect 25310 44380 25620 44400
rect 25880 44380 26120 44400
rect 26380 44380 26500 44400
rect 25310 44350 25600 44380
rect 25310 44150 25520 44350
rect 25590 44150 25600 44350
rect 25310 44120 25600 44150
rect 25900 44350 26100 44380
rect 25900 44150 25910 44350
rect 25980 44150 26020 44350
rect 26090 44150 26100 44350
rect 25900 44120 26100 44150
rect 26400 44350 26500 44380
rect 26400 44150 26410 44350
rect 26480 44150 26500 44350
rect 26400 44120 26500 44150
rect 25310 44100 25620 44120
rect 25880 44100 26120 44120
rect 26380 44100 26500 44120
rect 25310 44090 26500 44100
rect 25310 44020 25650 44090
rect 25850 44020 26150 44090
rect 26350 44020 26500 44090
rect 25310 43980 26500 44020
rect 25310 43910 25650 43980
rect 25850 43910 26150 43980
rect 26350 43910 26500 43980
rect 25310 43900 26500 43910
rect 25310 43880 25620 43900
rect 25880 43880 26120 43900
rect 26380 43880 26500 43900
rect 25310 43850 25600 43880
rect 25310 43650 25520 43850
rect 25590 43650 25600 43850
rect 25310 43620 25600 43650
rect 25900 43850 26100 43880
rect 25900 43650 25910 43850
rect 25980 43650 26020 43850
rect 26090 43650 26100 43850
rect 25900 43620 26100 43650
rect 26400 43850 26500 43880
rect 26400 43650 26410 43850
rect 26480 43650 26500 43850
rect 26400 43620 26500 43650
rect 25310 43600 25620 43620
rect 25880 43600 26120 43620
rect 26380 43600 26500 43620
rect 25310 43590 26500 43600
rect 25310 43520 25650 43590
rect 25850 43520 26150 43590
rect 26350 43520 26500 43590
rect 25310 43480 26500 43520
rect 25310 43410 25650 43480
rect 25850 43410 26150 43480
rect 26350 43410 26500 43480
rect 25310 43400 26500 43410
rect 25310 43380 25620 43400
rect 25880 43380 26120 43400
rect 26380 43380 26500 43400
rect 25310 43350 25600 43380
rect 25310 43150 25520 43350
rect 25590 43150 25600 43350
rect 25310 43120 25600 43150
rect 25900 43350 26100 43380
rect 25900 43150 25910 43350
rect 25980 43150 26020 43350
rect 26090 43150 26100 43350
rect 25900 43120 26100 43150
rect 26400 43350 26500 43380
rect 26400 43150 26410 43350
rect 26480 43150 26500 43350
rect 26400 43120 26500 43150
rect 25310 43100 25620 43120
rect 25880 43100 26120 43120
rect 26380 43100 26500 43120
rect 25310 43090 26500 43100
rect 25310 43020 25650 43090
rect 25850 43020 26150 43090
rect 26350 43020 26500 43090
rect 25310 42980 26500 43020
rect 25310 42910 25650 42980
rect 25850 42910 26150 42980
rect 26350 42910 26500 42980
rect 25310 42900 26500 42910
rect 25310 42880 25620 42900
rect 25880 42880 26120 42900
rect 26380 42880 26500 42900
rect 25310 42850 25600 42880
rect 25310 42650 25520 42850
rect 25590 42650 25600 42850
rect 25310 42620 25600 42650
rect 25900 42850 26100 42880
rect 25900 42650 25910 42850
rect 25980 42650 26020 42850
rect 26090 42650 26100 42850
rect 25900 42620 26100 42650
rect 26400 42850 26500 42880
rect 26400 42650 26410 42850
rect 26480 42650 26500 42850
rect 26400 42620 26500 42650
rect 25310 42600 25620 42620
rect 25880 42600 26120 42620
rect 26380 42600 26500 42620
rect 25310 42590 26500 42600
rect 25310 42520 25650 42590
rect 25850 42520 26150 42590
rect 26350 42520 26500 42590
rect 25310 42480 26500 42520
rect 25310 42410 25650 42480
rect 25850 42410 26150 42480
rect 26350 42410 26500 42480
rect 25310 42400 26500 42410
rect 25310 42380 25620 42400
rect 25880 42380 26120 42400
rect 26380 42380 26500 42400
rect 25310 42350 25600 42380
rect 25310 42150 25520 42350
rect 25590 42150 25600 42350
rect 25310 42120 25600 42150
rect 25900 42350 26100 42380
rect 25900 42150 25910 42350
rect 25980 42150 26020 42350
rect 26090 42150 26100 42350
rect 25900 42120 26100 42150
rect 26400 42350 26500 42380
rect 26400 42150 26410 42350
rect 26480 42150 26500 42350
rect 26400 42120 26500 42150
rect 25310 42100 25620 42120
rect 25880 42100 26120 42120
rect 26380 42100 26500 42120
rect 25310 42090 26500 42100
rect 25310 42020 25650 42090
rect 25850 42020 26150 42090
rect 26350 42020 26500 42090
rect 25310 41980 26500 42020
rect 25310 41910 25650 41980
rect 25850 41910 26150 41980
rect 26350 41910 26500 41980
rect 25310 41900 26500 41910
rect 25310 41880 25620 41900
rect 25880 41880 26120 41900
rect 26380 41880 26500 41900
rect 25310 41850 25600 41880
rect 25310 41650 25520 41850
rect 25590 41650 25600 41850
rect 25310 41620 25600 41650
rect 25900 41850 26100 41880
rect 25900 41650 25910 41850
rect 25980 41650 26020 41850
rect 26090 41650 26100 41850
rect 25900 41620 26100 41650
rect 26400 41850 26500 41880
rect 26400 41650 26410 41850
rect 26480 41650 26500 41850
rect 26400 41620 26500 41650
rect 25310 41600 25620 41620
rect 25880 41600 26120 41620
rect 26380 41600 26500 41620
rect 25310 41590 26500 41600
rect 25310 41520 25650 41590
rect 25850 41520 26150 41590
rect 26350 41520 26500 41590
rect 25310 41480 26500 41520
rect 25310 41410 25650 41480
rect 25850 41410 26150 41480
rect 26350 41410 26500 41480
rect 25310 41400 26500 41410
rect 25310 41380 25620 41400
rect 25880 41380 26120 41400
rect 26380 41380 26500 41400
rect 25310 41350 25600 41380
rect 25310 41150 25520 41350
rect 25590 41150 25600 41350
rect 25310 41120 25600 41150
rect 25900 41350 26100 41380
rect 25900 41150 25910 41350
rect 25980 41150 26020 41350
rect 26090 41150 26100 41350
rect 25900 41120 26100 41150
rect 26400 41350 26500 41380
rect 26400 41150 26410 41350
rect 26480 41150 26500 41350
rect 26400 41120 26500 41150
rect 25310 41100 25620 41120
rect 25880 41100 26120 41120
rect 26380 41100 26500 41120
rect 25310 41090 26500 41100
rect 25310 41020 25650 41090
rect 25850 41020 26150 41090
rect 26350 41020 26500 41090
rect 25310 40980 26500 41020
rect 25310 40910 25650 40980
rect 25850 40910 26150 40980
rect 26350 40910 26500 40980
rect 25310 40900 26500 40910
rect 25310 40880 25620 40900
rect 25880 40880 26120 40900
rect 26380 40880 26500 40900
rect 25310 40850 25600 40880
rect 25310 40650 25520 40850
rect 25590 40650 25600 40850
rect 25310 40620 25600 40650
rect 25900 40850 26100 40880
rect 25900 40650 25910 40850
rect 25980 40650 26020 40850
rect 26090 40650 26100 40850
rect 25900 40620 26100 40650
rect 26400 40850 26500 40880
rect 26400 40650 26410 40850
rect 26480 40650 26500 40850
rect 26400 40620 26500 40650
rect 25310 40600 25620 40620
rect 25880 40600 26120 40620
rect 26380 40600 26500 40620
rect 25310 40590 26500 40600
rect 25310 40520 25650 40590
rect 25850 40520 26150 40590
rect 26350 40520 26500 40590
rect 25310 40480 26500 40520
rect 25310 40410 25650 40480
rect 25850 40410 26150 40480
rect 26350 40410 26500 40480
rect 29900 40450 30100 40460
rect 25310 40400 26500 40410
rect 25310 40380 25620 40400
rect 25880 40380 26120 40400
rect 26380 40380 26500 40400
rect 25310 40350 25600 40380
rect 25310 40150 25520 40350
rect 25590 40150 25600 40350
rect 25310 40120 25600 40150
rect 25900 40350 26100 40380
rect 25900 40150 25910 40350
rect 25980 40150 26020 40350
rect 26090 40150 26100 40350
rect 25900 40120 26100 40150
rect 26400 40350 26500 40380
rect 26400 40150 26410 40350
rect 26480 40150 26500 40350
rect 26400 40120 26500 40150
rect 25310 40100 25620 40120
rect 25880 40100 26120 40120
rect 26380 40100 26500 40120
rect 25310 40090 26500 40100
rect 25310 40020 25650 40090
rect 25850 40020 26150 40090
rect 26350 40020 26500 40090
rect 25310 40000 26500 40020
rect 29780 40400 29860 40420
rect 29780 40000 29800 40400
rect 25310 39980 29800 40000
rect 20432 39920 20452 39926
rect 25086 39920 25106 39926
rect 20432 39886 20444 39920
rect 25094 39886 25106 39920
rect 20432 39826 20452 39886
rect 25086 39826 25106 39886
rect 20230 39794 20300 39800
rect 25310 39910 25650 39980
rect 25850 39910 26150 39980
rect 26350 39910 26650 39980
rect 26850 39910 27150 39980
rect 27350 39910 27650 39980
rect 27850 39910 28150 39980
rect 28350 39910 28650 39980
rect 28850 39910 29150 39980
rect 29350 39910 29800 39980
rect 25310 39900 29800 39910
rect 25310 39880 25620 39900
rect 25880 39880 26120 39900
rect 26380 39880 26620 39900
rect 26880 39880 27120 39900
rect 27380 39880 27620 39900
rect 27880 39880 28120 39900
rect 28380 39880 28620 39900
rect 28880 39880 29120 39900
rect 29380 39880 29800 39900
rect 25310 39850 25600 39880
rect 25310 39800 25520 39850
rect 25240 39794 25520 39800
rect 20230 39784 25520 39794
rect 20230 39746 20436 39784
rect 25102 39746 25520 39784
rect 20230 39730 25520 39746
rect 980 39650 1340 39730
rect 900 39620 1340 39650
rect -3000 39600 -2880 39620
rect -2620 39600 -2380 39620
rect -2120 39600 -1880 39620
rect -1620 39600 -1380 39620
rect -1120 39600 -880 39620
rect -620 39600 -380 39620
rect -120 39600 120 39620
rect 380 39600 620 39620
rect 880 39600 1340 39620
rect -3000 39590 1340 39600
rect -3000 39520 -2850 39590
rect -2650 39520 -2350 39590
rect -2150 39520 -1850 39590
rect -1650 39520 -1350 39590
rect -1150 39520 -850 39590
rect -650 39520 -350 39590
rect -150 39520 150 39590
rect 350 39520 650 39590
rect 850 39520 1340 39590
rect -3000 39480 1340 39520
rect -3000 39410 -2850 39480
rect -2650 39410 -2350 39480
rect -2150 39410 -1850 39480
rect -1650 39410 -1350 39480
rect -1150 39410 -850 39480
rect -650 39410 -350 39480
rect -150 39410 150 39480
rect 350 39410 650 39480
rect 850 39410 1340 39480
rect -3000 39400 1340 39410
rect -3000 39380 -2880 39400
rect -2620 39380 -2380 39400
rect -2120 39380 -1880 39400
rect -1620 39380 -1380 39400
rect -1120 39380 -880 39400
rect -620 39380 -380 39400
rect -120 39380 120 39400
rect 380 39380 620 39400
rect 880 39380 1340 39400
rect -3000 39350 -2900 39380
rect -3000 39150 -2980 39350
rect -2910 39150 -2900 39350
rect -3000 39120 -2900 39150
rect -2600 39350 -2400 39380
rect -2600 39150 -2590 39350
rect -2520 39150 -2480 39350
rect -2410 39150 -2400 39350
rect -2600 39120 -2400 39150
rect -2100 39350 -1900 39380
rect -2100 39150 -2090 39350
rect -2020 39150 -1980 39350
rect -1910 39150 -1900 39350
rect -2100 39120 -1900 39150
rect -1600 39350 -1400 39380
rect -1600 39150 -1590 39350
rect -1520 39150 -1480 39350
rect -1410 39150 -1400 39350
rect -1600 39120 -1400 39150
rect -1100 39350 -900 39380
rect -1100 39150 -1090 39350
rect -1020 39150 -980 39350
rect -910 39150 -900 39350
rect -1100 39120 -900 39150
rect -600 39350 -400 39380
rect -600 39150 -590 39350
rect -520 39150 -480 39350
rect -410 39150 -400 39350
rect -600 39120 -400 39150
rect -100 39350 100 39380
rect -100 39150 -90 39350
rect -20 39150 20 39350
rect 90 39150 100 39350
rect -100 39120 100 39150
rect 400 39350 600 39380
rect 400 39150 410 39350
rect 480 39150 520 39350
rect 590 39150 600 39350
rect 400 39120 600 39150
rect 900 39350 1340 39380
rect 900 39150 910 39350
rect 980 39180 1340 39350
rect 25260 39650 25520 39730
rect 25590 39650 25600 39850
rect 25260 39620 25600 39650
rect 25900 39850 26100 39880
rect 25900 39650 25910 39850
rect 25980 39650 26020 39850
rect 26090 39650 26100 39850
rect 25900 39620 26100 39650
rect 26400 39850 26600 39880
rect 26400 39650 26410 39850
rect 26480 39650 26520 39850
rect 26590 39650 26600 39850
rect 26400 39620 26600 39650
rect 26900 39850 27100 39880
rect 26900 39650 26910 39850
rect 26980 39650 27020 39850
rect 27090 39650 27100 39850
rect 26900 39620 27100 39650
rect 27400 39850 27600 39880
rect 27400 39650 27410 39850
rect 27480 39650 27520 39850
rect 27590 39650 27600 39850
rect 27400 39620 27600 39650
rect 27900 39850 28100 39880
rect 27900 39650 27910 39850
rect 27980 39650 28020 39850
rect 28090 39650 28100 39850
rect 27900 39620 28100 39650
rect 28400 39850 28600 39880
rect 28400 39650 28410 39850
rect 28480 39650 28520 39850
rect 28590 39650 28600 39850
rect 28400 39620 28600 39650
rect 28900 39850 29100 39880
rect 28900 39650 28910 39850
rect 28980 39650 29020 39850
rect 29090 39650 29100 39850
rect 28900 39620 29100 39650
rect 29400 39850 29800 39880
rect 29400 39650 29410 39850
rect 29480 39650 29800 39850
rect 29400 39620 29800 39650
rect 25260 39600 25620 39620
rect 25880 39600 26120 39620
rect 26380 39600 26620 39620
rect 26880 39600 27120 39620
rect 27380 39600 27620 39620
rect 27880 39600 28120 39620
rect 28380 39600 28620 39620
rect 28880 39600 29120 39620
rect 29380 39600 29800 39620
rect 25260 39590 29800 39600
rect 25260 39520 25650 39590
rect 25850 39520 26150 39590
rect 26350 39520 26650 39590
rect 26850 39520 27150 39590
rect 27350 39520 27650 39590
rect 27850 39520 28150 39590
rect 28350 39520 28650 39590
rect 28850 39520 29150 39590
rect 29350 39520 29800 39590
rect 25260 39480 29800 39520
rect 25260 39410 25650 39480
rect 25850 39410 26150 39480
rect 26350 39410 26650 39480
rect 26850 39410 27150 39480
rect 27350 39410 27650 39480
rect 27850 39410 28150 39480
rect 28350 39410 28650 39480
rect 28850 39410 29150 39480
rect 29350 39410 29800 39480
rect 25260 39400 29800 39410
rect 25260 39380 25620 39400
rect 25880 39380 26120 39400
rect 26380 39380 26620 39400
rect 26880 39380 27120 39400
rect 27380 39380 27620 39400
rect 27880 39380 28120 39400
rect 28380 39380 28620 39400
rect 28880 39380 29120 39400
rect 29380 39380 29800 39400
rect 25260 39350 25600 39380
rect 25260 39180 25520 39350
rect 980 39170 6410 39180
rect 980 39150 1536 39170
rect 900 39132 1536 39150
rect 6259 39132 6410 39170
rect 900 39122 6410 39132
rect 900 39120 1400 39122
rect -3000 39100 -2880 39120
rect -2620 39100 -2380 39120
rect -2120 39100 -1880 39120
rect -1620 39100 -1380 39120
rect -1120 39100 -880 39120
rect -620 39100 -380 39120
rect -120 39100 120 39120
rect 380 39100 620 39120
rect 880 39100 1330 39120
rect -3000 39090 1330 39100
rect -3000 39020 -2850 39090
rect -2650 39020 -2350 39090
rect -2150 39020 -1850 39090
rect -1650 39020 -1350 39090
rect -1150 39020 -850 39090
rect -650 39020 -350 39090
rect -150 39020 150 39090
rect 350 39020 650 39090
rect 850 39020 1330 39090
rect -3000 39000 1330 39020
rect -3000 38740 -2980 39000
rect -3060 38720 -2980 38740
rect 0 38980 1330 39000
rect 6340 39120 6410 39122
rect 1532 39030 1552 39090
rect 6186 39030 6206 39090
rect 1532 38996 1544 39030
rect 6194 38996 6206 39030
rect 1532 38990 1552 38996
rect 6186 38990 6206 38996
rect 0 38910 150 38980
rect 350 38910 650 38980
rect 850 38910 1330 38980
rect 0 38900 1330 38910
rect 0 38880 120 38900
rect 380 38880 620 38900
rect 880 38880 1330 38900
rect 0 38850 100 38880
rect -3300 38680 -3100 38690
rect 0 38650 20 38850
rect 90 38650 100 38850
rect 0 38620 100 38650
rect 400 38850 600 38880
rect 400 38650 410 38850
rect 480 38650 520 38850
rect 590 38650 600 38850
rect 400 38620 600 38650
rect 900 38850 1330 38880
rect 900 38650 910 38850
rect 980 38650 1330 38850
rect 900 38620 1330 38650
rect 0 38600 120 38620
rect 380 38600 620 38620
rect 880 38600 1330 38620
rect 0 38590 1330 38600
rect 0 38520 150 38590
rect 350 38520 650 38590
rect 850 38520 1330 38590
rect 0 38480 1330 38520
rect 0 38410 150 38480
rect 350 38410 650 38480
rect 850 38410 1330 38480
rect 0 38400 1330 38410
rect 0 38380 120 38400
rect 380 38380 620 38400
rect 880 38380 1330 38400
rect 0 38350 100 38380
rect 0 38150 20 38350
rect 90 38150 100 38350
rect 0 38120 100 38150
rect 400 38350 600 38380
rect 400 38150 410 38350
rect 480 38150 520 38350
rect 590 38150 600 38350
rect 400 38120 600 38150
rect 900 38350 1330 38380
rect 900 38150 910 38350
rect 980 38150 1330 38350
rect 900 38120 1330 38150
rect 0 38100 120 38120
rect 380 38100 620 38120
rect 880 38100 1330 38120
rect 0 38090 1330 38100
rect 0 38020 150 38090
rect 350 38020 650 38090
rect 850 38020 1330 38090
rect 0 37980 1330 38020
rect 0 37910 150 37980
rect 350 37910 650 37980
rect 850 37910 1330 37980
rect 0 37900 1330 37910
rect 0 37880 120 37900
rect 380 37880 620 37900
rect 880 37880 1330 37900
rect 0 37850 100 37880
rect 0 37650 20 37850
rect 90 37650 100 37850
rect 0 37620 100 37650
rect 400 37850 600 37880
rect 400 37650 410 37850
rect 480 37650 520 37850
rect 590 37650 600 37850
rect 400 37620 600 37650
rect 900 37850 1330 37880
rect 900 37650 910 37850
rect 980 37650 1330 37850
rect 900 37620 1330 37650
rect 0 37600 120 37620
rect 380 37600 620 37620
rect 880 37600 1330 37620
rect 0 37590 1330 37600
rect 0 37520 150 37590
rect 350 37520 650 37590
rect 850 37520 1330 37590
rect 0 37480 1330 37520
rect 0 37410 150 37480
rect 350 37410 650 37480
rect 850 37410 1330 37480
rect 0 37400 1330 37410
rect 0 37380 120 37400
rect 380 37380 620 37400
rect 880 37380 1330 37400
rect 0 37350 100 37380
rect 0 37150 20 37350
rect 90 37150 100 37350
rect 0 37120 100 37150
rect 400 37350 600 37380
rect 400 37150 410 37350
rect 480 37150 520 37350
rect 590 37150 600 37350
rect 400 37120 600 37150
rect 900 37350 1330 37380
rect 900 37150 910 37350
rect 980 37150 1330 37350
rect 900 37120 1330 37150
rect 0 37100 120 37120
rect 380 37100 620 37120
rect 880 37100 1330 37120
rect 0 37090 1330 37100
rect 0 37020 150 37090
rect 350 37020 650 37090
rect 850 37020 1330 37090
rect 0 36980 1330 37020
rect 0 36910 150 36980
rect 350 36910 650 36980
rect 850 36910 1330 36980
rect 0 36900 1330 36910
rect 0 36880 120 36900
rect 380 36880 620 36900
rect 880 36880 1330 36900
rect 0 36850 100 36880
rect 0 36650 20 36850
rect 90 36650 100 36850
rect 0 36620 100 36650
rect 400 36850 600 36880
rect 400 36650 410 36850
rect 480 36650 520 36850
rect 590 36650 600 36850
rect 400 36620 600 36650
rect 900 36850 1330 36880
rect 900 36650 910 36850
rect 980 36650 1330 36850
rect 900 36620 1330 36650
rect 0 36600 120 36620
rect 380 36600 620 36620
rect 880 36600 1330 36620
rect 0 36590 1330 36600
rect 0 36520 150 36590
rect 350 36520 650 36590
rect 850 36520 1330 36590
rect 0 36480 1330 36520
rect 0 36410 150 36480
rect 350 36410 650 36480
rect 850 36410 1330 36480
rect 0 36400 1330 36410
rect 0 36380 120 36400
rect 380 36380 620 36400
rect 880 36380 1330 36400
rect 0 36350 100 36380
rect 0 36150 20 36350
rect 90 36150 100 36350
rect 0 36120 100 36150
rect 400 36350 600 36380
rect 400 36150 410 36350
rect 480 36150 520 36350
rect 590 36150 600 36350
rect 400 36120 600 36150
rect 900 36350 1330 36380
rect 900 36150 910 36350
rect 980 36150 1330 36350
rect 900 36120 1330 36150
rect 0 36100 120 36120
rect 380 36100 620 36120
rect 880 36100 1330 36120
rect 0 36090 1330 36100
rect 0 36020 150 36090
rect 350 36020 650 36090
rect 850 36020 1330 36090
rect 0 35980 1330 36020
rect 0 35910 150 35980
rect 350 35910 650 35980
rect 850 35910 1330 35980
rect 0 35900 1330 35910
rect 0 35880 120 35900
rect 380 35880 620 35900
rect 880 35880 1330 35900
rect 0 35850 100 35880
rect 0 35650 20 35850
rect 90 35650 100 35850
rect 0 35620 100 35650
rect 400 35850 600 35880
rect 400 35650 410 35850
rect 480 35650 520 35850
rect 590 35650 600 35850
rect 400 35620 600 35650
rect 900 35850 1330 35880
rect 900 35650 910 35850
rect 980 35650 1330 35850
rect 900 35620 1330 35650
rect 0 35600 120 35620
rect 380 35600 620 35620
rect 880 35600 1330 35620
rect 0 35590 1330 35600
rect 0 35520 150 35590
rect 350 35520 650 35590
rect 850 35520 1330 35590
rect 0 35480 1330 35520
rect 0 35410 150 35480
rect 350 35410 650 35480
rect 850 35410 1330 35480
rect 0 35400 1330 35410
rect 0 35380 120 35400
rect 380 35380 620 35400
rect 880 35380 1330 35400
rect 0 35350 100 35380
rect 0 35150 20 35350
rect 90 35150 100 35350
rect 0 35120 100 35150
rect 400 35350 600 35380
rect 400 35150 410 35350
rect 480 35150 520 35350
rect 590 35150 600 35350
rect 400 35120 600 35150
rect 900 35350 1330 35380
rect 900 35150 910 35350
rect 980 35150 1330 35350
rect 900 35120 1330 35150
rect 0 35100 120 35120
rect 380 35100 620 35120
rect 880 35100 1330 35120
rect 0 35090 1330 35100
rect 0 35020 150 35090
rect 350 35020 650 35090
rect 850 35020 1330 35090
rect 0 34980 1330 35020
rect 0 34910 150 34980
rect 350 34910 650 34980
rect 850 34910 1330 34980
rect 0 34900 1330 34910
rect 0 34880 120 34900
rect 380 34880 620 34900
rect 880 34880 1330 34900
rect 0 34850 100 34880
rect 0 34650 20 34850
rect 90 34650 100 34850
rect 0 34620 100 34650
rect 400 34850 600 34880
rect 400 34650 410 34850
rect 480 34650 520 34850
rect 590 34650 600 34850
rect 400 34620 600 34650
rect 900 34850 1330 34880
rect 900 34650 910 34850
rect 980 34650 1330 34850
rect 900 34620 1330 34650
rect 0 34600 120 34620
rect 380 34600 620 34620
rect 880 34600 1330 34620
rect 0 34590 1330 34600
rect 0 34520 150 34590
rect 350 34520 650 34590
rect 850 34520 1330 34590
rect 0 34480 1330 34520
rect 0 34410 150 34480
rect 350 34410 650 34480
rect 850 34410 1330 34480
rect 0 34400 1330 34410
rect 0 34380 120 34400
rect 380 34380 620 34400
rect 880 34380 1330 34400
rect 0 34350 100 34380
rect 0 34150 20 34350
rect 90 34150 100 34350
rect 0 34120 100 34150
rect 400 34350 600 34380
rect 400 34150 410 34350
rect 480 34150 520 34350
rect 590 34150 600 34350
rect 400 34120 600 34150
rect 900 34350 1330 34380
rect 900 34150 910 34350
rect 980 34150 1330 34350
rect 900 34120 1330 34150
rect 0 34100 120 34120
rect 380 34100 620 34120
rect 880 34100 1330 34120
rect 0 34090 1330 34100
rect 0 34020 150 34090
rect 350 34020 650 34090
rect 850 34020 1330 34090
rect 0 33980 1330 34020
rect 0 33910 150 33980
rect 350 33910 650 33980
rect 850 33910 1330 33980
rect 0 33900 1330 33910
rect 0 33880 120 33900
rect 380 33880 620 33900
rect 880 33880 1330 33900
rect 0 33850 100 33880
rect 0 33650 20 33850
rect 90 33650 100 33850
rect 0 33620 100 33650
rect 400 33850 600 33880
rect 400 33650 410 33850
rect 480 33650 520 33850
rect 590 33650 600 33850
rect 400 33620 600 33650
rect 900 33850 1330 33880
rect 900 33650 910 33850
rect 980 33650 1330 33850
rect 900 33620 1330 33650
rect 0 33600 120 33620
rect 380 33600 620 33620
rect 880 33600 1330 33620
rect 0 33590 1330 33600
rect 0 33520 150 33590
rect 350 33520 650 33590
rect 850 33520 1330 33590
rect 0 33480 1330 33520
rect 0 33410 150 33480
rect 350 33410 650 33480
rect 850 33410 1330 33480
rect 0 33400 1330 33410
rect 0 33380 120 33400
rect 380 33380 620 33400
rect 880 33380 1330 33400
rect 0 33350 100 33380
rect 0 33150 20 33350
rect 90 33150 100 33350
rect 0 33120 100 33150
rect 400 33350 600 33380
rect 400 33150 410 33350
rect 480 33150 520 33350
rect 590 33150 600 33350
rect 400 33120 600 33150
rect 900 33350 1330 33380
rect 900 33150 910 33350
rect 980 33150 1330 33350
rect 900 33120 1330 33150
rect 0 33100 120 33120
rect 380 33100 620 33120
rect 880 33100 1330 33120
rect 0 33090 1330 33100
rect 0 33020 150 33090
rect 350 33020 650 33090
rect 850 33020 1330 33090
rect 0 32980 1330 33020
rect 0 32910 150 32980
rect 350 32910 650 32980
rect 850 32910 1330 32980
rect 1465 38946 1531 38958
rect 1465 38938 1482 38946
rect 1516 38938 1531 38946
rect 1465 32970 1482 32978
rect 1516 32970 1531 32978
rect 1465 32958 1531 32970
rect 1623 38946 1689 38958
rect 1623 38938 1640 38946
rect 1674 38938 1689 38946
rect 1623 32970 1640 32978
rect 1674 32970 1689 32978
rect 1623 32958 1689 32970
rect 1781 38946 1847 38958
rect 1781 38938 1798 38946
rect 1832 38938 1847 38946
rect 1781 32970 1798 32978
rect 1832 32970 1847 32978
rect 1781 32958 1847 32970
rect 1939 38946 2005 38958
rect 1939 38938 1956 38946
rect 1990 38938 2005 38946
rect 1939 32970 1956 32978
rect 1990 32970 2005 32978
rect 1939 32958 2005 32970
rect 2097 38946 2163 38958
rect 2097 38938 2114 38946
rect 2148 38938 2163 38946
rect 2097 32970 2114 32978
rect 2148 32970 2163 32978
rect 2097 32958 2163 32970
rect 2255 38946 2321 38958
rect 2255 38938 2272 38946
rect 2306 38938 2321 38946
rect 2255 32970 2272 32978
rect 2306 32970 2321 32978
rect 2255 32958 2321 32970
rect 2413 38946 2479 38958
rect 2413 38938 2430 38946
rect 2464 38938 2479 38946
rect 2413 32970 2430 32978
rect 2464 32970 2479 32978
rect 2413 32958 2479 32970
rect 2571 38946 2637 38958
rect 2571 38938 2588 38946
rect 2622 38938 2637 38946
rect 2571 32970 2588 32978
rect 2622 32970 2637 32978
rect 2571 32958 2637 32970
rect 2729 38946 2795 38958
rect 2729 38938 2746 38946
rect 2780 38938 2795 38946
rect 2729 32970 2746 32978
rect 2780 32970 2795 32978
rect 2729 32958 2795 32970
rect 2887 38946 2953 38958
rect 2887 38938 2904 38946
rect 2938 38938 2953 38946
rect 2887 32970 2904 32978
rect 2938 32970 2953 32978
rect 2887 32958 2953 32970
rect 3045 38946 3111 38958
rect 3045 38938 3062 38946
rect 3096 38938 3111 38946
rect 3045 32970 3062 32978
rect 3096 32970 3111 32978
rect 3045 32958 3111 32970
rect 3203 38946 3269 38958
rect 3203 38938 3220 38946
rect 3254 38938 3269 38946
rect 3203 32970 3220 32978
rect 3254 32970 3269 32978
rect 3203 32958 3269 32970
rect 3361 38946 3427 38958
rect 3361 38938 3378 38946
rect 3412 38938 3427 38946
rect 3361 32970 3378 32978
rect 3412 32970 3427 32978
rect 3361 32958 3427 32970
rect 3519 38946 3585 38958
rect 3519 38938 3536 38946
rect 3570 38938 3585 38946
rect 3519 32970 3536 32978
rect 3570 32970 3585 32978
rect 3519 32958 3585 32970
rect 3677 38946 3743 38958
rect 3677 38938 3694 38946
rect 3728 38938 3743 38946
rect 3677 32970 3694 32978
rect 3728 32970 3743 32978
rect 3677 32958 3743 32970
rect 3835 38946 3901 38958
rect 3835 38938 3852 38946
rect 3886 38938 3901 38946
rect 3835 32970 3852 32978
rect 3886 32970 3901 32978
rect 3835 32958 3901 32970
rect 3993 38946 4059 38958
rect 3993 38938 4010 38946
rect 4044 38938 4059 38946
rect 3993 32970 4010 32978
rect 4044 32970 4059 32978
rect 3993 32958 4059 32970
rect 4151 38946 4217 38958
rect 4151 38938 4168 38946
rect 4202 38938 4217 38946
rect 4151 32970 4168 32978
rect 4202 32970 4217 32978
rect 4151 32958 4217 32970
rect 4309 38946 4375 38958
rect 4309 38938 4326 38946
rect 4360 38938 4375 38946
rect 4309 32970 4326 32978
rect 4360 32970 4375 32978
rect 4309 32958 4375 32970
rect 4467 38946 4533 38958
rect 4467 38938 4484 38946
rect 4518 38938 4533 38946
rect 4467 32970 4484 32978
rect 4518 32970 4533 32978
rect 4467 32958 4533 32970
rect 4625 38946 4691 38958
rect 4625 38938 4642 38946
rect 4676 38938 4691 38946
rect 4625 32970 4642 32978
rect 4676 32970 4691 32978
rect 4625 32958 4691 32970
rect 4783 38946 4849 38958
rect 4783 38938 4800 38946
rect 4834 38938 4849 38946
rect 4783 32970 4800 32978
rect 4834 32970 4849 32978
rect 4783 32958 4849 32970
rect 4941 38946 5007 38958
rect 4941 38938 4958 38946
rect 4992 38938 5007 38946
rect 4941 32970 4958 32978
rect 4992 32970 5007 32978
rect 4941 32958 5007 32970
rect 5099 38946 5165 38958
rect 5099 38938 5116 38946
rect 5150 38938 5165 38946
rect 5099 32970 5116 32978
rect 5150 32970 5165 32978
rect 5099 32958 5165 32970
rect 5257 38946 5323 38958
rect 5257 38938 5274 38946
rect 5308 38938 5323 38946
rect 5257 32970 5274 32978
rect 5308 32970 5323 32978
rect 5257 32958 5323 32970
rect 5415 38946 5481 38958
rect 5415 38938 5432 38946
rect 5466 38938 5481 38946
rect 5415 32970 5432 32978
rect 5466 32970 5481 32978
rect 5415 32958 5481 32970
rect 5573 38946 5639 38958
rect 5573 38938 5590 38946
rect 5624 38938 5639 38946
rect 5573 32970 5590 32978
rect 5624 32970 5639 32978
rect 5573 32958 5639 32970
rect 5731 38946 5797 38958
rect 5731 38938 5748 38946
rect 5782 38938 5797 38946
rect 5731 32970 5748 32978
rect 5782 32970 5797 32978
rect 5731 32958 5797 32970
rect 5889 38946 5955 38958
rect 5889 38938 5906 38946
rect 5940 38938 5955 38946
rect 5889 32970 5906 32978
rect 5940 32970 5955 32978
rect 5889 32958 5955 32970
rect 6047 38946 6113 38958
rect 6047 38938 6064 38946
rect 6098 38938 6113 38946
rect 6047 32970 6064 32978
rect 6098 32970 6113 32978
rect 6047 32958 6113 32970
rect 6205 38946 6271 38958
rect 6205 38938 6222 38946
rect 6256 38938 6271 38946
rect 6205 32970 6222 32978
rect 6256 32970 6271 32978
rect 6205 32958 6271 32970
rect 0 32900 1330 32910
rect 0 32880 120 32900
rect 380 32880 620 32900
rect 880 32880 1330 32900
rect 0 32850 100 32880
rect 0 32650 20 32850
rect 90 32650 100 32850
rect 0 32620 100 32650
rect 400 32850 600 32880
rect 400 32650 410 32850
rect 480 32650 520 32850
rect 590 32650 600 32850
rect 400 32620 600 32650
rect 900 32850 1330 32880
rect 900 32650 910 32850
rect 980 32800 1330 32850
rect 7630 39170 12710 39180
rect 7630 39132 7836 39170
rect 12559 39132 12710 39170
rect 7630 39122 12710 39132
rect 7630 39120 7700 39122
rect 12640 39120 12710 39122
rect 7832 39030 7852 39090
rect 12486 39030 12506 39090
rect 7832 38996 7844 39030
rect 12494 38996 12506 39030
rect 7832 38990 7852 38996
rect 12486 38990 12506 38996
rect 1532 32920 1552 32926
rect 6186 32920 6206 32926
rect 1532 32886 1544 32920
rect 6194 32886 6206 32920
rect 1532 32826 1552 32886
rect 6186 32826 6206 32886
rect 980 32794 1400 32800
rect 6340 32794 6410 32800
rect 980 32784 6410 32794
rect 980 32746 1536 32784
rect 6202 32746 6410 32784
rect 980 32730 6410 32746
rect 6500 32980 7500 33000
rect 6500 32910 6650 32980
rect 6850 32910 7150 32980
rect 7350 32910 7500 32980
rect 6500 32900 7500 32910
rect 6500 32880 6620 32900
rect 6880 32880 7120 32900
rect 7380 32880 7500 32900
rect 6500 32850 6600 32880
rect 980 32650 1340 32730
rect 900 32620 1340 32650
rect 0 32600 120 32620
rect 380 32600 620 32620
rect 880 32600 1340 32620
rect 0 32590 1340 32600
rect 0 32520 150 32590
rect 350 32520 650 32590
rect 850 32520 1340 32590
rect 0 32500 1340 32520
rect 6500 32650 6520 32850
rect 6590 32650 6600 32850
rect 6500 32620 6600 32650
rect 6900 32850 7100 32880
rect 6900 32650 6910 32850
rect 6980 32650 7020 32850
rect 7090 32650 7100 32850
rect 6900 32620 7100 32650
rect 7400 32850 7500 32880
rect 7400 32650 7410 32850
rect 7480 32650 7500 32850
rect 7765 38946 7831 38958
rect 7765 38938 7782 38946
rect 7816 38938 7831 38946
rect 7765 32970 7782 32978
rect 7816 32970 7831 32978
rect 7765 32958 7831 32970
rect 7923 38946 7989 38958
rect 7923 38938 7940 38946
rect 7974 38938 7989 38946
rect 7923 32970 7940 32978
rect 7974 32970 7989 32978
rect 7923 32958 7989 32970
rect 8081 38946 8147 38958
rect 8081 38938 8098 38946
rect 8132 38938 8147 38946
rect 8081 32970 8098 32978
rect 8132 32970 8147 32978
rect 8081 32958 8147 32970
rect 8239 38946 8305 38958
rect 8239 38938 8256 38946
rect 8290 38938 8305 38946
rect 8239 32970 8256 32978
rect 8290 32970 8305 32978
rect 8239 32958 8305 32970
rect 8397 38946 8463 38958
rect 8397 38938 8414 38946
rect 8448 38938 8463 38946
rect 8397 32970 8414 32978
rect 8448 32970 8463 32978
rect 8397 32958 8463 32970
rect 8555 38946 8621 38958
rect 8555 38938 8572 38946
rect 8606 38938 8621 38946
rect 8555 32970 8572 32978
rect 8606 32970 8621 32978
rect 8555 32958 8621 32970
rect 8713 38946 8779 38958
rect 8713 38938 8730 38946
rect 8764 38938 8779 38946
rect 8713 32970 8730 32978
rect 8764 32970 8779 32978
rect 8713 32958 8779 32970
rect 8871 38946 8937 38958
rect 8871 38938 8888 38946
rect 8922 38938 8937 38946
rect 8871 32970 8888 32978
rect 8922 32970 8937 32978
rect 8871 32958 8937 32970
rect 9029 38946 9095 38958
rect 9029 38938 9046 38946
rect 9080 38938 9095 38946
rect 9029 32970 9046 32978
rect 9080 32970 9095 32978
rect 9029 32958 9095 32970
rect 9187 38946 9253 38958
rect 9187 38938 9204 38946
rect 9238 38938 9253 38946
rect 9187 32970 9204 32978
rect 9238 32970 9253 32978
rect 9187 32958 9253 32970
rect 9345 38946 9411 38958
rect 9345 38938 9362 38946
rect 9396 38938 9411 38946
rect 9345 32970 9362 32978
rect 9396 32970 9411 32978
rect 9345 32958 9411 32970
rect 9503 38946 9569 38958
rect 9503 38938 9520 38946
rect 9554 38938 9569 38946
rect 9503 32970 9520 32978
rect 9554 32970 9569 32978
rect 9503 32958 9569 32970
rect 9661 38946 9727 38958
rect 9661 38938 9678 38946
rect 9712 38938 9727 38946
rect 9661 32970 9678 32978
rect 9712 32970 9727 32978
rect 9661 32958 9727 32970
rect 9819 38946 9885 38958
rect 9819 38938 9836 38946
rect 9870 38938 9885 38946
rect 9819 32970 9836 32978
rect 9870 32970 9885 32978
rect 9819 32958 9885 32970
rect 9977 38946 10043 38958
rect 9977 38938 9994 38946
rect 10028 38938 10043 38946
rect 9977 32970 9994 32978
rect 10028 32970 10043 32978
rect 9977 32958 10043 32970
rect 10135 38946 10201 38958
rect 10135 38938 10152 38946
rect 10186 38938 10201 38946
rect 10135 32970 10152 32978
rect 10186 32970 10201 32978
rect 10135 32958 10201 32970
rect 10293 38946 10359 38958
rect 10293 38938 10310 38946
rect 10344 38938 10359 38946
rect 10293 32970 10310 32978
rect 10344 32970 10359 32978
rect 10293 32958 10359 32970
rect 10451 38946 10517 38958
rect 10451 38938 10468 38946
rect 10502 38938 10517 38946
rect 10451 32970 10468 32978
rect 10502 32970 10517 32978
rect 10451 32958 10517 32970
rect 10609 38946 10675 38958
rect 10609 38938 10626 38946
rect 10660 38938 10675 38946
rect 10609 32970 10626 32978
rect 10660 32970 10675 32978
rect 10609 32958 10675 32970
rect 10767 38946 10833 38958
rect 10767 38938 10784 38946
rect 10818 38938 10833 38946
rect 10767 32970 10784 32978
rect 10818 32970 10833 32978
rect 10767 32958 10833 32970
rect 10925 38946 10991 38958
rect 10925 38938 10942 38946
rect 10976 38938 10991 38946
rect 10925 32970 10942 32978
rect 10976 32970 10991 32978
rect 10925 32958 10991 32970
rect 11083 38946 11149 38958
rect 11083 38938 11100 38946
rect 11134 38938 11149 38946
rect 11083 32970 11100 32978
rect 11134 32970 11149 32978
rect 11083 32958 11149 32970
rect 11241 38946 11307 38958
rect 11241 38938 11258 38946
rect 11292 38938 11307 38946
rect 11241 32970 11258 32978
rect 11292 32970 11307 32978
rect 11241 32958 11307 32970
rect 11399 38946 11465 38958
rect 11399 38938 11416 38946
rect 11450 38938 11465 38946
rect 11399 32970 11416 32978
rect 11450 32970 11465 32978
rect 11399 32958 11465 32970
rect 11557 38946 11623 38958
rect 11557 38938 11574 38946
rect 11608 38938 11623 38946
rect 11557 32970 11574 32978
rect 11608 32970 11623 32978
rect 11557 32958 11623 32970
rect 11715 38946 11781 38958
rect 11715 38938 11732 38946
rect 11766 38938 11781 38946
rect 11715 32970 11732 32978
rect 11766 32970 11781 32978
rect 11715 32958 11781 32970
rect 11873 38946 11939 38958
rect 11873 38938 11890 38946
rect 11924 38938 11939 38946
rect 11873 32970 11890 32978
rect 11924 32970 11939 32978
rect 11873 32958 11939 32970
rect 12031 38946 12097 38958
rect 12031 38938 12048 38946
rect 12082 38938 12097 38946
rect 12031 32970 12048 32978
rect 12082 32970 12097 32978
rect 12031 32958 12097 32970
rect 12189 38946 12255 38958
rect 12189 38938 12206 38946
rect 12240 38938 12255 38946
rect 12189 32970 12206 32978
rect 12240 32970 12255 32978
rect 12189 32958 12255 32970
rect 12347 38946 12413 38958
rect 12347 38938 12364 38946
rect 12398 38938 12413 38946
rect 12347 32970 12364 32978
rect 12398 32970 12413 32978
rect 12347 32958 12413 32970
rect 12505 38946 12571 38958
rect 12505 38938 12522 38946
rect 12556 38938 12571 38946
rect 12505 32970 12522 32978
rect 12556 32970 12571 32978
rect 12505 32958 12571 32970
rect 13930 39170 19010 39180
rect 13930 39132 14136 39170
rect 18859 39132 19010 39170
rect 13930 39122 19010 39132
rect 13930 39120 14000 39122
rect 18940 39120 19010 39122
rect 14132 39030 14152 39090
rect 18786 39030 18806 39090
rect 14132 38996 14144 39030
rect 18794 38996 18806 39030
rect 14132 38990 14152 38996
rect 18786 38990 18806 38996
rect 7832 32920 7852 32926
rect 12486 32920 12506 32926
rect 7832 32886 7844 32920
rect 12494 32886 12506 32920
rect 7832 32826 7852 32886
rect 12486 32826 12506 32886
rect 7630 32794 7700 32800
rect 12640 32794 12710 32800
rect 7630 32784 12710 32794
rect 7630 32746 7836 32784
rect 12502 32746 12710 32784
rect 7630 32730 12710 32746
rect 13000 32980 13500 33000
rect 13000 32910 13150 32980
rect 13350 32910 13500 32980
rect 13000 32900 13500 32910
rect 13000 32880 13120 32900
rect 13380 32880 13500 32900
rect 13000 32850 13100 32880
rect 7400 32620 7500 32650
rect 6500 32600 6620 32620
rect 6880 32600 7120 32620
rect 7380 32600 7500 32620
rect 6500 32590 7500 32600
rect 6500 32520 6650 32590
rect 6850 32520 7150 32590
rect 7350 32520 7500 32590
rect 6500 32500 7500 32520
rect 13000 32650 13020 32850
rect 13090 32650 13100 32850
rect 13000 32620 13100 32650
rect 13400 32850 13500 32880
rect 13400 32650 13410 32850
rect 13480 32650 13500 32850
rect 14065 38946 14131 38958
rect 14065 38938 14082 38946
rect 14116 38938 14131 38946
rect 14065 32970 14082 32978
rect 14116 32970 14131 32978
rect 14065 32958 14131 32970
rect 14223 38946 14289 38958
rect 14223 38938 14240 38946
rect 14274 38938 14289 38946
rect 14223 32970 14240 32978
rect 14274 32970 14289 32978
rect 14223 32958 14289 32970
rect 14381 38946 14447 38958
rect 14381 38938 14398 38946
rect 14432 38938 14447 38946
rect 14381 32970 14398 32978
rect 14432 32970 14447 32978
rect 14381 32958 14447 32970
rect 14539 38946 14605 38958
rect 14539 38938 14556 38946
rect 14590 38938 14605 38946
rect 14539 32970 14556 32978
rect 14590 32970 14605 32978
rect 14539 32958 14605 32970
rect 14697 38946 14763 38958
rect 14697 38938 14714 38946
rect 14748 38938 14763 38946
rect 14697 32970 14714 32978
rect 14748 32970 14763 32978
rect 14697 32958 14763 32970
rect 14855 38946 14921 38958
rect 14855 38938 14872 38946
rect 14906 38938 14921 38946
rect 14855 32970 14872 32978
rect 14906 32970 14921 32978
rect 14855 32958 14921 32970
rect 15013 38946 15079 38958
rect 15013 38938 15030 38946
rect 15064 38938 15079 38946
rect 15013 32970 15030 32978
rect 15064 32970 15079 32978
rect 15013 32958 15079 32970
rect 15171 38946 15237 38958
rect 15171 38938 15188 38946
rect 15222 38938 15237 38946
rect 15171 32970 15188 32978
rect 15222 32970 15237 32978
rect 15171 32958 15237 32970
rect 15329 38946 15395 38958
rect 15329 38938 15346 38946
rect 15380 38938 15395 38946
rect 15329 32970 15346 32978
rect 15380 32970 15395 32978
rect 15329 32958 15395 32970
rect 15487 38946 15553 38958
rect 15487 38938 15504 38946
rect 15538 38938 15553 38946
rect 15487 32970 15504 32978
rect 15538 32970 15553 32978
rect 15487 32958 15553 32970
rect 15645 38946 15711 38958
rect 15645 38938 15662 38946
rect 15696 38938 15711 38946
rect 15645 32970 15662 32978
rect 15696 32970 15711 32978
rect 15645 32958 15711 32970
rect 15803 38946 15869 38958
rect 15803 38938 15820 38946
rect 15854 38938 15869 38946
rect 15803 32970 15820 32978
rect 15854 32970 15869 32978
rect 15803 32958 15869 32970
rect 15961 38946 16027 38958
rect 15961 38938 15978 38946
rect 16012 38938 16027 38946
rect 15961 32970 15978 32978
rect 16012 32970 16027 32978
rect 15961 32958 16027 32970
rect 16119 38946 16185 38958
rect 16119 38938 16136 38946
rect 16170 38938 16185 38946
rect 16119 32970 16136 32978
rect 16170 32970 16185 32978
rect 16119 32958 16185 32970
rect 16277 38946 16343 38958
rect 16277 38938 16294 38946
rect 16328 38938 16343 38946
rect 16277 32970 16294 32978
rect 16328 32970 16343 32978
rect 16277 32958 16343 32970
rect 16435 38946 16501 38958
rect 16435 38938 16452 38946
rect 16486 38938 16501 38946
rect 16435 32970 16452 32978
rect 16486 32970 16501 32978
rect 16435 32958 16501 32970
rect 16593 38946 16659 38958
rect 16593 38938 16610 38946
rect 16644 38938 16659 38946
rect 16593 32970 16610 32978
rect 16644 32970 16659 32978
rect 16593 32958 16659 32970
rect 16751 38946 16817 38958
rect 16751 38938 16768 38946
rect 16802 38938 16817 38946
rect 16751 32970 16768 32978
rect 16802 32970 16817 32978
rect 16751 32958 16817 32970
rect 16909 38946 16975 38958
rect 16909 38938 16926 38946
rect 16960 38938 16975 38946
rect 16909 32970 16926 32978
rect 16960 32970 16975 32978
rect 16909 32958 16975 32970
rect 17067 38946 17133 38958
rect 17067 38938 17084 38946
rect 17118 38938 17133 38946
rect 17067 32970 17084 32978
rect 17118 32970 17133 32978
rect 17067 32958 17133 32970
rect 17225 38946 17291 38958
rect 17225 38938 17242 38946
rect 17276 38938 17291 38946
rect 17225 32970 17242 32978
rect 17276 32970 17291 32978
rect 17225 32958 17291 32970
rect 17383 38946 17449 38958
rect 17383 38938 17400 38946
rect 17434 38938 17449 38946
rect 17383 32970 17400 32978
rect 17434 32970 17449 32978
rect 17383 32958 17449 32970
rect 17541 38946 17607 38958
rect 17541 38938 17558 38946
rect 17592 38938 17607 38946
rect 17541 32970 17558 32978
rect 17592 32970 17607 32978
rect 17541 32958 17607 32970
rect 17699 38946 17765 38958
rect 17699 38938 17716 38946
rect 17750 38938 17765 38946
rect 17699 32970 17716 32978
rect 17750 32970 17765 32978
rect 17699 32958 17765 32970
rect 17857 38946 17923 38958
rect 17857 38938 17874 38946
rect 17908 38938 17923 38946
rect 17857 32970 17874 32978
rect 17908 32970 17923 32978
rect 17857 32958 17923 32970
rect 18015 38946 18081 38958
rect 18015 38938 18032 38946
rect 18066 38938 18081 38946
rect 18015 32970 18032 32978
rect 18066 32970 18081 32978
rect 18015 32958 18081 32970
rect 18173 38946 18239 38958
rect 18173 38938 18190 38946
rect 18224 38938 18239 38946
rect 18173 32970 18190 32978
rect 18224 32970 18239 32978
rect 18173 32958 18239 32970
rect 18331 38946 18397 38958
rect 18331 38938 18348 38946
rect 18382 38938 18397 38946
rect 18331 32970 18348 32978
rect 18382 32970 18397 32978
rect 18331 32958 18397 32970
rect 18489 38946 18555 38958
rect 18489 38938 18506 38946
rect 18540 38938 18555 38946
rect 18489 32970 18506 32978
rect 18540 32970 18555 32978
rect 18489 32958 18555 32970
rect 18647 38946 18713 38958
rect 18647 38938 18664 38946
rect 18698 38938 18713 38946
rect 18647 32970 18664 32978
rect 18698 32970 18713 32978
rect 18647 32958 18713 32970
rect 18805 38946 18871 38958
rect 18805 38938 18822 38946
rect 18856 38938 18871 38946
rect 18805 32970 18822 32978
rect 18856 32970 18871 32978
rect 18805 32958 18871 32970
rect 20230 39170 25520 39180
rect 20230 39132 20436 39170
rect 25159 39150 25520 39170
rect 25590 39150 25600 39350
rect 25159 39132 25600 39150
rect 20230 39122 25600 39132
rect 20230 39120 20300 39122
rect 25240 39120 25600 39122
rect 25900 39350 26100 39380
rect 25900 39150 25910 39350
rect 25980 39150 26020 39350
rect 26090 39150 26100 39350
rect 25900 39120 26100 39150
rect 26400 39350 26600 39380
rect 26400 39150 26410 39350
rect 26480 39150 26520 39350
rect 26590 39150 26600 39350
rect 26400 39120 26600 39150
rect 26900 39350 27100 39380
rect 26900 39150 26910 39350
rect 26980 39150 27020 39350
rect 27090 39150 27100 39350
rect 26900 39120 27100 39150
rect 27400 39350 27600 39380
rect 27400 39150 27410 39350
rect 27480 39150 27520 39350
rect 27590 39150 27600 39350
rect 27400 39120 27600 39150
rect 27900 39350 28100 39380
rect 27900 39150 27910 39350
rect 27980 39150 28020 39350
rect 28090 39150 28100 39350
rect 27900 39120 28100 39150
rect 28400 39350 28600 39380
rect 28400 39150 28410 39350
rect 28480 39150 28520 39350
rect 28590 39150 28600 39350
rect 28400 39120 28600 39150
rect 28900 39350 29100 39380
rect 28900 39150 28910 39350
rect 28980 39150 29020 39350
rect 29090 39150 29100 39350
rect 28900 39120 29100 39150
rect 29400 39350 29800 39380
rect 29400 39150 29410 39350
rect 29480 39150 29800 39350
rect 29400 39120 29800 39150
rect 20432 39030 20452 39090
rect 25086 39030 25106 39090
rect 20432 38996 20444 39030
rect 25094 38996 25106 39030
rect 20432 38990 20452 38996
rect 25086 38990 25106 38996
rect 14132 32920 14152 32926
rect 18786 32920 18806 32926
rect 14132 32886 14144 32920
rect 18794 32886 18806 32920
rect 14132 32826 14152 32886
rect 18786 32826 18806 32886
rect 13930 32794 14000 32800
rect 18940 32794 19010 32800
rect 13930 32784 19010 32794
rect 13930 32746 14136 32784
rect 18802 32746 19010 32784
rect 13930 32730 19010 32746
rect 19500 32980 20000 33000
rect 19500 32910 19650 32980
rect 19850 32910 20000 32980
rect 19500 32900 20000 32910
rect 19500 32880 19620 32900
rect 19880 32880 20000 32900
rect 19500 32850 19600 32880
rect 13400 32620 13500 32650
rect 13000 32600 13120 32620
rect 13380 32600 13500 32620
rect 13000 32590 13500 32600
rect 13000 32520 13150 32590
rect 13350 32520 13500 32590
rect 13000 32500 13500 32520
rect 19500 32650 19520 32850
rect 19590 32650 19600 32850
rect 19500 32620 19600 32650
rect 19900 32850 20000 32880
rect 19900 32650 19910 32850
rect 19980 32650 20000 32850
rect 25310 39100 25620 39120
rect 25880 39100 26120 39120
rect 26380 39100 26620 39120
rect 26880 39100 27120 39120
rect 27380 39100 27620 39120
rect 27880 39100 28120 39120
rect 28380 39100 28620 39120
rect 28880 39100 29120 39120
rect 29380 39100 29800 39120
rect 25310 39090 29800 39100
rect 25310 39020 25650 39090
rect 25850 39020 26150 39090
rect 26350 39020 26650 39090
rect 26850 39020 27150 39090
rect 27350 39020 27650 39090
rect 27850 39020 28150 39090
rect 28350 39020 28650 39090
rect 28850 39020 29150 39090
rect 29350 39020 29800 39090
rect 25310 39000 29800 39020
rect 25310 38980 26500 39000
rect 20365 38946 20431 38958
rect 20365 38938 20382 38946
rect 20416 38938 20431 38946
rect 20365 32970 20382 32978
rect 20416 32970 20431 32978
rect 20365 32958 20431 32970
rect 20523 38946 20589 38958
rect 20523 38938 20540 38946
rect 20574 38938 20589 38946
rect 20523 32970 20540 32978
rect 20574 32970 20589 32978
rect 20523 32958 20589 32970
rect 20681 38946 20747 38958
rect 20681 38938 20698 38946
rect 20732 38938 20747 38946
rect 20681 32970 20698 32978
rect 20732 32970 20747 32978
rect 20681 32958 20747 32970
rect 20839 38946 20905 38958
rect 20839 38938 20856 38946
rect 20890 38938 20905 38946
rect 20839 32970 20856 32978
rect 20890 32970 20905 32978
rect 20839 32958 20905 32970
rect 20997 38946 21063 38958
rect 20997 38938 21014 38946
rect 21048 38938 21063 38946
rect 20997 32970 21014 32978
rect 21048 32970 21063 32978
rect 20997 32958 21063 32970
rect 21155 38946 21221 38958
rect 21155 38938 21172 38946
rect 21206 38938 21221 38946
rect 21155 32970 21172 32978
rect 21206 32970 21221 32978
rect 21155 32958 21221 32970
rect 21313 38946 21379 38958
rect 21313 38938 21330 38946
rect 21364 38938 21379 38946
rect 21313 32970 21330 32978
rect 21364 32970 21379 32978
rect 21313 32958 21379 32970
rect 21471 38946 21537 38958
rect 21471 38938 21488 38946
rect 21522 38938 21537 38946
rect 21471 32970 21488 32978
rect 21522 32970 21537 32978
rect 21471 32958 21537 32970
rect 21629 38946 21695 38958
rect 21629 38938 21646 38946
rect 21680 38938 21695 38946
rect 21629 32970 21646 32978
rect 21680 32970 21695 32978
rect 21629 32958 21695 32970
rect 21787 38946 21853 38958
rect 21787 38938 21804 38946
rect 21838 38938 21853 38946
rect 21787 32970 21804 32978
rect 21838 32970 21853 32978
rect 21787 32958 21853 32970
rect 21945 38946 22011 38958
rect 21945 38938 21962 38946
rect 21996 38938 22011 38946
rect 21945 32970 21962 32978
rect 21996 32970 22011 32978
rect 21945 32958 22011 32970
rect 22103 38946 22169 38958
rect 22103 38938 22120 38946
rect 22154 38938 22169 38946
rect 22103 32970 22120 32978
rect 22154 32970 22169 32978
rect 22103 32958 22169 32970
rect 22261 38946 22327 38958
rect 22261 38938 22278 38946
rect 22312 38938 22327 38946
rect 22261 32970 22278 32978
rect 22312 32970 22327 32978
rect 22261 32958 22327 32970
rect 22419 38946 22485 38958
rect 22419 38938 22436 38946
rect 22470 38938 22485 38946
rect 22419 32970 22436 32978
rect 22470 32970 22485 32978
rect 22419 32958 22485 32970
rect 22577 38946 22643 38958
rect 22577 38938 22594 38946
rect 22628 38938 22643 38946
rect 22577 32970 22594 32978
rect 22628 32970 22643 32978
rect 22577 32958 22643 32970
rect 22735 38946 22801 38958
rect 22735 38938 22752 38946
rect 22786 38938 22801 38946
rect 22735 32970 22752 32978
rect 22786 32970 22801 32978
rect 22735 32958 22801 32970
rect 22893 38946 22959 38958
rect 22893 38938 22910 38946
rect 22944 38938 22959 38946
rect 22893 32970 22910 32978
rect 22944 32970 22959 32978
rect 22893 32958 22959 32970
rect 23051 38946 23117 38958
rect 23051 38938 23068 38946
rect 23102 38938 23117 38946
rect 23051 32970 23068 32978
rect 23102 32970 23117 32978
rect 23051 32958 23117 32970
rect 23209 38946 23275 38958
rect 23209 38938 23226 38946
rect 23260 38938 23275 38946
rect 23209 32970 23226 32978
rect 23260 32970 23275 32978
rect 23209 32958 23275 32970
rect 23367 38946 23433 38958
rect 23367 38938 23384 38946
rect 23418 38938 23433 38946
rect 23367 32970 23384 32978
rect 23418 32970 23433 32978
rect 23367 32958 23433 32970
rect 23525 38946 23591 38958
rect 23525 38938 23542 38946
rect 23576 38938 23591 38946
rect 23525 32970 23542 32978
rect 23576 32970 23591 32978
rect 23525 32958 23591 32970
rect 23683 38946 23749 38958
rect 23683 38938 23700 38946
rect 23734 38938 23749 38946
rect 23683 32970 23700 32978
rect 23734 32970 23749 32978
rect 23683 32958 23749 32970
rect 23841 38946 23907 38958
rect 23841 38938 23858 38946
rect 23892 38938 23907 38946
rect 23841 32970 23858 32978
rect 23892 32970 23907 32978
rect 23841 32958 23907 32970
rect 23999 38946 24065 38958
rect 23999 38938 24016 38946
rect 24050 38938 24065 38946
rect 23999 32970 24016 32978
rect 24050 32970 24065 32978
rect 23999 32958 24065 32970
rect 24157 38946 24223 38958
rect 24157 38938 24174 38946
rect 24208 38938 24223 38946
rect 24157 32970 24174 32978
rect 24208 32970 24223 32978
rect 24157 32958 24223 32970
rect 24315 38946 24381 38958
rect 24315 38938 24332 38946
rect 24366 38938 24381 38946
rect 24315 32970 24332 32978
rect 24366 32970 24381 32978
rect 24315 32958 24381 32970
rect 24473 38946 24539 38958
rect 24473 38938 24490 38946
rect 24524 38938 24539 38946
rect 24473 32970 24490 32978
rect 24524 32970 24539 32978
rect 24473 32958 24539 32970
rect 24631 38946 24697 38958
rect 24631 38938 24648 38946
rect 24682 38938 24697 38946
rect 24631 32970 24648 32978
rect 24682 32970 24697 32978
rect 24631 32958 24697 32970
rect 24789 38946 24855 38958
rect 24789 38938 24806 38946
rect 24840 38938 24855 38946
rect 24789 32970 24806 32978
rect 24840 32970 24855 32978
rect 24789 32958 24855 32970
rect 24947 38946 25013 38958
rect 24947 38938 24964 38946
rect 24998 38938 25013 38946
rect 24947 32970 24964 32978
rect 24998 32970 25013 32978
rect 24947 32958 25013 32970
rect 25105 38946 25171 38958
rect 25105 38938 25122 38946
rect 25156 38938 25171 38946
rect 25105 32970 25122 32978
rect 25156 32970 25171 32978
rect 25105 32958 25171 32970
rect 25310 38910 25650 38980
rect 25850 38910 26150 38980
rect 26350 38910 26500 38980
rect 25310 38900 26500 38910
rect 25310 38880 25620 38900
rect 25880 38880 26120 38900
rect 26380 38880 26500 38900
rect 25310 38850 25600 38880
rect 25310 38650 25520 38850
rect 25590 38650 25600 38850
rect 25310 38620 25600 38650
rect 25900 38850 26100 38880
rect 25900 38650 25910 38850
rect 25980 38650 26020 38850
rect 26090 38650 26100 38850
rect 25900 38620 26100 38650
rect 26400 38850 26500 38880
rect 26400 38650 26410 38850
rect 26480 38650 26500 38850
rect 29780 38720 29800 39000
rect 29840 38720 29860 40400
rect 29900 40190 29910 40450
rect 30090 40190 30100 40450
rect 29900 40180 30100 40190
rect 29780 38700 29860 38720
rect 29900 38910 30100 38920
rect 29900 38690 29910 38910
rect 30090 38690 30100 38910
rect 29900 38680 30100 38690
rect 26400 38620 26500 38650
rect 25310 38600 25620 38620
rect 25880 38600 26120 38620
rect 26380 38600 26500 38620
rect 25310 38590 26500 38600
rect 25310 38520 25650 38590
rect 25850 38520 26150 38590
rect 26350 38520 26500 38590
rect 25310 38480 26500 38520
rect 25310 38410 25650 38480
rect 25850 38410 26150 38480
rect 26350 38410 26500 38480
rect 25310 38400 26500 38410
rect 25310 38380 25620 38400
rect 25880 38380 26120 38400
rect 26380 38380 26500 38400
rect 25310 38350 25600 38380
rect 25310 38150 25520 38350
rect 25590 38150 25600 38350
rect 25310 38120 25600 38150
rect 25900 38350 26100 38380
rect 25900 38150 25910 38350
rect 25980 38150 26020 38350
rect 26090 38150 26100 38350
rect 25900 38120 26100 38150
rect 26400 38350 26500 38380
rect 26400 38150 26410 38350
rect 26480 38150 26500 38350
rect 26400 38120 26500 38150
rect 25310 38100 25620 38120
rect 25880 38100 26120 38120
rect 26380 38100 26500 38120
rect 25310 38090 26500 38100
rect 25310 38020 25650 38090
rect 25850 38020 26150 38090
rect 26350 38020 26500 38090
rect 25310 37980 26500 38020
rect 25310 37910 25650 37980
rect 25850 37910 26150 37980
rect 26350 37910 26500 37980
rect 25310 37900 26500 37910
rect 25310 37880 25620 37900
rect 25880 37880 26120 37900
rect 26380 37880 26500 37900
rect 25310 37850 25600 37880
rect 25310 37650 25520 37850
rect 25590 37650 25600 37850
rect 25310 37620 25600 37650
rect 25900 37850 26100 37880
rect 25900 37650 25910 37850
rect 25980 37650 26020 37850
rect 26090 37650 26100 37850
rect 25900 37620 26100 37650
rect 26400 37850 26500 37880
rect 26400 37650 26410 37850
rect 26480 37650 26500 37850
rect 26400 37620 26500 37650
rect 25310 37600 25620 37620
rect 25880 37600 26120 37620
rect 26380 37600 26500 37620
rect 25310 37590 26500 37600
rect 25310 37520 25650 37590
rect 25850 37520 26150 37590
rect 26350 37520 26500 37590
rect 25310 37480 26500 37520
rect 25310 37410 25650 37480
rect 25850 37410 26150 37480
rect 26350 37410 26500 37480
rect 25310 37400 26500 37410
rect 25310 37380 25620 37400
rect 25880 37380 26120 37400
rect 26380 37380 26500 37400
rect 25310 37350 25600 37380
rect 25310 37150 25520 37350
rect 25590 37150 25600 37350
rect 25310 37120 25600 37150
rect 25900 37350 26100 37380
rect 25900 37150 25910 37350
rect 25980 37150 26020 37350
rect 26090 37150 26100 37350
rect 25900 37120 26100 37150
rect 26400 37350 26500 37380
rect 26400 37150 26410 37350
rect 26480 37150 26500 37350
rect 26400 37120 26500 37150
rect 25310 37100 25620 37120
rect 25880 37100 26120 37120
rect 26380 37100 26500 37120
rect 25310 37090 26500 37100
rect 25310 37020 25650 37090
rect 25850 37020 26150 37090
rect 26350 37020 26500 37090
rect 25310 36980 26500 37020
rect 25310 36910 25650 36980
rect 25850 36910 26150 36980
rect 26350 36910 26500 36980
rect 25310 36900 26500 36910
rect 25310 36880 25620 36900
rect 25880 36880 26120 36900
rect 26380 36880 26500 36900
rect 25310 36850 25600 36880
rect 25310 36650 25520 36850
rect 25590 36650 25600 36850
rect 25310 36620 25600 36650
rect 25900 36850 26100 36880
rect 25900 36650 25910 36850
rect 25980 36650 26020 36850
rect 26090 36650 26100 36850
rect 25900 36620 26100 36650
rect 26400 36850 26500 36880
rect 26400 36650 26410 36850
rect 26480 36650 26500 36850
rect 26400 36620 26500 36650
rect 25310 36600 25620 36620
rect 25880 36600 26120 36620
rect 26380 36600 26500 36620
rect 25310 36590 26500 36600
rect 25310 36520 25650 36590
rect 25850 36520 26150 36590
rect 26350 36520 26500 36590
rect 25310 36480 26500 36520
rect 25310 36410 25650 36480
rect 25850 36410 26150 36480
rect 26350 36410 26500 36480
rect 25310 36400 26500 36410
rect 25310 36380 25620 36400
rect 25880 36380 26120 36400
rect 26380 36380 26500 36400
rect 25310 36350 25600 36380
rect 25310 36150 25520 36350
rect 25590 36150 25600 36350
rect 25310 36120 25600 36150
rect 25900 36350 26100 36380
rect 25900 36150 25910 36350
rect 25980 36150 26020 36350
rect 26090 36150 26100 36350
rect 25900 36120 26100 36150
rect 26400 36350 26500 36380
rect 26400 36150 26410 36350
rect 26480 36150 26500 36350
rect 26400 36120 26500 36150
rect 25310 36100 25620 36120
rect 25880 36100 26120 36120
rect 26380 36100 26500 36120
rect 25310 36090 26500 36100
rect 25310 36020 25650 36090
rect 25850 36020 26150 36090
rect 26350 36020 26500 36090
rect 25310 35980 26500 36020
rect 25310 35910 25650 35980
rect 25850 35910 26150 35980
rect 26350 35910 26500 35980
rect 25310 35900 26500 35910
rect 25310 35880 25620 35900
rect 25880 35880 26120 35900
rect 26380 35880 26500 35900
rect 25310 35850 25600 35880
rect 25310 35650 25520 35850
rect 25590 35650 25600 35850
rect 25310 35620 25600 35650
rect 25900 35850 26100 35880
rect 25900 35650 25910 35850
rect 25980 35650 26020 35850
rect 26090 35650 26100 35850
rect 25900 35620 26100 35650
rect 26400 35850 26500 35880
rect 26400 35650 26410 35850
rect 26480 35650 26500 35850
rect 26400 35620 26500 35650
rect 25310 35600 25620 35620
rect 25880 35600 26120 35620
rect 26380 35600 26500 35620
rect 25310 35590 26500 35600
rect 25310 35520 25650 35590
rect 25850 35520 26150 35590
rect 26350 35520 26500 35590
rect 25310 35480 26500 35520
rect 25310 35410 25650 35480
rect 25850 35410 26150 35480
rect 26350 35410 26500 35480
rect 25310 35400 26500 35410
rect 25310 35380 25620 35400
rect 25880 35380 26120 35400
rect 26380 35380 26500 35400
rect 25310 35350 25600 35380
rect 25310 35150 25520 35350
rect 25590 35150 25600 35350
rect 25310 35120 25600 35150
rect 25900 35350 26100 35380
rect 25900 35150 25910 35350
rect 25980 35150 26020 35350
rect 26090 35150 26100 35350
rect 25900 35120 26100 35150
rect 26400 35350 26500 35380
rect 26400 35150 26410 35350
rect 26480 35150 26500 35350
rect 26400 35120 26500 35150
rect 25310 35100 25620 35120
rect 25880 35100 26120 35120
rect 26380 35100 26500 35120
rect 25310 35090 26500 35100
rect 25310 35020 25650 35090
rect 25850 35020 26150 35090
rect 26350 35020 26500 35090
rect 25310 34980 26500 35020
rect 25310 34910 25650 34980
rect 25850 34910 26150 34980
rect 26350 34910 26500 34980
rect 25310 34900 26500 34910
rect 25310 34880 25620 34900
rect 25880 34880 26120 34900
rect 26380 34880 26500 34900
rect 25310 34850 25600 34880
rect 25310 34650 25520 34850
rect 25590 34650 25600 34850
rect 25310 34620 25600 34650
rect 25900 34850 26100 34880
rect 25900 34650 25910 34850
rect 25980 34650 26020 34850
rect 26090 34650 26100 34850
rect 25900 34620 26100 34650
rect 26400 34850 26500 34880
rect 26400 34650 26410 34850
rect 26480 34650 26500 34850
rect 26400 34620 26500 34650
rect 25310 34600 25620 34620
rect 25880 34600 26120 34620
rect 26380 34600 26500 34620
rect 25310 34590 26500 34600
rect 25310 34520 25650 34590
rect 25850 34520 26150 34590
rect 26350 34520 26500 34590
rect 25310 34480 26500 34520
rect 25310 34410 25650 34480
rect 25850 34410 26150 34480
rect 26350 34410 26500 34480
rect 25310 34400 26500 34410
rect 25310 34380 25620 34400
rect 25880 34380 26120 34400
rect 26380 34380 26500 34400
rect 25310 34350 25600 34380
rect 25310 34150 25520 34350
rect 25590 34150 25600 34350
rect 25310 34120 25600 34150
rect 25900 34350 26100 34380
rect 25900 34150 25910 34350
rect 25980 34150 26020 34350
rect 26090 34150 26100 34350
rect 25900 34120 26100 34150
rect 26400 34350 26500 34380
rect 26400 34150 26410 34350
rect 26480 34150 26500 34350
rect 26400 34120 26500 34150
rect 25310 34100 25620 34120
rect 25880 34100 26120 34120
rect 26380 34100 26500 34120
rect 25310 34090 26500 34100
rect 25310 34020 25650 34090
rect 25850 34020 26150 34090
rect 26350 34020 26500 34090
rect 25310 33980 26500 34020
rect 25310 33910 25650 33980
rect 25850 33910 26150 33980
rect 26350 33910 26500 33980
rect 25310 33900 26500 33910
rect 25310 33880 25620 33900
rect 25880 33880 26120 33900
rect 26380 33880 26500 33900
rect 25310 33850 25600 33880
rect 25310 33650 25520 33850
rect 25590 33650 25600 33850
rect 25310 33620 25600 33650
rect 25900 33850 26100 33880
rect 25900 33650 25910 33850
rect 25980 33650 26020 33850
rect 26090 33650 26100 33850
rect 25900 33620 26100 33650
rect 26400 33850 26500 33880
rect 26400 33650 26410 33850
rect 26480 33650 26500 33850
rect 26400 33620 26500 33650
rect 25310 33600 25620 33620
rect 25880 33600 26120 33620
rect 26380 33600 26500 33620
rect 25310 33590 26500 33600
rect 25310 33520 25650 33590
rect 25850 33520 26150 33590
rect 26350 33520 26500 33590
rect 25310 33480 26500 33520
rect 25310 33410 25650 33480
rect 25850 33410 26150 33480
rect 26350 33410 26500 33480
rect 25310 33400 26500 33410
rect 25310 33380 25620 33400
rect 25880 33380 26120 33400
rect 26380 33380 26500 33400
rect 25310 33350 25600 33380
rect 25310 33150 25520 33350
rect 25590 33150 25600 33350
rect 25310 33120 25600 33150
rect 25900 33350 26100 33380
rect 25900 33150 25910 33350
rect 25980 33150 26020 33350
rect 26090 33150 26100 33350
rect 25900 33120 26100 33150
rect 26400 33350 26500 33380
rect 26400 33150 26410 33350
rect 26480 33150 26500 33350
rect 26400 33120 26500 33150
rect 25310 33100 25620 33120
rect 25880 33100 26120 33120
rect 26380 33100 26500 33120
rect 25310 33090 26500 33100
rect 25310 33020 25650 33090
rect 25850 33020 26150 33090
rect 26350 33020 26500 33090
rect 25310 32980 26500 33020
rect 20432 32920 20452 32926
rect 25086 32920 25106 32926
rect 20432 32886 20444 32920
rect 25094 32886 25106 32920
rect 20432 32826 20452 32886
rect 25086 32826 25106 32886
rect 20230 32794 20300 32800
rect 25310 32910 25650 32980
rect 25850 32910 26150 32980
rect 26350 32910 26500 32980
rect 25310 32900 26500 32910
rect 25310 32880 25620 32900
rect 25880 32880 26120 32900
rect 26380 32880 26500 32900
rect 25310 32850 25600 32880
rect 25310 32800 25520 32850
rect 25240 32794 25520 32800
rect 20230 32784 25520 32794
rect 20230 32746 20436 32784
rect 25102 32746 25520 32784
rect 20230 32730 25520 32746
rect 19900 32620 20000 32650
rect 19500 32600 19620 32620
rect 19880 32600 20000 32620
rect 19500 32590 20000 32600
rect 19500 32520 19650 32590
rect 19850 32520 20000 32590
rect 19500 32500 20000 32520
rect 25260 32650 25520 32730
rect 25590 32650 25600 32850
rect 25260 32620 25600 32650
rect 25900 32850 26100 32880
rect 25900 32650 25910 32850
rect 25980 32650 26020 32850
rect 26090 32650 26100 32850
rect 25900 32620 26100 32650
rect 26400 32850 26500 32880
rect 26400 32650 26410 32850
rect 26480 32650 26500 32850
rect 26400 32620 26500 32650
rect 25260 32600 25620 32620
rect 25880 32600 26120 32620
rect 26380 32600 26500 32620
rect 25260 32590 26500 32600
rect 25260 32520 25650 32590
rect 25850 32520 26150 32590
rect 26350 32520 26500 32590
rect 25260 32500 26500 32520
rect 0 32480 26500 32500
rect 0 32410 150 32480
rect 350 32410 650 32480
rect 850 32410 1150 32480
rect 1350 32410 1650 32480
rect 1850 32410 2150 32480
rect 2350 32410 2650 32480
rect 2850 32410 3150 32480
rect 3350 32410 3650 32480
rect 3850 32410 4150 32480
rect 4350 32410 4650 32480
rect 4850 32410 5150 32480
rect 5350 32410 5650 32480
rect 5850 32410 6150 32480
rect 6350 32410 6650 32480
rect 6850 32410 7150 32480
rect 7350 32410 7650 32480
rect 7850 32410 8150 32480
rect 8350 32410 8650 32480
rect 8850 32410 9150 32480
rect 9350 32410 9650 32480
rect 9850 32410 10150 32480
rect 10350 32410 10650 32480
rect 10850 32410 11150 32480
rect 11350 32410 11650 32480
rect 11850 32410 12150 32480
rect 12350 32410 12650 32480
rect 12850 32410 13150 32480
rect 13350 32410 13650 32480
rect 13850 32410 14150 32480
rect 14350 32410 14650 32480
rect 14850 32410 15150 32480
rect 15350 32410 15650 32480
rect 15850 32410 16150 32480
rect 16350 32410 16650 32480
rect 16850 32410 17150 32480
rect 17350 32410 17650 32480
rect 17850 32410 18150 32480
rect 18350 32410 18650 32480
rect 18850 32410 19150 32480
rect 19350 32410 19650 32480
rect 19850 32410 20150 32480
rect 20350 32410 20650 32480
rect 20850 32410 21150 32480
rect 21350 32410 21650 32480
rect 21850 32410 22150 32480
rect 22350 32410 22650 32480
rect 22850 32410 23150 32480
rect 23350 32410 23650 32480
rect 23850 32410 24150 32480
rect 24350 32410 24650 32480
rect 24850 32410 25150 32480
rect 25350 32410 25650 32480
rect 25850 32410 26150 32480
rect 26350 32410 26500 32480
rect 0 32400 26500 32410
rect 0 32380 120 32400
rect 380 32380 620 32400
rect 880 32380 1120 32400
rect 1380 32380 1620 32400
rect 1880 32380 2120 32400
rect 2380 32380 2620 32400
rect 2880 32380 3120 32400
rect 3380 32380 3620 32400
rect 3880 32380 4120 32400
rect 4380 32380 4620 32400
rect 4880 32380 5120 32400
rect 5380 32380 5620 32400
rect 5880 32380 6120 32400
rect 6380 32380 6620 32400
rect 6880 32380 7120 32400
rect 7380 32380 7620 32400
rect 7880 32380 8120 32400
rect 8380 32380 8620 32400
rect 8880 32380 9120 32400
rect 9380 32380 9620 32400
rect 9880 32380 10120 32400
rect 10380 32380 10620 32400
rect 10880 32380 11120 32400
rect 11380 32380 11620 32400
rect 11880 32380 12120 32400
rect 12380 32380 12620 32400
rect 12880 32380 13120 32400
rect 13380 32380 13620 32400
rect 13880 32380 14120 32400
rect 14380 32380 14620 32400
rect 14880 32380 15120 32400
rect 15380 32380 15620 32400
rect 15880 32380 16120 32400
rect 16380 32380 16620 32400
rect 16880 32380 17120 32400
rect 17380 32380 17620 32400
rect 17880 32380 18120 32400
rect 18380 32380 18620 32400
rect 18880 32380 19120 32400
rect 19380 32380 19620 32400
rect 19880 32380 20120 32400
rect 20380 32380 20620 32400
rect 20880 32380 21120 32400
rect 21380 32380 21620 32400
rect 21880 32380 22120 32400
rect 22380 32380 22620 32400
rect 22880 32380 23120 32400
rect 23380 32380 23620 32400
rect 23880 32380 24120 32400
rect 24380 32380 24620 32400
rect 24880 32380 25120 32400
rect 25380 32380 25620 32400
rect 25880 32380 26120 32400
rect 26380 32380 26500 32400
rect 0 32350 100 32380
rect 0 32150 20 32350
rect 90 32150 100 32350
rect 0 32120 100 32150
rect 400 32350 600 32380
rect 400 32150 410 32350
rect 480 32150 520 32350
rect 590 32150 600 32350
rect 400 32120 600 32150
rect 900 32350 1100 32380
rect 900 32150 910 32350
rect 980 32150 1020 32350
rect 1090 32150 1100 32350
rect 900 32120 1100 32150
rect 1400 32350 1600 32380
rect 1400 32150 1410 32350
rect 1480 32150 1520 32350
rect 1590 32150 1600 32350
rect 1400 32120 1600 32150
rect 1900 32350 2100 32380
rect 1900 32150 1910 32350
rect 1980 32150 2020 32350
rect 2090 32150 2100 32350
rect 1900 32120 2100 32150
rect 2400 32350 2600 32380
rect 2400 32150 2410 32350
rect 2480 32150 2520 32350
rect 2590 32150 2600 32350
rect 2400 32120 2600 32150
rect 2900 32350 3100 32380
rect 2900 32150 2910 32350
rect 2980 32150 3020 32350
rect 3090 32150 3100 32350
rect 2900 32120 3100 32150
rect 3400 32350 3600 32380
rect 3400 32150 3410 32350
rect 3480 32150 3520 32350
rect 3590 32150 3600 32350
rect 3400 32120 3600 32150
rect 3900 32350 4100 32380
rect 3900 32150 3910 32350
rect 3980 32150 4020 32350
rect 4090 32150 4100 32350
rect 3900 32120 4100 32150
rect 4400 32350 4600 32380
rect 4400 32150 4410 32350
rect 4480 32150 4520 32350
rect 4590 32150 4600 32350
rect 4400 32120 4600 32150
rect 4900 32350 5100 32380
rect 4900 32150 4910 32350
rect 4980 32150 5020 32350
rect 5090 32150 5100 32350
rect 4900 32120 5100 32150
rect 5400 32350 5600 32380
rect 5400 32150 5410 32350
rect 5480 32150 5520 32350
rect 5590 32150 5600 32350
rect 5400 32120 5600 32150
rect 5900 32350 6100 32380
rect 5900 32150 5910 32350
rect 5980 32150 6020 32350
rect 6090 32150 6100 32350
rect 5900 32120 6100 32150
rect 6400 32350 6600 32380
rect 6400 32150 6410 32350
rect 6480 32150 6520 32350
rect 6590 32150 6600 32350
rect 6400 32120 6600 32150
rect 6900 32350 7100 32380
rect 6900 32150 6910 32350
rect 6980 32150 7020 32350
rect 7090 32150 7100 32350
rect 6900 32120 7100 32150
rect 7400 32350 7600 32380
rect 7400 32150 7410 32350
rect 7480 32150 7520 32350
rect 7590 32150 7600 32350
rect 7400 32120 7600 32150
rect 7900 32350 8100 32380
rect 7900 32150 7910 32350
rect 7980 32150 8020 32350
rect 8090 32150 8100 32350
rect 7900 32120 8100 32150
rect 8400 32350 8600 32380
rect 8400 32150 8410 32350
rect 8480 32150 8520 32350
rect 8590 32150 8600 32350
rect 8400 32120 8600 32150
rect 8900 32350 9100 32380
rect 8900 32150 8910 32350
rect 8980 32150 9020 32350
rect 9090 32150 9100 32350
rect 8900 32120 9100 32150
rect 9400 32350 9600 32380
rect 9400 32150 9410 32350
rect 9480 32150 9520 32350
rect 9590 32150 9600 32350
rect 9400 32120 9600 32150
rect 9900 32350 10100 32380
rect 9900 32150 9910 32350
rect 9980 32150 10020 32350
rect 10090 32150 10100 32350
rect 9900 32120 10100 32150
rect 10400 32350 10600 32380
rect 10400 32150 10410 32350
rect 10480 32150 10520 32350
rect 10590 32150 10600 32350
rect 10400 32120 10600 32150
rect 10900 32350 11100 32380
rect 10900 32150 10910 32350
rect 10980 32150 11020 32350
rect 11090 32150 11100 32350
rect 10900 32120 11100 32150
rect 11400 32350 11600 32380
rect 11400 32150 11410 32350
rect 11480 32150 11520 32350
rect 11590 32150 11600 32350
rect 11400 32120 11600 32150
rect 11900 32350 12100 32380
rect 11900 32150 11910 32350
rect 11980 32150 12020 32350
rect 12090 32150 12100 32350
rect 11900 32120 12100 32150
rect 12400 32350 12600 32380
rect 12400 32150 12410 32350
rect 12480 32150 12520 32350
rect 12590 32150 12600 32350
rect 12400 32120 12600 32150
rect 12900 32350 13100 32380
rect 12900 32150 12910 32350
rect 12980 32150 13020 32350
rect 13090 32150 13100 32350
rect 12900 32120 13100 32150
rect 13400 32350 13600 32380
rect 13400 32150 13410 32350
rect 13480 32150 13520 32350
rect 13590 32150 13600 32350
rect 13400 32120 13600 32150
rect 13900 32350 14100 32380
rect 13900 32150 13910 32350
rect 13980 32150 14020 32350
rect 14090 32150 14100 32350
rect 13900 32120 14100 32150
rect 14400 32350 14600 32380
rect 14400 32150 14410 32350
rect 14480 32150 14520 32350
rect 14590 32150 14600 32350
rect 14400 32120 14600 32150
rect 14900 32350 15100 32380
rect 14900 32150 14910 32350
rect 14980 32150 15020 32350
rect 15090 32150 15100 32350
rect 14900 32120 15100 32150
rect 15400 32350 15600 32380
rect 15400 32150 15410 32350
rect 15480 32150 15520 32350
rect 15590 32150 15600 32350
rect 15400 32120 15600 32150
rect 15900 32350 16100 32380
rect 15900 32150 15910 32350
rect 15980 32150 16020 32350
rect 16090 32150 16100 32350
rect 15900 32120 16100 32150
rect 16400 32350 16600 32380
rect 16400 32150 16410 32350
rect 16480 32150 16520 32350
rect 16590 32150 16600 32350
rect 16400 32120 16600 32150
rect 16900 32350 17100 32380
rect 16900 32150 16910 32350
rect 16980 32150 17020 32350
rect 17090 32150 17100 32350
rect 16900 32120 17100 32150
rect 17400 32350 17600 32380
rect 17400 32150 17410 32350
rect 17480 32150 17520 32350
rect 17590 32150 17600 32350
rect 17400 32120 17600 32150
rect 17900 32350 18100 32380
rect 17900 32150 17910 32350
rect 17980 32150 18020 32350
rect 18090 32150 18100 32350
rect 17900 32120 18100 32150
rect 18400 32350 18600 32380
rect 18400 32150 18410 32350
rect 18480 32150 18520 32350
rect 18590 32150 18600 32350
rect 18400 32120 18600 32150
rect 18900 32350 19100 32380
rect 18900 32150 18910 32350
rect 18980 32150 19020 32350
rect 19090 32150 19100 32350
rect 18900 32120 19100 32150
rect 19400 32350 19600 32380
rect 19400 32150 19410 32350
rect 19480 32150 19520 32350
rect 19590 32150 19600 32350
rect 19400 32120 19600 32150
rect 19900 32350 20100 32380
rect 19900 32150 19910 32350
rect 19980 32150 20020 32350
rect 20090 32150 20100 32350
rect 19900 32120 20100 32150
rect 20400 32350 20600 32380
rect 20400 32150 20410 32350
rect 20480 32150 20520 32350
rect 20590 32150 20600 32350
rect 20400 32120 20600 32150
rect 20900 32350 21100 32380
rect 20900 32150 20910 32350
rect 20980 32150 21020 32350
rect 21090 32150 21100 32350
rect 20900 32120 21100 32150
rect 21400 32350 21600 32380
rect 21400 32150 21410 32350
rect 21480 32150 21520 32350
rect 21590 32150 21600 32350
rect 21400 32120 21600 32150
rect 21900 32350 22100 32380
rect 21900 32150 21910 32350
rect 21980 32150 22020 32350
rect 22090 32150 22100 32350
rect 21900 32120 22100 32150
rect 22400 32350 22600 32380
rect 22400 32150 22410 32350
rect 22480 32150 22520 32350
rect 22590 32150 22600 32350
rect 22400 32120 22600 32150
rect 22900 32350 23100 32380
rect 22900 32150 22910 32350
rect 22980 32150 23020 32350
rect 23090 32150 23100 32350
rect 22900 32120 23100 32150
rect 23400 32350 23600 32380
rect 23400 32150 23410 32350
rect 23480 32150 23520 32350
rect 23590 32150 23600 32350
rect 23400 32120 23600 32150
rect 23900 32350 24100 32380
rect 23900 32150 23910 32350
rect 23980 32150 24020 32350
rect 24090 32150 24100 32350
rect 23900 32120 24100 32150
rect 24400 32350 24600 32380
rect 24400 32150 24410 32350
rect 24480 32150 24520 32350
rect 24590 32150 24600 32350
rect 24400 32120 24600 32150
rect 24900 32350 25100 32380
rect 24900 32150 24910 32350
rect 24980 32150 25020 32350
rect 25090 32150 25100 32350
rect 24900 32120 25100 32150
rect 25400 32350 25600 32380
rect 25400 32150 25410 32350
rect 25480 32150 25520 32350
rect 25590 32150 25600 32350
rect 25400 32120 25600 32150
rect 25900 32350 26100 32380
rect 25900 32150 25910 32350
rect 25980 32150 26020 32350
rect 26090 32150 26100 32350
rect 25900 32120 26100 32150
rect 26400 32350 26500 32380
rect 26400 32150 26410 32350
rect 26480 32150 26500 32350
rect 26400 32120 26500 32150
rect 0 32100 120 32120
rect 380 32100 620 32120
rect 880 32100 1120 32120
rect 1380 32100 1620 32120
rect 1880 32100 2120 32120
rect 2380 32100 2620 32120
rect 2880 32100 3120 32120
rect 3380 32100 3620 32120
rect 3880 32100 4120 32120
rect 4380 32100 4620 32120
rect 4880 32100 5120 32120
rect 5380 32100 5620 32120
rect 5880 32100 6120 32120
rect 6380 32100 6620 32120
rect 6880 32100 7120 32120
rect 7380 32100 7620 32120
rect 7880 32100 8120 32120
rect 8380 32100 8620 32120
rect 8880 32100 9120 32120
rect 9380 32100 9620 32120
rect 9880 32100 10120 32120
rect 10380 32100 10620 32120
rect 10880 32100 11120 32120
rect 11380 32100 11620 32120
rect 11880 32100 12120 32120
rect 12380 32100 12620 32120
rect 12880 32100 13120 32120
rect 13380 32100 13620 32120
rect 13880 32100 14120 32120
rect 14380 32100 14620 32120
rect 14880 32100 15120 32120
rect 15380 32100 15620 32120
rect 15880 32100 16120 32120
rect 16380 32100 16620 32120
rect 16880 32100 17120 32120
rect 17380 32100 17620 32120
rect 17880 32100 18120 32120
rect 18380 32100 18620 32120
rect 18880 32100 19120 32120
rect 19380 32100 19620 32120
rect 19880 32100 20120 32120
rect 20380 32100 20620 32120
rect 20880 32100 21120 32120
rect 21380 32100 21620 32120
rect 21880 32100 22120 32120
rect 22380 32100 22620 32120
rect 22880 32100 23120 32120
rect 23380 32100 23620 32120
rect 23880 32100 24120 32120
rect 24380 32100 24620 32120
rect 24880 32100 25120 32120
rect 25380 32100 25620 32120
rect 25880 32100 26120 32120
rect 26380 32100 26500 32120
rect 0 32090 26500 32100
rect 0 32020 150 32090
rect 350 32020 650 32090
rect 850 32020 1150 32090
rect 1350 32020 1650 32090
rect 1850 32020 2150 32090
rect 2350 32020 2650 32090
rect 2850 32020 3150 32090
rect 3350 32020 3650 32090
rect 3850 32020 4150 32090
rect 4350 32020 4650 32090
rect 4850 32020 5150 32090
rect 5350 32020 5650 32090
rect 5850 32020 6150 32090
rect 6350 32020 6650 32090
rect 6850 32020 7150 32090
rect 7350 32020 7650 32090
rect 7850 32020 8150 32090
rect 8350 32020 8650 32090
rect 8850 32020 9150 32090
rect 9350 32020 9650 32090
rect 9850 32020 10150 32090
rect 10350 32020 10650 32090
rect 10850 32020 11150 32090
rect 11350 32020 11650 32090
rect 11850 32020 12150 32090
rect 12350 32020 12650 32090
rect 12850 32020 13150 32090
rect 13350 32020 13650 32090
rect 13850 32020 14150 32090
rect 14350 32020 14650 32090
rect 14850 32020 15150 32090
rect 15350 32020 15650 32090
rect 15850 32020 16150 32090
rect 16350 32020 16650 32090
rect 16850 32020 17150 32090
rect 17350 32020 17650 32090
rect 17850 32020 18150 32090
rect 18350 32020 18650 32090
rect 18850 32020 19150 32090
rect 19350 32020 19650 32090
rect 19850 32020 20150 32090
rect 20350 32020 20650 32090
rect 20850 32020 21150 32090
rect 21350 32020 21650 32090
rect 21850 32020 22150 32090
rect 22350 32020 22650 32090
rect 22850 32020 23150 32090
rect 23350 32020 23650 32090
rect 23850 32020 24150 32090
rect 24350 32020 24650 32090
rect 24850 32020 25150 32090
rect 25350 32020 25650 32090
rect 25850 32020 26150 32090
rect 26350 32020 26500 32090
rect 0 31980 26500 32020
rect 0 31910 150 31980
rect 350 31910 650 31980
rect 850 31910 1150 31980
rect 1350 31910 1650 31980
rect 1850 31910 2150 31980
rect 2350 31910 2650 31980
rect 2850 31910 3150 31980
rect 3350 31910 3650 31980
rect 3850 31910 4150 31980
rect 4350 31910 4650 31980
rect 4850 31910 5150 31980
rect 5350 31910 5650 31980
rect 5850 31910 6150 31980
rect 6350 31910 6650 31980
rect 6850 31910 7150 31980
rect 7350 31910 7650 31980
rect 7850 31910 8150 31980
rect 8350 31910 8650 31980
rect 8850 31910 9150 31980
rect 9350 31910 9650 31980
rect 9850 31910 10150 31980
rect 10350 31910 10650 31980
rect 10850 31910 11150 31980
rect 11350 31910 11650 31980
rect 11850 31910 12150 31980
rect 12350 31910 12650 31980
rect 12850 31910 13150 31980
rect 13350 31910 13650 31980
rect 13850 31910 14150 31980
rect 14350 31910 14650 31980
rect 14850 31910 15150 31980
rect 15350 31910 15650 31980
rect 15850 31910 16150 31980
rect 16350 31910 16650 31980
rect 16850 31910 17150 31980
rect 17350 31910 17650 31980
rect 17850 31910 18150 31980
rect 18350 31910 18650 31980
rect 18850 31910 19150 31980
rect 19350 31910 19650 31980
rect 19850 31910 20150 31980
rect 20350 31910 20650 31980
rect 20850 31910 21150 31980
rect 21350 31910 21650 31980
rect 21850 31910 22150 31980
rect 22350 31910 22650 31980
rect 22850 31910 23150 31980
rect 23350 31910 23650 31980
rect 23850 31910 24150 31980
rect 24350 31910 24650 31980
rect 24850 31910 25150 31980
rect 25350 31910 25650 31980
rect 25850 31910 26150 31980
rect 26350 31910 26500 31980
rect 0 31900 26500 31910
rect 0 31880 120 31900
rect 380 31880 620 31900
rect 880 31880 1120 31900
rect 1380 31880 1620 31900
rect 1880 31880 2120 31900
rect 2380 31880 2620 31900
rect 2880 31880 3120 31900
rect 3380 31880 3620 31900
rect 3880 31880 4120 31900
rect 4380 31880 4620 31900
rect 4880 31880 5120 31900
rect 5380 31880 5620 31900
rect 5880 31880 6120 31900
rect 6380 31880 6620 31900
rect 6880 31880 7120 31900
rect 7380 31880 7620 31900
rect 7880 31880 8120 31900
rect 8380 31880 8620 31900
rect 8880 31880 9120 31900
rect 9380 31880 9620 31900
rect 9880 31880 10120 31900
rect 10380 31880 10620 31900
rect 10880 31880 11120 31900
rect 11380 31880 11620 31900
rect 11880 31880 12120 31900
rect 12380 31880 12620 31900
rect 12880 31880 13120 31900
rect 13380 31880 13620 31900
rect 13880 31880 14120 31900
rect 14380 31880 14620 31900
rect 14880 31880 15120 31900
rect 15380 31880 15620 31900
rect 15880 31880 16120 31900
rect 16380 31880 16620 31900
rect 16880 31880 17120 31900
rect 17380 31880 17620 31900
rect 17880 31880 18120 31900
rect 18380 31880 18620 31900
rect 18880 31880 19120 31900
rect 19380 31880 19620 31900
rect 19880 31880 20120 31900
rect 20380 31880 20620 31900
rect 20880 31880 21120 31900
rect 21380 31880 21620 31900
rect 21880 31880 22120 31900
rect 22380 31880 22620 31900
rect 22880 31880 23120 31900
rect 23380 31880 23620 31900
rect 23880 31880 24120 31900
rect 24380 31880 24620 31900
rect 24880 31880 25120 31900
rect 25380 31880 25620 31900
rect 25880 31880 26120 31900
rect 26380 31880 26500 31900
rect 0 31850 100 31880
rect 0 31650 20 31850
rect 90 31650 100 31850
rect 0 31620 100 31650
rect 400 31850 600 31880
rect 400 31650 410 31850
rect 480 31650 520 31850
rect 590 31650 600 31850
rect 400 31620 600 31650
rect 900 31850 1100 31880
rect 900 31650 910 31850
rect 980 31650 1020 31850
rect 1090 31650 1100 31850
rect 900 31620 1100 31650
rect 1400 31850 1600 31880
rect 1400 31650 1410 31850
rect 1480 31650 1520 31850
rect 1590 31650 1600 31850
rect 1400 31620 1600 31650
rect 1900 31850 2100 31880
rect 1900 31650 1910 31850
rect 1980 31650 2020 31850
rect 2090 31650 2100 31850
rect 1900 31620 2100 31650
rect 2400 31850 2600 31880
rect 2400 31650 2410 31850
rect 2480 31650 2520 31850
rect 2590 31650 2600 31850
rect 2400 31620 2600 31650
rect 2900 31850 3100 31880
rect 2900 31650 2910 31850
rect 2980 31650 3020 31850
rect 3090 31650 3100 31850
rect 2900 31620 3100 31650
rect 3400 31850 3600 31880
rect 3400 31650 3410 31850
rect 3480 31650 3520 31850
rect 3590 31650 3600 31850
rect 3400 31620 3600 31650
rect 3900 31850 4100 31880
rect 3900 31650 3910 31850
rect 3980 31650 4020 31850
rect 4090 31650 4100 31850
rect 3900 31620 4100 31650
rect 4400 31850 4600 31880
rect 4400 31650 4410 31850
rect 4480 31650 4520 31850
rect 4590 31650 4600 31850
rect 4400 31620 4600 31650
rect 4900 31850 5100 31880
rect 4900 31650 4910 31850
rect 4980 31650 5020 31850
rect 5090 31650 5100 31850
rect 4900 31620 5100 31650
rect 5400 31850 5600 31880
rect 5400 31650 5410 31850
rect 5480 31650 5520 31850
rect 5590 31650 5600 31850
rect 5400 31620 5600 31650
rect 5900 31850 6100 31880
rect 5900 31650 5910 31850
rect 5980 31650 6020 31850
rect 6090 31650 6100 31850
rect 5900 31620 6100 31650
rect 6400 31850 6600 31880
rect 6400 31650 6410 31850
rect 6480 31650 6520 31850
rect 6590 31650 6600 31850
rect 6400 31620 6600 31650
rect 6900 31850 7100 31880
rect 6900 31650 6910 31850
rect 6980 31650 7020 31850
rect 7090 31650 7100 31850
rect 6900 31620 7100 31650
rect 7400 31850 7600 31880
rect 7400 31650 7410 31850
rect 7480 31650 7520 31850
rect 7590 31650 7600 31850
rect 7400 31620 7600 31650
rect 7900 31850 8100 31880
rect 7900 31650 7910 31850
rect 7980 31650 8020 31850
rect 8090 31650 8100 31850
rect 7900 31620 8100 31650
rect 8400 31850 8600 31880
rect 8400 31650 8410 31850
rect 8480 31650 8520 31850
rect 8590 31650 8600 31850
rect 8400 31620 8600 31650
rect 8900 31850 9100 31880
rect 8900 31650 8910 31850
rect 8980 31650 9020 31850
rect 9090 31650 9100 31850
rect 8900 31620 9100 31650
rect 9400 31850 9600 31880
rect 9400 31650 9410 31850
rect 9480 31650 9520 31850
rect 9590 31650 9600 31850
rect 9400 31620 9600 31650
rect 9900 31850 10100 31880
rect 9900 31650 9910 31850
rect 9980 31650 10020 31850
rect 10090 31650 10100 31850
rect 9900 31620 10100 31650
rect 10400 31850 10600 31880
rect 10400 31650 10410 31850
rect 10480 31650 10520 31850
rect 10590 31650 10600 31850
rect 10400 31620 10600 31650
rect 10900 31850 11100 31880
rect 10900 31650 10910 31850
rect 10980 31650 11020 31850
rect 11090 31650 11100 31850
rect 10900 31620 11100 31650
rect 11400 31850 11600 31880
rect 11400 31650 11410 31850
rect 11480 31650 11520 31850
rect 11590 31650 11600 31850
rect 11400 31620 11600 31650
rect 11900 31850 12100 31880
rect 11900 31650 11910 31850
rect 11980 31650 12020 31850
rect 12090 31650 12100 31850
rect 11900 31620 12100 31650
rect 12400 31850 12600 31880
rect 12400 31650 12410 31850
rect 12480 31650 12520 31850
rect 12590 31650 12600 31850
rect 12400 31620 12600 31650
rect 12900 31850 13100 31880
rect 12900 31650 12910 31850
rect 12980 31650 13020 31850
rect 13090 31650 13100 31850
rect 12900 31620 13100 31650
rect 13400 31850 13600 31880
rect 13400 31650 13410 31850
rect 13480 31650 13520 31850
rect 13590 31650 13600 31850
rect 13400 31620 13600 31650
rect 13900 31850 14100 31880
rect 13900 31650 13910 31850
rect 13980 31650 14020 31850
rect 14090 31650 14100 31850
rect 13900 31620 14100 31650
rect 14400 31850 14600 31880
rect 14400 31650 14410 31850
rect 14480 31650 14520 31850
rect 14590 31650 14600 31850
rect 14400 31620 14600 31650
rect 14900 31850 15100 31880
rect 14900 31650 14910 31850
rect 14980 31650 15020 31850
rect 15090 31650 15100 31850
rect 14900 31620 15100 31650
rect 15400 31850 15600 31880
rect 15400 31650 15410 31850
rect 15480 31650 15520 31850
rect 15590 31650 15600 31850
rect 15400 31620 15600 31650
rect 15900 31850 16100 31880
rect 15900 31650 15910 31850
rect 15980 31650 16020 31850
rect 16090 31650 16100 31850
rect 15900 31620 16100 31650
rect 16400 31850 16600 31880
rect 16400 31650 16410 31850
rect 16480 31650 16520 31850
rect 16590 31650 16600 31850
rect 16400 31620 16600 31650
rect 16900 31850 17100 31880
rect 16900 31650 16910 31850
rect 16980 31650 17020 31850
rect 17090 31650 17100 31850
rect 16900 31620 17100 31650
rect 17400 31850 17600 31880
rect 17400 31650 17410 31850
rect 17480 31650 17520 31850
rect 17590 31650 17600 31850
rect 17400 31620 17600 31650
rect 17900 31850 18100 31880
rect 17900 31650 17910 31850
rect 17980 31650 18020 31850
rect 18090 31650 18100 31850
rect 17900 31620 18100 31650
rect 18400 31850 18600 31880
rect 18400 31650 18410 31850
rect 18480 31650 18520 31850
rect 18590 31650 18600 31850
rect 18400 31620 18600 31650
rect 18900 31850 19100 31880
rect 18900 31650 18910 31850
rect 18980 31650 19020 31850
rect 19090 31650 19100 31850
rect 18900 31620 19100 31650
rect 19400 31850 19600 31880
rect 19400 31650 19410 31850
rect 19480 31650 19520 31850
rect 19590 31650 19600 31850
rect 19400 31620 19600 31650
rect 19900 31850 20100 31880
rect 19900 31650 19910 31850
rect 19980 31650 20020 31850
rect 20090 31650 20100 31850
rect 19900 31620 20100 31650
rect 20400 31850 20600 31880
rect 20400 31650 20410 31850
rect 20480 31650 20520 31850
rect 20590 31650 20600 31850
rect 20400 31620 20600 31650
rect 20900 31850 21100 31880
rect 20900 31650 20910 31850
rect 20980 31650 21020 31850
rect 21090 31650 21100 31850
rect 20900 31620 21100 31650
rect 21400 31850 21600 31880
rect 21400 31650 21410 31850
rect 21480 31650 21520 31850
rect 21590 31650 21600 31850
rect 21400 31620 21600 31650
rect 21900 31850 22100 31880
rect 21900 31650 21910 31850
rect 21980 31650 22020 31850
rect 22090 31650 22100 31850
rect 21900 31620 22100 31650
rect 22400 31850 22600 31880
rect 22400 31650 22410 31850
rect 22480 31650 22520 31850
rect 22590 31650 22600 31850
rect 22400 31620 22600 31650
rect 22900 31850 23100 31880
rect 22900 31650 22910 31850
rect 22980 31650 23020 31850
rect 23090 31650 23100 31850
rect 22900 31620 23100 31650
rect 23400 31850 23600 31880
rect 23400 31650 23410 31850
rect 23480 31650 23520 31850
rect 23590 31650 23600 31850
rect 23400 31620 23600 31650
rect 23900 31850 24100 31880
rect 23900 31650 23910 31850
rect 23980 31650 24020 31850
rect 24090 31650 24100 31850
rect 23900 31620 24100 31650
rect 24400 31850 24600 31880
rect 24400 31650 24410 31850
rect 24480 31650 24520 31850
rect 24590 31650 24600 31850
rect 24400 31620 24600 31650
rect 24900 31850 25100 31880
rect 24900 31650 24910 31850
rect 24980 31650 25020 31850
rect 25090 31650 25100 31850
rect 24900 31620 25100 31650
rect 25400 31850 25600 31880
rect 25400 31650 25410 31850
rect 25480 31650 25520 31850
rect 25590 31650 25600 31850
rect 25400 31620 25600 31650
rect 25900 31850 26100 31880
rect 25900 31650 25910 31850
rect 25980 31650 26020 31850
rect 26090 31650 26100 31850
rect 25900 31620 26100 31650
rect 26400 31850 26500 31880
rect 26400 31650 26410 31850
rect 26480 31650 26500 31850
rect 26400 31620 26500 31650
rect 0 31600 120 31620
rect 380 31600 620 31620
rect 880 31600 1120 31620
rect 1380 31600 1620 31620
rect 1880 31600 2120 31620
rect 2380 31600 2620 31620
rect 2880 31600 3120 31620
rect 3380 31600 3620 31620
rect 3880 31600 4120 31620
rect 4380 31600 4620 31620
rect 4880 31600 5120 31620
rect 5380 31600 5620 31620
rect 5880 31600 6120 31620
rect 6380 31600 6620 31620
rect 6880 31600 7120 31620
rect 7380 31600 7620 31620
rect 7880 31600 8120 31620
rect 8380 31600 8620 31620
rect 8880 31600 9120 31620
rect 9380 31600 9620 31620
rect 9880 31600 10120 31620
rect 10380 31600 10620 31620
rect 10880 31600 11120 31620
rect 11380 31600 11620 31620
rect 11880 31600 12120 31620
rect 12380 31600 12620 31620
rect 12880 31600 13120 31620
rect 13380 31600 13620 31620
rect 13880 31600 14120 31620
rect 14380 31600 14620 31620
rect 14880 31600 15120 31620
rect 15380 31600 15620 31620
rect 15880 31600 16120 31620
rect 16380 31600 16620 31620
rect 16880 31600 17120 31620
rect 17380 31600 17620 31620
rect 17880 31600 18120 31620
rect 18380 31600 18620 31620
rect 18880 31600 19120 31620
rect 19380 31600 19620 31620
rect 19880 31600 20120 31620
rect 20380 31600 20620 31620
rect 20880 31600 21120 31620
rect 21380 31600 21620 31620
rect 21880 31600 22120 31620
rect 22380 31600 22620 31620
rect 22880 31600 23120 31620
rect 23380 31600 23620 31620
rect 23880 31600 24120 31620
rect 24380 31600 24620 31620
rect 24880 31600 25120 31620
rect 25380 31600 25620 31620
rect 25880 31600 26120 31620
rect 26380 31600 26500 31620
rect 0 31590 26500 31600
rect 0 31520 150 31590
rect 350 31520 650 31590
rect 850 31520 1150 31590
rect 1350 31520 1650 31590
rect 1850 31520 2150 31590
rect 2350 31520 2650 31590
rect 2850 31520 3150 31590
rect 3350 31520 3650 31590
rect 3850 31520 4150 31590
rect 4350 31520 4650 31590
rect 4850 31520 5150 31590
rect 5350 31520 5650 31590
rect 5850 31520 6150 31590
rect 6350 31520 6650 31590
rect 6850 31520 7150 31590
rect 7350 31520 7650 31590
rect 7850 31520 8150 31590
rect 8350 31520 8650 31590
rect 8850 31520 9150 31590
rect 9350 31520 9650 31590
rect 9850 31520 10150 31590
rect 10350 31520 10650 31590
rect 10850 31520 11150 31590
rect 11350 31520 11650 31590
rect 11850 31520 12150 31590
rect 12350 31520 12650 31590
rect 12850 31520 13150 31590
rect 13350 31520 13650 31590
rect 13850 31520 14150 31590
rect 14350 31520 14650 31590
rect 14850 31520 15150 31590
rect 15350 31520 15650 31590
rect 15850 31520 16150 31590
rect 16350 31520 16650 31590
rect 16850 31520 17150 31590
rect 17350 31520 17650 31590
rect 17850 31520 18150 31590
rect 18350 31520 18650 31590
rect 18850 31520 19150 31590
rect 19350 31520 19650 31590
rect 19850 31520 20150 31590
rect 20350 31520 20650 31590
rect 20850 31520 21150 31590
rect 21350 31520 21650 31590
rect 21850 31520 22150 31590
rect 22350 31520 22650 31590
rect 22850 31520 23150 31590
rect 23350 31520 23650 31590
rect 23850 31520 24150 31590
rect 24350 31520 24650 31590
rect 24850 31520 25150 31590
rect 25350 31520 25650 31590
rect 25850 31520 26150 31590
rect 26350 31520 26500 31590
rect 0 31500 26500 31520
rect 0 31480 1340 31500
rect 0 31410 150 31480
rect 350 31410 650 31480
rect 850 31410 1340 31480
rect 0 31400 1340 31410
rect 0 31380 120 31400
rect 380 31380 620 31400
rect 880 31380 1340 31400
rect 0 31350 100 31380
rect 0 31150 20 31350
rect 90 31150 100 31350
rect 0 31120 100 31150
rect 400 31350 600 31380
rect 400 31150 410 31350
rect 480 31150 520 31350
rect 590 31150 600 31350
rect 400 31120 600 31150
rect 900 31350 1340 31380
rect 900 31150 910 31350
rect 980 31150 1340 31350
rect 900 31120 1340 31150
rect 0 31100 120 31120
rect 380 31100 620 31120
rect 880 31100 1340 31120
rect 0 31090 1340 31100
rect 0 31020 150 31090
rect 350 31020 650 31090
rect 850 31020 1340 31090
rect 0 30980 1340 31020
rect 0 30910 150 30980
rect 350 30910 650 30980
rect 850 30910 1340 30980
rect 0 30900 1340 30910
rect 0 30880 120 30900
rect 380 30880 620 30900
rect 880 30880 1340 30900
rect 6500 31480 7500 31500
rect 6500 31410 6650 31480
rect 6850 31410 7150 31480
rect 7350 31410 7500 31480
rect 6500 31400 7500 31410
rect 6500 31380 6620 31400
rect 6880 31380 7120 31400
rect 7380 31380 7500 31400
rect 6500 31350 6600 31380
rect 6500 31150 6520 31350
rect 6590 31150 6600 31350
rect 6500 31120 6600 31150
rect 6900 31350 7100 31380
rect 6900 31150 6910 31350
rect 6980 31150 7020 31350
rect 7090 31150 7100 31350
rect 6900 31120 7100 31150
rect 7400 31350 7500 31380
rect 7400 31150 7410 31350
rect 7480 31150 7500 31350
rect 7400 31120 7500 31150
rect 6500 31100 6620 31120
rect 6880 31100 7120 31120
rect 7380 31100 7500 31120
rect 6500 31090 7500 31100
rect 6500 31020 6650 31090
rect 6850 31020 7150 31090
rect 7350 31020 7500 31090
rect 6500 30980 7500 31020
rect 13000 31480 13500 31500
rect 13000 31410 13150 31480
rect 13350 31410 13500 31480
rect 13000 31400 13500 31410
rect 13000 31380 13120 31400
rect 13380 31380 13500 31400
rect 13000 31350 13100 31380
rect 13000 31150 13020 31350
rect 13090 31150 13100 31350
rect 13000 31120 13100 31150
rect 13400 31350 13500 31380
rect 13400 31150 13410 31350
rect 13480 31150 13500 31350
rect 13400 31120 13500 31150
rect 13000 31100 13120 31120
rect 13380 31100 13500 31120
rect 13000 31090 13500 31100
rect 13000 31020 13150 31090
rect 13350 31020 13500 31090
rect 13000 31000 13500 31020
rect 19500 31480 20000 31500
rect 19500 31410 19650 31480
rect 19850 31410 20000 31480
rect 19500 31400 20000 31410
rect 19500 31380 19620 31400
rect 19880 31380 20000 31400
rect 19500 31350 19600 31380
rect 19500 31150 19520 31350
rect 19590 31150 19600 31350
rect 19500 31120 19600 31150
rect 19900 31350 20000 31380
rect 19900 31150 19910 31350
rect 19980 31150 20000 31350
rect 19900 31120 20000 31150
rect 19500 31100 19620 31120
rect 19880 31100 20000 31120
rect 19500 31090 20000 31100
rect 19500 31020 19650 31090
rect 19850 31020 20000 31090
rect 6500 30910 6650 30980
rect 6850 30910 7150 30980
rect 7350 30910 7500 30980
rect 6500 30900 7500 30910
rect 6500 30880 6620 30900
rect 6880 30880 7120 30900
rect 7380 30880 7500 30900
rect 19500 30980 20000 31020
rect 19500 30910 19650 30980
rect 19850 30910 20000 30980
rect 19500 30900 20000 30910
rect 19500 30880 19620 30900
rect 19880 30880 20000 30900
rect 25260 31480 26500 31500
rect 25260 31410 25650 31480
rect 25850 31410 26150 31480
rect 26350 31410 26500 31480
rect 25260 31400 26500 31410
rect 25260 31380 25620 31400
rect 25880 31380 26120 31400
rect 26380 31380 26500 31400
rect 25260 31350 25600 31380
rect 25260 31150 25520 31350
rect 25590 31150 25600 31350
rect 25260 31120 25600 31150
rect 25900 31350 26100 31380
rect 25900 31150 25910 31350
rect 25980 31150 26020 31350
rect 26090 31150 26100 31350
rect 25900 31120 26100 31150
rect 26400 31350 26500 31380
rect 26400 31150 26410 31350
rect 26480 31150 26500 31350
rect 26400 31120 26500 31150
rect 25260 31100 25620 31120
rect 25880 31100 26120 31120
rect 26380 31100 26500 31120
rect 25260 31090 26500 31100
rect 25260 31020 25650 31090
rect 25850 31020 26150 31090
rect 26350 31020 26500 31090
rect 25260 30980 26500 31020
rect 25260 30910 25650 30980
rect 25850 30910 26150 30980
rect 26350 30910 26500 30980
rect 25260 30900 26500 30910
rect 25260 30880 25620 30900
rect 25880 30880 26120 30900
rect 26380 30880 26500 30900
rect 0 30850 100 30880
rect 0 30650 20 30850
rect 90 30650 100 30850
rect 0 30620 100 30650
rect 400 30850 600 30880
rect 400 30650 410 30850
rect 480 30650 520 30850
rect 590 30650 600 30850
rect 400 30620 600 30650
rect 900 30870 6410 30880
rect 900 30850 1536 30870
rect 900 30650 910 30850
rect 980 30832 1536 30850
rect 6259 30832 6410 30870
rect 980 30822 6410 30832
rect 980 30820 1400 30822
rect 980 30650 1330 30820
rect 6340 30820 6410 30822
rect 1532 30730 1552 30790
rect 6186 30730 6206 30790
rect 1532 30696 1544 30730
rect 6194 30696 6206 30730
rect 1532 30690 1552 30696
rect 6186 30690 6206 30696
rect 900 30620 1330 30650
rect 0 30600 120 30620
rect 380 30600 620 30620
rect 880 30600 1330 30620
rect 0 30590 1330 30600
rect 0 30520 150 30590
rect 350 30520 650 30590
rect 850 30520 1330 30590
rect 0 30480 1330 30520
rect 0 30410 150 30480
rect 350 30410 650 30480
rect 850 30410 1330 30480
rect 0 30400 1330 30410
rect 0 30380 120 30400
rect 380 30380 620 30400
rect 880 30380 1330 30400
rect 0 30350 100 30380
rect 0 30150 20 30350
rect 90 30150 100 30350
rect 0 30120 100 30150
rect 400 30350 600 30380
rect 400 30150 410 30350
rect 480 30150 520 30350
rect 590 30150 600 30350
rect 400 30120 600 30150
rect 900 30350 1330 30380
rect 900 30150 910 30350
rect 980 30150 1330 30350
rect 900 30120 1330 30150
rect 0 30100 120 30120
rect 380 30100 620 30120
rect 880 30100 1330 30120
rect 0 30090 1330 30100
rect 0 30020 150 30090
rect 350 30020 650 30090
rect 850 30020 1330 30090
rect 0 29980 1330 30020
rect 0 29910 150 29980
rect 350 29910 650 29980
rect 850 29910 1330 29980
rect 0 29900 1330 29910
rect 0 29880 120 29900
rect 380 29880 620 29900
rect 880 29880 1330 29900
rect 0 29850 100 29880
rect 0 29650 20 29850
rect 90 29650 100 29850
rect 0 29620 100 29650
rect 400 29850 600 29880
rect 400 29650 410 29850
rect 480 29650 520 29850
rect 590 29650 600 29850
rect 400 29620 600 29650
rect 900 29850 1330 29880
rect 900 29650 910 29850
rect 980 29650 1330 29850
rect 900 29620 1330 29650
rect 0 29600 120 29620
rect 380 29600 620 29620
rect 880 29600 1330 29620
rect 0 29590 1330 29600
rect 0 29520 150 29590
rect 350 29520 650 29590
rect 850 29520 1330 29590
rect 0 29480 1330 29520
rect 0 29410 150 29480
rect 350 29410 650 29480
rect 850 29410 1330 29480
rect 0 29400 1330 29410
rect 0 29380 120 29400
rect 380 29380 620 29400
rect 880 29380 1330 29400
rect 0 29350 100 29380
rect 0 29150 20 29350
rect 90 29150 100 29350
rect 0 29120 100 29150
rect 400 29350 600 29380
rect 400 29150 410 29350
rect 480 29150 520 29350
rect 590 29150 600 29350
rect 400 29120 600 29150
rect 900 29350 1330 29380
rect 900 29150 910 29350
rect 980 29150 1330 29350
rect 900 29120 1330 29150
rect 0 29100 120 29120
rect 380 29100 620 29120
rect 880 29100 1330 29120
rect 0 29090 1330 29100
rect 0 29020 150 29090
rect 350 29020 650 29090
rect 850 29020 1330 29090
rect 0 28980 1330 29020
rect 0 28910 150 28980
rect 350 28910 650 28980
rect 850 28910 1330 28980
rect 0 28900 1330 28910
rect 0 28880 120 28900
rect 380 28880 620 28900
rect 880 28880 1330 28900
rect 0 28850 100 28880
rect 0 28650 20 28850
rect 90 28650 100 28850
rect 0 28620 100 28650
rect 400 28850 600 28880
rect 400 28650 410 28850
rect 480 28650 520 28850
rect 590 28650 600 28850
rect 400 28620 600 28650
rect 900 28850 1330 28880
rect 900 28650 910 28850
rect 980 28650 1330 28850
rect 900 28620 1330 28650
rect 0 28600 120 28620
rect 380 28600 620 28620
rect 880 28600 1330 28620
rect 0 28590 1330 28600
rect 0 28520 150 28590
rect 350 28520 650 28590
rect 850 28520 1330 28590
rect 0 28480 1330 28520
rect 0 28410 150 28480
rect 350 28410 650 28480
rect 850 28410 1330 28480
rect 0 28400 1330 28410
rect 0 28380 120 28400
rect 380 28380 620 28400
rect 880 28380 1330 28400
rect 0 28350 100 28380
rect 0 28150 20 28350
rect 90 28150 100 28350
rect 0 28120 100 28150
rect 400 28350 600 28380
rect 400 28150 410 28350
rect 480 28150 520 28350
rect 590 28150 600 28350
rect 400 28120 600 28150
rect 900 28350 1330 28380
rect 900 28150 910 28350
rect 980 28150 1330 28350
rect 900 28120 1330 28150
rect 0 28100 120 28120
rect 380 28100 620 28120
rect 880 28100 1330 28120
rect 0 28090 1330 28100
rect 0 28020 150 28090
rect 350 28020 650 28090
rect 850 28020 1330 28090
rect 0 27980 1330 28020
rect 0 27910 150 27980
rect 350 27910 650 27980
rect 850 27910 1330 27980
rect 0 27900 1330 27910
rect 0 27880 120 27900
rect 380 27880 620 27900
rect 880 27880 1330 27900
rect 0 27850 100 27880
rect 0 27650 20 27850
rect 90 27650 100 27850
rect 0 27620 100 27650
rect 400 27850 600 27880
rect 400 27650 410 27850
rect 480 27650 520 27850
rect 590 27650 600 27850
rect 400 27620 600 27650
rect 900 27850 1330 27880
rect 900 27650 910 27850
rect 980 27650 1330 27850
rect 900 27620 1330 27650
rect 0 27600 120 27620
rect 380 27600 620 27620
rect 880 27600 1330 27620
rect 0 27590 1330 27600
rect 0 27520 150 27590
rect 350 27520 650 27590
rect 850 27520 1330 27590
rect 0 27480 1330 27520
rect 0 27410 150 27480
rect 350 27410 650 27480
rect 850 27410 1330 27480
rect 0 27400 1330 27410
rect 0 27380 120 27400
rect 380 27380 620 27400
rect 880 27380 1330 27400
rect 0 27350 100 27380
rect -4300 27250 -4100 27260
rect -4300 27030 -4290 27250
rect -4110 27030 -4100 27250
rect -4300 27020 -4100 27030
rect -4060 27200 -3980 27220
rect -4300 25710 -4100 25720
rect -4300 25490 -4290 25710
rect -4110 25490 -4100 25710
rect -4060 25540 -4040 27200
rect -4000 27000 -3980 27200
rect 0 27150 20 27350
rect 90 27150 100 27350
rect 0 27120 100 27150
rect 400 27350 600 27380
rect 400 27150 410 27350
rect 480 27150 520 27350
rect 590 27150 600 27350
rect 400 27120 600 27150
rect 900 27350 1330 27380
rect 900 27150 910 27350
rect 980 27150 1330 27350
rect 900 27120 1330 27150
rect 0 27100 120 27120
rect 380 27100 620 27120
rect 880 27100 1330 27120
rect 0 27090 1330 27100
rect 0 27020 150 27090
rect 350 27020 650 27090
rect 850 27020 1330 27090
rect 0 27000 1330 27020
rect -4000 26980 1330 27000
rect -4000 26910 -3850 26980
rect -3650 26910 -3350 26980
rect -3150 26910 -2850 26980
rect -2650 26910 -2350 26980
rect -2150 26910 -1850 26980
rect -1650 26910 -1350 26980
rect -1150 26910 -850 26980
rect -650 26910 -350 26980
rect -150 26910 150 26980
rect 350 26910 650 26980
rect 850 26910 1330 26980
rect -4000 26900 1330 26910
rect -4000 26880 -3880 26900
rect -3620 26880 -3380 26900
rect -3120 26880 -2880 26900
rect -2620 26880 -2380 26900
rect -2120 26880 -1880 26900
rect -1620 26880 -1380 26900
rect -1120 26880 -880 26900
rect -620 26880 -380 26900
rect -120 26880 120 26900
rect 380 26880 620 26900
rect 880 26880 1330 26900
rect -4000 26850 -3900 26880
rect -4000 26650 -3980 26850
rect -3910 26650 -3900 26850
rect -4000 26620 -3900 26650
rect -3600 26850 -3400 26880
rect -3600 26650 -3590 26850
rect -3520 26650 -3480 26850
rect -3410 26650 -3400 26850
rect -3600 26620 -3400 26650
rect -3100 26850 -2900 26880
rect -3100 26650 -3090 26850
rect -3020 26650 -2980 26850
rect -2910 26650 -2900 26850
rect -3100 26620 -2900 26650
rect -2600 26850 -2400 26880
rect -2600 26650 -2590 26850
rect -2520 26650 -2480 26850
rect -2410 26650 -2400 26850
rect -2600 26620 -2400 26650
rect -2100 26850 -1900 26880
rect -2100 26650 -2090 26850
rect -2020 26650 -1980 26850
rect -1910 26650 -1900 26850
rect -2100 26620 -1900 26650
rect -1600 26850 -1400 26880
rect -1600 26650 -1590 26850
rect -1520 26650 -1480 26850
rect -1410 26650 -1400 26850
rect -1600 26620 -1400 26650
rect -1100 26850 -900 26880
rect -1100 26650 -1090 26850
rect -1020 26650 -980 26850
rect -910 26650 -900 26850
rect -1100 26620 -900 26650
rect -600 26850 -400 26880
rect -600 26650 -590 26850
rect -520 26650 -480 26850
rect -410 26650 -400 26850
rect -600 26620 -400 26650
rect -100 26850 100 26880
rect -100 26650 -90 26850
rect -20 26650 20 26850
rect 90 26650 100 26850
rect -100 26620 100 26650
rect 400 26850 600 26880
rect 400 26650 410 26850
rect 480 26650 520 26850
rect 590 26650 600 26850
rect 400 26620 600 26650
rect 900 26850 1330 26880
rect 900 26650 910 26850
rect 980 26650 1330 26850
rect 900 26620 1330 26650
rect -4000 26600 -3880 26620
rect -3620 26600 -3380 26620
rect -3120 26600 -2880 26620
rect -2620 26600 -2380 26620
rect -2120 26600 -1880 26620
rect -1620 26600 -1380 26620
rect -1120 26600 -880 26620
rect -620 26600 -380 26620
rect -120 26600 120 26620
rect 380 26600 620 26620
rect 880 26600 1330 26620
rect -4000 26590 1330 26600
rect -4000 26520 -3850 26590
rect -3650 26520 -3350 26590
rect -3150 26520 -2850 26590
rect -2650 26520 -2350 26590
rect -2150 26520 -1850 26590
rect -1650 26520 -1350 26590
rect -1150 26520 -850 26590
rect -650 26520 -350 26590
rect -150 26520 150 26590
rect 350 26520 650 26590
rect 850 26520 1330 26590
rect -4000 26480 1330 26520
rect -4000 26410 -3850 26480
rect -3650 26410 -3350 26480
rect -3150 26410 -2850 26480
rect -2650 26410 -2350 26480
rect -2150 26410 -1850 26480
rect -1650 26410 -1350 26480
rect -1150 26410 -850 26480
rect -650 26410 -350 26480
rect -150 26410 150 26480
rect 350 26410 650 26480
rect 850 26410 1330 26480
rect -4000 26400 1330 26410
rect -4000 26380 -3880 26400
rect -3620 26380 -3380 26400
rect -3120 26380 -2880 26400
rect -2620 26380 -2380 26400
rect -2120 26380 -1880 26400
rect -1620 26380 -1380 26400
rect -1120 26380 -880 26400
rect -620 26380 -380 26400
rect -120 26380 120 26400
rect 380 26380 620 26400
rect 880 26380 1330 26400
rect -4000 26350 -3900 26380
rect -4000 26150 -3980 26350
rect -3910 26150 -3900 26350
rect -4000 26120 -3900 26150
rect -3600 26350 -3400 26380
rect -3600 26150 -3590 26350
rect -3520 26150 -3480 26350
rect -3410 26150 -3400 26350
rect -3600 26120 -3400 26150
rect -3100 26350 -2900 26380
rect -3100 26150 -3090 26350
rect -3020 26150 -2980 26350
rect -2910 26150 -2900 26350
rect -3100 26120 -2900 26150
rect -2600 26350 -2400 26380
rect -2600 26150 -2590 26350
rect -2520 26150 -2480 26350
rect -2410 26150 -2400 26350
rect -2600 26120 -2400 26150
rect -2100 26350 -1900 26380
rect -2100 26150 -2090 26350
rect -2020 26150 -1980 26350
rect -1910 26150 -1900 26350
rect -2100 26120 -1900 26150
rect -1600 26350 -1400 26380
rect -1600 26150 -1590 26350
rect -1520 26150 -1480 26350
rect -1410 26150 -1400 26350
rect -1600 26120 -1400 26150
rect -1100 26350 -900 26380
rect -1100 26150 -1090 26350
rect -1020 26150 -980 26350
rect -910 26150 -900 26350
rect -1100 26120 -900 26150
rect -600 26350 -400 26380
rect -600 26150 -590 26350
rect -520 26150 -480 26350
rect -410 26150 -400 26350
rect -600 26120 -400 26150
rect -100 26350 100 26380
rect -100 26150 -90 26350
rect -20 26150 20 26350
rect 90 26150 100 26350
rect -100 26120 100 26150
rect 400 26350 600 26380
rect 400 26150 410 26350
rect 480 26150 520 26350
rect 590 26150 600 26350
rect 400 26120 600 26150
rect 900 26350 1330 26380
rect 900 26150 910 26350
rect 980 26150 1330 26350
rect 900 26120 1330 26150
rect -4000 26100 -3880 26120
rect -3620 26100 -3380 26120
rect -3120 26100 -2880 26120
rect -2620 26100 -2380 26120
rect -2120 26100 -1880 26120
rect -1620 26100 -1380 26120
rect -1120 26100 -880 26120
rect -620 26100 -380 26120
rect -120 26100 120 26120
rect 380 26100 620 26120
rect 880 26100 1330 26120
rect -4000 26090 1330 26100
rect -4000 26020 -3850 26090
rect -3650 26020 -3350 26090
rect -3150 26020 -2850 26090
rect -2650 26020 -2350 26090
rect -2150 26020 -1850 26090
rect -1650 26020 -1350 26090
rect -1150 26020 -850 26090
rect -650 26020 -350 26090
rect -150 26020 150 26090
rect 350 26020 650 26090
rect 850 26020 1330 26090
rect -4000 26000 1330 26020
rect -4000 25540 -3980 26000
rect -4060 25520 -3980 25540
rect 0 25980 1330 26000
rect 0 25910 150 25980
rect 350 25910 650 25980
rect 850 25910 1330 25980
rect 0 25900 1330 25910
rect 0 25880 120 25900
rect 380 25880 620 25900
rect 880 25880 1330 25900
rect 0 25850 100 25880
rect 0 25650 20 25850
rect 90 25650 100 25850
rect 0 25620 100 25650
rect 400 25850 600 25880
rect 400 25650 410 25850
rect 480 25650 520 25850
rect 590 25650 600 25850
rect 400 25620 600 25650
rect 900 25850 1330 25880
rect 900 25650 910 25850
rect 980 25650 1330 25850
rect 900 25620 1330 25650
rect 0 25600 120 25620
rect 380 25600 620 25620
rect 880 25600 1330 25620
rect 0 25590 1330 25600
rect 0 25520 150 25590
rect 350 25520 650 25590
rect 850 25520 1330 25590
rect -4300 25480 -4100 25490
rect 0 25480 1330 25520
rect 0 25410 150 25480
rect 350 25410 650 25480
rect 850 25410 1330 25480
rect 0 25400 1330 25410
rect 0 25380 120 25400
rect 380 25380 620 25400
rect 880 25380 1330 25400
rect 0 25350 100 25380
rect 0 25150 20 25350
rect 90 25150 100 25350
rect 0 25120 100 25150
rect 400 25350 600 25380
rect 400 25150 410 25350
rect 480 25150 520 25350
rect 590 25150 600 25350
rect 400 25120 600 25150
rect 900 25350 1330 25380
rect 900 25150 910 25350
rect 980 25150 1330 25350
rect 900 25120 1330 25150
rect 0 25100 120 25120
rect 380 25100 620 25120
rect 880 25100 1330 25120
rect 0 25090 1330 25100
rect 0 25020 150 25090
rect 350 25020 650 25090
rect 850 25020 1330 25090
rect 0 24980 1330 25020
rect 0 24910 150 24980
rect 350 24910 650 24980
rect 850 24910 1330 24980
rect 0 24900 1330 24910
rect 0 24880 120 24900
rect 380 24880 620 24900
rect 880 24880 1330 24900
rect 0 24850 100 24880
rect 0 24650 20 24850
rect 90 24650 100 24850
rect 0 24620 100 24650
rect 400 24850 600 24880
rect 400 24650 410 24850
rect 480 24650 520 24850
rect 590 24650 600 24850
rect 400 24620 600 24650
rect 900 24850 1330 24880
rect 900 24650 910 24850
rect 980 24650 1330 24850
rect 900 24620 1330 24650
rect 1465 30646 1531 30658
rect 1465 30638 1482 30646
rect 1516 30638 1531 30646
rect 1465 24670 1482 24678
rect 1516 24670 1531 24678
rect 1465 24658 1531 24670
rect 1623 30646 1689 30658
rect 1623 30638 1640 30646
rect 1674 30638 1689 30646
rect 1623 24670 1640 24678
rect 1674 24670 1689 24678
rect 1623 24658 1689 24670
rect 1781 30646 1847 30658
rect 1781 30638 1798 30646
rect 1832 30638 1847 30646
rect 1781 24670 1798 24678
rect 1832 24670 1847 24678
rect 1781 24658 1847 24670
rect 1939 30646 2005 30658
rect 1939 30638 1956 30646
rect 1990 30638 2005 30646
rect 1939 24670 1956 24678
rect 1990 24670 2005 24678
rect 1939 24658 2005 24670
rect 2097 30646 2163 30658
rect 2097 30638 2114 30646
rect 2148 30638 2163 30646
rect 2097 24670 2114 24678
rect 2148 24670 2163 24678
rect 2097 24658 2163 24670
rect 2255 30646 2321 30658
rect 2255 30638 2272 30646
rect 2306 30638 2321 30646
rect 2255 24670 2272 24678
rect 2306 24670 2321 24678
rect 2255 24658 2321 24670
rect 2413 30646 2479 30658
rect 2413 30638 2430 30646
rect 2464 30638 2479 30646
rect 2413 24670 2430 24678
rect 2464 24670 2479 24678
rect 2413 24658 2479 24670
rect 2571 30646 2637 30658
rect 2571 30638 2588 30646
rect 2622 30638 2637 30646
rect 2571 24670 2588 24678
rect 2622 24670 2637 24678
rect 2571 24658 2637 24670
rect 2729 30646 2795 30658
rect 2729 30638 2746 30646
rect 2780 30638 2795 30646
rect 2729 24670 2746 24678
rect 2780 24670 2795 24678
rect 2729 24658 2795 24670
rect 2887 30646 2953 30658
rect 2887 30638 2904 30646
rect 2938 30638 2953 30646
rect 2887 24670 2904 24678
rect 2938 24670 2953 24678
rect 2887 24658 2953 24670
rect 3045 30646 3111 30658
rect 3045 30638 3062 30646
rect 3096 30638 3111 30646
rect 3045 24670 3062 24678
rect 3096 24670 3111 24678
rect 3045 24658 3111 24670
rect 3203 30646 3269 30658
rect 3203 30638 3220 30646
rect 3254 30638 3269 30646
rect 3203 24670 3220 24678
rect 3254 24670 3269 24678
rect 3203 24658 3269 24670
rect 3361 30646 3427 30658
rect 3361 30638 3378 30646
rect 3412 30638 3427 30646
rect 3361 24670 3378 24678
rect 3412 24670 3427 24678
rect 3361 24658 3427 24670
rect 3519 30646 3585 30658
rect 3519 30638 3536 30646
rect 3570 30638 3585 30646
rect 3519 24670 3536 24678
rect 3570 24670 3585 24678
rect 3519 24658 3585 24670
rect 3677 30646 3743 30658
rect 3677 30638 3694 30646
rect 3728 30638 3743 30646
rect 3677 24670 3694 24678
rect 3728 24670 3743 24678
rect 3677 24658 3743 24670
rect 3835 30646 3901 30658
rect 3835 30638 3852 30646
rect 3886 30638 3901 30646
rect 3835 24670 3852 24678
rect 3886 24670 3901 24678
rect 3835 24658 3901 24670
rect 3993 30646 4059 30658
rect 3993 30638 4010 30646
rect 4044 30638 4059 30646
rect 3993 24670 4010 24678
rect 4044 24670 4059 24678
rect 3993 24658 4059 24670
rect 4151 30646 4217 30658
rect 4151 30638 4168 30646
rect 4202 30638 4217 30646
rect 4151 24670 4168 24678
rect 4202 24670 4217 24678
rect 4151 24658 4217 24670
rect 4309 30646 4375 30658
rect 4309 30638 4326 30646
rect 4360 30638 4375 30646
rect 4309 24670 4326 24678
rect 4360 24670 4375 24678
rect 4309 24658 4375 24670
rect 4467 30646 4533 30658
rect 4467 30638 4484 30646
rect 4518 30638 4533 30646
rect 4467 24670 4484 24678
rect 4518 24670 4533 24678
rect 4467 24658 4533 24670
rect 4625 30646 4691 30658
rect 4625 30638 4642 30646
rect 4676 30638 4691 30646
rect 4625 24670 4642 24678
rect 4676 24670 4691 24678
rect 4625 24658 4691 24670
rect 4783 30646 4849 30658
rect 4783 30638 4800 30646
rect 4834 30638 4849 30646
rect 4783 24670 4800 24678
rect 4834 24670 4849 24678
rect 4783 24658 4849 24670
rect 4941 30646 5007 30658
rect 4941 30638 4958 30646
rect 4992 30638 5007 30646
rect 4941 24670 4958 24678
rect 4992 24670 5007 24678
rect 4941 24658 5007 24670
rect 5099 30646 5165 30658
rect 5099 30638 5116 30646
rect 5150 30638 5165 30646
rect 5099 24670 5116 24678
rect 5150 24670 5165 24678
rect 5099 24658 5165 24670
rect 5257 30646 5323 30658
rect 5257 30638 5274 30646
rect 5308 30638 5323 30646
rect 5257 24670 5274 24678
rect 5308 24670 5323 24678
rect 5257 24658 5323 24670
rect 5415 30646 5481 30658
rect 5415 30638 5432 30646
rect 5466 30638 5481 30646
rect 5415 24670 5432 24678
rect 5466 24670 5481 24678
rect 5415 24658 5481 24670
rect 5573 30646 5639 30658
rect 5573 30638 5590 30646
rect 5624 30638 5639 30646
rect 5573 24670 5590 24678
rect 5624 24670 5639 24678
rect 5573 24658 5639 24670
rect 5731 30646 5797 30658
rect 5731 30638 5748 30646
rect 5782 30638 5797 30646
rect 5731 24670 5748 24678
rect 5782 24670 5797 24678
rect 5731 24658 5797 24670
rect 5889 30646 5955 30658
rect 5889 30638 5906 30646
rect 5940 30638 5955 30646
rect 5889 24670 5906 24678
rect 5940 24670 5955 24678
rect 5889 24658 5955 24670
rect 6047 30646 6113 30658
rect 6047 30638 6064 30646
rect 6098 30638 6113 30646
rect 6047 24670 6064 24678
rect 6098 24670 6113 24678
rect 6047 24658 6113 24670
rect 6205 30646 6271 30658
rect 6205 30638 6222 30646
rect 6256 30638 6271 30646
rect 6205 24670 6222 24678
rect 6256 24670 6271 24678
rect 6205 24658 6271 24670
rect 0 24600 120 24620
rect 380 24600 620 24620
rect 880 24600 1330 24620
rect 0 24590 1330 24600
rect 0 24520 150 24590
rect 350 24520 650 24590
rect 850 24520 1330 24590
rect 0 24500 1330 24520
rect 6500 30850 6600 30880
rect 6500 30650 6520 30850
rect 6590 30650 6600 30850
rect 6500 30620 6600 30650
rect 6900 30850 7100 30880
rect 6900 30650 6910 30850
rect 6980 30650 7020 30850
rect 7090 30650 7100 30850
rect 6900 30620 7100 30650
rect 7400 30850 7500 30880
rect 7400 30650 7410 30850
rect 7480 30650 7500 30850
rect 7400 30620 7500 30650
rect 6500 30600 6620 30620
rect 6880 30600 7120 30620
rect 7380 30600 7500 30620
rect 6500 30590 7500 30600
rect 6500 30520 6650 30590
rect 6850 30520 7150 30590
rect 7350 30520 7500 30590
rect 6500 30500 7500 30520
rect 7630 30870 12710 30880
rect 7630 30832 7836 30870
rect 12559 30832 12710 30870
rect 7630 30822 12710 30832
rect 7630 30820 7700 30822
rect 12640 30820 12710 30822
rect 7832 30730 7852 30790
rect 12486 30730 12506 30790
rect 7832 30696 7844 30730
rect 12494 30696 12506 30730
rect 7832 30690 7852 30696
rect 12486 30690 12506 30696
rect 1532 24620 1552 24626
rect 6186 24620 6206 24626
rect 1532 24586 1544 24620
rect 6194 24586 6206 24620
rect 1532 24526 1552 24586
rect 6186 24526 6206 24586
rect 0 24494 1400 24500
rect 6340 24494 6410 24500
rect 0 24484 6410 24494
rect 0 24480 1536 24484
rect 0 24410 150 24480
rect 350 24410 650 24480
rect 850 24446 1536 24480
rect 6202 24446 6410 24484
rect 850 24430 6410 24446
rect 7765 30646 7831 30658
rect 7765 30638 7782 30646
rect 7816 30638 7831 30646
rect 7765 24670 7782 24678
rect 7816 24670 7831 24678
rect 7765 24658 7831 24670
rect 7923 30646 7989 30658
rect 7923 30638 7940 30646
rect 7974 30638 7989 30646
rect 7923 24670 7940 24678
rect 7974 24670 7989 24678
rect 7923 24658 7989 24670
rect 8081 30646 8147 30658
rect 8081 30638 8098 30646
rect 8132 30638 8147 30646
rect 8081 24670 8098 24678
rect 8132 24670 8147 24678
rect 8081 24658 8147 24670
rect 8239 30646 8305 30658
rect 8239 30638 8256 30646
rect 8290 30638 8305 30646
rect 8239 24670 8256 24678
rect 8290 24670 8305 24678
rect 8239 24658 8305 24670
rect 8397 30646 8463 30658
rect 8397 30638 8414 30646
rect 8448 30638 8463 30646
rect 8397 24670 8414 24678
rect 8448 24670 8463 24678
rect 8397 24658 8463 24670
rect 8555 30646 8621 30658
rect 8555 30638 8572 30646
rect 8606 30638 8621 30646
rect 8555 24670 8572 24678
rect 8606 24670 8621 24678
rect 8555 24658 8621 24670
rect 8713 30646 8779 30658
rect 8713 30638 8730 30646
rect 8764 30638 8779 30646
rect 8713 24670 8730 24678
rect 8764 24670 8779 24678
rect 8713 24658 8779 24670
rect 8871 30646 8937 30658
rect 8871 30638 8888 30646
rect 8922 30638 8937 30646
rect 8871 24670 8888 24678
rect 8922 24670 8937 24678
rect 8871 24658 8937 24670
rect 9029 30646 9095 30658
rect 9029 30638 9046 30646
rect 9080 30638 9095 30646
rect 9029 24670 9046 24678
rect 9080 24670 9095 24678
rect 9029 24658 9095 24670
rect 9187 30646 9253 30658
rect 9187 30638 9204 30646
rect 9238 30638 9253 30646
rect 9187 24670 9204 24678
rect 9238 24670 9253 24678
rect 9187 24658 9253 24670
rect 9345 30646 9411 30658
rect 9345 30638 9362 30646
rect 9396 30638 9411 30646
rect 9345 24670 9362 24678
rect 9396 24670 9411 24678
rect 9345 24658 9411 24670
rect 9503 30646 9569 30658
rect 9503 30638 9520 30646
rect 9554 30638 9569 30646
rect 9503 24670 9520 24678
rect 9554 24670 9569 24678
rect 9503 24658 9569 24670
rect 9661 30646 9727 30658
rect 9661 30638 9678 30646
rect 9712 30638 9727 30646
rect 9661 24670 9678 24678
rect 9712 24670 9727 24678
rect 9661 24658 9727 24670
rect 9819 30646 9885 30658
rect 9819 30638 9836 30646
rect 9870 30638 9885 30646
rect 9819 24670 9836 24678
rect 9870 24670 9885 24678
rect 9819 24658 9885 24670
rect 9977 30646 10043 30658
rect 9977 30638 9994 30646
rect 10028 30638 10043 30646
rect 9977 24670 9994 24678
rect 10028 24670 10043 24678
rect 9977 24658 10043 24670
rect 10135 30646 10201 30658
rect 10135 30638 10152 30646
rect 10186 30638 10201 30646
rect 10135 24670 10152 24678
rect 10186 24670 10201 24678
rect 10135 24658 10201 24670
rect 10293 30646 10359 30658
rect 10293 30638 10310 30646
rect 10344 30638 10359 30646
rect 10293 24670 10310 24678
rect 10344 24670 10359 24678
rect 10293 24658 10359 24670
rect 10451 30646 10517 30658
rect 10451 30638 10468 30646
rect 10502 30638 10517 30646
rect 10451 24670 10468 24678
rect 10502 24670 10517 24678
rect 10451 24658 10517 24670
rect 10609 30646 10675 30658
rect 10609 30638 10626 30646
rect 10660 30638 10675 30646
rect 10609 24670 10626 24678
rect 10660 24670 10675 24678
rect 10609 24658 10675 24670
rect 10767 30646 10833 30658
rect 10767 30638 10784 30646
rect 10818 30638 10833 30646
rect 10767 24670 10784 24678
rect 10818 24670 10833 24678
rect 10767 24658 10833 24670
rect 10925 30646 10991 30658
rect 10925 30638 10942 30646
rect 10976 30638 10991 30646
rect 10925 24670 10942 24678
rect 10976 24670 10991 24678
rect 10925 24658 10991 24670
rect 11083 30646 11149 30658
rect 11083 30638 11100 30646
rect 11134 30638 11149 30646
rect 11083 24670 11100 24678
rect 11134 24670 11149 24678
rect 11083 24658 11149 24670
rect 11241 30646 11307 30658
rect 11241 30638 11258 30646
rect 11292 30638 11307 30646
rect 11241 24670 11258 24678
rect 11292 24670 11307 24678
rect 11241 24658 11307 24670
rect 11399 30646 11465 30658
rect 11399 30638 11416 30646
rect 11450 30638 11465 30646
rect 11399 24670 11416 24678
rect 11450 24670 11465 24678
rect 11399 24658 11465 24670
rect 11557 30646 11623 30658
rect 11557 30638 11574 30646
rect 11608 30638 11623 30646
rect 11557 24670 11574 24678
rect 11608 24670 11623 24678
rect 11557 24658 11623 24670
rect 11715 30646 11781 30658
rect 11715 30638 11732 30646
rect 11766 30638 11781 30646
rect 11715 24670 11732 24678
rect 11766 24670 11781 24678
rect 11715 24658 11781 24670
rect 11873 30646 11939 30658
rect 11873 30638 11890 30646
rect 11924 30638 11939 30646
rect 11873 24670 11890 24678
rect 11924 24670 11939 24678
rect 11873 24658 11939 24670
rect 12031 30646 12097 30658
rect 12031 30638 12048 30646
rect 12082 30638 12097 30646
rect 12031 24670 12048 24678
rect 12082 24670 12097 24678
rect 12031 24658 12097 24670
rect 12189 30646 12255 30658
rect 12189 30638 12206 30646
rect 12240 30638 12255 30646
rect 12189 24670 12206 24678
rect 12240 24670 12255 24678
rect 12189 24658 12255 24670
rect 12347 30646 12413 30658
rect 12347 30638 12364 30646
rect 12398 30638 12413 30646
rect 12347 24670 12364 24678
rect 12398 24670 12413 24678
rect 12347 24658 12413 24670
rect 12505 30646 12571 30658
rect 12505 30638 12522 30646
rect 12556 30638 12571 30646
rect 12505 24670 12522 24678
rect 12556 24670 12571 24678
rect 12505 24658 12571 24670
rect 7832 24620 7852 24626
rect 12486 24620 12506 24626
rect 7832 24586 7844 24620
rect 12494 24586 12506 24620
rect 7832 24526 7852 24586
rect 12486 24526 12506 24586
rect 7630 24494 7700 24500
rect 12640 24494 12710 24500
rect 7630 24484 12710 24494
rect 7630 24446 7836 24484
rect 12502 24446 12710 24484
rect 7630 24430 12710 24446
rect 13930 30870 19010 30880
rect 13930 30832 14136 30870
rect 18859 30832 19010 30870
rect 13930 30822 19010 30832
rect 13930 30820 14000 30822
rect 18940 30820 19010 30822
rect 14132 30730 14152 30790
rect 18786 30730 18806 30790
rect 14132 30696 14144 30730
rect 18794 30696 18806 30730
rect 14132 30690 14152 30696
rect 18786 30690 18806 30696
rect 14065 30646 14131 30658
rect 14065 30638 14082 30646
rect 14116 30638 14131 30646
rect 14065 24670 14082 24678
rect 14116 24670 14131 24678
rect 14065 24658 14131 24670
rect 14223 30646 14289 30658
rect 14223 30638 14240 30646
rect 14274 30638 14289 30646
rect 14223 24670 14240 24678
rect 14274 24670 14289 24678
rect 14223 24658 14289 24670
rect 14381 30646 14447 30658
rect 14381 30638 14398 30646
rect 14432 30638 14447 30646
rect 14381 24670 14398 24678
rect 14432 24670 14447 24678
rect 14381 24658 14447 24670
rect 14539 30646 14605 30658
rect 14539 30638 14556 30646
rect 14590 30638 14605 30646
rect 14539 24670 14556 24678
rect 14590 24670 14605 24678
rect 14539 24658 14605 24670
rect 14697 30646 14763 30658
rect 14697 30638 14714 30646
rect 14748 30638 14763 30646
rect 14697 24670 14714 24678
rect 14748 24670 14763 24678
rect 14697 24658 14763 24670
rect 14855 30646 14921 30658
rect 14855 30638 14872 30646
rect 14906 30638 14921 30646
rect 14855 24670 14872 24678
rect 14906 24670 14921 24678
rect 14855 24658 14921 24670
rect 15013 30646 15079 30658
rect 15013 30638 15030 30646
rect 15064 30638 15079 30646
rect 15013 24670 15030 24678
rect 15064 24670 15079 24678
rect 15013 24658 15079 24670
rect 15171 30646 15237 30658
rect 15171 30638 15188 30646
rect 15222 30638 15237 30646
rect 15171 24670 15188 24678
rect 15222 24670 15237 24678
rect 15171 24658 15237 24670
rect 15329 30646 15395 30658
rect 15329 30638 15346 30646
rect 15380 30638 15395 30646
rect 15329 24670 15346 24678
rect 15380 24670 15395 24678
rect 15329 24658 15395 24670
rect 15487 30646 15553 30658
rect 15487 30638 15504 30646
rect 15538 30638 15553 30646
rect 15487 24670 15504 24678
rect 15538 24670 15553 24678
rect 15487 24658 15553 24670
rect 15645 30646 15711 30658
rect 15645 30638 15662 30646
rect 15696 30638 15711 30646
rect 15645 24670 15662 24678
rect 15696 24670 15711 24678
rect 15645 24658 15711 24670
rect 15803 30646 15869 30658
rect 15803 30638 15820 30646
rect 15854 30638 15869 30646
rect 15803 24670 15820 24678
rect 15854 24670 15869 24678
rect 15803 24658 15869 24670
rect 15961 30646 16027 30658
rect 15961 30638 15978 30646
rect 16012 30638 16027 30646
rect 15961 24670 15978 24678
rect 16012 24670 16027 24678
rect 15961 24658 16027 24670
rect 16119 30646 16185 30658
rect 16119 30638 16136 30646
rect 16170 30638 16185 30646
rect 16119 24670 16136 24678
rect 16170 24670 16185 24678
rect 16119 24658 16185 24670
rect 16277 30646 16343 30658
rect 16277 30638 16294 30646
rect 16328 30638 16343 30646
rect 16277 24670 16294 24678
rect 16328 24670 16343 24678
rect 16277 24658 16343 24670
rect 16435 30646 16501 30658
rect 16435 30638 16452 30646
rect 16486 30638 16501 30646
rect 16435 24670 16452 24678
rect 16486 24670 16501 24678
rect 16435 24658 16501 24670
rect 16593 30646 16659 30658
rect 16593 30638 16610 30646
rect 16644 30638 16659 30646
rect 16593 24670 16610 24678
rect 16644 24670 16659 24678
rect 16593 24658 16659 24670
rect 16751 30646 16817 30658
rect 16751 30638 16768 30646
rect 16802 30638 16817 30646
rect 16751 24670 16768 24678
rect 16802 24670 16817 24678
rect 16751 24658 16817 24670
rect 16909 30646 16975 30658
rect 16909 30638 16926 30646
rect 16960 30638 16975 30646
rect 16909 24670 16926 24678
rect 16960 24670 16975 24678
rect 16909 24658 16975 24670
rect 17067 30646 17133 30658
rect 17067 30638 17084 30646
rect 17118 30638 17133 30646
rect 17067 24670 17084 24678
rect 17118 24670 17133 24678
rect 17067 24658 17133 24670
rect 17225 30646 17291 30658
rect 17225 30638 17242 30646
rect 17276 30638 17291 30646
rect 17225 24670 17242 24678
rect 17276 24670 17291 24678
rect 17225 24658 17291 24670
rect 17383 30646 17449 30658
rect 17383 30638 17400 30646
rect 17434 30638 17449 30646
rect 17383 24670 17400 24678
rect 17434 24670 17449 24678
rect 17383 24658 17449 24670
rect 17541 30646 17607 30658
rect 17541 30638 17558 30646
rect 17592 30638 17607 30646
rect 17541 24670 17558 24678
rect 17592 24670 17607 24678
rect 17541 24658 17607 24670
rect 17699 30646 17765 30658
rect 17699 30638 17716 30646
rect 17750 30638 17765 30646
rect 17699 24670 17716 24678
rect 17750 24670 17765 24678
rect 17699 24658 17765 24670
rect 17857 30646 17923 30658
rect 17857 30638 17874 30646
rect 17908 30638 17923 30646
rect 17857 24670 17874 24678
rect 17908 24670 17923 24678
rect 17857 24658 17923 24670
rect 18015 30646 18081 30658
rect 18015 30638 18032 30646
rect 18066 30638 18081 30646
rect 18015 24670 18032 24678
rect 18066 24670 18081 24678
rect 18015 24658 18081 24670
rect 18173 30646 18239 30658
rect 18173 30638 18190 30646
rect 18224 30638 18239 30646
rect 18173 24670 18190 24678
rect 18224 24670 18239 24678
rect 18173 24658 18239 24670
rect 18331 30646 18397 30658
rect 18331 30638 18348 30646
rect 18382 30638 18397 30646
rect 18331 24670 18348 24678
rect 18382 24670 18397 24678
rect 18331 24658 18397 24670
rect 18489 30646 18555 30658
rect 18489 30638 18506 30646
rect 18540 30638 18555 30646
rect 18489 24670 18506 24678
rect 18540 24670 18555 24678
rect 18489 24658 18555 24670
rect 18647 30646 18713 30658
rect 18647 30638 18664 30646
rect 18698 30638 18713 30646
rect 18647 24670 18664 24678
rect 18698 24670 18713 24678
rect 18647 24658 18713 24670
rect 18805 30646 18871 30658
rect 18805 30638 18822 30646
rect 18856 30638 18871 30646
rect 18805 24670 18822 24678
rect 18856 24670 18871 24678
rect 18805 24658 18871 24670
rect 19500 30850 19600 30880
rect 19500 30650 19520 30850
rect 19590 30650 19600 30850
rect 19500 30620 19600 30650
rect 19900 30850 20000 30880
rect 19900 30650 19910 30850
rect 19980 30650 20000 30850
rect 19900 30620 20000 30650
rect 19500 30600 19620 30620
rect 19880 30600 20000 30620
rect 19500 30590 20000 30600
rect 19500 30520 19650 30590
rect 19850 30520 20000 30590
rect 19500 30500 20000 30520
rect 20230 30870 25600 30880
rect 20230 30832 20436 30870
rect 25159 30850 25600 30870
rect 25159 30832 25520 30850
rect 20230 30822 25520 30832
rect 20230 30820 20300 30822
rect 25240 30820 25520 30822
rect 20432 30730 20452 30790
rect 25086 30730 25106 30790
rect 20432 30696 20444 30730
rect 25094 30696 25106 30730
rect 20432 30690 20452 30696
rect 25086 30690 25106 30696
rect 14132 24620 14152 24626
rect 18786 24620 18806 24626
rect 14132 24586 14144 24620
rect 18794 24586 18806 24620
rect 14132 24526 14152 24586
rect 18786 24526 18806 24586
rect 13930 24494 14000 24500
rect 18940 24494 19010 24500
rect 13930 24484 19010 24494
rect 13930 24446 14136 24484
rect 18802 24446 19010 24484
rect 13930 24430 19010 24446
rect 20365 30646 20431 30658
rect 20365 30638 20382 30646
rect 20416 30638 20431 30646
rect 20365 24670 20382 24678
rect 20416 24670 20431 24678
rect 20365 24658 20431 24670
rect 20523 30646 20589 30658
rect 20523 30638 20540 30646
rect 20574 30638 20589 30646
rect 20523 24670 20540 24678
rect 20574 24670 20589 24678
rect 20523 24658 20589 24670
rect 20681 30646 20747 30658
rect 20681 30638 20698 30646
rect 20732 30638 20747 30646
rect 20681 24670 20698 24678
rect 20732 24670 20747 24678
rect 20681 24658 20747 24670
rect 20839 30646 20905 30658
rect 20839 30638 20856 30646
rect 20890 30638 20905 30646
rect 20839 24670 20856 24678
rect 20890 24670 20905 24678
rect 20839 24658 20905 24670
rect 20997 30646 21063 30658
rect 20997 30638 21014 30646
rect 21048 30638 21063 30646
rect 20997 24670 21014 24678
rect 21048 24670 21063 24678
rect 20997 24658 21063 24670
rect 21155 30646 21221 30658
rect 21155 30638 21172 30646
rect 21206 30638 21221 30646
rect 21155 24670 21172 24678
rect 21206 24670 21221 24678
rect 21155 24658 21221 24670
rect 21313 30646 21379 30658
rect 21313 30638 21330 30646
rect 21364 30638 21379 30646
rect 21313 24670 21330 24678
rect 21364 24670 21379 24678
rect 21313 24658 21379 24670
rect 21471 30646 21537 30658
rect 21471 30638 21488 30646
rect 21522 30638 21537 30646
rect 21471 24670 21488 24678
rect 21522 24670 21537 24678
rect 21471 24658 21537 24670
rect 21629 30646 21695 30658
rect 21629 30638 21646 30646
rect 21680 30638 21695 30646
rect 21629 24670 21646 24678
rect 21680 24670 21695 24678
rect 21629 24658 21695 24670
rect 21787 30646 21853 30658
rect 21787 30638 21804 30646
rect 21838 30638 21853 30646
rect 21787 24670 21804 24678
rect 21838 24670 21853 24678
rect 21787 24658 21853 24670
rect 21945 30646 22011 30658
rect 21945 30638 21962 30646
rect 21996 30638 22011 30646
rect 21945 24670 21962 24678
rect 21996 24670 22011 24678
rect 21945 24658 22011 24670
rect 22103 30646 22169 30658
rect 22103 30638 22120 30646
rect 22154 30638 22169 30646
rect 22103 24670 22120 24678
rect 22154 24670 22169 24678
rect 22103 24658 22169 24670
rect 22261 30646 22327 30658
rect 22261 30638 22278 30646
rect 22312 30638 22327 30646
rect 22261 24670 22278 24678
rect 22312 24670 22327 24678
rect 22261 24658 22327 24670
rect 22419 30646 22485 30658
rect 22419 30638 22436 30646
rect 22470 30638 22485 30646
rect 22419 24670 22436 24678
rect 22470 24670 22485 24678
rect 22419 24658 22485 24670
rect 22577 30646 22643 30658
rect 22577 30638 22594 30646
rect 22628 30638 22643 30646
rect 22577 24670 22594 24678
rect 22628 24670 22643 24678
rect 22577 24658 22643 24670
rect 22735 30646 22801 30658
rect 22735 30638 22752 30646
rect 22786 30638 22801 30646
rect 22735 24670 22752 24678
rect 22786 24670 22801 24678
rect 22735 24658 22801 24670
rect 22893 30646 22959 30658
rect 22893 30638 22910 30646
rect 22944 30638 22959 30646
rect 22893 24670 22910 24678
rect 22944 24670 22959 24678
rect 22893 24658 22959 24670
rect 23051 30646 23117 30658
rect 23051 30638 23068 30646
rect 23102 30638 23117 30646
rect 23051 24670 23068 24678
rect 23102 24670 23117 24678
rect 23051 24658 23117 24670
rect 23209 30646 23275 30658
rect 23209 30638 23226 30646
rect 23260 30638 23275 30646
rect 23209 24670 23226 24678
rect 23260 24670 23275 24678
rect 23209 24658 23275 24670
rect 23367 30646 23433 30658
rect 23367 30638 23384 30646
rect 23418 30638 23433 30646
rect 23367 24670 23384 24678
rect 23418 24670 23433 24678
rect 23367 24658 23433 24670
rect 23525 30646 23591 30658
rect 23525 30638 23542 30646
rect 23576 30638 23591 30646
rect 23525 24670 23542 24678
rect 23576 24670 23591 24678
rect 23525 24658 23591 24670
rect 23683 30646 23749 30658
rect 23683 30638 23700 30646
rect 23734 30638 23749 30646
rect 23683 24670 23700 24678
rect 23734 24670 23749 24678
rect 23683 24658 23749 24670
rect 23841 30646 23907 30658
rect 23841 30638 23858 30646
rect 23892 30638 23907 30646
rect 23841 24670 23858 24678
rect 23892 24670 23907 24678
rect 23841 24658 23907 24670
rect 23999 30646 24065 30658
rect 23999 30638 24016 30646
rect 24050 30638 24065 30646
rect 23999 24670 24016 24678
rect 24050 24670 24065 24678
rect 23999 24658 24065 24670
rect 24157 30646 24223 30658
rect 24157 30638 24174 30646
rect 24208 30638 24223 30646
rect 24157 24670 24174 24678
rect 24208 24670 24223 24678
rect 24157 24658 24223 24670
rect 24315 30646 24381 30658
rect 24315 30638 24332 30646
rect 24366 30638 24381 30646
rect 24315 24670 24332 24678
rect 24366 24670 24381 24678
rect 24315 24658 24381 24670
rect 24473 30646 24539 30658
rect 24473 30638 24490 30646
rect 24524 30638 24539 30646
rect 24473 24670 24490 24678
rect 24524 24670 24539 24678
rect 24473 24658 24539 24670
rect 24631 30646 24697 30658
rect 24631 30638 24648 30646
rect 24682 30638 24697 30646
rect 24631 24670 24648 24678
rect 24682 24670 24697 24678
rect 24631 24658 24697 24670
rect 24789 30646 24855 30658
rect 24789 30638 24806 30646
rect 24840 30638 24855 30646
rect 24789 24670 24806 24678
rect 24840 24670 24855 24678
rect 24789 24658 24855 24670
rect 24947 30646 25013 30658
rect 24947 30638 24964 30646
rect 24998 30638 25013 30646
rect 24947 24670 24964 24678
rect 24998 24670 25013 24678
rect 24947 24658 25013 24670
rect 25105 30646 25171 30658
rect 25105 30638 25122 30646
rect 25156 30638 25171 30646
rect 25105 24670 25122 24678
rect 25156 24670 25171 24678
rect 25105 24658 25171 24670
rect 25310 30650 25520 30820
rect 25590 30650 25600 30850
rect 25310 30620 25600 30650
rect 25900 30850 26100 30880
rect 25900 30650 25910 30850
rect 25980 30650 26020 30850
rect 26090 30650 26100 30850
rect 25900 30620 26100 30650
rect 26400 30850 26500 30880
rect 26400 30650 26410 30850
rect 26480 30650 26500 30850
rect 26400 30620 26500 30650
rect 25310 30600 25620 30620
rect 25880 30600 26120 30620
rect 26380 30600 26500 30620
rect 25310 30590 26500 30600
rect 25310 30520 25650 30590
rect 25850 30520 26150 30590
rect 26350 30520 26500 30590
rect 25310 30480 26500 30520
rect 25310 30410 25650 30480
rect 25850 30410 26150 30480
rect 26350 30410 26500 30480
rect 25310 30400 26500 30410
rect 25310 30380 25620 30400
rect 25880 30380 26120 30400
rect 26380 30380 26500 30400
rect 25310 30350 25600 30380
rect 25310 30150 25520 30350
rect 25590 30150 25600 30350
rect 25310 30120 25600 30150
rect 25900 30350 26100 30380
rect 25900 30150 25910 30350
rect 25980 30150 26020 30350
rect 26090 30150 26100 30350
rect 25900 30120 26100 30150
rect 26400 30350 26500 30380
rect 26400 30150 26410 30350
rect 26480 30150 26500 30350
rect 26400 30120 26500 30150
rect 25310 30100 25620 30120
rect 25880 30100 26120 30120
rect 26380 30100 26500 30120
rect 25310 30090 26500 30100
rect 25310 30020 25650 30090
rect 25850 30020 26150 30090
rect 26350 30020 26500 30090
rect 25310 29980 26500 30020
rect 25310 29910 25650 29980
rect 25850 29910 26150 29980
rect 26350 29910 26500 29980
rect 25310 29900 26500 29910
rect 25310 29880 25620 29900
rect 25880 29880 26120 29900
rect 26380 29880 26500 29900
rect 25310 29850 25600 29880
rect 25310 29650 25520 29850
rect 25590 29650 25600 29850
rect 25310 29620 25600 29650
rect 25900 29850 26100 29880
rect 25900 29650 25910 29850
rect 25980 29650 26020 29850
rect 26090 29650 26100 29850
rect 25900 29620 26100 29650
rect 26400 29850 26500 29880
rect 26400 29650 26410 29850
rect 26480 29650 26500 29850
rect 26400 29620 26500 29650
rect 25310 29600 25620 29620
rect 25880 29600 26120 29620
rect 26380 29600 26500 29620
rect 25310 29590 26500 29600
rect 25310 29520 25650 29590
rect 25850 29520 26150 29590
rect 26350 29520 26500 29590
rect 25310 29480 26500 29520
rect 25310 29410 25650 29480
rect 25850 29410 26150 29480
rect 26350 29410 26500 29480
rect 25310 29400 26500 29410
rect 25310 29380 25620 29400
rect 25880 29380 26120 29400
rect 26380 29380 26500 29400
rect 25310 29350 25600 29380
rect 25310 29150 25520 29350
rect 25590 29150 25600 29350
rect 25310 29120 25600 29150
rect 25900 29350 26100 29380
rect 25900 29150 25910 29350
rect 25980 29150 26020 29350
rect 26090 29150 26100 29350
rect 25900 29120 26100 29150
rect 26400 29350 26500 29380
rect 26400 29150 26410 29350
rect 26480 29150 26500 29350
rect 26400 29120 26500 29150
rect 25310 29100 25620 29120
rect 25880 29100 26120 29120
rect 26380 29100 26500 29120
rect 25310 29090 26500 29100
rect 25310 29020 25650 29090
rect 25850 29020 26150 29090
rect 26350 29020 26500 29090
rect 25310 28980 26500 29020
rect 25310 28910 25650 28980
rect 25850 28910 26150 28980
rect 26350 28910 26500 28980
rect 25310 28900 26500 28910
rect 25310 28880 25620 28900
rect 25880 28880 26120 28900
rect 26380 28880 26500 28900
rect 25310 28850 25600 28880
rect 25310 28650 25520 28850
rect 25590 28650 25600 28850
rect 25310 28620 25600 28650
rect 25900 28850 26100 28880
rect 25900 28650 25910 28850
rect 25980 28650 26020 28850
rect 26090 28650 26100 28850
rect 25900 28620 26100 28650
rect 26400 28850 26500 28880
rect 26400 28650 26410 28850
rect 26480 28650 26500 28850
rect 26400 28620 26500 28650
rect 25310 28600 25620 28620
rect 25880 28600 26120 28620
rect 26380 28600 26500 28620
rect 25310 28590 26500 28600
rect 25310 28520 25650 28590
rect 25850 28520 26150 28590
rect 26350 28520 26500 28590
rect 25310 28480 26500 28520
rect 25310 28410 25650 28480
rect 25850 28410 26150 28480
rect 26350 28410 26500 28480
rect 25310 28400 26500 28410
rect 25310 28380 25620 28400
rect 25880 28380 26120 28400
rect 26380 28380 26500 28400
rect 25310 28350 25600 28380
rect 25310 28150 25520 28350
rect 25590 28150 25600 28350
rect 25310 28120 25600 28150
rect 25900 28350 26100 28380
rect 25900 28150 25910 28350
rect 25980 28150 26020 28350
rect 26090 28150 26100 28350
rect 25900 28120 26100 28150
rect 26400 28350 26500 28380
rect 26400 28150 26410 28350
rect 26480 28150 26500 28350
rect 26400 28120 26500 28150
rect 25310 28100 25620 28120
rect 25880 28100 26120 28120
rect 26380 28100 26500 28120
rect 25310 28090 26500 28100
rect 25310 28020 25650 28090
rect 25850 28020 26150 28090
rect 26350 28020 26500 28090
rect 25310 27980 26500 28020
rect 25310 27910 25650 27980
rect 25850 27910 26150 27980
rect 26350 27910 26500 27980
rect 25310 27900 26500 27910
rect 25310 27880 25620 27900
rect 25880 27880 26120 27900
rect 26380 27880 26500 27900
rect 25310 27850 25600 27880
rect 25310 27650 25520 27850
rect 25590 27650 25600 27850
rect 25310 27620 25600 27650
rect 25900 27850 26100 27880
rect 25900 27650 25910 27850
rect 25980 27650 26020 27850
rect 26090 27650 26100 27850
rect 25900 27620 26100 27650
rect 26400 27850 26500 27880
rect 26400 27650 26410 27850
rect 26480 27650 26500 27850
rect 26400 27620 26500 27650
rect 25310 27600 25620 27620
rect 25880 27600 26120 27620
rect 26380 27600 26500 27620
rect 25310 27590 26500 27600
rect 25310 27520 25650 27590
rect 25850 27520 26150 27590
rect 26350 27520 26500 27590
rect 25310 27480 26500 27520
rect 25310 27410 25650 27480
rect 25850 27410 26150 27480
rect 26350 27410 26500 27480
rect 25310 27400 26500 27410
rect 25310 27380 25620 27400
rect 25880 27380 26120 27400
rect 26380 27380 26500 27400
rect 25310 27350 25600 27380
rect 25310 27150 25520 27350
rect 25590 27150 25600 27350
rect 25310 27120 25600 27150
rect 25900 27350 26100 27380
rect 25900 27150 25910 27350
rect 25980 27150 26020 27350
rect 26090 27150 26100 27350
rect 25900 27120 26100 27150
rect 26400 27350 26500 27380
rect 26400 27150 26410 27350
rect 26480 27150 26500 27350
rect 26400 27120 26500 27150
rect 25310 27100 25620 27120
rect 25880 27100 26120 27120
rect 26380 27100 26500 27120
rect 25310 27090 26500 27100
rect 25310 27020 25650 27090
rect 25850 27020 26150 27090
rect 26350 27020 26500 27090
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect 25310 27000 26500 27020
rect 25310 26980 30860 27000
rect 25310 26910 25650 26980
rect 25850 26910 26150 26980
rect 26350 26910 26650 26980
rect 26850 26910 27150 26980
rect 27350 26910 27650 26980
rect 27850 26910 28150 26980
rect 28350 26910 28650 26980
rect 28850 26910 29150 26980
rect 29350 26910 29650 26980
rect 29850 26910 30150 26980
rect 30350 26910 30800 26980
rect 25310 26900 30800 26910
rect 25310 26880 25620 26900
rect 25880 26880 26120 26900
rect 26380 26880 26620 26900
rect 26880 26880 27120 26900
rect 27380 26880 27620 26900
rect 27880 26880 28120 26900
rect 28380 26880 28620 26900
rect 28880 26880 29120 26900
rect 29380 26880 29620 26900
rect 29880 26880 30120 26900
rect 30380 26880 30800 26900
rect 25310 26850 25600 26880
rect 25310 26650 25520 26850
rect 25590 26650 25600 26850
rect 25310 26620 25600 26650
rect 25900 26850 26100 26880
rect 25900 26650 25910 26850
rect 25980 26650 26020 26850
rect 26090 26650 26100 26850
rect 25900 26620 26100 26650
rect 26400 26850 26600 26880
rect 26400 26650 26410 26850
rect 26480 26650 26520 26850
rect 26590 26650 26600 26850
rect 26400 26620 26600 26650
rect 26900 26850 27100 26880
rect 26900 26650 26910 26850
rect 26980 26650 27020 26850
rect 27090 26650 27100 26850
rect 26900 26620 27100 26650
rect 27400 26850 27600 26880
rect 27400 26650 27410 26850
rect 27480 26650 27520 26850
rect 27590 26650 27600 26850
rect 27400 26620 27600 26650
rect 27900 26850 28100 26880
rect 27900 26650 27910 26850
rect 27980 26650 28020 26850
rect 28090 26650 28100 26850
rect 27900 26620 28100 26650
rect 28400 26850 28600 26880
rect 28400 26650 28410 26850
rect 28480 26650 28520 26850
rect 28590 26650 28600 26850
rect 28400 26620 28600 26650
rect 28900 26850 29100 26880
rect 28900 26650 28910 26850
rect 28980 26650 29020 26850
rect 29090 26650 29100 26850
rect 28900 26620 29100 26650
rect 29400 26850 29600 26880
rect 29400 26650 29410 26850
rect 29480 26650 29520 26850
rect 29590 26650 29600 26850
rect 29400 26620 29600 26650
rect 29900 26850 30100 26880
rect 29900 26650 29910 26850
rect 29980 26650 30020 26850
rect 30090 26650 30100 26850
rect 29900 26620 30100 26650
rect 30400 26850 30800 26880
rect 30400 26650 30410 26850
rect 30480 26650 30800 26850
rect 30400 26620 30800 26650
rect 25310 26600 25620 26620
rect 25880 26600 26120 26620
rect 26380 26600 26620 26620
rect 26880 26600 27120 26620
rect 27380 26600 27620 26620
rect 27880 26600 28120 26620
rect 28380 26600 28620 26620
rect 28880 26600 29120 26620
rect 29380 26600 29620 26620
rect 29880 26600 30120 26620
rect 30380 26600 30800 26620
rect 25310 26590 30800 26600
rect 25310 26520 25650 26590
rect 25850 26520 26150 26590
rect 26350 26520 26650 26590
rect 26850 26520 27150 26590
rect 27350 26520 27650 26590
rect 27850 26520 28150 26590
rect 28350 26520 28650 26590
rect 28850 26520 29150 26590
rect 29350 26520 29650 26590
rect 29850 26520 30150 26590
rect 30350 26520 30800 26590
rect 25310 26480 30800 26520
rect 25310 26410 25650 26480
rect 25850 26410 26150 26480
rect 26350 26410 26650 26480
rect 26850 26410 27150 26480
rect 27350 26410 27650 26480
rect 27850 26410 28150 26480
rect 28350 26410 28650 26480
rect 28850 26410 29150 26480
rect 29350 26410 29650 26480
rect 29850 26410 30150 26480
rect 30350 26410 30800 26480
rect 25310 26400 30800 26410
rect 25310 26380 25620 26400
rect 25880 26380 26120 26400
rect 26380 26380 26620 26400
rect 26880 26380 27120 26400
rect 27380 26380 27620 26400
rect 27880 26380 28120 26400
rect 28380 26380 28620 26400
rect 28880 26380 29120 26400
rect 29380 26380 29620 26400
rect 29880 26380 30120 26400
rect 30380 26380 30800 26400
rect 25310 26350 25600 26380
rect 25310 26150 25520 26350
rect 25590 26150 25600 26350
rect 25310 26120 25600 26150
rect 25900 26350 26100 26380
rect 25900 26150 25910 26350
rect 25980 26150 26020 26350
rect 26090 26150 26100 26350
rect 25900 26120 26100 26150
rect 26400 26350 26600 26380
rect 26400 26150 26410 26350
rect 26480 26150 26520 26350
rect 26590 26150 26600 26350
rect 26400 26120 26600 26150
rect 26900 26350 27100 26380
rect 26900 26150 26910 26350
rect 26980 26150 27020 26350
rect 27090 26150 27100 26350
rect 26900 26120 27100 26150
rect 27400 26350 27600 26380
rect 27400 26150 27410 26350
rect 27480 26150 27520 26350
rect 27590 26150 27600 26350
rect 27400 26120 27600 26150
rect 27900 26350 28100 26380
rect 27900 26150 27910 26350
rect 27980 26150 28020 26350
rect 28090 26150 28100 26350
rect 27900 26120 28100 26150
rect 28400 26350 28600 26380
rect 28400 26150 28410 26350
rect 28480 26150 28520 26350
rect 28590 26150 28600 26350
rect 28400 26120 28600 26150
rect 28900 26350 29100 26380
rect 28900 26150 28910 26350
rect 28980 26150 29020 26350
rect 29090 26150 29100 26350
rect 28900 26120 29100 26150
rect 29400 26350 29600 26380
rect 29400 26150 29410 26350
rect 29480 26150 29520 26350
rect 29590 26150 29600 26350
rect 29400 26120 29600 26150
rect 29900 26350 30100 26380
rect 29900 26150 29910 26350
rect 29980 26150 30020 26350
rect 30090 26150 30100 26350
rect 29900 26120 30100 26150
rect 30400 26350 30800 26380
rect 30400 26150 30410 26350
rect 30480 26150 30800 26350
rect 30400 26120 30800 26150
rect 25310 26100 25620 26120
rect 25880 26100 26120 26120
rect 26380 26100 26620 26120
rect 26880 26100 27120 26120
rect 27380 26100 27620 26120
rect 27880 26100 28120 26120
rect 28380 26100 28620 26120
rect 28880 26100 29120 26120
rect 29380 26100 29620 26120
rect 29880 26100 30120 26120
rect 30380 26100 30800 26120
rect 25310 26090 30800 26100
rect 25310 26020 25650 26090
rect 25850 26020 26150 26090
rect 26350 26020 26650 26090
rect 26850 26020 27150 26090
rect 27350 26020 27650 26090
rect 27850 26020 28150 26090
rect 28350 26020 28650 26090
rect 28850 26020 29150 26090
rect 29350 26020 29650 26090
rect 29850 26020 30150 26090
rect 30350 26020 30800 26090
rect 30840 26020 30860 26980
rect 25310 26000 30860 26020
rect 25310 25980 26500 26000
rect 25310 25910 25650 25980
rect 25850 25910 26150 25980
rect 26350 25910 26500 25980
rect 25310 25900 26500 25910
rect 25310 25880 25620 25900
rect 25880 25880 26120 25900
rect 26380 25880 26500 25900
rect 25310 25850 25600 25880
rect 25310 25650 25520 25850
rect 25590 25650 25600 25850
rect 25310 25620 25600 25650
rect 25900 25850 26100 25880
rect 25900 25650 25910 25850
rect 25980 25650 26020 25850
rect 26090 25650 26100 25850
rect 25900 25620 26100 25650
rect 26400 25850 26500 25880
rect 26400 25650 26410 25850
rect 26480 25650 26500 25850
rect 26400 25620 26500 25650
rect 25310 25600 25620 25620
rect 25880 25600 26120 25620
rect 26380 25600 26500 25620
rect 25310 25590 26500 25600
rect 25310 25520 25650 25590
rect 25850 25520 26150 25590
rect 26350 25520 26500 25590
rect 25310 25480 26500 25520
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect 25310 25410 25650 25480
rect 25850 25410 26150 25480
rect 26350 25410 26500 25480
rect 25310 25400 26500 25410
rect 25310 25380 25620 25400
rect 25880 25380 26120 25400
rect 26380 25380 26500 25400
rect 25310 25350 25600 25380
rect 25310 25150 25520 25350
rect 25590 25150 25600 25350
rect 25310 25120 25600 25150
rect 25900 25350 26100 25380
rect 25900 25150 25910 25350
rect 25980 25150 26020 25350
rect 26090 25150 26100 25350
rect 25900 25120 26100 25150
rect 26400 25350 26500 25380
rect 26400 25150 26410 25350
rect 26480 25150 26500 25350
rect 26400 25120 26500 25150
rect 25310 25100 25620 25120
rect 25880 25100 26120 25120
rect 26380 25100 26500 25120
rect 25310 25090 26500 25100
rect 25310 25020 25650 25090
rect 25850 25020 26150 25090
rect 26350 25020 26500 25090
rect 25310 24980 26500 25020
rect 25310 24910 25650 24980
rect 25850 24910 26150 24980
rect 26350 24910 26500 24980
rect 25310 24900 26500 24910
rect 25310 24880 25620 24900
rect 25880 24880 26120 24900
rect 26380 24880 26500 24900
rect 25310 24850 25600 24880
rect 25310 24650 25520 24850
rect 25590 24650 25600 24850
rect 20432 24620 20452 24626
rect 25086 24620 25106 24626
rect 20432 24586 20444 24620
rect 25094 24586 25106 24620
rect 20432 24526 20452 24586
rect 25086 24526 25106 24586
rect 20230 24494 20300 24500
rect 25310 24620 25600 24650
rect 25900 24850 26100 24880
rect 25900 24650 25910 24850
rect 25980 24650 26020 24850
rect 26090 24650 26100 24850
rect 25900 24620 26100 24650
rect 26400 24850 26500 24880
rect 26400 24650 26410 24850
rect 26480 24650 26500 24850
rect 26400 24620 26500 24650
rect 25310 24600 25620 24620
rect 25880 24600 26120 24620
rect 26380 24600 26500 24620
rect 25310 24590 26500 24600
rect 25310 24520 25650 24590
rect 25850 24520 26150 24590
rect 26350 24520 26500 24590
rect 25310 24500 26500 24520
rect 25240 24494 26500 24500
rect 20230 24484 26500 24494
rect 20230 24446 20436 24484
rect 25102 24480 26500 24484
rect 25102 24446 25650 24480
rect 20230 24430 25650 24446
rect 850 24410 1340 24430
rect 0 24400 1340 24410
rect 0 24380 120 24400
rect 380 24380 620 24400
rect 880 24380 1340 24400
rect 0 24350 100 24380
rect 0 24150 20 24350
rect 90 24150 100 24350
rect 0 24120 100 24150
rect 400 24350 600 24380
rect 400 24150 410 24350
rect 480 24150 520 24350
rect 590 24150 600 24350
rect 400 24120 600 24150
rect 900 24350 1340 24380
rect 900 24150 910 24350
rect 980 24150 1340 24350
rect 900 24120 1340 24150
rect 0 24100 120 24120
rect 380 24100 620 24120
rect 880 24100 1340 24120
rect 0 24090 1340 24100
rect 0 24020 150 24090
rect 350 24020 650 24090
rect 850 24020 1340 24090
rect 0 23980 1340 24020
rect 0 23910 150 23980
rect 350 23910 650 23980
rect 850 23910 1340 23980
rect 0 23900 1340 23910
rect 0 23880 120 23900
rect 380 23880 620 23900
rect 880 23880 1340 23900
rect 25260 24410 25650 24430
rect 25850 24410 26150 24480
rect 26350 24410 26500 24480
rect 25260 24400 26500 24410
rect 25260 24380 25620 24400
rect 25880 24380 26120 24400
rect 26380 24380 26500 24400
rect 25260 24350 25600 24380
rect 25260 24150 25520 24350
rect 25590 24150 25600 24350
rect 25260 24120 25600 24150
rect 25900 24350 26100 24380
rect 25900 24150 25910 24350
rect 25980 24150 26020 24350
rect 26090 24150 26100 24350
rect 25900 24120 26100 24150
rect 26400 24350 26500 24380
rect 26400 24150 26410 24350
rect 26480 24150 26500 24350
rect 26400 24120 26500 24150
rect 25260 24100 25620 24120
rect 25880 24100 26120 24120
rect 26380 24100 26500 24120
rect 25260 24090 26500 24100
rect 25260 24020 25650 24090
rect 25850 24020 26150 24090
rect 26350 24020 26500 24090
rect 25260 23980 26500 24020
rect 25260 23910 25650 23980
rect 25850 23910 26150 23980
rect 26350 23910 26500 23980
rect 25260 23900 26500 23910
rect 25260 23880 25620 23900
rect 25880 23880 26120 23900
rect 26380 23880 26500 23900
rect 0 23850 100 23880
rect 0 23650 20 23850
rect 90 23650 100 23850
rect 0 23620 100 23650
rect 400 23850 600 23880
rect 400 23650 410 23850
rect 480 23650 520 23850
rect 590 23650 600 23850
rect 400 23620 600 23650
rect 900 23870 6410 23880
rect 900 23850 1536 23870
rect 900 23650 910 23850
rect 980 23832 1536 23850
rect 6259 23832 6410 23870
rect 980 23822 6410 23832
rect 980 23820 1400 23822
rect 980 23650 1330 23820
rect 6340 23820 6410 23822
rect 1532 23730 1552 23790
rect 6186 23730 6206 23790
rect 1532 23696 1544 23730
rect 6194 23696 6206 23730
rect 1532 23690 1552 23696
rect 6186 23690 6206 23696
rect 900 23620 1330 23650
rect 0 23600 120 23620
rect 380 23600 620 23620
rect 880 23600 1330 23620
rect 0 23590 1330 23600
rect 0 23520 150 23590
rect 350 23520 650 23590
rect 850 23520 1330 23590
rect 0 23480 1330 23520
rect 0 23410 150 23480
rect 350 23410 650 23480
rect 850 23410 1330 23480
rect 0 23400 1330 23410
rect 0 23380 120 23400
rect 380 23380 620 23400
rect 880 23380 1330 23400
rect 0 23350 100 23380
rect 0 23150 20 23350
rect 90 23150 100 23350
rect 0 23120 100 23150
rect 400 23350 600 23380
rect 400 23150 410 23350
rect 480 23150 520 23350
rect 590 23150 600 23350
rect 400 23120 600 23150
rect 900 23350 1330 23380
rect 900 23150 910 23350
rect 980 23150 1330 23350
rect 900 23120 1330 23150
rect 0 23100 120 23120
rect 380 23100 620 23120
rect 880 23100 1330 23120
rect 0 23090 1330 23100
rect 0 23020 150 23090
rect 350 23020 650 23090
rect 850 23020 1330 23090
rect 0 22980 1330 23020
rect 0 22910 150 22980
rect 350 22910 650 22980
rect 850 22910 1330 22980
rect 0 22900 1330 22910
rect 0 22880 120 22900
rect 380 22880 620 22900
rect 880 22880 1330 22900
rect 0 22850 100 22880
rect 0 22650 20 22850
rect 90 22650 100 22850
rect 0 22620 100 22650
rect 400 22850 600 22880
rect 400 22650 410 22850
rect 480 22650 520 22850
rect 590 22650 600 22850
rect 400 22620 600 22650
rect 900 22850 1330 22880
rect 900 22650 910 22850
rect 980 22650 1330 22850
rect 900 22620 1330 22650
rect 0 22600 120 22620
rect 380 22600 620 22620
rect 880 22600 1330 22620
rect 0 22590 1330 22600
rect 0 22520 150 22590
rect 350 22520 650 22590
rect 850 22520 1330 22590
rect 0 22480 1330 22520
rect 0 22410 150 22480
rect 350 22410 650 22480
rect 850 22410 1330 22480
rect 0 22400 1330 22410
rect 0 22380 120 22400
rect 380 22380 620 22400
rect 880 22380 1330 22400
rect 0 22350 100 22380
rect 0 22150 20 22350
rect 90 22150 100 22350
rect 0 22120 100 22150
rect 400 22350 600 22380
rect 400 22150 410 22350
rect 480 22150 520 22350
rect 590 22150 600 22350
rect 400 22120 600 22150
rect 900 22350 1330 22380
rect 900 22150 910 22350
rect 980 22150 1330 22350
rect 900 22120 1330 22150
rect 0 22100 120 22120
rect 380 22100 620 22120
rect 880 22100 1330 22120
rect 0 22090 1330 22100
rect 0 22020 150 22090
rect 350 22020 650 22090
rect 850 22020 1330 22090
rect 0 21980 1330 22020
rect 0 21910 150 21980
rect 350 21910 650 21980
rect 850 21910 1330 21980
rect 0 21900 1330 21910
rect 0 21880 120 21900
rect 380 21880 620 21900
rect 880 21880 1330 21900
rect 0 21850 100 21880
rect 0 21650 20 21850
rect 90 21650 100 21850
rect 0 21620 100 21650
rect 400 21850 600 21880
rect 400 21650 410 21850
rect 480 21650 520 21850
rect 590 21650 600 21850
rect 400 21620 600 21650
rect 900 21850 1330 21880
rect 900 21650 910 21850
rect 980 21650 1330 21850
rect 900 21620 1330 21650
rect 0 21600 120 21620
rect 380 21600 620 21620
rect 880 21600 1330 21620
rect 0 21590 1330 21600
rect 0 21520 150 21590
rect 350 21520 650 21590
rect 850 21520 1330 21590
rect 0 21480 1330 21520
rect 0 21410 150 21480
rect 350 21410 650 21480
rect 850 21410 1330 21480
rect 0 21400 1330 21410
rect 0 21380 120 21400
rect 380 21380 620 21400
rect 880 21380 1330 21400
rect 0 21350 100 21380
rect 0 21150 20 21350
rect 90 21150 100 21350
rect 0 21120 100 21150
rect 400 21350 600 21380
rect 400 21150 410 21350
rect 480 21150 520 21350
rect 590 21150 600 21350
rect 400 21120 600 21150
rect 900 21350 1330 21380
rect 900 21150 910 21350
rect 980 21150 1330 21350
rect 900 21120 1330 21150
rect 0 21100 120 21120
rect 380 21100 620 21120
rect 880 21100 1330 21120
rect 0 21090 1330 21100
rect 0 21020 150 21090
rect 350 21020 650 21090
rect 850 21020 1330 21090
rect 0 20980 1330 21020
rect 0 20910 150 20980
rect 350 20910 650 20980
rect 850 20910 1330 20980
rect 0 20900 1330 20910
rect 0 20880 120 20900
rect 380 20880 620 20900
rect 880 20880 1330 20900
rect 0 20850 100 20880
rect 0 20650 20 20850
rect 90 20650 100 20850
rect 0 20620 100 20650
rect 400 20850 600 20880
rect 400 20650 410 20850
rect 480 20650 520 20850
rect 590 20650 600 20850
rect 400 20620 600 20650
rect 900 20850 1330 20880
rect 900 20650 910 20850
rect 980 20650 1330 20850
rect 900 20620 1330 20650
rect 0 20600 120 20620
rect 380 20600 620 20620
rect 880 20600 1330 20620
rect 0 20590 1330 20600
rect 0 20520 150 20590
rect 350 20520 650 20590
rect 850 20520 1330 20590
rect 0 20480 1330 20520
rect 0 20410 150 20480
rect 350 20410 650 20480
rect 850 20410 1330 20480
rect 0 20400 1330 20410
rect 0 20380 120 20400
rect 380 20380 620 20400
rect 880 20380 1330 20400
rect 0 20350 100 20380
rect 0 20150 20 20350
rect 90 20150 100 20350
rect 0 20120 100 20150
rect 400 20350 600 20380
rect 400 20150 410 20350
rect 480 20150 520 20350
rect 590 20150 600 20350
rect 400 20120 600 20150
rect 900 20350 1330 20380
rect 900 20150 910 20350
rect 980 20150 1330 20350
rect 900 20120 1330 20150
rect 0 20100 120 20120
rect 380 20100 620 20120
rect 880 20100 1330 20120
rect 0 20090 1330 20100
rect 0 20020 150 20090
rect 350 20020 650 20090
rect 850 20020 1330 20090
rect 0 19980 1330 20020
rect 0 19910 150 19980
rect 350 19910 650 19980
rect 850 19910 1330 19980
rect 0 19900 1330 19910
rect 0 19880 120 19900
rect 380 19880 620 19900
rect 880 19880 1330 19900
rect 0 19850 100 19880
rect 0 19650 20 19850
rect 90 19650 100 19850
rect 0 19620 100 19650
rect 400 19850 600 19880
rect 400 19650 410 19850
rect 480 19650 520 19850
rect 590 19650 600 19850
rect 400 19620 600 19650
rect 900 19850 1330 19880
rect 900 19650 910 19850
rect 980 19650 1330 19850
rect 900 19620 1330 19650
rect 0 19600 120 19620
rect 380 19600 620 19620
rect 880 19600 1330 19620
rect 0 19590 1330 19600
rect 0 19520 150 19590
rect 350 19520 650 19590
rect 850 19520 1330 19590
rect 0 19480 1330 19520
rect 0 19410 150 19480
rect 350 19410 650 19480
rect 850 19410 1330 19480
rect 0 19400 1330 19410
rect 0 19380 120 19400
rect 380 19380 620 19400
rect 880 19380 1330 19400
rect 0 19350 100 19380
rect 0 19150 20 19350
rect 90 19150 100 19350
rect 0 19120 100 19150
rect 400 19350 600 19380
rect 400 19150 410 19350
rect 480 19150 520 19350
rect 590 19150 600 19350
rect 400 19120 600 19150
rect 900 19350 1330 19380
rect 900 19150 910 19350
rect 980 19150 1330 19350
rect 900 19120 1330 19150
rect 0 19100 120 19120
rect 380 19100 620 19120
rect 880 19100 1330 19120
rect 0 19090 1330 19100
rect 0 19020 150 19090
rect 350 19020 650 19090
rect 850 19020 1330 19090
rect 0 18980 1330 19020
rect 0 18910 150 18980
rect 350 18910 650 18980
rect 850 18910 1330 18980
rect 0 18900 1330 18910
rect 0 18880 120 18900
rect 380 18880 620 18900
rect 880 18880 1330 18900
rect 0 18850 100 18880
rect 0 18650 20 18850
rect 90 18650 100 18850
rect 0 18620 100 18650
rect 400 18850 600 18880
rect 400 18650 410 18850
rect 480 18650 520 18850
rect 590 18650 600 18850
rect 400 18620 600 18650
rect 900 18850 1330 18880
rect 900 18650 910 18850
rect 980 18650 1330 18850
rect 900 18620 1330 18650
rect 0 18600 120 18620
rect 380 18600 620 18620
rect 880 18600 1330 18620
rect 0 18590 1330 18600
rect 0 18520 150 18590
rect 350 18520 650 18590
rect 850 18520 1330 18590
rect 0 18480 1330 18520
rect 0 18410 150 18480
rect 350 18410 650 18480
rect 850 18410 1330 18480
rect 0 18400 1330 18410
rect 0 18380 120 18400
rect 380 18380 620 18400
rect 880 18380 1330 18400
rect 0 18350 100 18380
rect 0 18150 20 18350
rect 90 18150 100 18350
rect 0 18120 100 18150
rect 400 18350 600 18380
rect 400 18150 410 18350
rect 480 18150 520 18350
rect 590 18150 600 18350
rect 400 18120 600 18150
rect 900 18350 1330 18380
rect 900 18150 910 18350
rect 980 18150 1330 18350
rect 900 18120 1330 18150
rect 0 18100 120 18120
rect 380 18100 620 18120
rect 880 18100 1330 18120
rect 0 18090 1330 18100
rect 0 18020 150 18090
rect 350 18020 650 18090
rect 850 18020 1330 18090
rect 0 17980 1330 18020
rect 0 17910 150 17980
rect 350 17910 650 17980
rect 850 17910 1330 17980
rect 0 17900 1330 17910
rect 0 17880 120 17900
rect 380 17880 620 17900
rect 880 17880 1330 17900
rect 0 17850 100 17880
rect 0 17650 20 17850
rect 90 17650 100 17850
rect 0 17620 100 17650
rect 400 17850 600 17880
rect 400 17650 410 17850
rect 480 17650 520 17850
rect 590 17650 600 17850
rect 400 17620 600 17650
rect 900 17850 1330 17880
rect 900 17650 910 17850
rect 980 17650 1330 17850
rect 900 17620 1330 17650
rect 1465 23646 1531 23658
rect 1465 23638 1482 23646
rect 1516 23638 1531 23646
rect 1465 17670 1482 17678
rect 1516 17670 1531 17678
rect 1465 17658 1531 17670
rect 1623 23646 1689 23658
rect 1623 23638 1640 23646
rect 1674 23638 1689 23646
rect 1623 17670 1640 17678
rect 1674 17670 1689 17678
rect 1623 17658 1689 17670
rect 1781 23646 1847 23658
rect 1781 23638 1798 23646
rect 1832 23638 1847 23646
rect 1781 17670 1798 17678
rect 1832 17670 1847 17678
rect 1781 17658 1847 17670
rect 1939 23646 2005 23658
rect 1939 23638 1956 23646
rect 1990 23638 2005 23646
rect 1939 17670 1956 17678
rect 1990 17670 2005 17678
rect 1939 17658 2005 17670
rect 2097 23646 2163 23658
rect 2097 23638 2114 23646
rect 2148 23638 2163 23646
rect 2097 17670 2114 17678
rect 2148 17670 2163 17678
rect 2097 17658 2163 17670
rect 2255 23646 2321 23658
rect 2255 23638 2272 23646
rect 2306 23638 2321 23646
rect 2255 17670 2272 17678
rect 2306 17670 2321 17678
rect 2255 17658 2321 17670
rect 2413 23646 2479 23658
rect 2413 23638 2430 23646
rect 2464 23638 2479 23646
rect 2413 17670 2430 17678
rect 2464 17670 2479 17678
rect 2413 17658 2479 17670
rect 2571 23646 2637 23658
rect 2571 23638 2588 23646
rect 2622 23638 2637 23646
rect 2571 17670 2588 17678
rect 2622 17670 2637 17678
rect 2571 17658 2637 17670
rect 2729 23646 2795 23658
rect 2729 23638 2746 23646
rect 2780 23638 2795 23646
rect 2729 17670 2746 17678
rect 2780 17670 2795 17678
rect 2729 17658 2795 17670
rect 2887 23646 2953 23658
rect 2887 23638 2904 23646
rect 2938 23638 2953 23646
rect 2887 17670 2904 17678
rect 2938 17670 2953 17678
rect 2887 17658 2953 17670
rect 3045 23646 3111 23658
rect 3045 23638 3062 23646
rect 3096 23638 3111 23646
rect 3045 17670 3062 17678
rect 3096 17670 3111 17678
rect 3045 17658 3111 17670
rect 3203 23646 3269 23658
rect 3203 23638 3220 23646
rect 3254 23638 3269 23646
rect 3203 17670 3220 17678
rect 3254 17670 3269 17678
rect 3203 17658 3269 17670
rect 3361 23646 3427 23658
rect 3361 23638 3378 23646
rect 3412 23638 3427 23646
rect 3361 17670 3378 17678
rect 3412 17670 3427 17678
rect 3361 17658 3427 17670
rect 3519 23646 3585 23658
rect 3519 23638 3536 23646
rect 3570 23638 3585 23646
rect 3519 17670 3536 17678
rect 3570 17670 3585 17678
rect 3519 17658 3585 17670
rect 3677 23646 3743 23658
rect 3677 23638 3694 23646
rect 3728 23638 3743 23646
rect 3677 17670 3694 17678
rect 3728 17670 3743 17678
rect 3677 17658 3743 17670
rect 3835 23646 3901 23658
rect 3835 23638 3852 23646
rect 3886 23638 3901 23646
rect 3835 17670 3852 17678
rect 3886 17670 3901 17678
rect 3835 17658 3901 17670
rect 3993 23646 4059 23658
rect 3993 23638 4010 23646
rect 4044 23638 4059 23646
rect 3993 17670 4010 17678
rect 4044 17670 4059 17678
rect 3993 17658 4059 17670
rect 4151 23646 4217 23658
rect 4151 23638 4168 23646
rect 4202 23638 4217 23646
rect 4151 17670 4168 17678
rect 4202 17670 4217 17678
rect 4151 17658 4217 17670
rect 4309 23646 4375 23658
rect 4309 23638 4326 23646
rect 4360 23638 4375 23646
rect 4309 17670 4326 17678
rect 4360 17670 4375 17678
rect 4309 17658 4375 17670
rect 4467 23646 4533 23658
rect 4467 23638 4484 23646
rect 4518 23638 4533 23646
rect 4467 17670 4484 17678
rect 4518 17670 4533 17678
rect 4467 17658 4533 17670
rect 4625 23646 4691 23658
rect 4625 23638 4642 23646
rect 4676 23638 4691 23646
rect 4625 17670 4642 17678
rect 4676 17670 4691 17678
rect 4625 17658 4691 17670
rect 4783 23646 4849 23658
rect 4783 23638 4800 23646
rect 4834 23638 4849 23646
rect 4783 17670 4800 17678
rect 4834 17670 4849 17678
rect 4783 17658 4849 17670
rect 4941 23646 5007 23658
rect 4941 23638 4958 23646
rect 4992 23638 5007 23646
rect 4941 17670 4958 17678
rect 4992 17670 5007 17678
rect 4941 17658 5007 17670
rect 5099 23646 5165 23658
rect 5099 23638 5116 23646
rect 5150 23638 5165 23646
rect 5099 17670 5116 17678
rect 5150 17670 5165 17678
rect 5099 17658 5165 17670
rect 5257 23646 5323 23658
rect 5257 23638 5274 23646
rect 5308 23638 5323 23646
rect 5257 17670 5274 17678
rect 5308 17670 5323 17678
rect 5257 17658 5323 17670
rect 5415 23646 5481 23658
rect 5415 23638 5432 23646
rect 5466 23638 5481 23646
rect 5415 17670 5432 17678
rect 5466 17670 5481 17678
rect 5415 17658 5481 17670
rect 5573 23646 5639 23658
rect 5573 23638 5590 23646
rect 5624 23638 5639 23646
rect 5573 17670 5590 17678
rect 5624 17670 5639 17678
rect 5573 17658 5639 17670
rect 5731 23646 5797 23658
rect 5731 23638 5748 23646
rect 5782 23638 5797 23646
rect 5731 17670 5748 17678
rect 5782 17670 5797 17678
rect 5731 17658 5797 17670
rect 5889 23646 5955 23658
rect 5889 23638 5906 23646
rect 5940 23638 5955 23646
rect 5889 17670 5906 17678
rect 5940 17670 5955 17678
rect 5889 17658 5955 17670
rect 6047 23646 6113 23658
rect 6047 23638 6064 23646
rect 6098 23638 6113 23646
rect 6047 17670 6064 17678
rect 6098 17670 6113 17678
rect 6047 17658 6113 17670
rect 6205 23646 6271 23658
rect 6205 23638 6222 23646
rect 6256 23638 6271 23646
rect 6205 17670 6222 17678
rect 6256 17670 6271 17678
rect 6205 17658 6271 17670
rect 0 17600 120 17620
rect 380 17600 620 17620
rect 880 17600 1330 17620
rect 0 17590 1330 17600
rect 0 17520 150 17590
rect 350 17520 650 17590
rect 850 17520 1330 17590
rect 0 17500 1330 17520
rect 1532 17620 1552 17626
rect 6186 17620 6206 17626
rect 1532 17586 1544 17620
rect 6194 17586 6206 17620
rect 1532 17526 1552 17586
rect 6186 17526 6206 17586
rect 0 17494 1400 17500
rect 7630 23870 12710 23880
rect 7630 23832 7836 23870
rect 12559 23832 12710 23870
rect 7630 23822 12710 23832
rect 7630 23820 7700 23822
rect 12640 23820 12710 23822
rect 7832 23730 7852 23790
rect 12486 23730 12506 23790
rect 7832 23696 7844 23730
rect 12494 23696 12506 23730
rect 7832 23690 7852 23696
rect 12486 23690 12506 23696
rect 7765 23646 7831 23658
rect 7765 23638 7782 23646
rect 7816 23638 7831 23646
rect 7765 17670 7782 17678
rect 7816 17670 7831 17678
rect 7765 17658 7831 17670
rect 7923 23646 7989 23658
rect 7923 23638 7940 23646
rect 7974 23638 7989 23646
rect 7923 17670 7940 17678
rect 7974 17670 7989 17678
rect 7923 17658 7989 17670
rect 8081 23646 8147 23658
rect 8081 23638 8098 23646
rect 8132 23638 8147 23646
rect 8081 17670 8098 17678
rect 8132 17670 8147 17678
rect 8081 17658 8147 17670
rect 8239 23646 8305 23658
rect 8239 23638 8256 23646
rect 8290 23638 8305 23646
rect 8239 17670 8256 17678
rect 8290 17670 8305 17678
rect 8239 17658 8305 17670
rect 8397 23646 8463 23658
rect 8397 23638 8414 23646
rect 8448 23638 8463 23646
rect 8397 17670 8414 17678
rect 8448 17670 8463 17678
rect 8397 17658 8463 17670
rect 8555 23646 8621 23658
rect 8555 23638 8572 23646
rect 8606 23638 8621 23646
rect 8555 17670 8572 17678
rect 8606 17670 8621 17678
rect 8555 17658 8621 17670
rect 8713 23646 8779 23658
rect 8713 23638 8730 23646
rect 8764 23638 8779 23646
rect 8713 17670 8730 17678
rect 8764 17670 8779 17678
rect 8713 17658 8779 17670
rect 8871 23646 8937 23658
rect 8871 23638 8888 23646
rect 8922 23638 8937 23646
rect 8871 17670 8888 17678
rect 8922 17670 8937 17678
rect 8871 17658 8937 17670
rect 9029 23646 9095 23658
rect 9029 23638 9046 23646
rect 9080 23638 9095 23646
rect 9029 17670 9046 17678
rect 9080 17670 9095 17678
rect 9029 17658 9095 17670
rect 9187 23646 9253 23658
rect 9187 23638 9204 23646
rect 9238 23638 9253 23646
rect 9187 17670 9204 17678
rect 9238 17670 9253 17678
rect 9187 17658 9253 17670
rect 9345 23646 9411 23658
rect 9345 23638 9362 23646
rect 9396 23638 9411 23646
rect 9345 17670 9362 17678
rect 9396 17670 9411 17678
rect 9345 17658 9411 17670
rect 9503 23646 9569 23658
rect 9503 23638 9520 23646
rect 9554 23638 9569 23646
rect 9503 17670 9520 17678
rect 9554 17670 9569 17678
rect 9503 17658 9569 17670
rect 9661 23646 9727 23658
rect 9661 23638 9678 23646
rect 9712 23638 9727 23646
rect 9661 17670 9678 17678
rect 9712 17670 9727 17678
rect 9661 17658 9727 17670
rect 9819 23646 9885 23658
rect 9819 23638 9836 23646
rect 9870 23638 9885 23646
rect 9819 17670 9836 17678
rect 9870 17670 9885 17678
rect 9819 17658 9885 17670
rect 9977 23646 10043 23658
rect 9977 23638 9994 23646
rect 10028 23638 10043 23646
rect 9977 17670 9994 17678
rect 10028 17670 10043 17678
rect 9977 17658 10043 17670
rect 10135 23646 10201 23658
rect 10135 23638 10152 23646
rect 10186 23638 10201 23646
rect 10135 17670 10152 17678
rect 10186 17670 10201 17678
rect 10135 17658 10201 17670
rect 10293 23646 10359 23658
rect 10293 23638 10310 23646
rect 10344 23638 10359 23646
rect 10293 17670 10310 17678
rect 10344 17670 10359 17678
rect 10293 17658 10359 17670
rect 10451 23646 10517 23658
rect 10451 23638 10468 23646
rect 10502 23638 10517 23646
rect 10451 17670 10468 17678
rect 10502 17670 10517 17678
rect 10451 17658 10517 17670
rect 10609 23646 10675 23658
rect 10609 23638 10626 23646
rect 10660 23638 10675 23646
rect 10609 17670 10626 17678
rect 10660 17670 10675 17678
rect 10609 17658 10675 17670
rect 10767 23646 10833 23658
rect 10767 23638 10784 23646
rect 10818 23638 10833 23646
rect 10767 17670 10784 17678
rect 10818 17670 10833 17678
rect 10767 17658 10833 17670
rect 10925 23646 10991 23658
rect 10925 23638 10942 23646
rect 10976 23638 10991 23646
rect 10925 17670 10942 17678
rect 10976 17670 10991 17678
rect 10925 17658 10991 17670
rect 11083 23646 11149 23658
rect 11083 23638 11100 23646
rect 11134 23638 11149 23646
rect 11083 17670 11100 17678
rect 11134 17670 11149 17678
rect 11083 17658 11149 17670
rect 11241 23646 11307 23658
rect 11241 23638 11258 23646
rect 11292 23638 11307 23646
rect 11241 17670 11258 17678
rect 11292 17670 11307 17678
rect 11241 17658 11307 17670
rect 11399 23646 11465 23658
rect 11399 23638 11416 23646
rect 11450 23638 11465 23646
rect 11399 17670 11416 17678
rect 11450 17670 11465 17678
rect 11399 17658 11465 17670
rect 11557 23646 11623 23658
rect 11557 23638 11574 23646
rect 11608 23638 11623 23646
rect 11557 17670 11574 17678
rect 11608 17670 11623 17678
rect 11557 17658 11623 17670
rect 11715 23646 11781 23658
rect 11715 23638 11732 23646
rect 11766 23638 11781 23646
rect 11715 17670 11732 17678
rect 11766 17670 11781 17678
rect 11715 17658 11781 17670
rect 11873 23646 11939 23658
rect 11873 23638 11890 23646
rect 11924 23638 11939 23646
rect 11873 17670 11890 17678
rect 11924 17670 11939 17678
rect 11873 17658 11939 17670
rect 12031 23646 12097 23658
rect 12031 23638 12048 23646
rect 12082 23638 12097 23646
rect 12031 17670 12048 17678
rect 12082 17670 12097 17678
rect 12031 17658 12097 17670
rect 12189 23646 12255 23658
rect 12189 23638 12206 23646
rect 12240 23638 12255 23646
rect 12189 17670 12206 17678
rect 12240 17670 12255 17678
rect 12189 17658 12255 17670
rect 12347 23646 12413 23658
rect 12347 23638 12364 23646
rect 12398 23638 12413 23646
rect 12347 17670 12364 17678
rect 12398 17670 12413 17678
rect 12347 17658 12413 17670
rect 12505 23646 12571 23658
rect 12505 23638 12522 23646
rect 12556 23638 12571 23646
rect 12505 17670 12522 17678
rect 12556 17670 12571 17678
rect 12505 17658 12571 17670
rect 7832 17620 7852 17626
rect 12486 17620 12506 17626
rect 7832 17586 7844 17620
rect 12494 17586 12506 17620
rect 7832 17526 7852 17586
rect 12486 17526 12506 17586
rect 6340 17494 6410 17500
rect 0 17484 6410 17494
rect 0 17480 1536 17484
rect 0 17410 150 17480
rect 350 17410 650 17480
rect 850 17446 1536 17480
rect 6202 17446 6410 17484
rect 850 17430 6410 17446
rect 6500 17480 7500 17500
rect 850 17410 1340 17430
rect 0 17400 1340 17410
rect 0 17380 120 17400
rect 380 17380 620 17400
rect 880 17380 1340 17400
rect 0 17350 100 17380
rect 0 17150 20 17350
rect 90 17150 100 17350
rect 0 17120 100 17150
rect 400 17350 600 17380
rect 400 17150 410 17350
rect 480 17150 520 17350
rect 590 17150 600 17350
rect 400 17120 600 17150
rect 900 17350 1340 17380
rect 900 17150 910 17350
rect 980 17150 1340 17350
rect 900 17120 1340 17150
rect 0 17100 120 17120
rect 380 17100 620 17120
rect 880 17100 1340 17120
rect 0 17090 1340 17100
rect 0 17020 150 17090
rect 350 17020 650 17090
rect 850 17020 1340 17090
rect 0 17000 1340 17020
rect 6500 17410 6650 17480
rect 6850 17410 7150 17480
rect 7350 17410 7500 17480
rect 7630 17494 7700 17500
rect 13930 23870 19010 23880
rect 13930 23832 14136 23870
rect 18859 23832 19010 23870
rect 13930 23822 19010 23832
rect 13930 23820 14000 23822
rect 18940 23820 19010 23822
rect 14132 23730 14152 23790
rect 18786 23730 18806 23790
rect 14132 23696 14144 23730
rect 18794 23696 18806 23730
rect 14132 23690 14152 23696
rect 18786 23690 18806 23696
rect 14065 23646 14131 23658
rect 14065 23638 14082 23646
rect 14116 23638 14131 23646
rect 14065 17670 14082 17678
rect 14116 17670 14131 17678
rect 14065 17658 14131 17670
rect 14223 23646 14289 23658
rect 14223 23638 14240 23646
rect 14274 23638 14289 23646
rect 14223 17670 14240 17678
rect 14274 17670 14289 17678
rect 14223 17658 14289 17670
rect 14381 23646 14447 23658
rect 14381 23638 14398 23646
rect 14432 23638 14447 23646
rect 14381 17670 14398 17678
rect 14432 17670 14447 17678
rect 14381 17658 14447 17670
rect 14539 23646 14605 23658
rect 14539 23638 14556 23646
rect 14590 23638 14605 23646
rect 14539 17670 14556 17678
rect 14590 17670 14605 17678
rect 14539 17658 14605 17670
rect 14697 23646 14763 23658
rect 14697 23638 14714 23646
rect 14748 23638 14763 23646
rect 14697 17670 14714 17678
rect 14748 17670 14763 17678
rect 14697 17658 14763 17670
rect 14855 23646 14921 23658
rect 14855 23638 14872 23646
rect 14906 23638 14921 23646
rect 14855 17670 14872 17678
rect 14906 17670 14921 17678
rect 14855 17658 14921 17670
rect 15013 23646 15079 23658
rect 15013 23638 15030 23646
rect 15064 23638 15079 23646
rect 15013 17670 15030 17678
rect 15064 17670 15079 17678
rect 15013 17658 15079 17670
rect 15171 23646 15237 23658
rect 15171 23638 15188 23646
rect 15222 23638 15237 23646
rect 15171 17670 15188 17678
rect 15222 17670 15237 17678
rect 15171 17658 15237 17670
rect 15329 23646 15395 23658
rect 15329 23638 15346 23646
rect 15380 23638 15395 23646
rect 15329 17670 15346 17678
rect 15380 17670 15395 17678
rect 15329 17658 15395 17670
rect 15487 23646 15553 23658
rect 15487 23638 15504 23646
rect 15538 23638 15553 23646
rect 15487 17670 15504 17678
rect 15538 17670 15553 17678
rect 15487 17658 15553 17670
rect 15645 23646 15711 23658
rect 15645 23638 15662 23646
rect 15696 23638 15711 23646
rect 15645 17670 15662 17678
rect 15696 17670 15711 17678
rect 15645 17658 15711 17670
rect 15803 23646 15869 23658
rect 15803 23638 15820 23646
rect 15854 23638 15869 23646
rect 15803 17670 15820 17678
rect 15854 17670 15869 17678
rect 15803 17658 15869 17670
rect 15961 23646 16027 23658
rect 15961 23638 15978 23646
rect 16012 23638 16027 23646
rect 15961 17670 15978 17678
rect 16012 17670 16027 17678
rect 15961 17658 16027 17670
rect 16119 23646 16185 23658
rect 16119 23638 16136 23646
rect 16170 23638 16185 23646
rect 16119 17670 16136 17678
rect 16170 17670 16185 17678
rect 16119 17658 16185 17670
rect 16277 23646 16343 23658
rect 16277 23638 16294 23646
rect 16328 23638 16343 23646
rect 16277 17670 16294 17678
rect 16328 17670 16343 17678
rect 16277 17658 16343 17670
rect 16435 23646 16501 23658
rect 16435 23638 16452 23646
rect 16486 23638 16501 23646
rect 16435 17670 16452 17678
rect 16486 17670 16501 17678
rect 16435 17658 16501 17670
rect 16593 23646 16659 23658
rect 16593 23638 16610 23646
rect 16644 23638 16659 23646
rect 16593 17670 16610 17678
rect 16644 17670 16659 17678
rect 16593 17658 16659 17670
rect 16751 23646 16817 23658
rect 16751 23638 16768 23646
rect 16802 23638 16817 23646
rect 16751 17670 16768 17678
rect 16802 17670 16817 17678
rect 16751 17658 16817 17670
rect 16909 23646 16975 23658
rect 16909 23638 16926 23646
rect 16960 23638 16975 23646
rect 16909 17670 16926 17678
rect 16960 17670 16975 17678
rect 16909 17658 16975 17670
rect 17067 23646 17133 23658
rect 17067 23638 17084 23646
rect 17118 23638 17133 23646
rect 17067 17670 17084 17678
rect 17118 17670 17133 17678
rect 17067 17658 17133 17670
rect 17225 23646 17291 23658
rect 17225 23638 17242 23646
rect 17276 23638 17291 23646
rect 17225 17670 17242 17678
rect 17276 17670 17291 17678
rect 17225 17658 17291 17670
rect 17383 23646 17449 23658
rect 17383 23638 17400 23646
rect 17434 23638 17449 23646
rect 17383 17670 17400 17678
rect 17434 17670 17449 17678
rect 17383 17658 17449 17670
rect 17541 23646 17607 23658
rect 17541 23638 17558 23646
rect 17592 23638 17607 23646
rect 17541 17670 17558 17678
rect 17592 17670 17607 17678
rect 17541 17658 17607 17670
rect 17699 23646 17765 23658
rect 17699 23638 17716 23646
rect 17750 23638 17765 23646
rect 17699 17670 17716 17678
rect 17750 17670 17765 17678
rect 17699 17658 17765 17670
rect 17857 23646 17923 23658
rect 17857 23638 17874 23646
rect 17908 23638 17923 23646
rect 17857 17670 17874 17678
rect 17908 17670 17923 17678
rect 17857 17658 17923 17670
rect 18015 23646 18081 23658
rect 18015 23638 18032 23646
rect 18066 23638 18081 23646
rect 18015 17670 18032 17678
rect 18066 17670 18081 17678
rect 18015 17658 18081 17670
rect 18173 23646 18239 23658
rect 18173 23638 18190 23646
rect 18224 23638 18239 23646
rect 18173 17670 18190 17678
rect 18224 17670 18239 17678
rect 18173 17658 18239 17670
rect 18331 23646 18397 23658
rect 18331 23638 18348 23646
rect 18382 23638 18397 23646
rect 18331 17670 18348 17678
rect 18382 17670 18397 17678
rect 18331 17658 18397 17670
rect 18489 23646 18555 23658
rect 18489 23638 18506 23646
rect 18540 23638 18555 23646
rect 18489 17670 18506 17678
rect 18540 17670 18555 17678
rect 18489 17658 18555 17670
rect 18647 23646 18713 23658
rect 18647 23638 18664 23646
rect 18698 23638 18713 23646
rect 18647 17670 18664 17678
rect 18698 17670 18713 17678
rect 18647 17658 18713 17670
rect 18805 23646 18871 23658
rect 18805 23638 18822 23646
rect 18856 23638 18871 23646
rect 18805 17670 18822 17678
rect 18856 17670 18871 17678
rect 18805 17658 18871 17670
rect 14132 17620 14152 17626
rect 18786 17620 18806 17626
rect 14132 17586 14144 17620
rect 18794 17586 18806 17620
rect 14132 17526 14152 17586
rect 18786 17526 18806 17586
rect 12640 17494 12710 17500
rect 7630 17484 12710 17494
rect 7630 17446 7836 17484
rect 12502 17446 12710 17484
rect 7630 17430 12710 17446
rect 13000 17494 14000 17500
rect 20230 23870 25600 23880
rect 20230 23832 20436 23870
rect 25159 23850 25600 23870
rect 25159 23832 25520 23850
rect 20230 23822 25520 23832
rect 20230 23820 20300 23822
rect 25240 23820 25520 23822
rect 20432 23730 20452 23790
rect 25086 23730 25106 23790
rect 20432 23696 20444 23730
rect 25094 23696 25106 23730
rect 20432 23690 20452 23696
rect 25086 23690 25106 23696
rect 20365 23646 20431 23658
rect 20365 23638 20382 23646
rect 20416 23638 20431 23646
rect 20365 17670 20382 17678
rect 20416 17670 20431 17678
rect 20365 17658 20431 17670
rect 20523 23646 20589 23658
rect 20523 23638 20540 23646
rect 20574 23638 20589 23646
rect 20523 17670 20540 17678
rect 20574 17670 20589 17678
rect 20523 17658 20589 17670
rect 20681 23646 20747 23658
rect 20681 23638 20698 23646
rect 20732 23638 20747 23646
rect 20681 17670 20698 17678
rect 20732 17670 20747 17678
rect 20681 17658 20747 17670
rect 20839 23646 20905 23658
rect 20839 23638 20856 23646
rect 20890 23638 20905 23646
rect 20839 17670 20856 17678
rect 20890 17670 20905 17678
rect 20839 17658 20905 17670
rect 20997 23646 21063 23658
rect 20997 23638 21014 23646
rect 21048 23638 21063 23646
rect 20997 17670 21014 17678
rect 21048 17670 21063 17678
rect 20997 17658 21063 17670
rect 21155 23646 21221 23658
rect 21155 23638 21172 23646
rect 21206 23638 21221 23646
rect 21155 17670 21172 17678
rect 21206 17670 21221 17678
rect 21155 17658 21221 17670
rect 21313 23646 21379 23658
rect 21313 23638 21330 23646
rect 21364 23638 21379 23646
rect 21313 17670 21330 17678
rect 21364 17670 21379 17678
rect 21313 17658 21379 17670
rect 21471 23646 21537 23658
rect 21471 23638 21488 23646
rect 21522 23638 21537 23646
rect 21471 17670 21488 17678
rect 21522 17670 21537 17678
rect 21471 17658 21537 17670
rect 21629 23646 21695 23658
rect 21629 23638 21646 23646
rect 21680 23638 21695 23646
rect 21629 17670 21646 17678
rect 21680 17670 21695 17678
rect 21629 17658 21695 17670
rect 21787 23646 21853 23658
rect 21787 23638 21804 23646
rect 21838 23638 21853 23646
rect 21787 17670 21804 17678
rect 21838 17670 21853 17678
rect 21787 17658 21853 17670
rect 21945 23646 22011 23658
rect 21945 23638 21962 23646
rect 21996 23638 22011 23646
rect 21945 17670 21962 17678
rect 21996 17670 22011 17678
rect 21945 17658 22011 17670
rect 22103 23646 22169 23658
rect 22103 23638 22120 23646
rect 22154 23638 22169 23646
rect 22103 17670 22120 17678
rect 22154 17670 22169 17678
rect 22103 17658 22169 17670
rect 22261 23646 22327 23658
rect 22261 23638 22278 23646
rect 22312 23638 22327 23646
rect 22261 17670 22278 17678
rect 22312 17670 22327 17678
rect 22261 17658 22327 17670
rect 22419 23646 22485 23658
rect 22419 23638 22436 23646
rect 22470 23638 22485 23646
rect 22419 17670 22436 17678
rect 22470 17670 22485 17678
rect 22419 17658 22485 17670
rect 22577 23646 22643 23658
rect 22577 23638 22594 23646
rect 22628 23638 22643 23646
rect 22577 17670 22594 17678
rect 22628 17670 22643 17678
rect 22577 17658 22643 17670
rect 22735 23646 22801 23658
rect 22735 23638 22752 23646
rect 22786 23638 22801 23646
rect 22735 17670 22752 17678
rect 22786 17670 22801 17678
rect 22735 17658 22801 17670
rect 22893 23646 22959 23658
rect 22893 23638 22910 23646
rect 22944 23638 22959 23646
rect 22893 17670 22910 17678
rect 22944 17670 22959 17678
rect 22893 17658 22959 17670
rect 23051 23646 23117 23658
rect 23051 23638 23068 23646
rect 23102 23638 23117 23646
rect 23051 17670 23068 17678
rect 23102 17670 23117 17678
rect 23051 17658 23117 17670
rect 23209 23646 23275 23658
rect 23209 23638 23226 23646
rect 23260 23638 23275 23646
rect 23209 17670 23226 17678
rect 23260 17670 23275 17678
rect 23209 17658 23275 17670
rect 23367 23646 23433 23658
rect 23367 23638 23384 23646
rect 23418 23638 23433 23646
rect 23367 17670 23384 17678
rect 23418 17670 23433 17678
rect 23367 17658 23433 17670
rect 23525 23646 23591 23658
rect 23525 23638 23542 23646
rect 23576 23638 23591 23646
rect 23525 17670 23542 17678
rect 23576 17670 23591 17678
rect 23525 17658 23591 17670
rect 23683 23646 23749 23658
rect 23683 23638 23700 23646
rect 23734 23638 23749 23646
rect 23683 17670 23700 17678
rect 23734 17670 23749 17678
rect 23683 17658 23749 17670
rect 23841 23646 23907 23658
rect 23841 23638 23858 23646
rect 23892 23638 23907 23646
rect 23841 17670 23858 17678
rect 23892 17670 23907 17678
rect 23841 17658 23907 17670
rect 23999 23646 24065 23658
rect 23999 23638 24016 23646
rect 24050 23638 24065 23646
rect 23999 17670 24016 17678
rect 24050 17670 24065 17678
rect 23999 17658 24065 17670
rect 24157 23646 24223 23658
rect 24157 23638 24174 23646
rect 24208 23638 24223 23646
rect 24157 17670 24174 17678
rect 24208 17670 24223 17678
rect 24157 17658 24223 17670
rect 24315 23646 24381 23658
rect 24315 23638 24332 23646
rect 24366 23638 24381 23646
rect 24315 17670 24332 17678
rect 24366 17670 24381 17678
rect 24315 17658 24381 17670
rect 24473 23646 24539 23658
rect 24473 23638 24490 23646
rect 24524 23638 24539 23646
rect 24473 17670 24490 17678
rect 24524 17670 24539 17678
rect 24473 17658 24539 17670
rect 24631 23646 24697 23658
rect 24631 23638 24648 23646
rect 24682 23638 24697 23646
rect 24631 17670 24648 17678
rect 24682 17670 24697 17678
rect 24631 17658 24697 17670
rect 24789 23646 24855 23658
rect 24789 23638 24806 23646
rect 24840 23638 24855 23646
rect 24789 17670 24806 17678
rect 24840 17670 24855 17678
rect 24789 17658 24855 17670
rect 24947 23646 25013 23658
rect 24947 23638 24964 23646
rect 24998 23638 25013 23646
rect 24947 17670 24964 17678
rect 24998 17670 25013 17678
rect 24947 17658 25013 17670
rect 25105 23646 25171 23658
rect 25105 23638 25122 23646
rect 25156 23638 25171 23646
rect 25105 17670 25122 17678
rect 25156 17670 25171 17678
rect 25105 17658 25171 17670
rect 25310 23650 25520 23820
rect 25590 23650 25600 23850
rect 25310 23620 25600 23650
rect 25900 23850 26100 23880
rect 25900 23650 25910 23850
rect 25980 23650 26020 23850
rect 26090 23650 26100 23850
rect 25900 23620 26100 23650
rect 26400 23850 26500 23880
rect 26400 23650 26410 23850
rect 26480 23650 26500 23850
rect 26400 23620 26500 23650
rect 25310 23600 25620 23620
rect 25880 23600 26120 23620
rect 26380 23600 26500 23620
rect 25310 23590 26500 23600
rect 25310 23520 25650 23590
rect 25850 23520 26150 23590
rect 26350 23520 26500 23590
rect 25310 23480 26500 23520
rect 25310 23410 25650 23480
rect 25850 23410 26150 23480
rect 26350 23410 26500 23480
rect 25310 23400 26500 23410
rect 25310 23380 25620 23400
rect 25880 23380 26120 23400
rect 26380 23380 26500 23400
rect 25310 23350 25600 23380
rect 25310 23150 25520 23350
rect 25590 23150 25600 23350
rect 25310 23120 25600 23150
rect 25900 23350 26100 23380
rect 25900 23150 25910 23350
rect 25980 23150 26020 23350
rect 26090 23150 26100 23350
rect 25900 23120 26100 23150
rect 26400 23350 26500 23380
rect 26400 23150 26410 23350
rect 26480 23150 26500 23350
rect 26400 23120 26500 23150
rect 25310 23100 25620 23120
rect 25880 23100 26120 23120
rect 26380 23100 26500 23120
rect 25310 23090 26500 23100
rect 25310 23020 25650 23090
rect 25850 23020 26150 23090
rect 26350 23020 26500 23090
rect 25310 22980 26500 23020
rect 25310 22910 25650 22980
rect 25850 22910 26150 22980
rect 26350 22910 26500 22980
rect 25310 22900 26500 22910
rect 25310 22880 25620 22900
rect 25880 22880 26120 22900
rect 26380 22880 26500 22900
rect 25310 22850 25600 22880
rect 25310 22650 25520 22850
rect 25590 22650 25600 22850
rect 25310 22620 25600 22650
rect 25900 22850 26100 22880
rect 25900 22650 25910 22850
rect 25980 22650 26020 22850
rect 26090 22650 26100 22850
rect 25900 22620 26100 22650
rect 26400 22850 26500 22880
rect 26400 22650 26410 22850
rect 26480 22650 26500 22850
rect 26400 22620 26500 22650
rect 25310 22600 25620 22620
rect 25880 22600 26120 22620
rect 26380 22600 26500 22620
rect 25310 22590 26500 22600
rect 25310 22520 25650 22590
rect 25850 22520 26150 22590
rect 26350 22520 26500 22590
rect 25310 22480 26500 22520
rect 25310 22410 25650 22480
rect 25850 22410 26150 22480
rect 26350 22410 26500 22480
rect 25310 22400 26500 22410
rect 25310 22380 25620 22400
rect 25880 22380 26120 22400
rect 26380 22380 26500 22400
rect 25310 22350 25600 22380
rect 25310 22150 25520 22350
rect 25590 22150 25600 22350
rect 25310 22120 25600 22150
rect 25900 22350 26100 22380
rect 25900 22150 25910 22350
rect 25980 22150 26020 22350
rect 26090 22150 26100 22350
rect 25900 22120 26100 22150
rect 26400 22350 26500 22380
rect 26400 22150 26410 22350
rect 26480 22150 26500 22350
rect 26400 22120 26500 22150
rect 25310 22100 25620 22120
rect 25880 22100 26120 22120
rect 26380 22100 26500 22120
rect 25310 22090 26500 22100
rect 25310 22020 25650 22090
rect 25850 22020 26150 22090
rect 26350 22020 26500 22090
rect 25310 21980 26500 22020
rect 25310 21910 25650 21980
rect 25850 21910 26150 21980
rect 26350 21910 26500 21980
rect 25310 21900 26500 21910
rect 25310 21880 25620 21900
rect 25880 21880 26120 21900
rect 26380 21880 26500 21900
rect 25310 21850 25600 21880
rect 25310 21650 25520 21850
rect 25590 21650 25600 21850
rect 25310 21620 25600 21650
rect 25900 21850 26100 21880
rect 25900 21650 25910 21850
rect 25980 21650 26020 21850
rect 26090 21650 26100 21850
rect 25900 21620 26100 21650
rect 26400 21850 26500 21880
rect 26400 21650 26410 21850
rect 26480 21650 26500 21850
rect 26400 21620 26500 21650
rect 25310 21600 25620 21620
rect 25880 21600 26120 21620
rect 26380 21600 26500 21620
rect 25310 21590 26500 21600
rect 25310 21520 25650 21590
rect 25850 21520 26150 21590
rect 26350 21520 26500 21590
rect 25310 21480 26500 21520
rect 25310 21410 25650 21480
rect 25850 21410 26150 21480
rect 26350 21410 26500 21480
rect 25310 21400 26500 21410
rect 25310 21380 25620 21400
rect 25880 21380 26120 21400
rect 26380 21380 26500 21400
rect 25310 21350 25600 21380
rect 25310 21150 25520 21350
rect 25590 21150 25600 21350
rect 25310 21120 25600 21150
rect 25900 21350 26100 21380
rect 25900 21150 25910 21350
rect 25980 21150 26020 21350
rect 26090 21150 26100 21350
rect 25900 21120 26100 21150
rect 26400 21350 26500 21380
rect 26400 21150 26410 21350
rect 26480 21150 26500 21350
rect 26400 21120 26500 21150
rect 25310 21100 25620 21120
rect 25880 21100 26120 21120
rect 26380 21100 26500 21120
rect 25310 21090 26500 21100
rect 25310 21020 25650 21090
rect 25850 21020 26150 21090
rect 26350 21020 26500 21090
rect 25310 20980 26500 21020
rect 25310 20910 25650 20980
rect 25850 20910 26150 20980
rect 26350 20910 26500 20980
rect 25310 20900 26500 20910
rect 25310 20880 25620 20900
rect 25880 20880 26120 20900
rect 26380 20880 26500 20900
rect 25310 20850 25600 20880
rect 25310 20650 25520 20850
rect 25590 20650 25600 20850
rect 25310 20620 25600 20650
rect 25900 20850 26100 20880
rect 25900 20650 25910 20850
rect 25980 20650 26020 20850
rect 26090 20650 26100 20850
rect 25900 20620 26100 20650
rect 26400 20850 26500 20880
rect 26400 20650 26410 20850
rect 26480 20650 26500 20850
rect 26400 20620 26500 20650
rect 25310 20600 25620 20620
rect 25880 20600 26120 20620
rect 26380 20600 26500 20620
rect 25310 20590 26500 20600
rect 25310 20520 25650 20590
rect 25850 20520 26150 20590
rect 26350 20520 26500 20590
rect 25310 20480 26500 20520
rect 25310 20410 25650 20480
rect 25850 20410 26150 20480
rect 26350 20410 26500 20480
rect 25310 20400 26500 20410
rect 25310 20380 25620 20400
rect 25880 20380 26120 20400
rect 26380 20380 26500 20400
rect 25310 20350 25600 20380
rect 25310 20150 25520 20350
rect 25590 20150 25600 20350
rect 25310 20120 25600 20150
rect 25900 20350 26100 20380
rect 25900 20150 25910 20350
rect 25980 20150 26020 20350
rect 26090 20150 26100 20350
rect 25900 20120 26100 20150
rect 26400 20350 26500 20380
rect 26400 20150 26410 20350
rect 26480 20150 26500 20350
rect 26400 20120 26500 20150
rect 25310 20100 25620 20120
rect 25880 20100 26120 20120
rect 26380 20100 26500 20120
rect 25310 20090 26500 20100
rect 25310 20020 25650 20090
rect 25850 20020 26150 20090
rect 26350 20020 26500 20090
rect 25310 19980 26500 20020
rect 25310 19910 25650 19980
rect 25850 19910 26150 19980
rect 26350 19910 26500 19980
rect 25310 19900 26500 19910
rect 25310 19880 25620 19900
rect 25880 19880 26120 19900
rect 26380 19880 26500 19900
rect 25310 19850 25600 19880
rect 25310 19650 25520 19850
rect 25590 19650 25600 19850
rect 25310 19620 25600 19650
rect 25900 19850 26100 19880
rect 25900 19650 25910 19850
rect 25980 19650 26020 19850
rect 26090 19650 26100 19850
rect 25900 19620 26100 19650
rect 26400 19850 26500 19880
rect 26400 19650 26410 19850
rect 26480 19650 26500 19850
rect 26400 19620 26500 19650
rect 25310 19600 25620 19620
rect 25880 19600 26120 19620
rect 26380 19600 26500 19620
rect 25310 19590 26500 19600
rect 25310 19520 25650 19590
rect 25850 19520 26150 19590
rect 26350 19520 26500 19590
rect 25310 19480 26500 19520
rect 25310 19410 25650 19480
rect 25850 19410 26150 19480
rect 26350 19410 26500 19480
rect 25310 19400 26500 19410
rect 25310 19380 25620 19400
rect 25880 19380 26120 19400
rect 26380 19380 26500 19400
rect 25310 19350 25600 19380
rect 25310 19150 25520 19350
rect 25590 19150 25600 19350
rect 25310 19120 25600 19150
rect 25900 19350 26100 19380
rect 25900 19150 25910 19350
rect 25980 19150 26020 19350
rect 26090 19150 26100 19350
rect 25900 19120 26100 19150
rect 26400 19350 26500 19380
rect 26400 19150 26410 19350
rect 26480 19150 26500 19350
rect 26400 19120 26500 19150
rect 25310 19100 25620 19120
rect 25880 19100 26120 19120
rect 26380 19100 26500 19120
rect 25310 19090 26500 19100
rect 25310 19020 25650 19090
rect 25850 19020 26150 19090
rect 26350 19020 26500 19090
rect 25310 18980 26500 19020
rect 25310 18910 25650 18980
rect 25850 18910 26150 18980
rect 26350 18910 26500 18980
rect 25310 18900 26500 18910
rect 25310 18880 25620 18900
rect 25880 18880 26120 18900
rect 26380 18880 26500 18900
rect 25310 18850 25600 18880
rect 25310 18650 25520 18850
rect 25590 18650 25600 18850
rect 25310 18620 25600 18650
rect 25900 18850 26100 18880
rect 25900 18650 25910 18850
rect 25980 18650 26020 18850
rect 26090 18650 26100 18850
rect 25900 18620 26100 18650
rect 26400 18850 26500 18880
rect 26400 18650 26410 18850
rect 26480 18650 26500 18850
rect 26400 18620 26500 18650
rect 25310 18600 25620 18620
rect 25880 18600 26120 18620
rect 26380 18600 26500 18620
rect 25310 18590 26500 18600
rect 25310 18520 25650 18590
rect 25850 18520 26150 18590
rect 26350 18520 26500 18590
rect 25310 18480 26500 18520
rect 25310 18410 25650 18480
rect 25850 18410 26150 18480
rect 26350 18410 26500 18480
rect 25310 18400 26500 18410
rect 25310 18380 25620 18400
rect 25880 18380 26120 18400
rect 26380 18380 26500 18400
rect 25310 18350 25600 18380
rect 25310 18150 25520 18350
rect 25590 18150 25600 18350
rect 25310 18120 25600 18150
rect 25900 18350 26100 18380
rect 25900 18150 25910 18350
rect 25980 18150 26020 18350
rect 26090 18150 26100 18350
rect 25900 18120 26100 18150
rect 26400 18350 26500 18380
rect 26400 18150 26410 18350
rect 26480 18150 26500 18350
rect 26400 18120 26500 18150
rect 25310 18100 25620 18120
rect 25880 18100 26120 18120
rect 26380 18100 26500 18120
rect 25310 18090 26500 18100
rect 25310 18020 25650 18090
rect 25850 18020 26150 18090
rect 26350 18020 26500 18090
rect 25310 17980 26500 18020
rect 25310 17910 25650 17980
rect 25850 17910 26150 17980
rect 26350 17910 26500 17980
rect 25310 17900 26500 17910
rect 25310 17880 25620 17900
rect 25880 17880 26120 17900
rect 26380 17880 26500 17900
rect 25310 17850 25600 17880
rect 25310 17650 25520 17850
rect 25590 17650 25600 17850
rect 20432 17620 20452 17626
rect 25086 17620 25106 17626
rect 20432 17586 20444 17620
rect 25094 17586 25106 17620
rect 20432 17526 20452 17586
rect 25086 17526 25106 17586
rect 18940 17494 20000 17500
rect 13000 17484 20000 17494
rect 13000 17480 14136 17484
rect 6500 17400 7500 17410
rect 6500 17380 6620 17400
rect 6880 17380 7120 17400
rect 7380 17380 7500 17400
rect 6500 17350 6600 17380
rect 6500 17150 6520 17350
rect 6590 17150 6600 17350
rect 6500 17120 6600 17150
rect 6900 17350 7100 17380
rect 6900 17150 6910 17350
rect 6980 17150 7020 17350
rect 7090 17150 7100 17350
rect 6900 17120 7100 17150
rect 7400 17350 7500 17380
rect 7400 17150 7410 17350
rect 7480 17150 7500 17350
rect 7400 17120 7500 17150
rect 6500 17100 6620 17120
rect 6880 17100 7120 17120
rect 7380 17100 7500 17120
rect 6500 17090 7500 17100
rect 6500 17020 6650 17090
rect 6850 17020 7150 17090
rect 7350 17020 7500 17090
rect 6500 17000 7500 17020
rect 13000 17410 13150 17480
rect 13350 17410 13650 17480
rect 13850 17446 14136 17480
rect 18802 17480 20000 17484
rect 18802 17446 19150 17480
rect 13850 17430 19150 17446
rect 13850 17410 14000 17430
rect 13000 17400 14000 17410
rect 13000 17380 13120 17400
rect 13380 17380 13620 17400
rect 13880 17380 14000 17400
rect 13000 17350 13100 17380
rect 13000 17150 13020 17350
rect 13090 17150 13100 17350
rect 13000 17120 13100 17150
rect 13400 17350 13600 17380
rect 13400 17150 13410 17350
rect 13480 17150 13520 17350
rect 13590 17150 13600 17350
rect 13400 17120 13600 17150
rect 13900 17350 14000 17380
rect 13900 17150 13910 17350
rect 13980 17150 14000 17350
rect 13900 17120 14000 17150
rect 13000 17100 13120 17120
rect 13380 17100 13620 17120
rect 13880 17100 14000 17120
rect 13000 17090 14000 17100
rect 13000 17020 13150 17090
rect 13350 17020 13650 17090
rect 13850 17020 14000 17090
rect 13000 17000 14000 17020
rect 19000 17410 19150 17430
rect 19350 17410 19650 17480
rect 19850 17410 20000 17480
rect 20230 17494 20300 17500
rect 25310 17620 25600 17650
rect 25900 17850 26100 17880
rect 25900 17650 25910 17850
rect 25980 17650 26020 17850
rect 26090 17650 26100 17850
rect 25900 17620 26100 17650
rect 26400 17850 26500 17880
rect 26400 17650 26410 17850
rect 26480 17650 26500 17850
rect 26400 17620 26500 17650
rect 25310 17600 25620 17620
rect 25880 17600 26120 17620
rect 26380 17600 26500 17620
rect 25310 17590 26500 17600
rect 25310 17520 25650 17590
rect 25850 17520 26150 17590
rect 26350 17520 26500 17590
rect 25310 17500 26500 17520
rect 25240 17494 26500 17500
rect 20230 17484 26500 17494
rect 20230 17446 20436 17484
rect 25102 17480 26500 17484
rect 25102 17446 25650 17480
rect 20230 17430 25650 17446
rect 19000 17400 20000 17410
rect 19000 17380 19120 17400
rect 19380 17380 19620 17400
rect 19880 17380 20000 17400
rect 19000 17350 19100 17380
rect 19000 17150 19020 17350
rect 19090 17150 19100 17350
rect 19000 17120 19100 17150
rect 19400 17350 19600 17380
rect 19400 17150 19410 17350
rect 19480 17150 19520 17350
rect 19590 17150 19600 17350
rect 19400 17120 19600 17150
rect 19900 17350 20000 17380
rect 19900 17150 19910 17350
rect 19980 17150 20000 17350
rect 19900 17120 20000 17150
rect 19000 17100 19120 17120
rect 19380 17100 19620 17120
rect 19880 17100 20000 17120
rect 19000 17090 20000 17100
rect 19000 17020 19150 17090
rect 19350 17020 19650 17090
rect 19850 17020 20000 17090
rect 19000 17000 20000 17020
rect 25260 17410 25650 17430
rect 25850 17410 26150 17480
rect 26350 17410 26500 17480
rect 25260 17400 26500 17410
rect 25260 17380 25620 17400
rect 25880 17380 26120 17400
rect 26380 17380 26500 17400
rect 25260 17350 25600 17380
rect 25260 17150 25520 17350
rect 25590 17150 25600 17350
rect 25260 17120 25600 17150
rect 25900 17350 26100 17380
rect 25900 17150 25910 17350
rect 25980 17150 26020 17350
rect 26090 17150 26100 17350
rect 25900 17120 26100 17150
rect 26400 17350 26500 17380
rect 26400 17150 26410 17350
rect 26480 17150 26500 17350
rect 26400 17120 26500 17150
rect 25260 17100 25620 17120
rect 25880 17100 26120 17120
rect 26380 17100 26500 17120
rect 25260 17090 26500 17100
rect 25260 17020 25650 17090
rect 25850 17020 26150 17090
rect 26350 17020 26500 17090
rect 25260 17000 26500 17020
rect 0 16980 26500 17000
rect 0 16910 150 16980
rect 350 16910 650 16980
rect 850 16910 1150 16980
rect 1350 16910 1650 16980
rect 1850 16910 2150 16980
rect 2350 16910 2650 16980
rect 2850 16910 3150 16980
rect 3350 16910 3650 16980
rect 3850 16910 4150 16980
rect 4350 16910 4650 16980
rect 4850 16910 5150 16980
rect 5350 16910 5650 16980
rect 5850 16910 6150 16980
rect 6350 16910 6650 16980
rect 6850 16910 7150 16980
rect 7350 16910 7650 16980
rect 7850 16910 8150 16980
rect 8350 16910 8650 16980
rect 8850 16910 9150 16980
rect 9350 16910 9650 16980
rect 9850 16910 10150 16980
rect 10350 16910 10650 16980
rect 10850 16910 11150 16980
rect 11350 16910 11650 16980
rect 11850 16910 12150 16980
rect 12350 16910 12650 16980
rect 12850 16910 13150 16980
rect 13350 16910 13650 16980
rect 13850 16910 14150 16980
rect 14350 16910 14650 16980
rect 14850 16910 15150 16980
rect 15350 16910 15650 16980
rect 15850 16910 16150 16980
rect 16350 16910 16650 16980
rect 16850 16910 17150 16980
rect 17350 16910 17650 16980
rect 17850 16910 18150 16980
rect 18350 16910 18650 16980
rect 18850 16910 19150 16980
rect 19350 16910 19650 16980
rect 19850 16910 20150 16980
rect 20350 16910 20650 16980
rect 20850 16910 21150 16980
rect 21350 16910 21650 16980
rect 21850 16910 22150 16980
rect 22350 16910 22650 16980
rect 22850 16910 23150 16980
rect 23350 16910 23650 16980
rect 23850 16910 24150 16980
rect 24350 16910 24650 16980
rect 24850 16910 25150 16980
rect 25350 16910 25650 16980
rect 25850 16910 26150 16980
rect 26350 16910 26500 16980
rect 0 16900 26500 16910
rect 0 16880 120 16900
rect 380 16880 620 16900
rect 880 16880 1120 16900
rect 1380 16880 1620 16900
rect 1880 16880 2120 16900
rect 2380 16880 2620 16900
rect 2880 16880 3120 16900
rect 3380 16880 3620 16900
rect 3880 16880 4120 16900
rect 4380 16880 4620 16900
rect 4880 16880 5120 16900
rect 5380 16880 5620 16900
rect 5880 16880 6120 16900
rect 6380 16880 6620 16900
rect 6880 16880 7120 16900
rect 7380 16880 7620 16900
rect 7880 16880 8120 16900
rect 8380 16880 8620 16900
rect 8880 16880 9120 16900
rect 9380 16880 9620 16900
rect 9880 16880 10120 16900
rect 10380 16880 10620 16900
rect 10880 16880 11120 16900
rect 11380 16880 11620 16900
rect 11880 16880 12120 16900
rect 12380 16880 12620 16900
rect 12880 16880 13120 16900
rect 13380 16880 13620 16900
rect 13880 16880 14120 16900
rect 14380 16880 14620 16900
rect 14880 16880 15120 16900
rect 15380 16880 15620 16900
rect 15880 16880 16120 16900
rect 16380 16880 16620 16900
rect 16880 16880 17120 16900
rect 17380 16880 17620 16900
rect 17880 16880 18120 16900
rect 18380 16880 18620 16900
rect 18880 16880 19120 16900
rect 19380 16880 19620 16900
rect 19880 16880 20120 16900
rect 20380 16880 20620 16900
rect 20880 16880 21120 16900
rect 21380 16880 21620 16900
rect 21880 16880 22120 16900
rect 22380 16880 22620 16900
rect 22880 16880 23120 16900
rect 23380 16880 23620 16900
rect 23880 16880 24120 16900
rect 24380 16880 24620 16900
rect 24880 16880 25120 16900
rect 25380 16880 25620 16900
rect 25880 16880 26120 16900
rect 26380 16880 26500 16900
rect 0 16850 100 16880
rect 0 16650 20 16850
rect 90 16650 100 16850
rect 0 16620 100 16650
rect 400 16850 600 16880
rect 400 16650 410 16850
rect 480 16650 520 16850
rect 590 16650 600 16850
rect 400 16620 600 16650
rect 900 16850 1100 16880
rect 900 16650 910 16850
rect 980 16650 1020 16850
rect 1090 16650 1100 16850
rect 900 16620 1100 16650
rect 1400 16850 1600 16880
rect 1400 16650 1410 16850
rect 1480 16650 1520 16850
rect 1590 16650 1600 16850
rect 1400 16620 1600 16650
rect 1900 16850 2100 16880
rect 1900 16650 1910 16850
rect 1980 16650 2020 16850
rect 2090 16650 2100 16850
rect 1900 16620 2100 16650
rect 2400 16850 2600 16880
rect 2400 16650 2410 16850
rect 2480 16650 2520 16850
rect 2590 16650 2600 16850
rect 2400 16620 2600 16650
rect 2900 16850 3100 16880
rect 2900 16650 2910 16850
rect 2980 16650 3020 16850
rect 3090 16650 3100 16850
rect 2900 16620 3100 16650
rect 3400 16850 3600 16880
rect 3400 16650 3410 16850
rect 3480 16650 3520 16850
rect 3590 16650 3600 16850
rect 3400 16620 3600 16650
rect 3900 16850 4100 16880
rect 3900 16650 3910 16850
rect 3980 16650 4020 16850
rect 4090 16650 4100 16850
rect 3900 16620 4100 16650
rect 4400 16850 4600 16880
rect 4400 16650 4410 16850
rect 4480 16650 4520 16850
rect 4590 16650 4600 16850
rect 4400 16620 4600 16650
rect 4900 16850 5100 16880
rect 4900 16650 4910 16850
rect 4980 16650 5020 16850
rect 5090 16650 5100 16850
rect 4900 16620 5100 16650
rect 5400 16850 5600 16880
rect 5400 16650 5410 16850
rect 5480 16650 5520 16850
rect 5590 16650 5600 16850
rect 5400 16620 5600 16650
rect 5900 16850 6100 16880
rect 5900 16650 5910 16850
rect 5980 16650 6020 16850
rect 6090 16650 6100 16850
rect 5900 16620 6100 16650
rect 6400 16850 6600 16880
rect 6400 16650 6410 16850
rect 6480 16650 6520 16850
rect 6590 16650 6600 16850
rect 6400 16620 6600 16650
rect 6900 16850 7100 16880
rect 6900 16650 6910 16850
rect 6980 16650 7020 16850
rect 7090 16650 7100 16850
rect 6900 16620 7100 16650
rect 7400 16850 7600 16880
rect 7400 16650 7410 16850
rect 7480 16650 7520 16850
rect 7590 16650 7600 16850
rect 7400 16620 7600 16650
rect 7900 16850 8100 16880
rect 7900 16650 7910 16850
rect 7980 16650 8020 16850
rect 8090 16650 8100 16850
rect 7900 16620 8100 16650
rect 8400 16850 8600 16880
rect 8400 16650 8410 16850
rect 8480 16650 8520 16850
rect 8590 16650 8600 16850
rect 8400 16620 8600 16650
rect 8900 16850 9100 16880
rect 8900 16650 8910 16850
rect 8980 16650 9020 16850
rect 9090 16650 9100 16850
rect 8900 16620 9100 16650
rect 9400 16850 9600 16880
rect 9400 16650 9410 16850
rect 9480 16650 9520 16850
rect 9590 16650 9600 16850
rect 9400 16620 9600 16650
rect 9900 16850 10100 16880
rect 9900 16650 9910 16850
rect 9980 16650 10020 16850
rect 10090 16650 10100 16850
rect 9900 16620 10100 16650
rect 10400 16850 10600 16880
rect 10400 16650 10410 16850
rect 10480 16650 10520 16850
rect 10590 16650 10600 16850
rect 10400 16620 10600 16650
rect 10900 16850 11100 16880
rect 10900 16650 10910 16850
rect 10980 16650 11020 16850
rect 11090 16650 11100 16850
rect 10900 16620 11100 16650
rect 11400 16850 11600 16880
rect 11400 16650 11410 16850
rect 11480 16650 11520 16850
rect 11590 16650 11600 16850
rect 11400 16620 11600 16650
rect 11900 16850 12100 16880
rect 11900 16650 11910 16850
rect 11980 16650 12020 16850
rect 12090 16650 12100 16850
rect 11900 16620 12100 16650
rect 12400 16850 12600 16880
rect 12400 16650 12410 16850
rect 12480 16650 12520 16850
rect 12590 16650 12600 16850
rect 12400 16620 12600 16650
rect 12900 16850 13100 16880
rect 12900 16650 12910 16850
rect 12980 16650 13020 16850
rect 13090 16650 13100 16850
rect 12900 16620 13100 16650
rect 13400 16850 13600 16880
rect 13400 16650 13410 16850
rect 13480 16650 13520 16850
rect 13590 16650 13600 16850
rect 13400 16620 13600 16650
rect 13900 16850 14100 16880
rect 13900 16650 13910 16850
rect 13980 16650 14020 16850
rect 14090 16650 14100 16850
rect 13900 16620 14100 16650
rect 14400 16850 14600 16880
rect 14400 16650 14410 16850
rect 14480 16650 14520 16850
rect 14590 16650 14600 16850
rect 14400 16620 14600 16650
rect 14900 16850 15100 16880
rect 14900 16650 14910 16850
rect 14980 16650 15020 16850
rect 15090 16650 15100 16850
rect 14900 16620 15100 16650
rect 15400 16850 15600 16880
rect 15400 16650 15410 16850
rect 15480 16650 15520 16850
rect 15590 16650 15600 16850
rect 15400 16620 15600 16650
rect 15900 16850 16100 16880
rect 15900 16650 15910 16850
rect 15980 16650 16020 16850
rect 16090 16650 16100 16850
rect 15900 16620 16100 16650
rect 16400 16850 16600 16880
rect 16400 16650 16410 16850
rect 16480 16650 16520 16850
rect 16590 16650 16600 16850
rect 16400 16620 16600 16650
rect 16900 16850 17100 16880
rect 16900 16650 16910 16850
rect 16980 16650 17020 16850
rect 17090 16650 17100 16850
rect 16900 16620 17100 16650
rect 17400 16850 17600 16880
rect 17400 16650 17410 16850
rect 17480 16650 17520 16850
rect 17590 16650 17600 16850
rect 17400 16620 17600 16650
rect 17900 16850 18100 16880
rect 17900 16650 17910 16850
rect 17980 16650 18020 16850
rect 18090 16650 18100 16850
rect 17900 16620 18100 16650
rect 18400 16850 18600 16880
rect 18400 16650 18410 16850
rect 18480 16650 18520 16850
rect 18590 16650 18600 16850
rect 18400 16620 18600 16650
rect 18900 16850 19100 16880
rect 18900 16650 18910 16850
rect 18980 16650 19020 16850
rect 19090 16650 19100 16850
rect 18900 16620 19100 16650
rect 19400 16850 19600 16880
rect 19400 16650 19410 16850
rect 19480 16650 19520 16850
rect 19590 16650 19600 16850
rect 19400 16620 19600 16650
rect 19900 16850 20100 16880
rect 19900 16650 19910 16850
rect 19980 16650 20020 16850
rect 20090 16650 20100 16850
rect 19900 16620 20100 16650
rect 20400 16850 20600 16880
rect 20400 16650 20410 16850
rect 20480 16650 20520 16850
rect 20590 16650 20600 16850
rect 20400 16620 20600 16650
rect 20900 16850 21100 16880
rect 20900 16650 20910 16850
rect 20980 16650 21020 16850
rect 21090 16650 21100 16850
rect 20900 16620 21100 16650
rect 21400 16850 21600 16880
rect 21400 16650 21410 16850
rect 21480 16650 21520 16850
rect 21590 16650 21600 16850
rect 21400 16620 21600 16650
rect 21900 16850 22100 16880
rect 21900 16650 21910 16850
rect 21980 16650 22020 16850
rect 22090 16650 22100 16850
rect 21900 16620 22100 16650
rect 22400 16850 22600 16880
rect 22400 16650 22410 16850
rect 22480 16650 22520 16850
rect 22590 16650 22600 16850
rect 22400 16620 22600 16650
rect 22900 16850 23100 16880
rect 22900 16650 22910 16850
rect 22980 16650 23020 16850
rect 23090 16650 23100 16850
rect 22900 16620 23100 16650
rect 23400 16850 23600 16880
rect 23400 16650 23410 16850
rect 23480 16650 23520 16850
rect 23590 16650 23600 16850
rect 23400 16620 23600 16650
rect 23900 16850 24100 16880
rect 23900 16650 23910 16850
rect 23980 16650 24020 16850
rect 24090 16650 24100 16850
rect 23900 16620 24100 16650
rect 24400 16850 24600 16880
rect 24400 16650 24410 16850
rect 24480 16650 24520 16850
rect 24590 16650 24600 16850
rect 24400 16620 24600 16650
rect 24900 16850 25100 16880
rect 24900 16650 24910 16850
rect 24980 16650 25020 16850
rect 25090 16650 25100 16850
rect 24900 16620 25100 16650
rect 25400 16850 25600 16880
rect 25400 16650 25410 16850
rect 25480 16650 25520 16850
rect 25590 16650 25600 16850
rect 25400 16620 25600 16650
rect 25900 16850 26100 16880
rect 25900 16650 25910 16850
rect 25980 16650 26020 16850
rect 26090 16650 26100 16850
rect 25900 16620 26100 16650
rect 26400 16850 26500 16880
rect 26400 16650 26410 16850
rect 26480 16650 26500 16850
rect 26400 16620 26500 16650
rect 0 16600 120 16620
rect 380 16600 620 16620
rect 880 16600 1120 16620
rect 1380 16600 1620 16620
rect 1880 16600 2120 16620
rect 2380 16600 2620 16620
rect 2880 16600 3120 16620
rect 3380 16600 3620 16620
rect 3880 16600 4120 16620
rect 4380 16600 4620 16620
rect 4880 16600 5120 16620
rect 5380 16600 5620 16620
rect 5880 16600 6120 16620
rect 6380 16600 6620 16620
rect 6880 16600 7120 16620
rect 7380 16600 7620 16620
rect 7880 16600 8120 16620
rect 8380 16600 8620 16620
rect 8880 16600 9120 16620
rect 9380 16600 9620 16620
rect 9880 16600 10120 16620
rect 10380 16600 10620 16620
rect 10880 16600 11120 16620
rect 11380 16600 11620 16620
rect 11880 16600 12120 16620
rect 12380 16600 12620 16620
rect 12880 16600 13120 16620
rect 13380 16600 13620 16620
rect 13880 16600 14120 16620
rect 14380 16600 14620 16620
rect 14880 16600 15120 16620
rect 15380 16600 15620 16620
rect 15880 16600 16120 16620
rect 16380 16600 16620 16620
rect 16880 16600 17120 16620
rect 17380 16600 17620 16620
rect 17880 16600 18120 16620
rect 18380 16600 18620 16620
rect 18880 16600 19120 16620
rect 19380 16600 19620 16620
rect 19880 16600 20120 16620
rect 20380 16600 20620 16620
rect 20880 16600 21120 16620
rect 21380 16600 21620 16620
rect 21880 16600 22120 16620
rect 22380 16600 22620 16620
rect 22880 16600 23120 16620
rect 23380 16600 23620 16620
rect 23880 16600 24120 16620
rect 24380 16600 24620 16620
rect 24880 16600 25120 16620
rect 25380 16600 25620 16620
rect 25880 16600 26120 16620
rect 26380 16600 26500 16620
rect 0 16590 26500 16600
rect 0 16520 150 16590
rect 350 16520 650 16590
rect 850 16520 1150 16590
rect 1350 16520 1650 16590
rect 1850 16520 2150 16590
rect 2350 16520 2650 16590
rect 2850 16520 3150 16590
rect 3350 16520 3650 16590
rect 3850 16520 4150 16590
rect 4350 16520 4650 16590
rect 4850 16520 5150 16590
rect 5350 16520 5650 16590
rect 5850 16520 6150 16590
rect 6350 16520 6650 16590
rect 6850 16520 7150 16590
rect 7350 16520 7650 16590
rect 7850 16520 8150 16590
rect 8350 16520 8650 16590
rect 8850 16520 9150 16590
rect 9350 16520 9650 16590
rect 9850 16520 10150 16590
rect 10350 16520 10650 16590
rect 10850 16520 11150 16590
rect 11350 16520 11650 16590
rect 11850 16520 12150 16590
rect 12350 16520 12650 16590
rect 12850 16520 13150 16590
rect 13350 16520 13650 16590
rect 13850 16520 14150 16590
rect 14350 16520 14650 16590
rect 14850 16520 15150 16590
rect 15350 16520 15650 16590
rect 15850 16520 16150 16590
rect 16350 16520 16650 16590
rect 16850 16520 17150 16590
rect 17350 16520 17650 16590
rect 17850 16520 18150 16590
rect 18350 16520 18650 16590
rect 18850 16520 19150 16590
rect 19350 16520 19650 16590
rect 19850 16520 20150 16590
rect 20350 16520 20650 16590
rect 20850 16520 21150 16590
rect 21350 16520 21650 16590
rect 21850 16520 22150 16590
rect 22350 16520 22650 16590
rect 22850 16520 23150 16590
rect 23350 16520 23650 16590
rect 23850 16520 24150 16590
rect 24350 16520 24650 16590
rect 24850 16520 25150 16590
rect 25350 16520 25650 16590
rect 25850 16520 26150 16590
rect 26350 16520 26500 16590
rect 0 16480 26500 16520
rect 0 16410 150 16480
rect 350 16410 650 16480
rect 850 16410 1150 16480
rect 1350 16410 1650 16480
rect 1850 16410 2150 16480
rect 2350 16410 2650 16480
rect 2850 16410 3150 16480
rect 3350 16410 3650 16480
rect 3850 16410 4150 16480
rect 4350 16410 4650 16480
rect 4850 16410 5150 16480
rect 5350 16410 5650 16480
rect 5850 16410 6150 16480
rect 6350 16410 6650 16480
rect 6850 16410 7150 16480
rect 7350 16410 7650 16480
rect 7850 16410 8150 16480
rect 8350 16410 8650 16480
rect 8850 16410 9150 16480
rect 9350 16410 9650 16480
rect 9850 16410 10150 16480
rect 10350 16410 10650 16480
rect 10850 16410 11150 16480
rect 11350 16410 11650 16480
rect 11850 16410 12150 16480
rect 12350 16410 12650 16480
rect 12850 16410 13150 16480
rect 13350 16410 13650 16480
rect 13850 16410 14150 16480
rect 14350 16410 14650 16480
rect 14850 16410 15150 16480
rect 15350 16410 15650 16480
rect 15850 16410 16150 16480
rect 16350 16410 16650 16480
rect 16850 16410 17150 16480
rect 17350 16410 17650 16480
rect 17850 16410 18150 16480
rect 18350 16410 18650 16480
rect 18850 16410 19150 16480
rect 19350 16410 19650 16480
rect 19850 16410 20150 16480
rect 20350 16410 20650 16480
rect 20850 16410 21150 16480
rect 21350 16410 21650 16480
rect 21850 16410 22150 16480
rect 22350 16410 22650 16480
rect 22850 16410 23150 16480
rect 23350 16410 23650 16480
rect 23850 16410 24150 16480
rect 24350 16410 24650 16480
rect 24850 16410 25150 16480
rect 25350 16410 25650 16480
rect 25850 16410 26150 16480
rect 26350 16410 26500 16480
rect 0 16400 26500 16410
rect 0 16380 120 16400
rect 380 16380 620 16400
rect 880 16380 1120 16400
rect 1380 16380 1620 16400
rect 1880 16380 2120 16400
rect 2380 16380 2620 16400
rect 2880 16380 3120 16400
rect 3380 16380 3620 16400
rect 3880 16380 4120 16400
rect 4380 16380 4620 16400
rect 4880 16380 5120 16400
rect 5380 16380 5620 16400
rect 5880 16380 6120 16400
rect 6380 16380 6620 16400
rect 6880 16380 7120 16400
rect 7380 16380 7620 16400
rect 7880 16380 8120 16400
rect 8380 16380 8620 16400
rect 8880 16380 9120 16400
rect 9380 16380 9620 16400
rect 9880 16380 10120 16400
rect 10380 16380 10620 16400
rect 10880 16380 11120 16400
rect 11380 16380 11620 16400
rect 11880 16380 12120 16400
rect 12380 16380 12620 16400
rect 12880 16380 13120 16400
rect 13380 16380 13620 16400
rect 13880 16380 14120 16400
rect 14380 16380 14620 16400
rect 14880 16380 15120 16400
rect 15380 16380 15620 16400
rect 15880 16380 16120 16400
rect 16380 16380 16620 16400
rect 16880 16380 17120 16400
rect 17380 16380 17620 16400
rect 17880 16380 18120 16400
rect 18380 16380 18620 16400
rect 18880 16380 19120 16400
rect 19380 16380 19620 16400
rect 19880 16380 20120 16400
rect 20380 16380 20620 16400
rect 20880 16380 21120 16400
rect 21380 16380 21620 16400
rect 21880 16380 22120 16400
rect 22380 16380 22620 16400
rect 22880 16380 23120 16400
rect 23380 16380 23620 16400
rect 23880 16380 24120 16400
rect 24380 16380 24620 16400
rect 24880 16380 25120 16400
rect 25380 16380 25620 16400
rect 25880 16380 26120 16400
rect 26380 16380 26500 16400
rect 0 16350 100 16380
rect 0 16150 20 16350
rect 90 16150 100 16350
rect 0 16120 100 16150
rect 400 16350 600 16380
rect 400 16150 410 16350
rect 480 16150 520 16350
rect 590 16150 600 16350
rect 400 16120 600 16150
rect 900 16350 1100 16380
rect 900 16150 910 16350
rect 980 16150 1020 16350
rect 1090 16150 1100 16350
rect 900 16120 1100 16150
rect 1400 16350 1600 16380
rect 1400 16150 1410 16350
rect 1480 16150 1520 16350
rect 1590 16150 1600 16350
rect 1400 16120 1600 16150
rect 1900 16350 2100 16380
rect 1900 16150 1910 16350
rect 1980 16150 2020 16350
rect 2090 16150 2100 16350
rect 1900 16120 2100 16150
rect 2400 16350 2600 16380
rect 2400 16150 2410 16350
rect 2480 16150 2520 16350
rect 2590 16150 2600 16350
rect 2400 16120 2600 16150
rect 2900 16350 3100 16380
rect 2900 16150 2910 16350
rect 2980 16150 3020 16350
rect 3090 16150 3100 16350
rect 2900 16120 3100 16150
rect 3400 16350 3600 16380
rect 3400 16150 3410 16350
rect 3480 16150 3520 16350
rect 3590 16150 3600 16350
rect 3400 16120 3600 16150
rect 3900 16350 4100 16380
rect 3900 16150 3910 16350
rect 3980 16150 4020 16350
rect 4090 16150 4100 16350
rect 3900 16120 4100 16150
rect 4400 16350 4600 16380
rect 4400 16150 4410 16350
rect 4480 16150 4520 16350
rect 4590 16150 4600 16350
rect 4400 16120 4600 16150
rect 4900 16350 5100 16380
rect 4900 16150 4910 16350
rect 4980 16150 5020 16350
rect 5090 16150 5100 16350
rect 4900 16120 5100 16150
rect 5400 16350 5600 16380
rect 5400 16150 5410 16350
rect 5480 16150 5520 16350
rect 5590 16150 5600 16350
rect 5400 16120 5600 16150
rect 5900 16350 6100 16380
rect 5900 16150 5910 16350
rect 5980 16150 6020 16350
rect 6090 16150 6100 16350
rect 5900 16120 6100 16150
rect 6400 16350 6600 16380
rect 6400 16150 6410 16350
rect 6480 16150 6520 16350
rect 6590 16150 6600 16350
rect 6400 16120 6600 16150
rect 6900 16350 7100 16380
rect 6900 16150 6910 16350
rect 6980 16150 7020 16350
rect 7090 16150 7100 16350
rect 6900 16120 7100 16150
rect 7400 16350 7600 16380
rect 7400 16150 7410 16350
rect 7480 16150 7520 16350
rect 7590 16150 7600 16350
rect 7400 16120 7600 16150
rect 7900 16350 8100 16380
rect 7900 16150 7910 16350
rect 7980 16150 8020 16350
rect 8090 16150 8100 16350
rect 7900 16120 8100 16150
rect 8400 16350 8600 16380
rect 8400 16150 8410 16350
rect 8480 16150 8520 16350
rect 8590 16150 8600 16350
rect 8400 16120 8600 16150
rect 8900 16350 9100 16380
rect 8900 16150 8910 16350
rect 8980 16150 9020 16350
rect 9090 16150 9100 16350
rect 8900 16120 9100 16150
rect 9400 16350 9600 16380
rect 9400 16150 9410 16350
rect 9480 16150 9520 16350
rect 9590 16150 9600 16350
rect 9400 16120 9600 16150
rect 9900 16350 10100 16380
rect 9900 16150 9910 16350
rect 9980 16150 10020 16350
rect 10090 16150 10100 16350
rect 9900 16120 10100 16150
rect 10400 16350 10600 16380
rect 10400 16150 10410 16350
rect 10480 16150 10520 16350
rect 10590 16150 10600 16350
rect 10400 16120 10600 16150
rect 10900 16350 11100 16380
rect 10900 16150 10910 16350
rect 10980 16150 11020 16350
rect 11090 16150 11100 16350
rect 10900 16120 11100 16150
rect 11400 16350 11600 16380
rect 11400 16150 11410 16350
rect 11480 16150 11520 16350
rect 11590 16150 11600 16350
rect 11400 16120 11600 16150
rect 11900 16350 12100 16380
rect 11900 16150 11910 16350
rect 11980 16150 12020 16350
rect 12090 16150 12100 16350
rect 11900 16120 12100 16150
rect 12400 16350 12600 16380
rect 12400 16150 12410 16350
rect 12480 16150 12520 16350
rect 12590 16150 12600 16350
rect 12400 16120 12600 16150
rect 12900 16350 13100 16380
rect 12900 16150 12910 16350
rect 12980 16150 13020 16350
rect 13090 16150 13100 16350
rect 12900 16120 13100 16150
rect 13400 16350 13600 16380
rect 13400 16150 13410 16350
rect 13480 16150 13520 16350
rect 13590 16150 13600 16350
rect 13400 16120 13600 16150
rect 13900 16350 14100 16380
rect 13900 16150 13910 16350
rect 13980 16150 14020 16350
rect 14090 16150 14100 16350
rect 13900 16120 14100 16150
rect 14400 16350 14600 16380
rect 14400 16150 14410 16350
rect 14480 16150 14520 16350
rect 14590 16150 14600 16350
rect 14400 16120 14600 16150
rect 14900 16350 15100 16380
rect 14900 16150 14910 16350
rect 14980 16150 15020 16350
rect 15090 16150 15100 16350
rect 14900 16120 15100 16150
rect 15400 16350 15600 16380
rect 15400 16150 15410 16350
rect 15480 16150 15520 16350
rect 15590 16150 15600 16350
rect 15400 16120 15600 16150
rect 15900 16350 16100 16380
rect 15900 16150 15910 16350
rect 15980 16150 16020 16350
rect 16090 16150 16100 16350
rect 15900 16120 16100 16150
rect 16400 16350 16600 16380
rect 16400 16150 16410 16350
rect 16480 16150 16520 16350
rect 16590 16150 16600 16350
rect 16400 16120 16600 16150
rect 16900 16350 17100 16380
rect 16900 16150 16910 16350
rect 16980 16150 17020 16350
rect 17090 16150 17100 16350
rect 16900 16120 17100 16150
rect 17400 16350 17600 16380
rect 17400 16150 17410 16350
rect 17480 16150 17520 16350
rect 17590 16150 17600 16350
rect 17400 16120 17600 16150
rect 17900 16350 18100 16380
rect 17900 16150 17910 16350
rect 17980 16150 18020 16350
rect 18090 16150 18100 16350
rect 17900 16120 18100 16150
rect 18400 16350 18600 16380
rect 18400 16150 18410 16350
rect 18480 16150 18520 16350
rect 18590 16150 18600 16350
rect 18400 16120 18600 16150
rect 18900 16350 19100 16380
rect 18900 16150 18910 16350
rect 18980 16150 19020 16350
rect 19090 16150 19100 16350
rect 18900 16120 19100 16150
rect 19400 16350 19600 16380
rect 19400 16150 19410 16350
rect 19480 16150 19520 16350
rect 19590 16150 19600 16350
rect 19400 16120 19600 16150
rect 19900 16350 20100 16380
rect 19900 16150 19910 16350
rect 19980 16150 20020 16350
rect 20090 16150 20100 16350
rect 19900 16120 20100 16150
rect 20400 16350 20600 16380
rect 20400 16150 20410 16350
rect 20480 16150 20520 16350
rect 20590 16150 20600 16350
rect 20400 16120 20600 16150
rect 20900 16350 21100 16380
rect 20900 16150 20910 16350
rect 20980 16150 21020 16350
rect 21090 16150 21100 16350
rect 20900 16120 21100 16150
rect 21400 16350 21600 16380
rect 21400 16150 21410 16350
rect 21480 16150 21520 16350
rect 21590 16150 21600 16350
rect 21400 16120 21600 16150
rect 21900 16350 22100 16380
rect 21900 16150 21910 16350
rect 21980 16150 22020 16350
rect 22090 16150 22100 16350
rect 21900 16120 22100 16150
rect 22400 16350 22600 16380
rect 22400 16150 22410 16350
rect 22480 16150 22520 16350
rect 22590 16150 22600 16350
rect 22400 16120 22600 16150
rect 22900 16350 23100 16380
rect 22900 16150 22910 16350
rect 22980 16150 23020 16350
rect 23090 16150 23100 16350
rect 22900 16120 23100 16150
rect 23400 16350 23600 16380
rect 23400 16150 23410 16350
rect 23480 16150 23520 16350
rect 23590 16150 23600 16350
rect 23400 16120 23600 16150
rect 23900 16350 24100 16380
rect 23900 16150 23910 16350
rect 23980 16150 24020 16350
rect 24090 16150 24100 16350
rect 23900 16120 24100 16150
rect 24400 16350 24600 16380
rect 24400 16150 24410 16350
rect 24480 16150 24520 16350
rect 24590 16150 24600 16350
rect 24400 16120 24600 16150
rect 24900 16350 25100 16380
rect 24900 16150 24910 16350
rect 24980 16150 25020 16350
rect 25090 16150 25100 16350
rect 24900 16120 25100 16150
rect 25400 16350 25600 16380
rect 25400 16150 25410 16350
rect 25480 16150 25520 16350
rect 25590 16150 25600 16350
rect 25400 16120 25600 16150
rect 25900 16350 26100 16380
rect 25900 16150 25910 16350
rect 25980 16150 26020 16350
rect 26090 16150 26100 16350
rect 25900 16120 26100 16150
rect 26400 16350 26500 16380
rect 26400 16150 26410 16350
rect 26480 16150 26500 16350
rect 26400 16120 26500 16150
rect 0 16100 120 16120
rect 380 16100 620 16120
rect 880 16100 1120 16120
rect 1380 16100 1620 16120
rect 1880 16100 2120 16120
rect 2380 16100 2620 16120
rect 2880 16100 3120 16120
rect 3380 16100 3620 16120
rect 3880 16100 4120 16120
rect 4380 16100 4620 16120
rect 4880 16100 5120 16120
rect 5380 16100 5620 16120
rect 5880 16100 6120 16120
rect 6380 16100 6620 16120
rect 6880 16100 7120 16120
rect 7380 16100 7620 16120
rect 7880 16100 8120 16120
rect 8380 16100 8620 16120
rect 8880 16100 9120 16120
rect 9380 16100 9620 16120
rect 9880 16100 10120 16120
rect 10380 16100 10620 16120
rect 10880 16100 11120 16120
rect 11380 16100 11620 16120
rect 11880 16100 12120 16120
rect 12380 16100 12620 16120
rect 12880 16100 13120 16120
rect 13380 16100 13620 16120
rect 13880 16100 14120 16120
rect 14380 16100 14620 16120
rect 14880 16100 15120 16120
rect 15380 16100 15620 16120
rect 15880 16100 16120 16120
rect 16380 16100 16620 16120
rect 16880 16100 17120 16120
rect 17380 16100 17620 16120
rect 17880 16100 18120 16120
rect 18380 16100 18620 16120
rect 18880 16100 19120 16120
rect 19380 16100 19620 16120
rect 19880 16100 20120 16120
rect 20380 16100 20620 16120
rect 20880 16100 21120 16120
rect 21380 16100 21620 16120
rect 21880 16100 22120 16120
rect 22380 16100 22620 16120
rect 22880 16100 23120 16120
rect 23380 16100 23620 16120
rect 23880 16100 24120 16120
rect 24380 16100 24620 16120
rect 24880 16100 25120 16120
rect 25380 16100 25620 16120
rect 25880 16100 26120 16120
rect 26380 16100 26500 16120
rect 0 16090 26500 16100
rect 0 16020 150 16090
rect 350 16020 650 16090
rect 850 16020 1150 16090
rect 1350 16020 1650 16090
rect 1850 16020 2150 16090
rect 2350 16020 2650 16090
rect 2850 16020 3150 16090
rect 3350 16020 3650 16090
rect 3850 16020 4150 16090
rect 4350 16020 4650 16090
rect 4850 16020 5150 16090
rect 5350 16020 5650 16090
rect 5850 16020 6150 16090
rect 6350 16020 6650 16090
rect 6850 16020 7150 16090
rect 7350 16020 7650 16090
rect 7850 16020 8150 16090
rect 8350 16020 8650 16090
rect 8850 16020 9150 16090
rect 9350 16020 9650 16090
rect 9850 16020 10150 16090
rect 10350 16020 10650 16090
rect 10850 16020 11150 16090
rect 11350 16020 11650 16090
rect 11850 16020 12150 16090
rect 12350 16020 12650 16090
rect 12850 16020 13150 16090
rect 13350 16020 13650 16090
rect 13850 16020 14150 16090
rect 14350 16020 14650 16090
rect 14850 16020 15150 16090
rect 15350 16020 15650 16090
rect 15850 16020 16150 16090
rect 16350 16020 16650 16090
rect 16850 16020 17150 16090
rect 17350 16020 17650 16090
rect 17850 16020 18150 16090
rect 18350 16020 18650 16090
rect 18850 16020 19150 16090
rect 19350 16020 19650 16090
rect 19850 16020 20150 16090
rect 20350 16020 20650 16090
rect 20850 16020 21150 16090
rect 21350 16020 21650 16090
rect 21850 16020 22150 16090
rect 22350 16020 22650 16090
rect 22850 16020 23150 16090
rect 23350 16020 23650 16090
rect 23850 16020 24150 16090
rect 24350 16020 24650 16090
rect 24850 16020 25150 16090
rect 25350 16020 25650 16090
rect 25850 16020 26150 16090
rect 26350 16020 26500 16090
rect 0 16000 26500 16020
rect 0 15980 1340 16000
rect 0 15910 150 15980
rect 350 15910 650 15980
rect 850 15910 1340 15980
rect 0 15900 1340 15910
rect 0 15880 120 15900
rect 380 15880 620 15900
rect 880 15880 1340 15900
rect 0 15850 100 15880
rect 0 15650 20 15850
rect 90 15650 100 15850
rect 0 15620 100 15650
rect 400 15850 600 15880
rect 400 15650 410 15850
rect 480 15650 520 15850
rect 590 15650 600 15850
rect 400 15620 600 15650
rect 900 15850 1340 15880
rect 900 15650 910 15850
rect 980 15650 1340 15850
rect 900 15620 1340 15650
rect 0 15600 120 15620
rect 380 15600 620 15620
rect 880 15600 1340 15620
rect 0 15590 1340 15600
rect 0 15520 150 15590
rect 350 15520 650 15590
rect 850 15580 1340 15590
rect 6500 15980 7500 16000
rect 6500 15910 6650 15980
rect 6850 15910 7150 15980
rect 7350 15910 7500 15980
rect 6500 15900 7500 15910
rect 6500 15880 6620 15900
rect 6880 15880 7120 15900
rect 7380 15880 7500 15900
rect 6500 15850 6600 15880
rect 6500 15650 6520 15850
rect 6590 15650 6600 15850
rect 6500 15620 6600 15650
rect 6900 15850 7100 15880
rect 6900 15650 6910 15850
rect 6980 15650 7020 15850
rect 7090 15650 7100 15850
rect 6900 15620 7100 15650
rect 7400 15850 7500 15880
rect 7400 15650 7410 15850
rect 7480 15650 7500 15850
rect 7400 15620 7500 15650
rect 6500 15600 6620 15620
rect 6880 15600 7120 15620
rect 7380 15600 7500 15620
rect 6500 15590 7500 15600
rect 850 15570 6410 15580
rect 850 15532 1536 15570
rect 6259 15532 6410 15570
rect 850 15522 6410 15532
rect 850 15520 1400 15522
rect 0 15480 1330 15520
rect 0 15410 150 15480
rect 350 15410 650 15480
rect 850 15410 1330 15480
rect 0 15400 1330 15410
rect 0 15380 120 15400
rect 380 15380 620 15400
rect 880 15380 1330 15400
rect 6340 15520 6410 15522
rect 1532 15430 1552 15490
rect 6186 15430 6206 15490
rect 1532 15396 1544 15430
rect 6194 15396 6206 15430
rect 1532 15390 1552 15396
rect 6186 15390 6206 15396
rect 0 15350 100 15380
rect 0 15150 20 15350
rect 90 15150 100 15350
rect 0 15120 100 15150
rect 400 15350 600 15380
rect 400 15150 410 15350
rect 480 15150 520 15350
rect 590 15150 600 15350
rect 400 15120 600 15150
rect 900 15350 1330 15380
rect 900 15150 910 15350
rect 980 15150 1330 15350
rect 900 15120 1330 15150
rect 0 15100 120 15120
rect 380 15100 620 15120
rect 880 15100 1330 15120
rect 0 15090 1330 15100
rect 0 15020 150 15090
rect 350 15020 650 15090
rect 850 15020 1330 15090
rect 0 14980 1330 15020
rect 0 14910 150 14980
rect 350 14910 650 14980
rect 850 14910 1330 14980
rect 0 14900 1330 14910
rect 0 14880 120 14900
rect 380 14880 620 14900
rect 880 14880 1330 14900
rect 0 14850 100 14880
rect 0 14650 20 14850
rect 90 14650 100 14850
rect 0 14620 100 14650
rect 400 14850 600 14880
rect 400 14650 410 14850
rect 480 14650 520 14850
rect 590 14650 600 14850
rect 400 14620 600 14650
rect 900 14850 1330 14880
rect 900 14650 910 14850
rect 980 14650 1330 14850
rect 900 14620 1330 14650
rect 0 14600 120 14620
rect 380 14600 620 14620
rect 880 14600 1330 14620
rect 0 14590 1330 14600
rect 0 14520 150 14590
rect 350 14520 650 14590
rect 850 14520 1330 14590
rect 0 14480 1330 14520
rect 0 14410 150 14480
rect 350 14410 650 14480
rect 850 14410 1330 14480
rect 0 14400 1330 14410
rect 0 14380 120 14400
rect 380 14380 620 14400
rect 880 14380 1330 14400
rect 0 14350 100 14380
rect 0 14150 20 14350
rect 90 14150 100 14350
rect 0 14120 100 14150
rect 400 14350 600 14380
rect 400 14150 410 14350
rect 480 14150 520 14350
rect 590 14150 600 14350
rect 400 14120 600 14150
rect 900 14350 1330 14380
rect 900 14150 910 14350
rect 980 14150 1330 14350
rect 900 14120 1330 14150
rect 0 14100 120 14120
rect 380 14100 620 14120
rect 880 14100 1330 14120
rect 0 14090 1330 14100
rect 0 14020 150 14090
rect 350 14020 650 14090
rect 850 14020 1330 14090
rect 0 14000 1330 14020
rect -4000 13980 1330 14000
rect -4000 13960 -3850 13980
rect -4060 13940 -3850 13960
rect -4300 13900 -4100 13910
rect -4300 13420 -4290 13900
rect -4110 13420 -4100 13900
rect -4300 13410 -4100 13420
rect -4300 13090 -4100 13100
rect -4300 12610 -4290 13090
rect -4110 12610 -4100 13090
rect -4300 12600 -4100 12610
rect -4060 12560 -4040 13940
rect -4000 13910 -3850 13940
rect -3650 13910 -3350 13980
rect -3150 13910 -2850 13980
rect -2650 13910 -2350 13980
rect -2150 13910 -1850 13980
rect -1650 13910 -1350 13980
rect -1150 13910 -850 13980
rect -650 13910 -350 13980
rect -150 13910 150 13980
rect 350 13910 650 13980
rect 850 13910 1330 13980
rect -4000 13900 1330 13910
rect -4000 13880 -3880 13900
rect -3620 13880 -3380 13900
rect -3120 13880 -2880 13900
rect -2620 13880 -2380 13900
rect -2120 13880 -1880 13900
rect -1620 13880 -1380 13900
rect -1120 13880 -880 13900
rect -620 13880 -380 13900
rect -120 13880 120 13900
rect 380 13880 620 13900
rect 880 13880 1330 13900
rect -4000 13850 -3900 13880
rect -4000 13650 -3980 13850
rect -3910 13650 -3900 13850
rect -4000 13620 -3900 13650
rect -3600 13850 -3400 13880
rect -3600 13650 -3590 13850
rect -3520 13650 -3480 13850
rect -3410 13650 -3400 13850
rect -3600 13620 -3400 13650
rect -3100 13850 -2900 13880
rect -3100 13650 -3090 13850
rect -3020 13650 -2980 13850
rect -2910 13650 -2900 13850
rect -3100 13620 -2900 13650
rect -2600 13850 -2400 13880
rect -2600 13650 -2590 13850
rect -2520 13650 -2480 13850
rect -2410 13650 -2400 13850
rect -2600 13620 -2400 13650
rect -2100 13850 -1900 13880
rect -2100 13650 -2090 13850
rect -2020 13650 -1980 13850
rect -1910 13650 -1900 13850
rect -2100 13620 -1900 13650
rect -1600 13850 -1400 13880
rect -1600 13650 -1590 13850
rect -1520 13650 -1480 13850
rect -1410 13650 -1400 13850
rect -1600 13620 -1400 13650
rect -1100 13850 -900 13880
rect -1100 13650 -1090 13850
rect -1020 13650 -980 13850
rect -910 13650 -900 13850
rect -1100 13620 -900 13650
rect -600 13850 -400 13880
rect -600 13650 -590 13850
rect -520 13650 -480 13850
rect -410 13650 -400 13850
rect -600 13620 -400 13650
rect -100 13850 100 13880
rect -100 13650 -90 13850
rect -20 13650 20 13850
rect 90 13650 100 13850
rect -100 13620 100 13650
rect 400 13850 600 13880
rect 400 13650 410 13850
rect 480 13650 520 13850
rect 590 13650 600 13850
rect 400 13620 600 13650
rect 900 13850 1330 13880
rect 900 13650 910 13850
rect 980 13650 1330 13850
rect 900 13620 1330 13650
rect -4000 13600 -3880 13620
rect -3620 13600 -3380 13620
rect -3120 13600 -2880 13620
rect -2620 13600 -2380 13620
rect -2120 13600 -1880 13620
rect -1620 13600 -1380 13620
rect -1120 13600 -880 13620
rect -620 13600 -380 13620
rect -120 13600 120 13620
rect 380 13600 620 13620
rect 880 13600 1330 13620
rect -4000 13590 1330 13600
rect -4000 13520 -3850 13590
rect -3650 13520 -3350 13590
rect -3150 13520 -2850 13590
rect -2650 13520 -2350 13590
rect -2150 13520 -1850 13590
rect -1650 13520 -1350 13590
rect -1150 13520 -850 13590
rect -650 13520 -350 13590
rect -150 13520 150 13590
rect 350 13520 650 13590
rect 850 13520 1330 13590
rect -4000 13480 1330 13520
rect -4000 13410 -3850 13480
rect -3650 13410 -3350 13480
rect -3150 13410 -2850 13480
rect -2650 13410 -2350 13480
rect -2150 13410 -1850 13480
rect -1650 13410 -1350 13480
rect -1150 13410 -850 13480
rect -650 13410 -350 13480
rect -150 13410 150 13480
rect 350 13410 650 13480
rect 850 13410 1330 13480
rect -4000 13400 1330 13410
rect -4000 13380 -3880 13400
rect -3620 13380 -3380 13400
rect -3120 13380 -2880 13400
rect -2620 13380 -2380 13400
rect -2120 13380 -1880 13400
rect -1620 13380 -1380 13400
rect -1120 13380 -880 13400
rect -620 13380 -380 13400
rect -120 13380 120 13400
rect 380 13380 620 13400
rect 880 13380 1330 13400
rect -4000 13350 -3900 13380
rect -4000 13150 -3980 13350
rect -3910 13150 -3900 13350
rect -4000 13120 -3900 13150
rect -3600 13350 -3400 13380
rect -3600 13150 -3590 13350
rect -3520 13150 -3480 13350
rect -3410 13150 -3400 13350
rect -3600 13120 -3400 13150
rect -3100 13350 -2900 13380
rect -3100 13150 -3090 13350
rect -3020 13150 -2980 13350
rect -2910 13150 -2900 13350
rect -3100 13120 -2900 13150
rect -2600 13350 -2400 13380
rect -2600 13150 -2590 13350
rect -2520 13150 -2480 13350
rect -2410 13150 -2400 13350
rect -2600 13120 -2400 13150
rect -2100 13350 -1900 13380
rect -2100 13150 -2090 13350
rect -2020 13150 -1980 13350
rect -1910 13150 -1900 13350
rect -2100 13120 -1900 13150
rect -1600 13350 -1400 13380
rect -1600 13150 -1590 13350
rect -1520 13150 -1480 13350
rect -1410 13150 -1400 13350
rect -1600 13120 -1400 13150
rect -1100 13350 -900 13380
rect -1100 13150 -1090 13350
rect -1020 13150 -980 13350
rect -910 13150 -900 13350
rect -1100 13120 -900 13150
rect -600 13350 -400 13380
rect -600 13150 -590 13350
rect -520 13150 -480 13350
rect -410 13150 -400 13350
rect -600 13120 -400 13150
rect -100 13350 100 13380
rect -100 13150 -90 13350
rect -20 13150 20 13350
rect 90 13150 100 13350
rect -100 13120 100 13150
rect 400 13350 600 13380
rect 400 13150 410 13350
rect 480 13150 520 13350
rect 590 13150 600 13350
rect 400 13120 600 13150
rect 900 13350 1330 13380
rect 900 13150 910 13350
rect 980 13150 1330 13350
rect 900 13120 1330 13150
rect -4000 13100 -3880 13120
rect -3620 13100 -3380 13120
rect -3120 13100 -2880 13120
rect -2620 13100 -2380 13120
rect -2120 13100 -1880 13120
rect -1620 13100 -1380 13120
rect -1120 13100 -880 13120
rect -620 13100 -380 13120
rect -120 13100 120 13120
rect 380 13100 620 13120
rect 880 13100 1330 13120
rect -4000 13090 1330 13100
rect -4000 13020 -3850 13090
rect -3650 13020 -3350 13090
rect -3150 13020 -2850 13090
rect -2650 13020 -2350 13090
rect -2150 13020 -1850 13090
rect -1650 13020 -1350 13090
rect -1150 13020 -850 13090
rect -650 13020 -350 13090
rect -150 13020 150 13090
rect 350 13020 650 13090
rect 850 13020 1330 13090
rect -4000 13000 1330 13020
rect -4000 12560 -3980 13000
rect -4060 12540 -3980 12560
rect 0 12980 1330 13000
rect 0 12910 150 12980
rect 350 12910 650 12980
rect 850 12910 1330 12980
rect 0 12900 1330 12910
rect 0 12880 120 12900
rect 380 12880 620 12900
rect 880 12880 1330 12900
rect 0 12850 100 12880
rect 0 12650 20 12850
rect 90 12650 100 12850
rect 0 12620 100 12650
rect 400 12850 600 12880
rect 400 12650 410 12850
rect 480 12650 520 12850
rect 590 12650 600 12850
rect 400 12620 600 12650
rect 900 12850 1330 12880
rect 900 12650 910 12850
rect 980 12650 1330 12850
rect 900 12620 1330 12650
rect 0 12600 120 12620
rect 380 12600 620 12620
rect 880 12600 1330 12620
rect 0 12590 1330 12600
rect 0 12520 150 12590
rect 350 12520 650 12590
rect 850 12520 1330 12590
rect 0 12480 1330 12520
rect 0 12410 150 12480
rect 350 12410 650 12480
rect 850 12410 1330 12480
rect 0 12400 1330 12410
rect 0 12380 120 12400
rect 380 12380 620 12400
rect 880 12380 1330 12400
rect 0 12350 100 12380
rect 0 12150 20 12350
rect 90 12150 100 12350
rect 0 12120 100 12150
rect 400 12350 600 12380
rect 400 12150 410 12350
rect 480 12150 520 12350
rect 590 12150 600 12350
rect 400 12120 600 12150
rect 900 12350 1330 12380
rect 900 12150 910 12350
rect 980 12150 1330 12350
rect 900 12120 1330 12150
rect 0 12100 120 12120
rect 380 12100 620 12120
rect 880 12100 1330 12120
rect 0 12090 1330 12100
rect 0 12020 150 12090
rect 350 12020 650 12090
rect 850 12020 1330 12090
rect 0 11980 1330 12020
rect 0 11910 150 11980
rect 350 11910 650 11980
rect 850 11910 1330 11980
rect 0 11900 1330 11910
rect 0 11880 120 11900
rect 380 11880 620 11900
rect 880 11880 1330 11900
rect 0 11850 100 11880
rect 0 11650 20 11850
rect 90 11650 100 11850
rect 0 11620 100 11650
rect 400 11850 600 11880
rect 400 11650 410 11850
rect 480 11650 520 11850
rect 590 11650 600 11850
rect 400 11620 600 11650
rect 900 11850 1330 11880
rect 900 11650 910 11850
rect 980 11650 1330 11850
rect 900 11620 1330 11650
rect 0 11600 120 11620
rect 380 11600 620 11620
rect 880 11600 1330 11620
rect 0 11590 1330 11600
rect 0 11520 150 11590
rect 350 11520 650 11590
rect 850 11520 1330 11590
rect 0 11480 1330 11520
rect 0 11410 150 11480
rect 350 11410 650 11480
rect 850 11410 1330 11480
rect 0 11400 1330 11410
rect 0 11380 120 11400
rect 380 11380 620 11400
rect 880 11380 1330 11400
rect 0 11350 100 11380
rect 0 11150 20 11350
rect 90 11150 100 11350
rect 0 11120 100 11150
rect 400 11350 600 11380
rect 400 11150 410 11350
rect 480 11150 520 11350
rect 590 11150 600 11350
rect 400 11120 600 11150
rect 900 11350 1330 11380
rect 900 11150 910 11350
rect 980 11150 1330 11350
rect 900 11120 1330 11150
rect 0 11100 120 11120
rect 380 11100 620 11120
rect 880 11100 1330 11120
rect 0 11090 1330 11100
rect 0 11020 150 11090
rect 350 11020 650 11090
rect 850 11020 1330 11090
rect 0 10980 1330 11020
rect 0 10910 150 10980
rect 350 10910 650 10980
rect 850 10910 1330 10980
rect 0 10900 1330 10910
rect 0 10880 120 10900
rect 380 10880 620 10900
rect 880 10880 1330 10900
rect 0 10850 100 10880
rect 0 10650 20 10850
rect 90 10650 100 10850
rect 0 10620 100 10650
rect 400 10850 600 10880
rect 400 10650 410 10850
rect 480 10650 520 10850
rect 590 10650 600 10850
rect 400 10620 600 10650
rect 900 10850 1330 10880
rect 900 10650 910 10850
rect 980 10650 1330 10850
rect 900 10620 1330 10650
rect 0 10600 120 10620
rect 380 10600 620 10620
rect 880 10600 1330 10620
rect 0 10590 1330 10600
rect 0 10520 150 10590
rect 350 10520 650 10590
rect 850 10520 1330 10590
rect 0 10480 1330 10520
rect 0 10410 150 10480
rect 350 10410 650 10480
rect 850 10410 1330 10480
rect 0 10400 1330 10410
rect 0 10380 120 10400
rect 380 10380 620 10400
rect 880 10380 1330 10400
rect 0 10350 100 10380
rect 0 10150 20 10350
rect 90 10150 100 10350
rect 0 10120 100 10150
rect 400 10350 600 10380
rect 400 10150 410 10350
rect 480 10150 520 10350
rect 590 10150 600 10350
rect 400 10120 600 10150
rect 900 10350 1330 10380
rect 900 10150 910 10350
rect 980 10150 1330 10350
rect 900 10120 1330 10150
rect 0 10100 120 10120
rect 380 10100 620 10120
rect 880 10100 1330 10120
rect 0 10090 1330 10100
rect 0 10020 150 10090
rect 350 10020 650 10090
rect 850 10020 1330 10090
rect 0 9980 1330 10020
rect 0 9910 150 9980
rect 350 9910 650 9980
rect 850 9910 1330 9980
rect 0 9900 1330 9910
rect 0 9880 120 9900
rect 380 9880 620 9900
rect 880 9880 1330 9900
rect 0 9850 100 9880
rect 0 9650 20 9850
rect 90 9650 100 9850
rect 0 9620 100 9650
rect 400 9850 600 9880
rect 400 9650 410 9850
rect 480 9650 520 9850
rect 590 9650 600 9850
rect 400 9620 600 9650
rect 900 9850 1330 9880
rect 900 9650 910 9850
rect 980 9650 1330 9850
rect 900 9620 1330 9650
rect 0 9600 120 9620
rect 380 9600 620 9620
rect 880 9600 1330 9620
rect 0 9590 1330 9600
rect 0 9520 150 9590
rect 350 9520 650 9590
rect 850 9520 1330 9590
rect 0 9480 1330 9520
rect 0 9410 150 9480
rect 350 9410 650 9480
rect 850 9410 1330 9480
rect 0 9400 1330 9410
rect 0 9380 120 9400
rect 380 9380 620 9400
rect 880 9380 1330 9400
rect 0 9350 100 9380
rect 0 9150 20 9350
rect 90 9150 100 9350
rect 0 9120 100 9150
rect 400 9350 600 9380
rect 400 9150 410 9350
rect 480 9150 520 9350
rect 590 9150 600 9350
rect 400 9120 600 9150
rect 900 9350 1330 9380
rect 900 9150 910 9350
rect 980 9200 1330 9350
rect 6500 15520 6650 15590
rect 6850 15520 7150 15590
rect 7350 15520 7500 15590
rect 13000 15980 14000 16000
rect 13000 15910 13150 15980
rect 13350 15910 13650 15980
rect 13850 15910 14000 15980
rect 13000 15900 14000 15910
rect 13000 15880 13120 15900
rect 13380 15880 13620 15900
rect 13880 15880 14000 15900
rect 13000 15850 13100 15880
rect 13000 15650 13020 15850
rect 13090 15650 13100 15850
rect 13000 15620 13100 15650
rect 13400 15850 13600 15880
rect 13400 15650 13410 15850
rect 13480 15650 13520 15850
rect 13590 15650 13600 15850
rect 13400 15620 13600 15650
rect 13900 15850 14000 15880
rect 13900 15650 13910 15850
rect 13980 15650 14000 15850
rect 13900 15620 14000 15650
rect 13000 15600 13120 15620
rect 13380 15600 13620 15620
rect 13880 15600 14000 15620
rect 13000 15590 14000 15600
rect 6500 15500 7500 15520
rect 7630 15570 12710 15580
rect 7630 15532 7836 15570
rect 12559 15532 12710 15570
rect 7630 15522 12710 15532
rect 7630 15520 7700 15522
rect 1465 15346 1531 15358
rect 1465 15338 1482 15346
rect 1516 15338 1531 15346
rect 1465 9370 1482 9378
rect 1516 9370 1531 9378
rect 1465 9358 1531 9370
rect 1623 15346 1689 15358
rect 1623 15338 1640 15346
rect 1674 15338 1689 15346
rect 1623 9370 1640 9378
rect 1674 9370 1689 9378
rect 1623 9358 1689 9370
rect 1781 15346 1847 15358
rect 1781 15338 1798 15346
rect 1832 15338 1847 15346
rect 1781 9370 1798 9378
rect 1832 9370 1847 9378
rect 1781 9358 1847 9370
rect 1939 15346 2005 15358
rect 1939 15338 1956 15346
rect 1990 15338 2005 15346
rect 1939 9370 1956 9378
rect 1990 9370 2005 9378
rect 1939 9358 2005 9370
rect 2097 15346 2163 15358
rect 2097 15338 2114 15346
rect 2148 15338 2163 15346
rect 2097 9370 2114 9378
rect 2148 9370 2163 9378
rect 2097 9358 2163 9370
rect 2255 15346 2321 15358
rect 2255 15338 2272 15346
rect 2306 15338 2321 15346
rect 2255 9370 2272 9378
rect 2306 9370 2321 9378
rect 2255 9358 2321 9370
rect 2413 15346 2479 15358
rect 2413 15338 2430 15346
rect 2464 15338 2479 15346
rect 2413 9370 2430 9378
rect 2464 9370 2479 9378
rect 2413 9358 2479 9370
rect 2571 15346 2637 15358
rect 2571 15338 2588 15346
rect 2622 15338 2637 15346
rect 2571 9370 2588 9378
rect 2622 9370 2637 9378
rect 2571 9358 2637 9370
rect 2729 15346 2795 15358
rect 2729 15338 2746 15346
rect 2780 15338 2795 15346
rect 2729 9370 2746 9378
rect 2780 9370 2795 9378
rect 2729 9358 2795 9370
rect 2887 15346 2953 15358
rect 2887 15338 2904 15346
rect 2938 15338 2953 15346
rect 2887 9370 2904 9378
rect 2938 9370 2953 9378
rect 2887 9358 2953 9370
rect 3045 15346 3111 15358
rect 3045 15338 3062 15346
rect 3096 15338 3111 15346
rect 3045 9370 3062 9378
rect 3096 9370 3111 9378
rect 3045 9358 3111 9370
rect 3203 15346 3269 15358
rect 3203 15338 3220 15346
rect 3254 15338 3269 15346
rect 3203 9370 3220 9378
rect 3254 9370 3269 9378
rect 3203 9358 3269 9370
rect 3361 15346 3427 15358
rect 3361 15338 3378 15346
rect 3412 15338 3427 15346
rect 3361 9370 3378 9378
rect 3412 9370 3427 9378
rect 3361 9358 3427 9370
rect 3519 15346 3585 15358
rect 3519 15338 3536 15346
rect 3570 15338 3585 15346
rect 3519 9370 3536 9378
rect 3570 9370 3585 9378
rect 3519 9358 3585 9370
rect 3677 15346 3743 15358
rect 3677 15338 3694 15346
rect 3728 15338 3743 15346
rect 3677 9370 3694 9378
rect 3728 9370 3743 9378
rect 3677 9358 3743 9370
rect 3835 15346 3901 15358
rect 3835 15338 3852 15346
rect 3886 15338 3901 15346
rect 3835 9370 3852 9378
rect 3886 9370 3901 9378
rect 3835 9358 3901 9370
rect 3993 15346 4059 15358
rect 3993 15338 4010 15346
rect 4044 15338 4059 15346
rect 3993 9370 4010 9378
rect 4044 9370 4059 9378
rect 3993 9358 4059 9370
rect 4151 15346 4217 15358
rect 4151 15338 4168 15346
rect 4202 15338 4217 15346
rect 4151 9370 4168 9378
rect 4202 9370 4217 9378
rect 4151 9358 4217 9370
rect 4309 15346 4375 15358
rect 4309 15338 4326 15346
rect 4360 15338 4375 15346
rect 4309 9370 4326 9378
rect 4360 9370 4375 9378
rect 4309 9358 4375 9370
rect 4467 15346 4533 15358
rect 4467 15338 4484 15346
rect 4518 15338 4533 15346
rect 4467 9370 4484 9378
rect 4518 9370 4533 9378
rect 4467 9358 4533 9370
rect 4625 15346 4691 15358
rect 4625 15338 4642 15346
rect 4676 15338 4691 15346
rect 4625 9370 4642 9378
rect 4676 9370 4691 9378
rect 4625 9358 4691 9370
rect 4783 15346 4849 15358
rect 4783 15338 4800 15346
rect 4834 15338 4849 15346
rect 4783 9370 4800 9378
rect 4834 9370 4849 9378
rect 4783 9358 4849 9370
rect 4941 15346 5007 15358
rect 4941 15338 4958 15346
rect 4992 15338 5007 15346
rect 4941 9370 4958 9378
rect 4992 9370 5007 9378
rect 4941 9358 5007 9370
rect 5099 15346 5165 15358
rect 5099 15338 5116 15346
rect 5150 15338 5165 15346
rect 5099 9370 5116 9378
rect 5150 9370 5165 9378
rect 5099 9358 5165 9370
rect 5257 15346 5323 15358
rect 5257 15338 5274 15346
rect 5308 15338 5323 15346
rect 5257 9370 5274 9378
rect 5308 9370 5323 9378
rect 5257 9358 5323 9370
rect 5415 15346 5481 15358
rect 5415 15338 5432 15346
rect 5466 15338 5481 15346
rect 5415 9370 5432 9378
rect 5466 9370 5481 9378
rect 5415 9358 5481 9370
rect 5573 15346 5639 15358
rect 5573 15338 5590 15346
rect 5624 15338 5639 15346
rect 5573 9370 5590 9378
rect 5624 9370 5639 9378
rect 5573 9358 5639 9370
rect 5731 15346 5797 15358
rect 5731 15338 5748 15346
rect 5782 15338 5797 15346
rect 5731 9370 5748 9378
rect 5782 9370 5797 9378
rect 5731 9358 5797 9370
rect 5889 15346 5955 15358
rect 5889 15338 5906 15346
rect 5940 15338 5955 15346
rect 5889 9370 5906 9378
rect 5940 9370 5955 9378
rect 5889 9358 5955 9370
rect 6047 15346 6113 15358
rect 6047 15338 6064 15346
rect 6098 15338 6113 15346
rect 6047 9370 6064 9378
rect 6098 9370 6113 9378
rect 6047 9358 6113 9370
rect 6205 15346 6271 15358
rect 6205 15338 6222 15346
rect 6256 15338 6271 15346
rect 6205 9370 6222 9378
rect 6256 9370 6271 9378
rect 6205 9358 6271 9370
rect 1532 9320 1552 9326
rect 6186 9320 6206 9326
rect 1532 9286 1544 9320
rect 6194 9286 6206 9320
rect 1532 9226 1552 9286
rect 6186 9226 6206 9286
rect 980 9194 1400 9200
rect 6340 9194 6410 9200
rect 980 9184 6410 9194
rect 980 9150 1536 9184
rect 900 9146 1536 9150
rect 6202 9146 6410 9184
rect 900 9130 6410 9146
rect 12640 15520 12710 15522
rect 7832 15430 7852 15490
rect 12486 15430 12506 15490
rect 7832 15396 7844 15430
rect 12494 15396 12506 15430
rect 7832 15390 7852 15396
rect 12486 15390 12506 15396
rect 13000 15520 13150 15590
rect 13350 15520 13650 15590
rect 13850 15580 14000 15590
rect 19000 15980 20000 16000
rect 19000 15910 19150 15980
rect 19350 15910 19650 15980
rect 19850 15910 20000 15980
rect 19000 15900 20000 15910
rect 19000 15880 19120 15900
rect 19380 15880 19620 15900
rect 19880 15880 20000 15900
rect 19000 15850 19100 15880
rect 19000 15650 19020 15850
rect 19090 15650 19100 15850
rect 19000 15620 19100 15650
rect 19400 15850 19600 15880
rect 19400 15650 19410 15850
rect 19480 15650 19520 15850
rect 19590 15650 19600 15850
rect 19400 15620 19600 15650
rect 19900 15850 20000 15880
rect 19900 15650 19910 15850
rect 19980 15650 20000 15850
rect 19900 15620 20000 15650
rect 19000 15600 19120 15620
rect 19380 15600 19620 15620
rect 19880 15600 20000 15620
rect 19000 15590 20000 15600
rect 19000 15580 19150 15590
rect 13850 15570 19150 15580
rect 13850 15532 14136 15570
rect 18859 15532 19150 15570
rect 13850 15522 19150 15532
rect 13850 15520 14000 15522
rect 13000 15500 13930 15520
rect 7765 15346 7831 15358
rect 7765 15338 7782 15346
rect 7816 15338 7831 15346
rect 7765 9370 7782 9378
rect 7816 9370 7831 9378
rect 7765 9358 7831 9370
rect 7923 15346 7989 15358
rect 7923 15338 7940 15346
rect 7974 15338 7989 15346
rect 7923 9370 7940 9378
rect 7974 9370 7989 9378
rect 7923 9358 7989 9370
rect 8081 15346 8147 15358
rect 8081 15338 8098 15346
rect 8132 15338 8147 15346
rect 8081 9370 8098 9378
rect 8132 9370 8147 9378
rect 8081 9358 8147 9370
rect 8239 15346 8305 15358
rect 8239 15338 8256 15346
rect 8290 15338 8305 15346
rect 8239 9370 8256 9378
rect 8290 9370 8305 9378
rect 8239 9358 8305 9370
rect 8397 15346 8463 15358
rect 8397 15338 8414 15346
rect 8448 15338 8463 15346
rect 8397 9370 8414 9378
rect 8448 9370 8463 9378
rect 8397 9358 8463 9370
rect 8555 15346 8621 15358
rect 8555 15338 8572 15346
rect 8606 15338 8621 15346
rect 8555 9370 8572 9378
rect 8606 9370 8621 9378
rect 8555 9358 8621 9370
rect 8713 15346 8779 15358
rect 8713 15338 8730 15346
rect 8764 15338 8779 15346
rect 8713 9370 8730 9378
rect 8764 9370 8779 9378
rect 8713 9358 8779 9370
rect 8871 15346 8937 15358
rect 8871 15338 8888 15346
rect 8922 15338 8937 15346
rect 8871 9370 8888 9378
rect 8922 9370 8937 9378
rect 8871 9358 8937 9370
rect 9029 15346 9095 15358
rect 9029 15338 9046 15346
rect 9080 15338 9095 15346
rect 9029 9370 9046 9378
rect 9080 9370 9095 9378
rect 9029 9358 9095 9370
rect 9187 15346 9253 15358
rect 9187 15338 9204 15346
rect 9238 15338 9253 15346
rect 9187 9370 9204 9378
rect 9238 9370 9253 9378
rect 9187 9358 9253 9370
rect 9345 15346 9411 15358
rect 9345 15338 9362 15346
rect 9396 15338 9411 15346
rect 9345 9370 9362 9378
rect 9396 9370 9411 9378
rect 9345 9358 9411 9370
rect 9503 15346 9569 15358
rect 9503 15338 9520 15346
rect 9554 15338 9569 15346
rect 9503 9370 9520 9378
rect 9554 9370 9569 9378
rect 9503 9358 9569 9370
rect 9661 15346 9727 15358
rect 9661 15338 9678 15346
rect 9712 15338 9727 15346
rect 9661 9370 9678 9378
rect 9712 9370 9727 9378
rect 9661 9358 9727 9370
rect 9819 15346 9885 15358
rect 9819 15338 9836 15346
rect 9870 15338 9885 15346
rect 9819 9370 9836 9378
rect 9870 9370 9885 9378
rect 9819 9358 9885 9370
rect 9977 15346 10043 15358
rect 9977 15338 9994 15346
rect 10028 15338 10043 15346
rect 9977 9370 9994 9378
rect 10028 9370 10043 9378
rect 9977 9358 10043 9370
rect 10135 15346 10201 15358
rect 10135 15338 10152 15346
rect 10186 15338 10201 15346
rect 10135 9370 10152 9378
rect 10186 9370 10201 9378
rect 10135 9358 10201 9370
rect 10293 15346 10359 15358
rect 10293 15338 10310 15346
rect 10344 15338 10359 15346
rect 10293 9370 10310 9378
rect 10344 9370 10359 9378
rect 10293 9358 10359 9370
rect 10451 15346 10517 15358
rect 10451 15338 10468 15346
rect 10502 15338 10517 15346
rect 10451 9370 10468 9378
rect 10502 9370 10517 9378
rect 10451 9358 10517 9370
rect 10609 15346 10675 15358
rect 10609 15338 10626 15346
rect 10660 15338 10675 15346
rect 10609 9370 10626 9378
rect 10660 9370 10675 9378
rect 10609 9358 10675 9370
rect 10767 15346 10833 15358
rect 10767 15338 10784 15346
rect 10818 15338 10833 15346
rect 10767 9370 10784 9378
rect 10818 9370 10833 9378
rect 10767 9358 10833 9370
rect 10925 15346 10991 15358
rect 10925 15338 10942 15346
rect 10976 15338 10991 15346
rect 10925 9370 10942 9378
rect 10976 9370 10991 9378
rect 10925 9358 10991 9370
rect 11083 15346 11149 15358
rect 11083 15338 11100 15346
rect 11134 15338 11149 15346
rect 11083 9370 11100 9378
rect 11134 9370 11149 9378
rect 11083 9358 11149 9370
rect 11241 15346 11307 15358
rect 11241 15338 11258 15346
rect 11292 15338 11307 15346
rect 11241 9370 11258 9378
rect 11292 9370 11307 9378
rect 11241 9358 11307 9370
rect 11399 15346 11465 15358
rect 11399 15338 11416 15346
rect 11450 15338 11465 15346
rect 11399 9370 11416 9378
rect 11450 9370 11465 9378
rect 11399 9358 11465 9370
rect 11557 15346 11623 15358
rect 11557 15338 11574 15346
rect 11608 15338 11623 15346
rect 11557 9370 11574 9378
rect 11608 9370 11623 9378
rect 11557 9358 11623 9370
rect 11715 15346 11781 15358
rect 11715 15338 11732 15346
rect 11766 15338 11781 15346
rect 11715 9370 11732 9378
rect 11766 9370 11781 9378
rect 11715 9358 11781 9370
rect 11873 15346 11939 15358
rect 11873 15338 11890 15346
rect 11924 15338 11939 15346
rect 11873 9370 11890 9378
rect 11924 9370 11939 9378
rect 11873 9358 11939 9370
rect 12031 15346 12097 15358
rect 12031 15338 12048 15346
rect 12082 15338 12097 15346
rect 12031 9370 12048 9378
rect 12082 9370 12097 9378
rect 12031 9358 12097 9370
rect 12189 15346 12255 15358
rect 12189 15338 12206 15346
rect 12240 15338 12255 15346
rect 12189 9370 12206 9378
rect 12240 9370 12255 9378
rect 12189 9358 12255 9370
rect 12347 15346 12413 15358
rect 12347 15338 12364 15346
rect 12398 15338 12413 15346
rect 12347 9370 12364 9378
rect 12398 9370 12413 9378
rect 12347 9358 12413 9370
rect 12505 15346 12571 15358
rect 12505 15338 12522 15346
rect 12556 15338 12571 15346
rect 12505 9370 12522 9378
rect 12556 9370 12571 9378
rect 12505 9358 12571 9370
rect 7832 9320 7852 9326
rect 12486 9320 12506 9326
rect 7832 9286 7844 9320
rect 12494 9286 12506 9320
rect 7832 9226 7852 9286
rect 12486 9226 12506 9286
rect 7630 9194 7700 9200
rect 12640 9194 12710 9200
rect 7630 9184 12710 9194
rect 7630 9146 7836 9184
rect 12502 9146 12710 9184
rect 7630 9130 12710 9146
rect 18940 15520 19150 15522
rect 19350 15520 19650 15590
rect 19850 15520 20000 15590
rect 25260 15980 26500 16000
rect 25260 15910 25650 15980
rect 25850 15910 26150 15980
rect 26350 15910 26500 15980
rect 25260 15900 26500 15910
rect 25260 15880 25620 15900
rect 25880 15880 26120 15900
rect 26380 15880 26500 15900
rect 25260 15850 25600 15880
rect 25260 15650 25520 15850
rect 25590 15650 25600 15850
rect 25260 15620 25600 15650
rect 25900 15850 26100 15880
rect 25900 15650 25910 15850
rect 25980 15650 26020 15850
rect 26090 15650 26100 15850
rect 25900 15620 26100 15650
rect 26400 15850 26500 15880
rect 26400 15650 26410 15850
rect 26480 15650 26500 15850
rect 26400 15620 26500 15650
rect 25260 15600 25620 15620
rect 25880 15600 26120 15620
rect 26380 15600 26500 15620
rect 25260 15590 26500 15600
rect 25260 15580 25650 15590
rect 14132 15430 14152 15490
rect 18786 15430 18806 15490
rect 14132 15396 14144 15430
rect 18794 15396 18806 15430
rect 14132 15390 14152 15396
rect 18786 15390 18806 15396
rect 19010 15500 20000 15520
rect 20230 15570 25650 15580
rect 20230 15532 20436 15570
rect 25159 15532 25650 15570
rect 20230 15522 25650 15532
rect 20230 15520 20300 15522
rect 14065 15346 14131 15358
rect 14065 15338 14082 15346
rect 14116 15338 14131 15346
rect 14065 9370 14082 9378
rect 14116 9370 14131 9378
rect 14065 9358 14131 9370
rect 14223 15346 14289 15358
rect 14223 15338 14240 15346
rect 14274 15338 14289 15346
rect 14223 9370 14240 9378
rect 14274 9370 14289 9378
rect 14223 9358 14289 9370
rect 14381 15346 14447 15358
rect 14381 15338 14398 15346
rect 14432 15338 14447 15346
rect 14381 9370 14398 9378
rect 14432 9370 14447 9378
rect 14381 9358 14447 9370
rect 14539 15346 14605 15358
rect 14539 15338 14556 15346
rect 14590 15338 14605 15346
rect 14539 9370 14556 9378
rect 14590 9370 14605 9378
rect 14539 9358 14605 9370
rect 14697 15346 14763 15358
rect 14697 15338 14714 15346
rect 14748 15338 14763 15346
rect 14697 9370 14714 9378
rect 14748 9370 14763 9378
rect 14697 9358 14763 9370
rect 14855 15346 14921 15358
rect 14855 15338 14872 15346
rect 14906 15338 14921 15346
rect 14855 9370 14872 9378
rect 14906 9370 14921 9378
rect 14855 9358 14921 9370
rect 15013 15346 15079 15358
rect 15013 15338 15030 15346
rect 15064 15338 15079 15346
rect 15013 9370 15030 9378
rect 15064 9370 15079 9378
rect 15013 9358 15079 9370
rect 15171 15346 15237 15358
rect 15171 15338 15188 15346
rect 15222 15338 15237 15346
rect 15171 9370 15188 9378
rect 15222 9370 15237 9378
rect 15171 9358 15237 9370
rect 15329 15346 15395 15358
rect 15329 15338 15346 15346
rect 15380 15338 15395 15346
rect 15329 9370 15346 9378
rect 15380 9370 15395 9378
rect 15329 9358 15395 9370
rect 15487 15346 15553 15358
rect 15487 15338 15504 15346
rect 15538 15338 15553 15346
rect 15487 9370 15504 9378
rect 15538 9370 15553 9378
rect 15487 9358 15553 9370
rect 15645 15346 15711 15358
rect 15645 15338 15662 15346
rect 15696 15338 15711 15346
rect 15645 9370 15662 9378
rect 15696 9370 15711 9378
rect 15645 9358 15711 9370
rect 15803 15346 15869 15358
rect 15803 15338 15820 15346
rect 15854 15338 15869 15346
rect 15803 9370 15820 9378
rect 15854 9370 15869 9378
rect 15803 9358 15869 9370
rect 15961 15346 16027 15358
rect 15961 15338 15978 15346
rect 16012 15338 16027 15346
rect 15961 9370 15978 9378
rect 16012 9370 16027 9378
rect 15961 9358 16027 9370
rect 16119 15346 16185 15358
rect 16119 15338 16136 15346
rect 16170 15338 16185 15346
rect 16119 9370 16136 9378
rect 16170 9370 16185 9378
rect 16119 9358 16185 9370
rect 16277 15346 16343 15358
rect 16277 15338 16294 15346
rect 16328 15338 16343 15346
rect 16277 9370 16294 9378
rect 16328 9370 16343 9378
rect 16277 9358 16343 9370
rect 16435 15346 16501 15358
rect 16435 15338 16452 15346
rect 16486 15338 16501 15346
rect 16435 9370 16452 9378
rect 16486 9370 16501 9378
rect 16435 9358 16501 9370
rect 16593 15346 16659 15358
rect 16593 15338 16610 15346
rect 16644 15338 16659 15346
rect 16593 9370 16610 9378
rect 16644 9370 16659 9378
rect 16593 9358 16659 9370
rect 16751 15346 16817 15358
rect 16751 15338 16768 15346
rect 16802 15338 16817 15346
rect 16751 9370 16768 9378
rect 16802 9370 16817 9378
rect 16751 9358 16817 9370
rect 16909 15346 16975 15358
rect 16909 15338 16926 15346
rect 16960 15338 16975 15346
rect 16909 9370 16926 9378
rect 16960 9370 16975 9378
rect 16909 9358 16975 9370
rect 17067 15346 17133 15358
rect 17067 15338 17084 15346
rect 17118 15338 17133 15346
rect 17067 9370 17084 9378
rect 17118 9370 17133 9378
rect 17067 9358 17133 9370
rect 17225 15346 17291 15358
rect 17225 15338 17242 15346
rect 17276 15338 17291 15346
rect 17225 9370 17242 9378
rect 17276 9370 17291 9378
rect 17225 9358 17291 9370
rect 17383 15346 17449 15358
rect 17383 15338 17400 15346
rect 17434 15338 17449 15346
rect 17383 9370 17400 9378
rect 17434 9370 17449 9378
rect 17383 9358 17449 9370
rect 17541 15346 17607 15358
rect 17541 15338 17558 15346
rect 17592 15338 17607 15346
rect 17541 9370 17558 9378
rect 17592 9370 17607 9378
rect 17541 9358 17607 9370
rect 17699 15346 17765 15358
rect 17699 15338 17716 15346
rect 17750 15338 17765 15346
rect 17699 9370 17716 9378
rect 17750 9370 17765 9378
rect 17699 9358 17765 9370
rect 17857 15346 17923 15358
rect 17857 15338 17874 15346
rect 17908 15338 17923 15346
rect 17857 9370 17874 9378
rect 17908 9370 17923 9378
rect 17857 9358 17923 9370
rect 18015 15346 18081 15358
rect 18015 15338 18032 15346
rect 18066 15338 18081 15346
rect 18015 9370 18032 9378
rect 18066 9370 18081 9378
rect 18015 9358 18081 9370
rect 18173 15346 18239 15358
rect 18173 15338 18190 15346
rect 18224 15338 18239 15346
rect 18173 9370 18190 9378
rect 18224 9370 18239 9378
rect 18173 9358 18239 9370
rect 18331 15346 18397 15358
rect 18331 15338 18348 15346
rect 18382 15338 18397 15346
rect 18331 9370 18348 9378
rect 18382 9370 18397 9378
rect 18331 9358 18397 9370
rect 18489 15346 18555 15358
rect 18489 15338 18506 15346
rect 18540 15338 18555 15346
rect 18489 9370 18506 9378
rect 18540 9370 18555 9378
rect 18489 9358 18555 9370
rect 18647 15346 18713 15358
rect 18647 15338 18664 15346
rect 18698 15338 18713 15346
rect 18647 9370 18664 9378
rect 18698 9370 18713 9378
rect 18647 9358 18713 9370
rect 18805 15346 18871 15358
rect 18805 15338 18822 15346
rect 18856 15338 18871 15346
rect 18805 9370 18822 9378
rect 18856 9370 18871 9378
rect 18805 9358 18871 9370
rect 14132 9320 14152 9326
rect 18786 9320 18806 9326
rect 14132 9286 14144 9320
rect 18794 9286 18806 9320
rect 14132 9226 14152 9286
rect 18786 9226 18806 9286
rect 13930 9194 14000 9200
rect 18940 9194 19010 9200
rect 13930 9184 19010 9194
rect 13930 9146 14136 9184
rect 18802 9146 19010 9184
rect 13930 9130 19010 9146
rect 25240 15520 25650 15522
rect 25850 15520 26150 15590
rect 26350 15520 26500 15590
rect 20432 15430 20452 15490
rect 25086 15430 25106 15490
rect 20432 15396 20444 15430
rect 25094 15396 25106 15430
rect 20432 15390 20452 15396
rect 25086 15390 25106 15396
rect 25310 15480 26500 15520
rect 25310 15410 25650 15480
rect 25850 15410 26150 15480
rect 26350 15410 26500 15480
rect 25310 15400 26500 15410
rect 25310 15380 25620 15400
rect 25880 15380 26120 15400
rect 26380 15380 26500 15400
rect 20365 15346 20431 15358
rect 20365 15338 20382 15346
rect 20416 15338 20431 15346
rect 20365 9370 20382 9378
rect 20416 9370 20431 9378
rect 20365 9358 20431 9370
rect 20523 15346 20589 15358
rect 20523 15338 20540 15346
rect 20574 15338 20589 15346
rect 20523 9370 20540 9378
rect 20574 9370 20589 9378
rect 20523 9358 20589 9370
rect 20681 15346 20747 15358
rect 20681 15338 20698 15346
rect 20732 15338 20747 15346
rect 20681 9370 20698 9378
rect 20732 9370 20747 9378
rect 20681 9358 20747 9370
rect 20839 15346 20905 15358
rect 20839 15338 20856 15346
rect 20890 15338 20905 15346
rect 20839 9370 20856 9378
rect 20890 9370 20905 9378
rect 20839 9358 20905 9370
rect 20997 15346 21063 15358
rect 20997 15338 21014 15346
rect 21048 15338 21063 15346
rect 20997 9370 21014 9378
rect 21048 9370 21063 9378
rect 20997 9358 21063 9370
rect 21155 15346 21221 15358
rect 21155 15338 21172 15346
rect 21206 15338 21221 15346
rect 21155 9370 21172 9378
rect 21206 9370 21221 9378
rect 21155 9358 21221 9370
rect 21313 15346 21379 15358
rect 21313 15338 21330 15346
rect 21364 15338 21379 15346
rect 21313 9370 21330 9378
rect 21364 9370 21379 9378
rect 21313 9358 21379 9370
rect 21471 15346 21537 15358
rect 21471 15338 21488 15346
rect 21522 15338 21537 15346
rect 21471 9370 21488 9378
rect 21522 9370 21537 9378
rect 21471 9358 21537 9370
rect 21629 15346 21695 15358
rect 21629 15338 21646 15346
rect 21680 15338 21695 15346
rect 21629 9370 21646 9378
rect 21680 9370 21695 9378
rect 21629 9358 21695 9370
rect 21787 15346 21853 15358
rect 21787 15338 21804 15346
rect 21838 15338 21853 15346
rect 21787 9370 21804 9378
rect 21838 9370 21853 9378
rect 21787 9358 21853 9370
rect 21945 15346 22011 15358
rect 21945 15338 21962 15346
rect 21996 15338 22011 15346
rect 21945 9370 21962 9378
rect 21996 9370 22011 9378
rect 21945 9358 22011 9370
rect 22103 15346 22169 15358
rect 22103 15338 22120 15346
rect 22154 15338 22169 15346
rect 22103 9370 22120 9378
rect 22154 9370 22169 9378
rect 22103 9358 22169 9370
rect 22261 15346 22327 15358
rect 22261 15338 22278 15346
rect 22312 15338 22327 15346
rect 22261 9370 22278 9378
rect 22312 9370 22327 9378
rect 22261 9358 22327 9370
rect 22419 15346 22485 15358
rect 22419 15338 22436 15346
rect 22470 15338 22485 15346
rect 22419 9370 22436 9378
rect 22470 9370 22485 9378
rect 22419 9358 22485 9370
rect 22577 15346 22643 15358
rect 22577 15338 22594 15346
rect 22628 15338 22643 15346
rect 22577 9370 22594 9378
rect 22628 9370 22643 9378
rect 22577 9358 22643 9370
rect 22735 15346 22801 15358
rect 22735 15338 22752 15346
rect 22786 15338 22801 15346
rect 22735 9370 22752 9378
rect 22786 9370 22801 9378
rect 22735 9358 22801 9370
rect 22893 15346 22959 15358
rect 22893 15338 22910 15346
rect 22944 15338 22959 15346
rect 22893 9370 22910 9378
rect 22944 9370 22959 9378
rect 22893 9358 22959 9370
rect 23051 15346 23117 15358
rect 23051 15338 23068 15346
rect 23102 15338 23117 15346
rect 23051 9370 23068 9378
rect 23102 9370 23117 9378
rect 23051 9358 23117 9370
rect 23209 15346 23275 15358
rect 23209 15338 23226 15346
rect 23260 15338 23275 15346
rect 23209 9370 23226 9378
rect 23260 9370 23275 9378
rect 23209 9358 23275 9370
rect 23367 15346 23433 15358
rect 23367 15338 23384 15346
rect 23418 15338 23433 15346
rect 23367 9370 23384 9378
rect 23418 9370 23433 9378
rect 23367 9358 23433 9370
rect 23525 15346 23591 15358
rect 23525 15338 23542 15346
rect 23576 15338 23591 15346
rect 23525 9370 23542 9378
rect 23576 9370 23591 9378
rect 23525 9358 23591 9370
rect 23683 15346 23749 15358
rect 23683 15338 23700 15346
rect 23734 15338 23749 15346
rect 23683 9370 23700 9378
rect 23734 9370 23749 9378
rect 23683 9358 23749 9370
rect 23841 15346 23907 15358
rect 23841 15338 23858 15346
rect 23892 15338 23907 15346
rect 23841 9370 23858 9378
rect 23892 9370 23907 9378
rect 23841 9358 23907 9370
rect 23999 15346 24065 15358
rect 23999 15338 24016 15346
rect 24050 15338 24065 15346
rect 23999 9370 24016 9378
rect 24050 9370 24065 9378
rect 23999 9358 24065 9370
rect 24157 15346 24223 15358
rect 24157 15338 24174 15346
rect 24208 15338 24223 15346
rect 24157 9370 24174 9378
rect 24208 9370 24223 9378
rect 24157 9358 24223 9370
rect 24315 15346 24381 15358
rect 24315 15338 24332 15346
rect 24366 15338 24381 15346
rect 24315 9370 24332 9378
rect 24366 9370 24381 9378
rect 24315 9358 24381 9370
rect 24473 15346 24539 15358
rect 24473 15338 24490 15346
rect 24524 15338 24539 15346
rect 24473 9370 24490 9378
rect 24524 9370 24539 9378
rect 24473 9358 24539 9370
rect 24631 15346 24697 15358
rect 24631 15338 24648 15346
rect 24682 15338 24697 15346
rect 24631 9370 24648 9378
rect 24682 9370 24697 9378
rect 24631 9358 24697 9370
rect 24789 15346 24855 15358
rect 24789 15338 24806 15346
rect 24840 15338 24855 15346
rect 24789 9370 24806 9378
rect 24840 9370 24855 9378
rect 24789 9358 24855 9370
rect 24947 15346 25013 15358
rect 24947 15338 24964 15346
rect 24998 15338 25013 15346
rect 24947 9370 24964 9378
rect 24998 9370 25013 9378
rect 24947 9358 25013 9370
rect 25105 15346 25171 15358
rect 25105 15338 25122 15346
rect 25156 15338 25171 15346
rect 25105 9370 25122 9378
rect 25156 9370 25171 9378
rect 25105 9358 25171 9370
rect 25310 15350 25600 15380
rect 25310 15150 25520 15350
rect 25590 15150 25600 15350
rect 25310 15120 25600 15150
rect 25900 15350 26100 15380
rect 25900 15150 25910 15350
rect 25980 15150 26020 15350
rect 26090 15150 26100 15350
rect 25900 15120 26100 15150
rect 26400 15350 26500 15380
rect 26400 15150 26410 15350
rect 26480 15150 26500 15350
rect 26400 15120 26500 15150
rect 25310 15100 25620 15120
rect 25880 15100 26120 15120
rect 26380 15100 26500 15120
rect 25310 15090 26500 15100
rect 25310 15020 25650 15090
rect 25850 15020 26150 15090
rect 26350 15020 26500 15090
rect 25310 14980 26500 15020
rect 25310 14910 25650 14980
rect 25850 14910 26150 14980
rect 26350 14910 26500 14980
rect 25310 14900 26500 14910
rect 25310 14880 25620 14900
rect 25880 14880 26120 14900
rect 26380 14880 26500 14900
rect 25310 14850 25600 14880
rect 25310 14650 25520 14850
rect 25590 14650 25600 14850
rect 25310 14620 25600 14650
rect 25900 14850 26100 14880
rect 25900 14650 25910 14850
rect 25980 14650 26020 14850
rect 26090 14650 26100 14850
rect 25900 14620 26100 14650
rect 26400 14850 26500 14880
rect 26400 14650 26410 14850
rect 26480 14650 26500 14850
rect 26400 14620 26500 14650
rect 25310 14600 25620 14620
rect 25880 14600 26120 14620
rect 26380 14600 26500 14620
rect 25310 14590 26500 14600
rect 25310 14520 25650 14590
rect 25850 14520 26150 14590
rect 26350 14520 26500 14590
rect 25310 14480 26500 14520
rect 25310 14410 25650 14480
rect 25850 14410 26150 14480
rect 26350 14410 26500 14480
rect 25310 14400 26500 14410
rect 25310 14380 25620 14400
rect 25880 14380 26120 14400
rect 26380 14380 26500 14400
rect 25310 14350 25600 14380
rect 25310 14150 25520 14350
rect 25590 14150 25600 14350
rect 25310 14120 25600 14150
rect 25900 14350 26100 14380
rect 25900 14150 25910 14350
rect 25980 14150 26020 14350
rect 26090 14150 26100 14350
rect 25900 14120 26100 14150
rect 26400 14350 26500 14380
rect 26400 14150 26410 14350
rect 26480 14150 26500 14350
rect 26400 14120 26500 14150
rect 25310 14100 25620 14120
rect 25880 14100 26120 14120
rect 26380 14100 26500 14120
rect 25310 14090 26500 14100
rect 25310 14020 25650 14090
rect 25850 14020 26150 14090
rect 26350 14020 26500 14090
rect 25310 14000 26500 14020
rect 25310 13980 30860 14000
rect 25310 13910 25650 13980
rect 25850 13910 26150 13980
rect 26350 13910 26650 13980
rect 26850 13910 27150 13980
rect 27350 13910 27650 13980
rect 27850 13910 28150 13980
rect 28350 13910 28650 13980
rect 28850 13910 29150 13980
rect 29350 13910 29650 13980
rect 29850 13910 30150 13980
rect 30350 13910 30800 13980
rect 25310 13900 30800 13910
rect 25310 13880 25620 13900
rect 25880 13880 26120 13900
rect 26380 13880 26620 13900
rect 26880 13880 27120 13900
rect 27380 13880 27620 13900
rect 27880 13880 28120 13900
rect 28380 13880 28620 13900
rect 28880 13880 29120 13900
rect 29380 13880 29620 13900
rect 29880 13880 30120 13900
rect 30380 13880 30800 13900
rect 25310 13850 25600 13880
rect 25310 13650 25520 13850
rect 25590 13650 25600 13850
rect 25310 13620 25600 13650
rect 25900 13850 26100 13880
rect 25900 13650 25910 13850
rect 25980 13650 26020 13850
rect 26090 13650 26100 13850
rect 25900 13620 26100 13650
rect 26400 13850 26600 13880
rect 26400 13650 26410 13850
rect 26480 13650 26520 13850
rect 26590 13650 26600 13850
rect 26400 13620 26600 13650
rect 26900 13850 27100 13880
rect 26900 13650 26910 13850
rect 26980 13650 27020 13850
rect 27090 13650 27100 13850
rect 26900 13620 27100 13650
rect 27400 13850 27600 13880
rect 27400 13650 27410 13850
rect 27480 13650 27520 13850
rect 27590 13650 27600 13850
rect 27400 13620 27600 13650
rect 27900 13850 28100 13880
rect 27900 13650 27910 13850
rect 27980 13650 28020 13850
rect 28090 13650 28100 13850
rect 27900 13620 28100 13650
rect 28400 13850 28600 13880
rect 28400 13650 28410 13850
rect 28480 13650 28520 13850
rect 28590 13650 28600 13850
rect 28400 13620 28600 13650
rect 28900 13850 29100 13880
rect 28900 13650 28910 13850
rect 28980 13650 29020 13850
rect 29090 13650 29100 13850
rect 28900 13620 29100 13650
rect 29400 13850 29600 13880
rect 29400 13650 29410 13850
rect 29480 13650 29520 13850
rect 29590 13650 29600 13850
rect 29400 13620 29600 13650
rect 29900 13850 30100 13880
rect 29900 13650 29910 13850
rect 29980 13650 30020 13850
rect 30090 13650 30100 13850
rect 29900 13620 30100 13650
rect 30400 13850 30800 13880
rect 30400 13650 30410 13850
rect 30480 13650 30800 13850
rect 30400 13620 30800 13650
rect 25310 13600 25620 13620
rect 25880 13600 26120 13620
rect 26380 13600 26620 13620
rect 26880 13600 27120 13620
rect 27380 13600 27620 13620
rect 27880 13600 28120 13620
rect 28380 13600 28620 13620
rect 28880 13600 29120 13620
rect 29380 13600 29620 13620
rect 29880 13600 30120 13620
rect 30380 13600 30800 13620
rect 25310 13590 30800 13600
rect 25310 13520 25650 13590
rect 25850 13520 26150 13590
rect 26350 13520 26650 13590
rect 26850 13520 27150 13590
rect 27350 13520 27650 13590
rect 27850 13520 28150 13590
rect 28350 13520 28650 13590
rect 28850 13520 29150 13590
rect 29350 13520 29650 13590
rect 29850 13520 30150 13590
rect 30350 13520 30800 13590
rect 25310 13480 30800 13520
rect 25310 13410 25650 13480
rect 25850 13410 26150 13480
rect 26350 13410 26650 13480
rect 26850 13410 27150 13480
rect 27350 13410 27650 13480
rect 27850 13410 28150 13480
rect 28350 13410 28650 13480
rect 28850 13410 29150 13480
rect 29350 13410 29650 13480
rect 29850 13410 30150 13480
rect 30350 13410 30800 13480
rect 25310 13400 30800 13410
rect 25310 13380 25620 13400
rect 25880 13380 26120 13400
rect 26380 13380 26620 13400
rect 26880 13380 27120 13400
rect 27380 13380 27620 13400
rect 27880 13380 28120 13400
rect 28380 13380 28620 13400
rect 28880 13380 29120 13400
rect 29380 13380 29620 13400
rect 29880 13380 30120 13400
rect 30380 13380 30800 13400
rect 25310 13350 25600 13380
rect 25310 13150 25520 13350
rect 25590 13150 25600 13350
rect 25310 13120 25600 13150
rect 25900 13350 26100 13380
rect 25900 13150 25910 13350
rect 25980 13150 26020 13350
rect 26090 13150 26100 13350
rect 25900 13120 26100 13150
rect 26400 13350 26600 13380
rect 26400 13150 26410 13350
rect 26480 13150 26520 13350
rect 26590 13150 26600 13350
rect 26400 13120 26600 13150
rect 26900 13350 27100 13380
rect 26900 13150 26910 13350
rect 26980 13150 27020 13350
rect 27090 13150 27100 13350
rect 26900 13120 27100 13150
rect 27400 13350 27600 13380
rect 27400 13150 27410 13350
rect 27480 13150 27520 13350
rect 27590 13150 27600 13350
rect 27400 13120 27600 13150
rect 27900 13350 28100 13380
rect 27900 13150 27910 13350
rect 27980 13150 28020 13350
rect 28090 13150 28100 13350
rect 27900 13120 28100 13150
rect 28400 13350 28600 13380
rect 28400 13150 28410 13350
rect 28480 13150 28520 13350
rect 28590 13150 28600 13350
rect 28400 13120 28600 13150
rect 28900 13350 29100 13380
rect 28900 13150 28910 13350
rect 28980 13150 29020 13350
rect 29090 13150 29100 13350
rect 28900 13120 29100 13150
rect 29400 13350 29600 13380
rect 29400 13150 29410 13350
rect 29480 13150 29520 13350
rect 29590 13150 29600 13350
rect 29400 13120 29600 13150
rect 29900 13350 30100 13380
rect 29900 13150 29910 13350
rect 29980 13150 30020 13350
rect 30090 13150 30100 13350
rect 29900 13120 30100 13150
rect 30400 13350 30800 13380
rect 30400 13150 30410 13350
rect 30480 13150 30800 13350
rect 30400 13120 30800 13150
rect 25310 13100 25620 13120
rect 25880 13100 26120 13120
rect 26380 13100 26620 13120
rect 26880 13100 27120 13120
rect 27380 13100 27620 13120
rect 27880 13100 28120 13120
rect 28380 13100 28620 13120
rect 28880 13100 29120 13120
rect 29380 13100 29620 13120
rect 29880 13100 30120 13120
rect 30380 13100 30800 13120
rect 25310 13090 30800 13100
rect 25310 13020 25650 13090
rect 25850 13020 26150 13090
rect 26350 13020 26650 13090
rect 26850 13020 27150 13090
rect 27350 13020 27650 13090
rect 27850 13020 28150 13090
rect 28350 13020 28650 13090
rect 28850 13020 29150 13090
rect 29350 13020 29650 13090
rect 29850 13020 30150 13090
rect 30350 13020 30800 13090
rect 25310 13000 30800 13020
rect 25310 12980 26500 13000
rect 25310 12910 25650 12980
rect 25850 12910 26150 12980
rect 26350 12910 26500 12980
rect 25310 12900 26500 12910
rect 25310 12880 25620 12900
rect 25880 12880 26120 12900
rect 26380 12880 26500 12900
rect 25310 12850 25600 12880
rect 25310 12650 25520 12850
rect 25590 12650 25600 12850
rect 25310 12620 25600 12650
rect 25900 12850 26100 12880
rect 25900 12650 25910 12850
rect 25980 12650 26020 12850
rect 26090 12650 26100 12850
rect 25900 12620 26100 12650
rect 26400 12850 26500 12880
rect 26400 12650 26410 12850
rect 26480 12650 26500 12850
rect 26400 12620 26500 12650
rect 25310 12600 25620 12620
rect 25880 12600 26120 12620
rect 26380 12600 26500 12620
rect 25310 12590 26500 12600
rect 25310 12520 25650 12590
rect 25850 12520 26150 12590
rect 26350 12520 26500 12590
rect 25310 12480 26500 12520
rect 30780 12520 30800 13000
rect 30840 12520 30860 13980
rect 30900 13900 31100 13910
rect 30900 13420 30910 13900
rect 31090 13420 31100 13900
rect 30900 13410 31100 13420
rect 30900 13090 31100 13100
rect 30900 12610 30910 13090
rect 31090 12610 31100 13090
rect 30900 12600 31100 12610
rect 30780 12500 30860 12520
rect 25310 12410 25650 12480
rect 25850 12410 26150 12480
rect 26350 12410 26500 12480
rect 25310 12400 26500 12410
rect 25310 12380 25620 12400
rect 25880 12380 26120 12400
rect 26380 12380 26500 12400
rect 25310 12350 25600 12380
rect 25310 12150 25520 12350
rect 25590 12150 25600 12350
rect 25310 12120 25600 12150
rect 25900 12350 26100 12380
rect 25900 12150 25910 12350
rect 25980 12150 26020 12350
rect 26090 12150 26100 12350
rect 25900 12120 26100 12150
rect 26400 12350 26500 12380
rect 26400 12150 26410 12350
rect 26480 12150 26500 12350
rect 26400 12120 26500 12150
rect 25310 12100 25620 12120
rect 25880 12100 26120 12120
rect 26380 12100 26500 12120
rect 25310 12090 26500 12100
rect 25310 12020 25650 12090
rect 25850 12020 26150 12090
rect 26350 12020 26500 12090
rect 25310 11980 26500 12020
rect 25310 11910 25650 11980
rect 25850 11910 26150 11980
rect 26350 11910 26500 11980
rect 25310 11900 26500 11910
rect 25310 11880 25620 11900
rect 25880 11880 26120 11900
rect 26380 11880 26500 11900
rect 25310 11850 25600 11880
rect 25310 11650 25520 11850
rect 25590 11650 25600 11850
rect 25310 11620 25600 11650
rect 25900 11850 26100 11880
rect 25900 11650 25910 11850
rect 25980 11650 26020 11850
rect 26090 11650 26100 11850
rect 25900 11620 26100 11650
rect 26400 11850 26500 11880
rect 26400 11650 26410 11850
rect 26480 11650 26500 11850
rect 26400 11620 26500 11650
rect 25310 11600 25620 11620
rect 25880 11600 26120 11620
rect 26380 11600 26500 11620
rect 25310 11590 26500 11600
rect 25310 11520 25650 11590
rect 25850 11520 26150 11590
rect 26350 11520 26500 11590
rect 25310 11480 26500 11520
rect 25310 11410 25650 11480
rect 25850 11410 26150 11480
rect 26350 11410 26500 11480
rect 25310 11400 26500 11410
rect 25310 11380 25620 11400
rect 25880 11380 26120 11400
rect 26380 11380 26500 11400
rect 25310 11350 25600 11380
rect 25310 11150 25520 11350
rect 25590 11150 25600 11350
rect 25310 11120 25600 11150
rect 25900 11350 26100 11380
rect 25900 11150 25910 11350
rect 25980 11150 26020 11350
rect 26090 11150 26100 11350
rect 25900 11120 26100 11150
rect 26400 11350 26500 11380
rect 26400 11150 26410 11350
rect 26480 11150 26500 11350
rect 26400 11120 26500 11150
rect 25310 11100 25620 11120
rect 25880 11100 26120 11120
rect 26380 11100 26500 11120
rect 25310 11090 26500 11100
rect 25310 11020 25650 11090
rect 25850 11020 26150 11090
rect 26350 11020 26500 11090
rect 25310 10980 26500 11020
rect 25310 10910 25650 10980
rect 25850 10910 26150 10980
rect 26350 10910 26500 10980
rect 25310 10900 26500 10910
rect 25310 10880 25620 10900
rect 25880 10880 26120 10900
rect 26380 10880 26500 10900
rect 25310 10850 25600 10880
rect 25310 10650 25520 10850
rect 25590 10650 25600 10850
rect 25310 10620 25600 10650
rect 25900 10850 26100 10880
rect 25900 10650 25910 10850
rect 25980 10650 26020 10850
rect 26090 10650 26100 10850
rect 25900 10620 26100 10650
rect 26400 10850 26500 10880
rect 26400 10650 26410 10850
rect 26480 10650 26500 10850
rect 26400 10620 26500 10650
rect 25310 10600 25620 10620
rect 25880 10600 26120 10620
rect 26380 10600 26500 10620
rect 25310 10590 26500 10600
rect 25310 10520 25650 10590
rect 25850 10520 26150 10590
rect 26350 10520 26500 10590
rect 25310 10480 26500 10520
rect 25310 10410 25650 10480
rect 25850 10410 26150 10480
rect 26350 10410 26500 10480
rect 25310 10400 26500 10410
rect 25310 10380 25620 10400
rect 25880 10380 26120 10400
rect 26380 10380 26500 10400
rect 25310 10350 25600 10380
rect 25310 10150 25520 10350
rect 25590 10150 25600 10350
rect 25310 10120 25600 10150
rect 25900 10350 26100 10380
rect 25900 10150 25910 10350
rect 25980 10150 26020 10350
rect 26090 10150 26100 10350
rect 25900 10120 26100 10150
rect 26400 10350 26500 10380
rect 26400 10150 26410 10350
rect 26480 10150 26500 10350
rect 26400 10120 26500 10150
rect 25310 10100 25620 10120
rect 25880 10100 26120 10120
rect 26380 10100 26500 10120
rect 25310 10090 26500 10100
rect 25310 10020 25650 10090
rect 25850 10020 26150 10090
rect 26350 10020 26500 10090
rect 25310 9980 26500 10020
rect 25310 9910 25650 9980
rect 25850 9910 26150 9980
rect 26350 9910 26500 9980
rect 25310 9900 26500 9910
rect 25310 9880 25620 9900
rect 25880 9880 26120 9900
rect 26380 9880 26500 9900
rect 25310 9850 25600 9880
rect 25310 9650 25520 9850
rect 25590 9650 25600 9850
rect 25310 9620 25600 9650
rect 25900 9850 26100 9880
rect 25900 9650 25910 9850
rect 25980 9650 26020 9850
rect 26090 9650 26100 9850
rect 25900 9620 26100 9650
rect 26400 9850 26500 9880
rect 26400 9650 26410 9850
rect 26480 9650 26500 9850
rect 26400 9620 26500 9650
rect 25310 9600 25620 9620
rect 25880 9600 26120 9620
rect 26380 9600 26500 9620
rect 25310 9590 26500 9600
rect 25310 9520 25650 9590
rect 25850 9520 26150 9590
rect 26350 9520 26500 9590
rect 25310 9480 26500 9520
rect 25310 9410 25650 9480
rect 25850 9410 26150 9480
rect 26350 9410 26500 9480
rect 25310 9400 26500 9410
rect 25310 9380 25620 9400
rect 25880 9380 26120 9400
rect 26380 9380 26500 9400
rect 25310 9350 25600 9380
rect 20432 9320 20452 9326
rect 25086 9320 25106 9326
rect 20432 9286 20444 9320
rect 25094 9286 25106 9320
rect 20432 9226 20452 9286
rect 25086 9226 25106 9286
rect 20230 9194 20300 9200
rect 25310 9200 25520 9350
rect 25240 9194 25520 9200
rect 20230 9184 25520 9194
rect 20230 9146 20436 9184
rect 25102 9150 25520 9184
rect 25590 9150 25600 9350
rect 25102 9146 25600 9150
rect 20230 9130 25600 9146
rect 900 9120 1340 9130
rect 0 9100 120 9120
rect 380 9100 620 9120
rect 880 9100 1340 9120
rect 0 9090 1340 9100
rect 0 9020 150 9090
rect 350 9020 650 9090
rect 850 9020 1340 9090
rect 0 8980 1340 9020
rect 0 8910 150 8980
rect 350 8910 650 8980
rect 850 8910 1340 8980
rect 0 8900 1340 8910
rect 0 8880 120 8900
rect 380 8880 620 8900
rect 880 8880 1340 8900
rect 0 8850 100 8880
rect 0 8650 20 8850
rect 90 8650 100 8850
rect 0 8620 100 8650
rect 400 8850 600 8880
rect 400 8650 410 8850
rect 480 8650 520 8850
rect 590 8650 600 8850
rect 400 8620 600 8650
rect 900 8850 1340 8880
rect 900 8650 910 8850
rect 980 8650 1340 8850
rect 900 8620 1340 8650
rect 0 8600 120 8620
rect 380 8600 620 8620
rect 880 8600 1340 8620
rect 0 8590 1340 8600
rect 0 8520 150 8590
rect 350 8520 650 8590
rect 850 8580 1340 8590
rect 25260 9120 25600 9130
rect 25900 9350 26100 9380
rect 25900 9150 25910 9350
rect 25980 9150 26020 9350
rect 26090 9150 26100 9350
rect 25900 9120 26100 9150
rect 26400 9350 26500 9380
rect 26400 9150 26410 9350
rect 26480 9150 26500 9350
rect 26400 9120 26500 9150
rect 25260 9100 25620 9120
rect 25880 9100 26120 9120
rect 26380 9100 26500 9120
rect 25260 9090 26500 9100
rect 25260 9020 25650 9090
rect 25850 9020 26150 9090
rect 26350 9020 26500 9090
rect 25260 8980 26500 9020
rect 25260 8910 25650 8980
rect 25850 8910 26150 8980
rect 26350 8910 26500 8980
rect 25260 8900 26500 8910
rect 25260 8880 25620 8900
rect 25880 8880 26120 8900
rect 26380 8880 26500 8900
rect 25260 8850 25600 8880
rect 25260 8650 25520 8850
rect 25590 8650 25600 8850
rect 25260 8620 25600 8650
rect 25900 8850 26100 8880
rect 25900 8650 25910 8850
rect 25980 8650 26020 8850
rect 26090 8650 26100 8850
rect 25900 8620 26100 8650
rect 26400 8850 26500 8880
rect 26400 8650 26410 8850
rect 26480 8650 26500 8850
rect 26400 8620 26500 8650
rect 25260 8600 25620 8620
rect 25880 8600 26120 8620
rect 26380 8600 26500 8620
rect 25260 8590 26500 8600
rect 25260 8580 25650 8590
rect 850 8570 6410 8580
rect 850 8532 1536 8570
rect 6259 8532 6410 8570
rect 850 8522 6410 8532
rect 850 8520 1400 8522
rect 0 8480 1330 8520
rect 0 8410 150 8480
rect 350 8410 650 8480
rect 850 8410 1330 8480
rect 0 8400 1330 8410
rect 0 8380 120 8400
rect 380 8380 620 8400
rect 880 8380 1330 8400
rect 6340 8520 6410 8522
rect 1532 8430 1552 8490
rect 6186 8430 6206 8490
rect 1532 8396 1544 8430
rect 6194 8396 6206 8430
rect 1532 8390 1552 8396
rect 6186 8390 6206 8396
rect 0 8350 100 8380
rect 0 8150 20 8350
rect 90 8150 100 8350
rect 0 8120 100 8150
rect 400 8350 600 8380
rect 400 8150 410 8350
rect 480 8150 520 8350
rect 590 8150 600 8350
rect 400 8120 600 8150
rect 900 8350 1330 8380
rect 900 8150 910 8350
rect 980 8150 1330 8350
rect 900 8120 1330 8150
rect 0 8100 120 8120
rect 380 8100 620 8120
rect 880 8100 1330 8120
rect 0 8090 1330 8100
rect 0 8020 150 8090
rect 350 8020 650 8090
rect 850 8020 1330 8090
rect 0 7980 1330 8020
rect 0 7910 150 7980
rect 350 7910 650 7980
rect 850 7910 1330 7980
rect 0 7900 1330 7910
rect 0 7880 120 7900
rect 380 7880 620 7900
rect 880 7880 1330 7900
rect 0 7850 100 7880
rect 0 7650 20 7850
rect 90 7650 100 7850
rect 0 7620 100 7650
rect 400 7850 600 7880
rect 400 7650 410 7850
rect 480 7650 520 7850
rect 590 7650 600 7850
rect 400 7620 600 7650
rect 900 7850 1330 7880
rect 900 7650 910 7850
rect 980 7650 1330 7850
rect 900 7620 1330 7650
rect 0 7600 120 7620
rect 380 7600 620 7620
rect 880 7600 1330 7620
rect 0 7590 1330 7600
rect 0 7520 150 7590
rect 350 7520 650 7590
rect 850 7520 1330 7590
rect 0 7480 1330 7520
rect 0 7410 150 7480
rect 350 7410 650 7480
rect 850 7410 1330 7480
rect 0 7400 1330 7410
rect 0 7380 120 7400
rect 380 7380 620 7400
rect 880 7380 1330 7400
rect 0 7350 100 7380
rect 0 7150 20 7350
rect 90 7150 100 7350
rect 0 7120 100 7150
rect 400 7350 600 7380
rect 400 7150 410 7350
rect 480 7150 520 7350
rect 590 7150 600 7350
rect 400 7120 600 7150
rect 900 7350 1330 7380
rect 900 7150 910 7350
rect 980 7150 1330 7350
rect 900 7120 1330 7150
rect 0 7100 120 7120
rect 380 7100 620 7120
rect 880 7100 1330 7120
rect 0 7090 1330 7100
rect 0 7020 150 7090
rect 350 7020 650 7090
rect 850 7020 1330 7090
rect 0 6980 1330 7020
rect 0 6910 150 6980
rect 350 6910 650 6980
rect 850 6910 1330 6980
rect 0 6900 1330 6910
rect 0 6880 120 6900
rect 380 6880 620 6900
rect 880 6880 1330 6900
rect 0 6850 100 6880
rect 0 6650 20 6850
rect 90 6650 100 6850
rect 0 6620 100 6650
rect 400 6850 600 6880
rect 400 6650 410 6850
rect 480 6650 520 6850
rect 590 6650 600 6850
rect 400 6620 600 6650
rect 900 6850 1330 6880
rect 900 6650 910 6850
rect 980 6650 1330 6850
rect 900 6620 1330 6650
rect 0 6600 120 6620
rect 380 6600 620 6620
rect 880 6600 1330 6620
rect 0 6590 1330 6600
rect 0 6520 150 6590
rect 350 6520 650 6590
rect 850 6520 1330 6590
rect 0 6480 1330 6520
rect 0 6410 150 6480
rect 350 6410 650 6480
rect 850 6410 1330 6480
rect 0 6400 1330 6410
rect 0 6380 120 6400
rect 380 6380 620 6400
rect 880 6380 1330 6400
rect 0 6350 100 6380
rect 0 6150 20 6350
rect 90 6150 100 6350
rect 0 6120 100 6150
rect 400 6350 600 6380
rect 400 6150 410 6350
rect 480 6150 520 6350
rect 590 6150 600 6350
rect 400 6120 600 6150
rect 900 6350 1330 6380
rect 900 6150 910 6350
rect 980 6150 1330 6350
rect 900 6120 1330 6150
rect 0 6100 120 6120
rect 380 6100 620 6120
rect 880 6100 1330 6120
rect 0 6090 1330 6100
rect 0 6020 150 6090
rect 350 6020 650 6090
rect 850 6020 1330 6090
rect 0 5980 1330 6020
rect 0 5910 150 5980
rect 350 5910 650 5980
rect 850 5910 1330 5980
rect 0 5900 1330 5910
rect 0 5880 120 5900
rect 380 5880 620 5900
rect 880 5880 1330 5900
rect 0 5850 100 5880
rect 0 5650 20 5850
rect 90 5650 100 5850
rect 0 5620 100 5650
rect 400 5850 600 5880
rect 400 5650 410 5850
rect 480 5650 520 5850
rect 590 5650 600 5850
rect 400 5620 600 5650
rect 900 5850 1330 5880
rect 900 5650 910 5850
rect 980 5650 1330 5850
rect 900 5620 1330 5650
rect 0 5600 120 5620
rect 380 5600 620 5620
rect 880 5600 1330 5620
rect 0 5590 1330 5600
rect 0 5520 150 5590
rect 350 5520 650 5590
rect 850 5520 1330 5590
rect 0 5480 1330 5520
rect 0 5410 150 5480
rect 350 5410 650 5480
rect 850 5410 1330 5480
rect 0 5400 1330 5410
rect 0 5380 120 5400
rect 380 5380 620 5400
rect 880 5380 1330 5400
rect 0 5350 100 5380
rect 0 5150 20 5350
rect 90 5150 100 5350
rect 0 5120 100 5150
rect 400 5350 600 5380
rect 400 5150 410 5350
rect 480 5150 520 5350
rect 590 5150 600 5350
rect 400 5120 600 5150
rect 900 5350 1330 5380
rect 900 5150 910 5350
rect 980 5150 1330 5350
rect 900 5120 1330 5150
rect 0 5100 120 5120
rect 380 5100 620 5120
rect 880 5100 1330 5120
rect 0 5090 1330 5100
rect 0 5020 150 5090
rect 350 5020 650 5090
rect 850 5020 1330 5090
rect 0 4980 1330 5020
rect 0 4910 150 4980
rect 350 4910 650 4980
rect 850 4910 1330 4980
rect 0 4900 1330 4910
rect 0 4880 120 4900
rect 380 4880 620 4900
rect 880 4880 1330 4900
rect 0 4850 100 4880
rect 0 4650 20 4850
rect 90 4650 100 4850
rect 0 4620 100 4650
rect 400 4850 600 4880
rect 400 4650 410 4850
rect 480 4650 520 4850
rect 590 4650 600 4850
rect 400 4620 600 4650
rect 900 4850 1330 4880
rect 900 4650 910 4850
rect 980 4650 1330 4850
rect 900 4620 1330 4650
rect 0 4600 120 4620
rect 380 4600 620 4620
rect 880 4600 1330 4620
rect 0 4590 1330 4600
rect 0 4520 150 4590
rect 350 4520 650 4590
rect 850 4520 1330 4590
rect 0 4480 1330 4520
rect 0 4410 150 4480
rect 350 4410 650 4480
rect 850 4410 1330 4480
rect 0 4400 1330 4410
rect 0 4380 120 4400
rect 380 4380 620 4400
rect 880 4380 1330 4400
rect 0 4350 100 4380
rect 0 4150 20 4350
rect 90 4150 100 4350
rect 0 4120 100 4150
rect 400 4350 600 4380
rect 400 4150 410 4350
rect 480 4150 520 4350
rect 590 4150 600 4350
rect 400 4120 600 4150
rect 900 4350 1330 4380
rect 900 4150 910 4350
rect 980 4150 1330 4350
rect 900 4120 1330 4150
rect 0 4100 120 4120
rect 380 4100 620 4120
rect 880 4100 1330 4120
rect 0 4090 1330 4100
rect 0 4020 150 4090
rect 350 4020 650 4090
rect 850 4020 1330 4090
rect 0 3980 1330 4020
rect 0 3910 150 3980
rect 350 3910 650 3980
rect 850 3910 1330 3980
rect 0 3900 1330 3910
rect 0 3880 120 3900
rect 380 3880 620 3900
rect 880 3880 1330 3900
rect 0 3850 100 3880
rect 0 3650 20 3850
rect 90 3650 100 3850
rect 0 3620 100 3650
rect 400 3850 600 3880
rect 400 3650 410 3850
rect 480 3650 520 3850
rect 590 3650 600 3850
rect 400 3620 600 3650
rect 900 3850 1330 3880
rect 900 3650 910 3850
rect 980 3650 1330 3850
rect 900 3620 1330 3650
rect 0 3600 120 3620
rect 380 3600 620 3620
rect 880 3600 1330 3620
rect 0 3590 1330 3600
rect 0 3520 150 3590
rect 350 3520 650 3590
rect 850 3520 1330 3590
rect 0 3480 1330 3520
rect 0 3410 150 3480
rect 350 3410 650 3480
rect 850 3410 1330 3480
rect 0 3400 1330 3410
rect 0 3380 120 3400
rect 380 3380 620 3400
rect 880 3380 1330 3400
rect 0 3350 100 3380
rect 0 3150 20 3350
rect 90 3150 100 3350
rect 0 3120 100 3150
rect 400 3350 600 3380
rect 400 3150 410 3350
rect 480 3150 520 3350
rect 590 3150 600 3350
rect 400 3120 600 3150
rect 900 3350 1330 3380
rect 900 3150 910 3350
rect 980 3150 1330 3350
rect 900 3120 1330 3150
rect 0 3100 120 3120
rect 380 3100 620 3120
rect 880 3100 1330 3120
rect 0 3090 1330 3100
rect 0 3020 150 3090
rect 350 3020 650 3090
rect 850 3020 1330 3090
rect 0 2980 1330 3020
rect 0 2910 150 2980
rect 350 2910 650 2980
rect 850 2910 1330 2980
rect 0 2900 1330 2910
rect 0 2880 120 2900
rect 380 2880 620 2900
rect 880 2880 1330 2900
rect 0 2850 100 2880
rect 0 2650 20 2850
rect 90 2650 100 2850
rect 0 2620 100 2650
rect 400 2850 600 2880
rect 400 2650 410 2850
rect 480 2650 520 2850
rect 590 2650 600 2850
rect 400 2620 600 2650
rect 900 2850 1330 2880
rect 900 2650 910 2850
rect 980 2650 1330 2850
rect 900 2620 1330 2650
rect 0 2600 120 2620
rect 380 2600 620 2620
rect 880 2600 1330 2620
rect 0 2590 1330 2600
rect 0 2520 150 2590
rect 350 2520 650 2590
rect 850 2520 1330 2590
rect 0 2480 1330 2520
rect 0 2410 150 2480
rect 350 2410 650 2480
rect 850 2410 1330 2480
rect 0 2400 1330 2410
rect 0 2380 120 2400
rect 380 2380 620 2400
rect 880 2380 1330 2400
rect 0 2350 100 2380
rect 0 2150 20 2350
rect 90 2150 100 2350
rect 0 2120 100 2150
rect 400 2350 600 2380
rect 400 2150 410 2350
rect 480 2150 520 2350
rect 590 2150 600 2350
rect 400 2120 600 2150
rect 900 2350 1330 2380
rect 900 2150 910 2350
rect 980 2200 1330 2350
rect 1465 8346 1531 8358
rect 1465 8338 1482 8346
rect 1516 8338 1531 8346
rect 1465 2370 1482 2378
rect 1516 2370 1531 2378
rect 1465 2358 1531 2370
rect 1623 8346 1689 8358
rect 1623 8338 1640 8346
rect 1674 8338 1689 8346
rect 1623 2370 1640 2378
rect 1674 2370 1689 2378
rect 1623 2358 1689 2370
rect 1781 8346 1847 8358
rect 1781 8338 1798 8346
rect 1832 8338 1847 8346
rect 1781 2370 1798 2378
rect 1832 2370 1847 2378
rect 1781 2358 1847 2370
rect 1939 8346 2005 8358
rect 1939 8338 1956 8346
rect 1990 8338 2005 8346
rect 1939 2370 1956 2378
rect 1990 2370 2005 2378
rect 1939 2358 2005 2370
rect 2097 8346 2163 8358
rect 2097 8338 2114 8346
rect 2148 8338 2163 8346
rect 2097 2370 2114 2378
rect 2148 2370 2163 2378
rect 2097 2358 2163 2370
rect 2255 8346 2321 8358
rect 2255 8338 2272 8346
rect 2306 8338 2321 8346
rect 2255 2370 2272 2378
rect 2306 2370 2321 2378
rect 2255 2358 2321 2370
rect 2413 8346 2479 8358
rect 2413 8338 2430 8346
rect 2464 8338 2479 8346
rect 2413 2370 2430 2378
rect 2464 2370 2479 2378
rect 2413 2358 2479 2370
rect 2571 8346 2637 8358
rect 2571 8338 2588 8346
rect 2622 8338 2637 8346
rect 2571 2370 2588 2378
rect 2622 2370 2637 2378
rect 2571 2358 2637 2370
rect 2729 8346 2795 8358
rect 2729 8338 2746 8346
rect 2780 8338 2795 8346
rect 2729 2370 2746 2378
rect 2780 2370 2795 2378
rect 2729 2358 2795 2370
rect 2887 8346 2953 8358
rect 2887 8338 2904 8346
rect 2938 8338 2953 8346
rect 2887 2370 2904 2378
rect 2938 2370 2953 2378
rect 2887 2358 2953 2370
rect 3045 8346 3111 8358
rect 3045 8338 3062 8346
rect 3096 8338 3111 8346
rect 3045 2370 3062 2378
rect 3096 2370 3111 2378
rect 3045 2358 3111 2370
rect 3203 8346 3269 8358
rect 3203 8338 3220 8346
rect 3254 8338 3269 8346
rect 3203 2370 3220 2378
rect 3254 2370 3269 2378
rect 3203 2358 3269 2370
rect 3361 8346 3427 8358
rect 3361 8338 3378 8346
rect 3412 8338 3427 8346
rect 3361 2370 3378 2378
rect 3412 2370 3427 2378
rect 3361 2358 3427 2370
rect 3519 8346 3585 8358
rect 3519 8338 3536 8346
rect 3570 8338 3585 8346
rect 3519 2370 3536 2378
rect 3570 2370 3585 2378
rect 3519 2358 3585 2370
rect 3677 8346 3743 8358
rect 3677 8338 3694 8346
rect 3728 8338 3743 8346
rect 3677 2370 3694 2378
rect 3728 2370 3743 2378
rect 3677 2358 3743 2370
rect 3835 8346 3901 8358
rect 3835 8338 3852 8346
rect 3886 8338 3901 8346
rect 3835 2370 3852 2378
rect 3886 2370 3901 2378
rect 3835 2358 3901 2370
rect 3993 8346 4059 8358
rect 3993 8338 4010 8346
rect 4044 8338 4059 8346
rect 3993 2370 4010 2378
rect 4044 2370 4059 2378
rect 3993 2358 4059 2370
rect 4151 8346 4217 8358
rect 4151 8338 4168 8346
rect 4202 8338 4217 8346
rect 4151 2370 4168 2378
rect 4202 2370 4217 2378
rect 4151 2358 4217 2370
rect 4309 8346 4375 8358
rect 4309 8338 4326 8346
rect 4360 8338 4375 8346
rect 4309 2370 4326 2378
rect 4360 2370 4375 2378
rect 4309 2358 4375 2370
rect 4467 8346 4533 8358
rect 4467 8338 4484 8346
rect 4518 8338 4533 8346
rect 4467 2370 4484 2378
rect 4518 2370 4533 2378
rect 4467 2358 4533 2370
rect 4625 8346 4691 8358
rect 4625 8338 4642 8346
rect 4676 8338 4691 8346
rect 4625 2370 4642 2378
rect 4676 2370 4691 2378
rect 4625 2358 4691 2370
rect 4783 8346 4849 8358
rect 4783 8338 4800 8346
rect 4834 8338 4849 8346
rect 4783 2370 4800 2378
rect 4834 2370 4849 2378
rect 4783 2358 4849 2370
rect 4941 8346 5007 8358
rect 4941 8338 4958 8346
rect 4992 8338 5007 8346
rect 4941 2370 4958 2378
rect 4992 2370 5007 2378
rect 4941 2358 5007 2370
rect 5099 8346 5165 8358
rect 5099 8338 5116 8346
rect 5150 8338 5165 8346
rect 5099 2370 5116 2378
rect 5150 2370 5165 2378
rect 5099 2358 5165 2370
rect 5257 8346 5323 8358
rect 5257 8338 5274 8346
rect 5308 8338 5323 8346
rect 5257 2370 5274 2378
rect 5308 2370 5323 2378
rect 5257 2358 5323 2370
rect 5415 8346 5481 8358
rect 5415 8338 5432 8346
rect 5466 8338 5481 8346
rect 5415 2370 5432 2378
rect 5466 2370 5481 2378
rect 5415 2358 5481 2370
rect 5573 8346 5639 8358
rect 5573 8338 5590 8346
rect 5624 8338 5639 8346
rect 5573 2370 5590 2378
rect 5624 2370 5639 2378
rect 5573 2358 5639 2370
rect 5731 8346 5797 8358
rect 5731 8338 5748 8346
rect 5782 8338 5797 8346
rect 5731 2370 5748 2378
rect 5782 2370 5797 2378
rect 5731 2358 5797 2370
rect 5889 8346 5955 8358
rect 5889 8338 5906 8346
rect 5940 8338 5955 8346
rect 5889 2370 5906 2378
rect 5940 2370 5955 2378
rect 5889 2358 5955 2370
rect 6047 8346 6113 8358
rect 6047 8338 6064 8346
rect 6098 8338 6113 8346
rect 6047 2370 6064 2378
rect 6098 2370 6113 2378
rect 6047 2358 6113 2370
rect 6205 8346 6271 8358
rect 6205 8338 6222 8346
rect 6256 8338 6271 8346
rect 6205 2370 6222 2378
rect 6256 2370 6271 2378
rect 6205 2358 6271 2370
rect 7630 8570 12710 8580
rect 7630 8532 7836 8570
rect 12559 8532 12710 8570
rect 7630 8522 12710 8532
rect 7630 8520 7700 8522
rect 12640 8520 12710 8522
rect 7832 8430 7852 8490
rect 12486 8430 12506 8490
rect 7832 8396 7844 8430
rect 12494 8396 12506 8430
rect 7832 8390 7852 8396
rect 12486 8390 12506 8396
rect 6410 2480 7630 2500
rect 6410 2410 6650 2480
rect 6850 2410 7150 2480
rect 7350 2410 7630 2480
rect 6410 2400 7630 2410
rect 6410 2380 6620 2400
rect 6880 2380 7120 2400
rect 7380 2380 7630 2400
rect 6410 2350 6600 2380
rect 1532 2320 1552 2326
rect 6186 2320 6206 2326
rect 1532 2286 1544 2320
rect 6194 2286 6206 2320
rect 1532 2226 1552 2286
rect 6186 2226 6206 2286
rect 980 2194 1400 2200
rect 6410 2200 6520 2350
rect 6340 2194 6520 2200
rect 980 2184 6520 2194
rect 980 2150 1536 2184
rect 900 2146 1536 2150
rect 6202 2150 6520 2184
rect 6590 2150 6600 2350
rect 6202 2146 6600 2150
rect 900 2120 6600 2146
rect 6900 2350 7100 2380
rect 6900 2150 6910 2350
rect 6980 2150 7020 2350
rect 7090 2150 7100 2350
rect 6900 2120 7100 2150
rect 7400 2350 7630 2380
rect 7400 2150 7410 2350
rect 7480 2200 7630 2350
rect 7765 8346 7831 8358
rect 7765 8338 7782 8346
rect 7816 8338 7831 8346
rect 7765 2370 7782 2378
rect 7816 2370 7831 2378
rect 7765 2358 7831 2370
rect 7923 8346 7989 8358
rect 7923 8338 7940 8346
rect 7974 8338 7989 8346
rect 7923 2370 7940 2378
rect 7974 2370 7989 2378
rect 7923 2358 7989 2370
rect 8081 8346 8147 8358
rect 8081 8338 8098 8346
rect 8132 8338 8147 8346
rect 8081 2370 8098 2378
rect 8132 2370 8147 2378
rect 8081 2358 8147 2370
rect 8239 8346 8305 8358
rect 8239 8338 8256 8346
rect 8290 8338 8305 8346
rect 8239 2370 8256 2378
rect 8290 2370 8305 2378
rect 8239 2358 8305 2370
rect 8397 8346 8463 8358
rect 8397 8338 8414 8346
rect 8448 8338 8463 8346
rect 8397 2370 8414 2378
rect 8448 2370 8463 2378
rect 8397 2358 8463 2370
rect 8555 8346 8621 8358
rect 8555 8338 8572 8346
rect 8606 8338 8621 8346
rect 8555 2370 8572 2378
rect 8606 2370 8621 2378
rect 8555 2358 8621 2370
rect 8713 8346 8779 8358
rect 8713 8338 8730 8346
rect 8764 8338 8779 8346
rect 8713 2370 8730 2378
rect 8764 2370 8779 2378
rect 8713 2358 8779 2370
rect 8871 8346 8937 8358
rect 8871 8338 8888 8346
rect 8922 8338 8937 8346
rect 8871 2370 8888 2378
rect 8922 2370 8937 2378
rect 8871 2358 8937 2370
rect 9029 8346 9095 8358
rect 9029 8338 9046 8346
rect 9080 8338 9095 8346
rect 9029 2370 9046 2378
rect 9080 2370 9095 2378
rect 9029 2358 9095 2370
rect 9187 8346 9253 8358
rect 9187 8338 9204 8346
rect 9238 8338 9253 8346
rect 9187 2370 9204 2378
rect 9238 2370 9253 2378
rect 9187 2358 9253 2370
rect 9345 8346 9411 8358
rect 9345 8338 9362 8346
rect 9396 8338 9411 8346
rect 9345 2370 9362 2378
rect 9396 2370 9411 2378
rect 9345 2358 9411 2370
rect 9503 8346 9569 8358
rect 9503 8338 9520 8346
rect 9554 8338 9569 8346
rect 9503 2370 9520 2378
rect 9554 2370 9569 2378
rect 9503 2358 9569 2370
rect 9661 8346 9727 8358
rect 9661 8338 9678 8346
rect 9712 8338 9727 8346
rect 9661 2370 9678 2378
rect 9712 2370 9727 2378
rect 9661 2358 9727 2370
rect 9819 8346 9885 8358
rect 9819 8338 9836 8346
rect 9870 8338 9885 8346
rect 9819 2370 9836 2378
rect 9870 2370 9885 2378
rect 9819 2358 9885 2370
rect 9977 8346 10043 8358
rect 9977 8338 9994 8346
rect 10028 8338 10043 8346
rect 9977 2370 9994 2378
rect 10028 2370 10043 2378
rect 9977 2358 10043 2370
rect 10135 8346 10201 8358
rect 10135 8338 10152 8346
rect 10186 8338 10201 8346
rect 10135 2370 10152 2378
rect 10186 2370 10201 2378
rect 10135 2358 10201 2370
rect 10293 8346 10359 8358
rect 10293 8338 10310 8346
rect 10344 8338 10359 8346
rect 10293 2370 10310 2378
rect 10344 2370 10359 2378
rect 10293 2358 10359 2370
rect 10451 8346 10517 8358
rect 10451 8338 10468 8346
rect 10502 8338 10517 8346
rect 10451 2370 10468 2378
rect 10502 2370 10517 2378
rect 10451 2358 10517 2370
rect 10609 8346 10675 8358
rect 10609 8338 10626 8346
rect 10660 8338 10675 8346
rect 10609 2370 10626 2378
rect 10660 2370 10675 2378
rect 10609 2358 10675 2370
rect 10767 8346 10833 8358
rect 10767 8338 10784 8346
rect 10818 8338 10833 8346
rect 10767 2370 10784 2378
rect 10818 2370 10833 2378
rect 10767 2358 10833 2370
rect 10925 8346 10991 8358
rect 10925 8338 10942 8346
rect 10976 8338 10991 8346
rect 10925 2370 10942 2378
rect 10976 2370 10991 2378
rect 10925 2358 10991 2370
rect 11083 8346 11149 8358
rect 11083 8338 11100 8346
rect 11134 8338 11149 8346
rect 11083 2370 11100 2378
rect 11134 2370 11149 2378
rect 11083 2358 11149 2370
rect 11241 8346 11307 8358
rect 11241 8338 11258 8346
rect 11292 8338 11307 8346
rect 11241 2370 11258 2378
rect 11292 2370 11307 2378
rect 11241 2358 11307 2370
rect 11399 8346 11465 8358
rect 11399 8338 11416 8346
rect 11450 8338 11465 8346
rect 11399 2370 11416 2378
rect 11450 2370 11465 2378
rect 11399 2358 11465 2370
rect 11557 8346 11623 8358
rect 11557 8338 11574 8346
rect 11608 8338 11623 8346
rect 11557 2370 11574 2378
rect 11608 2370 11623 2378
rect 11557 2358 11623 2370
rect 11715 8346 11781 8358
rect 11715 8338 11732 8346
rect 11766 8338 11781 8346
rect 11715 2370 11732 2378
rect 11766 2370 11781 2378
rect 11715 2358 11781 2370
rect 11873 8346 11939 8358
rect 11873 8338 11890 8346
rect 11924 8338 11939 8346
rect 11873 2370 11890 2378
rect 11924 2370 11939 2378
rect 11873 2358 11939 2370
rect 12031 8346 12097 8358
rect 12031 8338 12048 8346
rect 12082 8338 12097 8346
rect 12031 2370 12048 2378
rect 12082 2370 12097 2378
rect 12031 2358 12097 2370
rect 12189 8346 12255 8358
rect 12189 8338 12206 8346
rect 12240 8338 12255 8346
rect 12189 2370 12206 2378
rect 12240 2370 12255 2378
rect 12189 2358 12255 2370
rect 12347 8346 12413 8358
rect 12347 8338 12364 8346
rect 12398 8338 12413 8346
rect 12347 2370 12364 2378
rect 12398 2370 12413 2378
rect 12347 2358 12413 2370
rect 12505 8346 12571 8358
rect 12505 8338 12522 8346
rect 12556 8338 12571 8346
rect 12505 2370 12522 2378
rect 12556 2370 12571 2378
rect 12505 2358 12571 2370
rect 13930 8570 19010 8580
rect 13930 8532 14136 8570
rect 18859 8532 19010 8570
rect 13930 8522 19010 8532
rect 13930 8520 14000 8522
rect 18940 8520 19010 8522
rect 14132 8430 14152 8490
rect 18786 8430 18806 8490
rect 14132 8396 14144 8430
rect 18794 8396 18806 8430
rect 14132 8390 14152 8396
rect 18786 8390 18806 8396
rect 12710 2480 13930 2500
rect 12710 2410 13150 2480
rect 13350 2410 13930 2480
rect 12710 2400 13930 2410
rect 12710 2380 13120 2400
rect 13380 2380 13930 2400
rect 12710 2350 13100 2380
rect 7832 2320 7852 2326
rect 12486 2320 12506 2326
rect 7832 2286 7844 2320
rect 12494 2286 12506 2320
rect 7832 2226 7852 2286
rect 12486 2226 12506 2286
rect 7480 2194 7700 2200
rect 12710 2200 13020 2350
rect 12640 2194 13020 2200
rect 7480 2184 13020 2194
rect 7480 2150 7836 2184
rect 7400 2146 7836 2150
rect 12502 2150 13020 2184
rect 13090 2150 13100 2350
rect 12502 2146 13100 2150
rect 7400 2120 13100 2146
rect 13400 2350 13930 2380
rect 13400 2150 13410 2350
rect 13480 2200 13930 2350
rect 14065 8346 14131 8358
rect 14065 8338 14082 8346
rect 14116 8338 14131 8346
rect 14065 2370 14082 2378
rect 14116 2370 14131 2378
rect 14065 2358 14131 2370
rect 14223 8346 14289 8358
rect 14223 8338 14240 8346
rect 14274 8338 14289 8346
rect 14223 2370 14240 2378
rect 14274 2370 14289 2378
rect 14223 2358 14289 2370
rect 14381 8346 14447 8358
rect 14381 8338 14398 8346
rect 14432 8338 14447 8346
rect 14381 2370 14398 2378
rect 14432 2370 14447 2378
rect 14381 2358 14447 2370
rect 14539 8346 14605 8358
rect 14539 8338 14556 8346
rect 14590 8338 14605 8346
rect 14539 2370 14556 2378
rect 14590 2370 14605 2378
rect 14539 2358 14605 2370
rect 14697 8346 14763 8358
rect 14697 8338 14714 8346
rect 14748 8338 14763 8346
rect 14697 2370 14714 2378
rect 14748 2370 14763 2378
rect 14697 2358 14763 2370
rect 14855 8346 14921 8358
rect 14855 8338 14872 8346
rect 14906 8338 14921 8346
rect 14855 2370 14872 2378
rect 14906 2370 14921 2378
rect 14855 2358 14921 2370
rect 15013 8346 15079 8358
rect 15013 8338 15030 8346
rect 15064 8338 15079 8346
rect 15013 2370 15030 2378
rect 15064 2370 15079 2378
rect 15013 2358 15079 2370
rect 15171 8346 15237 8358
rect 15171 8338 15188 8346
rect 15222 8338 15237 8346
rect 15171 2370 15188 2378
rect 15222 2370 15237 2378
rect 15171 2358 15237 2370
rect 15329 8346 15395 8358
rect 15329 8338 15346 8346
rect 15380 8338 15395 8346
rect 15329 2370 15346 2378
rect 15380 2370 15395 2378
rect 15329 2358 15395 2370
rect 15487 8346 15553 8358
rect 15487 8338 15504 8346
rect 15538 8338 15553 8346
rect 15487 2370 15504 2378
rect 15538 2370 15553 2378
rect 15487 2358 15553 2370
rect 15645 8346 15711 8358
rect 15645 8338 15662 8346
rect 15696 8338 15711 8346
rect 15645 2370 15662 2378
rect 15696 2370 15711 2378
rect 15645 2358 15711 2370
rect 15803 8346 15869 8358
rect 15803 8338 15820 8346
rect 15854 8338 15869 8346
rect 15803 2370 15820 2378
rect 15854 2370 15869 2378
rect 15803 2358 15869 2370
rect 15961 8346 16027 8358
rect 15961 8338 15978 8346
rect 16012 8338 16027 8346
rect 15961 2370 15978 2378
rect 16012 2370 16027 2378
rect 15961 2358 16027 2370
rect 16119 8346 16185 8358
rect 16119 8338 16136 8346
rect 16170 8338 16185 8346
rect 16119 2370 16136 2378
rect 16170 2370 16185 2378
rect 16119 2358 16185 2370
rect 16277 8346 16343 8358
rect 16277 8338 16294 8346
rect 16328 8338 16343 8346
rect 16277 2370 16294 2378
rect 16328 2370 16343 2378
rect 16277 2358 16343 2370
rect 16435 8346 16501 8358
rect 16435 8338 16452 8346
rect 16486 8338 16501 8346
rect 16435 2370 16452 2378
rect 16486 2370 16501 2378
rect 16435 2358 16501 2370
rect 16593 8346 16659 8358
rect 16593 8338 16610 8346
rect 16644 8338 16659 8346
rect 16593 2370 16610 2378
rect 16644 2370 16659 2378
rect 16593 2358 16659 2370
rect 16751 8346 16817 8358
rect 16751 8338 16768 8346
rect 16802 8338 16817 8346
rect 16751 2370 16768 2378
rect 16802 2370 16817 2378
rect 16751 2358 16817 2370
rect 16909 8346 16975 8358
rect 16909 8338 16926 8346
rect 16960 8338 16975 8346
rect 16909 2370 16926 2378
rect 16960 2370 16975 2378
rect 16909 2358 16975 2370
rect 17067 8346 17133 8358
rect 17067 8338 17084 8346
rect 17118 8338 17133 8346
rect 17067 2370 17084 2378
rect 17118 2370 17133 2378
rect 17067 2358 17133 2370
rect 17225 8346 17291 8358
rect 17225 8338 17242 8346
rect 17276 8338 17291 8346
rect 17225 2370 17242 2378
rect 17276 2370 17291 2378
rect 17225 2358 17291 2370
rect 17383 8346 17449 8358
rect 17383 8338 17400 8346
rect 17434 8338 17449 8346
rect 17383 2370 17400 2378
rect 17434 2370 17449 2378
rect 17383 2358 17449 2370
rect 17541 8346 17607 8358
rect 17541 8338 17558 8346
rect 17592 8338 17607 8346
rect 17541 2370 17558 2378
rect 17592 2370 17607 2378
rect 17541 2358 17607 2370
rect 17699 8346 17765 8358
rect 17699 8338 17716 8346
rect 17750 8338 17765 8346
rect 17699 2370 17716 2378
rect 17750 2370 17765 2378
rect 17699 2358 17765 2370
rect 17857 8346 17923 8358
rect 17857 8338 17874 8346
rect 17908 8338 17923 8346
rect 17857 2370 17874 2378
rect 17908 2370 17923 2378
rect 17857 2358 17923 2370
rect 18015 8346 18081 8358
rect 18015 8338 18032 8346
rect 18066 8338 18081 8346
rect 18015 2370 18032 2378
rect 18066 2370 18081 2378
rect 18015 2358 18081 2370
rect 18173 8346 18239 8358
rect 18173 8338 18190 8346
rect 18224 8338 18239 8346
rect 18173 2370 18190 2378
rect 18224 2370 18239 2378
rect 18173 2358 18239 2370
rect 18331 8346 18397 8358
rect 18331 8338 18348 8346
rect 18382 8338 18397 8346
rect 18331 2370 18348 2378
rect 18382 2370 18397 2378
rect 18331 2358 18397 2370
rect 18489 8346 18555 8358
rect 18489 8338 18506 8346
rect 18540 8338 18555 8346
rect 18489 2370 18506 2378
rect 18540 2370 18555 2378
rect 18489 2358 18555 2370
rect 18647 8346 18713 8358
rect 18647 8338 18664 8346
rect 18698 8338 18713 8346
rect 18647 2370 18664 2378
rect 18698 2370 18713 2378
rect 18647 2358 18713 2370
rect 18805 8346 18871 8358
rect 18805 8338 18822 8346
rect 18856 8338 18871 8346
rect 18805 2370 18822 2378
rect 18856 2370 18871 2378
rect 18805 2358 18871 2370
rect 20230 8570 25650 8580
rect 20230 8532 20436 8570
rect 25159 8532 25650 8570
rect 20230 8522 25650 8532
rect 20230 8520 20300 8522
rect 25240 8520 25650 8522
rect 25850 8520 26150 8590
rect 26350 8520 26500 8590
rect 20432 8430 20452 8490
rect 25086 8430 25106 8490
rect 20432 8396 20444 8430
rect 25094 8396 25106 8430
rect 20432 8390 20452 8396
rect 25086 8390 25106 8396
rect 19010 2480 20230 2500
rect 19010 2410 19650 2480
rect 19850 2410 20230 2480
rect 19010 2400 20230 2410
rect 19010 2380 19620 2400
rect 19880 2380 20230 2400
rect 19010 2350 19600 2380
rect 14132 2320 14152 2326
rect 18786 2320 18806 2326
rect 14132 2286 14144 2320
rect 18794 2286 18806 2320
rect 14132 2226 14152 2286
rect 18786 2226 18806 2286
rect 13480 2194 14000 2200
rect 19010 2200 19520 2350
rect 18940 2194 19520 2200
rect 13480 2184 19520 2194
rect 13480 2150 14136 2184
rect 13400 2146 14136 2150
rect 18802 2150 19520 2184
rect 19590 2150 19600 2350
rect 18802 2146 19600 2150
rect 13400 2120 19600 2146
rect 19900 2350 20230 2380
rect 19900 2150 19910 2350
rect 19980 2200 20230 2350
rect 25310 8480 26500 8520
rect 25310 8410 25650 8480
rect 25850 8410 26150 8480
rect 26350 8410 26500 8480
rect 25310 8400 26500 8410
rect 25310 8380 25620 8400
rect 25880 8380 26120 8400
rect 26380 8380 26500 8400
rect 20365 8346 20431 8358
rect 20365 8338 20382 8346
rect 20416 8338 20431 8346
rect 20365 2370 20382 2378
rect 20416 2370 20431 2378
rect 20365 2358 20431 2370
rect 20523 8346 20589 8358
rect 20523 8338 20540 8346
rect 20574 8338 20589 8346
rect 20523 2370 20540 2378
rect 20574 2370 20589 2378
rect 20523 2358 20589 2370
rect 20681 8346 20747 8358
rect 20681 8338 20698 8346
rect 20732 8338 20747 8346
rect 20681 2370 20698 2378
rect 20732 2370 20747 2378
rect 20681 2358 20747 2370
rect 20839 8346 20905 8358
rect 20839 8338 20856 8346
rect 20890 8338 20905 8346
rect 20839 2370 20856 2378
rect 20890 2370 20905 2378
rect 20839 2358 20905 2370
rect 20997 8346 21063 8358
rect 20997 8338 21014 8346
rect 21048 8338 21063 8346
rect 20997 2370 21014 2378
rect 21048 2370 21063 2378
rect 20997 2358 21063 2370
rect 21155 8346 21221 8358
rect 21155 8338 21172 8346
rect 21206 8338 21221 8346
rect 21155 2370 21172 2378
rect 21206 2370 21221 2378
rect 21155 2358 21221 2370
rect 21313 8346 21379 8358
rect 21313 8338 21330 8346
rect 21364 8338 21379 8346
rect 21313 2370 21330 2378
rect 21364 2370 21379 2378
rect 21313 2358 21379 2370
rect 21471 8346 21537 8358
rect 21471 8338 21488 8346
rect 21522 8338 21537 8346
rect 21471 2370 21488 2378
rect 21522 2370 21537 2378
rect 21471 2358 21537 2370
rect 21629 8346 21695 8358
rect 21629 8338 21646 8346
rect 21680 8338 21695 8346
rect 21629 2370 21646 2378
rect 21680 2370 21695 2378
rect 21629 2358 21695 2370
rect 21787 8346 21853 8358
rect 21787 8338 21804 8346
rect 21838 8338 21853 8346
rect 21787 2370 21804 2378
rect 21838 2370 21853 2378
rect 21787 2358 21853 2370
rect 21945 8346 22011 8358
rect 21945 8338 21962 8346
rect 21996 8338 22011 8346
rect 21945 2370 21962 2378
rect 21996 2370 22011 2378
rect 21945 2358 22011 2370
rect 22103 8346 22169 8358
rect 22103 8338 22120 8346
rect 22154 8338 22169 8346
rect 22103 2370 22120 2378
rect 22154 2370 22169 2378
rect 22103 2358 22169 2370
rect 22261 8346 22327 8358
rect 22261 8338 22278 8346
rect 22312 8338 22327 8346
rect 22261 2370 22278 2378
rect 22312 2370 22327 2378
rect 22261 2358 22327 2370
rect 22419 8346 22485 8358
rect 22419 8338 22436 8346
rect 22470 8338 22485 8346
rect 22419 2370 22436 2378
rect 22470 2370 22485 2378
rect 22419 2358 22485 2370
rect 22577 8346 22643 8358
rect 22577 8338 22594 8346
rect 22628 8338 22643 8346
rect 22577 2370 22594 2378
rect 22628 2370 22643 2378
rect 22577 2358 22643 2370
rect 22735 8346 22801 8358
rect 22735 8338 22752 8346
rect 22786 8338 22801 8346
rect 22735 2370 22752 2378
rect 22786 2370 22801 2378
rect 22735 2358 22801 2370
rect 22893 8346 22959 8358
rect 22893 8338 22910 8346
rect 22944 8338 22959 8346
rect 22893 2370 22910 2378
rect 22944 2370 22959 2378
rect 22893 2358 22959 2370
rect 23051 8346 23117 8358
rect 23051 8338 23068 8346
rect 23102 8338 23117 8346
rect 23051 2370 23068 2378
rect 23102 2370 23117 2378
rect 23051 2358 23117 2370
rect 23209 8346 23275 8358
rect 23209 8338 23226 8346
rect 23260 8338 23275 8346
rect 23209 2370 23226 2378
rect 23260 2370 23275 2378
rect 23209 2358 23275 2370
rect 23367 8346 23433 8358
rect 23367 8338 23384 8346
rect 23418 8338 23433 8346
rect 23367 2370 23384 2378
rect 23418 2370 23433 2378
rect 23367 2358 23433 2370
rect 23525 8346 23591 8358
rect 23525 8338 23542 8346
rect 23576 8338 23591 8346
rect 23525 2370 23542 2378
rect 23576 2370 23591 2378
rect 23525 2358 23591 2370
rect 23683 8346 23749 8358
rect 23683 8338 23700 8346
rect 23734 8338 23749 8346
rect 23683 2370 23700 2378
rect 23734 2370 23749 2378
rect 23683 2358 23749 2370
rect 23841 8346 23907 8358
rect 23841 8338 23858 8346
rect 23892 8338 23907 8346
rect 23841 2370 23858 2378
rect 23892 2370 23907 2378
rect 23841 2358 23907 2370
rect 23999 8346 24065 8358
rect 23999 8338 24016 8346
rect 24050 8338 24065 8346
rect 23999 2370 24016 2378
rect 24050 2370 24065 2378
rect 23999 2358 24065 2370
rect 24157 8346 24223 8358
rect 24157 8338 24174 8346
rect 24208 8338 24223 8346
rect 24157 2370 24174 2378
rect 24208 2370 24223 2378
rect 24157 2358 24223 2370
rect 24315 8346 24381 8358
rect 24315 8338 24332 8346
rect 24366 8338 24381 8346
rect 24315 2370 24332 2378
rect 24366 2370 24381 2378
rect 24315 2358 24381 2370
rect 24473 8346 24539 8358
rect 24473 8338 24490 8346
rect 24524 8338 24539 8346
rect 24473 2370 24490 2378
rect 24524 2370 24539 2378
rect 24473 2358 24539 2370
rect 24631 8346 24697 8358
rect 24631 8338 24648 8346
rect 24682 8338 24697 8346
rect 24631 2370 24648 2378
rect 24682 2370 24697 2378
rect 24631 2358 24697 2370
rect 24789 8346 24855 8358
rect 24789 8338 24806 8346
rect 24840 8338 24855 8346
rect 24789 2370 24806 2378
rect 24840 2370 24855 2378
rect 24789 2358 24855 2370
rect 24947 8346 25013 8358
rect 24947 8338 24964 8346
rect 24998 8338 25013 8346
rect 24947 2370 24964 2378
rect 24998 2370 25013 2378
rect 24947 2358 25013 2370
rect 25105 8346 25171 8358
rect 25105 8338 25122 8346
rect 25156 8338 25171 8346
rect 25105 2370 25122 2378
rect 25156 2370 25171 2378
rect 25105 2358 25171 2370
rect 25310 8350 25600 8380
rect 25310 8150 25520 8350
rect 25590 8150 25600 8350
rect 25310 8120 25600 8150
rect 25900 8350 26100 8380
rect 25900 8150 25910 8350
rect 25980 8150 26020 8350
rect 26090 8150 26100 8350
rect 25900 8120 26100 8150
rect 26400 8350 26500 8380
rect 26400 8150 26410 8350
rect 26480 8150 26500 8350
rect 26400 8120 26500 8150
rect 25310 8100 25620 8120
rect 25880 8100 26120 8120
rect 26380 8100 26500 8120
rect 25310 8090 26500 8100
rect 25310 8020 25650 8090
rect 25850 8020 26150 8090
rect 26350 8020 26500 8090
rect 25310 7980 26500 8020
rect 25310 7910 25650 7980
rect 25850 7910 26150 7980
rect 26350 7910 26500 7980
rect 25310 7900 26500 7910
rect 25310 7880 25620 7900
rect 25880 7880 26120 7900
rect 26380 7880 26500 7900
rect 25310 7850 25600 7880
rect 25310 7650 25520 7850
rect 25590 7650 25600 7850
rect 25310 7620 25600 7650
rect 25900 7850 26100 7880
rect 25900 7650 25910 7850
rect 25980 7650 26020 7850
rect 26090 7650 26100 7850
rect 25900 7620 26100 7650
rect 26400 7850 26500 7880
rect 26400 7650 26410 7850
rect 26480 7650 26500 7850
rect 26400 7620 26500 7650
rect 25310 7600 25620 7620
rect 25880 7600 26120 7620
rect 26380 7600 26500 7620
rect 25310 7590 26500 7600
rect 25310 7520 25650 7590
rect 25850 7520 26150 7590
rect 26350 7520 26500 7590
rect 25310 7480 26500 7520
rect 25310 7410 25650 7480
rect 25850 7410 26150 7480
rect 26350 7410 26500 7480
rect 25310 7400 26500 7410
rect 25310 7380 25620 7400
rect 25880 7380 26120 7400
rect 26380 7380 26500 7400
rect 25310 7350 25600 7380
rect 25310 7150 25520 7350
rect 25590 7150 25600 7350
rect 25310 7120 25600 7150
rect 25900 7350 26100 7380
rect 25900 7150 25910 7350
rect 25980 7150 26020 7350
rect 26090 7150 26100 7350
rect 25900 7120 26100 7150
rect 26400 7350 26500 7380
rect 26400 7150 26410 7350
rect 26480 7150 26500 7350
rect 26400 7120 26500 7150
rect 25310 7100 25620 7120
rect 25880 7100 26120 7120
rect 26380 7100 26500 7120
rect 25310 7090 26500 7100
rect 25310 7020 25650 7090
rect 25850 7020 26150 7090
rect 26350 7020 26500 7090
rect 25310 6980 26500 7020
rect 25310 6910 25650 6980
rect 25850 6910 26150 6980
rect 26350 6910 26500 6980
rect 25310 6900 26500 6910
rect 25310 6880 25620 6900
rect 25880 6880 26120 6900
rect 26380 6880 26500 6900
rect 25310 6850 25600 6880
rect 25310 6650 25520 6850
rect 25590 6650 25600 6850
rect 25310 6620 25600 6650
rect 25900 6850 26100 6880
rect 25900 6650 25910 6850
rect 25980 6650 26020 6850
rect 26090 6650 26100 6850
rect 25900 6620 26100 6650
rect 26400 6850 26500 6880
rect 26400 6650 26410 6850
rect 26480 6650 26500 6850
rect 26400 6620 26500 6650
rect 25310 6600 25620 6620
rect 25880 6600 26120 6620
rect 26380 6600 26500 6620
rect 25310 6590 26500 6600
rect 25310 6520 25650 6590
rect 25850 6520 26150 6590
rect 26350 6520 26500 6590
rect 25310 6480 26500 6520
rect 25310 6410 25650 6480
rect 25850 6410 26150 6480
rect 26350 6410 26500 6480
rect 25310 6400 26500 6410
rect 25310 6380 25620 6400
rect 25880 6380 26120 6400
rect 26380 6380 26500 6400
rect 25310 6350 25600 6380
rect 25310 6150 25520 6350
rect 25590 6150 25600 6350
rect 25310 6120 25600 6150
rect 25900 6350 26100 6380
rect 25900 6150 25910 6350
rect 25980 6150 26020 6350
rect 26090 6150 26100 6350
rect 25900 6120 26100 6150
rect 26400 6350 26500 6380
rect 26400 6150 26410 6350
rect 26480 6150 26500 6350
rect 26400 6120 26500 6150
rect 25310 6100 25620 6120
rect 25880 6100 26120 6120
rect 26380 6100 26500 6120
rect 25310 6090 26500 6100
rect 25310 6020 25650 6090
rect 25850 6020 26150 6090
rect 26350 6020 26500 6090
rect 25310 5980 26500 6020
rect 25310 5910 25650 5980
rect 25850 5910 26150 5980
rect 26350 5910 26500 5980
rect 25310 5900 26500 5910
rect 25310 5880 25620 5900
rect 25880 5880 26120 5900
rect 26380 5880 26500 5900
rect 25310 5850 25600 5880
rect 25310 5650 25520 5850
rect 25590 5650 25600 5850
rect 25310 5620 25600 5650
rect 25900 5850 26100 5880
rect 25900 5650 25910 5850
rect 25980 5650 26020 5850
rect 26090 5650 26100 5850
rect 25900 5620 26100 5650
rect 26400 5850 26500 5880
rect 26400 5650 26410 5850
rect 26480 5650 26500 5850
rect 26400 5620 26500 5650
rect 25310 5600 25620 5620
rect 25880 5600 26120 5620
rect 26380 5600 26500 5620
rect 25310 5590 26500 5600
rect 25310 5520 25650 5590
rect 25850 5520 26150 5590
rect 26350 5520 26500 5590
rect 25310 5480 26500 5520
rect 25310 5410 25650 5480
rect 25850 5410 26150 5480
rect 26350 5410 26500 5480
rect 25310 5400 26500 5410
rect 25310 5380 25620 5400
rect 25880 5380 26120 5400
rect 26380 5380 26500 5400
rect 25310 5350 25600 5380
rect 25310 5150 25520 5350
rect 25590 5150 25600 5350
rect 25310 5120 25600 5150
rect 25900 5350 26100 5380
rect 25900 5150 25910 5350
rect 25980 5150 26020 5350
rect 26090 5150 26100 5350
rect 25900 5120 26100 5150
rect 26400 5350 26500 5380
rect 26400 5150 26410 5350
rect 26480 5150 26500 5350
rect 26400 5120 26500 5150
rect 25310 5100 25620 5120
rect 25880 5100 26120 5120
rect 26380 5100 26500 5120
rect 25310 5090 26500 5100
rect 25310 5020 25650 5090
rect 25850 5020 26150 5090
rect 26350 5020 26500 5090
rect 25310 4980 26500 5020
rect 25310 4910 25650 4980
rect 25850 4910 26150 4980
rect 26350 4910 26500 4980
rect 25310 4900 26500 4910
rect 25310 4880 25620 4900
rect 25880 4880 26120 4900
rect 26380 4880 26500 4900
rect 25310 4850 25600 4880
rect 25310 4650 25520 4850
rect 25590 4650 25600 4850
rect 25310 4620 25600 4650
rect 25900 4850 26100 4880
rect 25900 4650 25910 4850
rect 25980 4650 26020 4850
rect 26090 4650 26100 4850
rect 25900 4620 26100 4650
rect 26400 4850 26500 4880
rect 26400 4650 26410 4850
rect 26480 4650 26500 4850
rect 26400 4620 26500 4650
rect 25310 4600 25620 4620
rect 25880 4600 26120 4620
rect 26380 4600 26500 4620
rect 25310 4590 26500 4600
rect 25310 4520 25650 4590
rect 25850 4520 26150 4590
rect 26350 4520 26500 4590
rect 25310 4480 26500 4520
rect 25310 4410 25650 4480
rect 25850 4410 26150 4480
rect 26350 4410 26500 4480
rect 25310 4400 26500 4410
rect 25310 4380 25620 4400
rect 25880 4380 26120 4400
rect 26380 4380 26500 4400
rect 25310 4350 25600 4380
rect 25310 4150 25520 4350
rect 25590 4150 25600 4350
rect 25310 4120 25600 4150
rect 25900 4350 26100 4380
rect 25900 4150 25910 4350
rect 25980 4150 26020 4350
rect 26090 4150 26100 4350
rect 25900 4120 26100 4150
rect 26400 4350 26500 4380
rect 26400 4150 26410 4350
rect 26480 4150 26500 4350
rect 26400 4120 26500 4150
rect 25310 4100 25620 4120
rect 25880 4100 26120 4120
rect 26380 4100 26500 4120
rect 25310 4090 26500 4100
rect 25310 4020 25650 4090
rect 25850 4020 26150 4090
rect 26350 4020 26500 4090
rect 25310 3980 26500 4020
rect 25310 3910 25650 3980
rect 25850 3910 26150 3980
rect 26350 3910 26500 3980
rect 25310 3900 26500 3910
rect 25310 3880 25620 3900
rect 25880 3880 26120 3900
rect 26380 3880 26500 3900
rect 25310 3850 25600 3880
rect 25310 3650 25520 3850
rect 25590 3650 25600 3850
rect 25310 3620 25600 3650
rect 25900 3850 26100 3880
rect 25900 3650 25910 3850
rect 25980 3650 26020 3850
rect 26090 3650 26100 3850
rect 25900 3620 26100 3650
rect 26400 3850 26500 3880
rect 26400 3650 26410 3850
rect 26480 3650 26500 3850
rect 26400 3620 26500 3650
rect 25310 3600 25620 3620
rect 25880 3600 26120 3620
rect 26380 3600 26500 3620
rect 25310 3590 26500 3600
rect 25310 3520 25650 3590
rect 25850 3520 26150 3590
rect 26350 3520 26500 3590
rect 25310 3480 26500 3520
rect 25310 3410 25650 3480
rect 25850 3410 26150 3480
rect 26350 3410 26500 3480
rect 25310 3400 26500 3410
rect 25310 3380 25620 3400
rect 25880 3380 26120 3400
rect 26380 3380 26500 3400
rect 25310 3350 25600 3380
rect 25310 3150 25520 3350
rect 25590 3150 25600 3350
rect 25310 3120 25600 3150
rect 25900 3350 26100 3380
rect 25900 3150 25910 3350
rect 25980 3150 26020 3350
rect 26090 3150 26100 3350
rect 25900 3120 26100 3150
rect 26400 3350 26500 3380
rect 26400 3150 26410 3350
rect 26480 3150 26500 3350
rect 26400 3120 26500 3150
rect 25310 3100 25620 3120
rect 25880 3100 26120 3120
rect 26380 3100 26500 3120
rect 25310 3090 26500 3100
rect 25310 3020 25650 3090
rect 25850 3020 26150 3090
rect 26350 3020 26500 3090
rect 25310 2980 26500 3020
rect 25310 2910 25650 2980
rect 25850 2910 26150 2980
rect 26350 2910 26500 2980
rect 25310 2900 26500 2910
rect 25310 2880 25620 2900
rect 25880 2880 26120 2900
rect 26380 2880 26500 2900
rect 25310 2850 25600 2880
rect 25310 2650 25520 2850
rect 25590 2650 25600 2850
rect 25310 2620 25600 2650
rect 25900 2850 26100 2880
rect 25900 2650 25910 2850
rect 25980 2650 26020 2850
rect 26090 2650 26100 2850
rect 25900 2620 26100 2650
rect 26400 2850 26500 2880
rect 26400 2650 26410 2850
rect 26480 2650 26500 2850
rect 26400 2620 26500 2650
rect 25310 2600 25620 2620
rect 25880 2600 26120 2620
rect 26380 2600 26500 2620
rect 25310 2590 26500 2600
rect 25310 2520 25650 2590
rect 25850 2520 26150 2590
rect 26350 2520 26500 2590
rect 25310 2480 26500 2520
rect 25310 2410 25650 2480
rect 25850 2410 26150 2480
rect 26350 2410 26500 2480
rect 25310 2400 26500 2410
rect 25310 2380 25620 2400
rect 25880 2380 26120 2400
rect 26380 2380 26500 2400
rect 25310 2350 25600 2380
rect 20432 2320 20452 2326
rect 25086 2320 25106 2326
rect 20432 2286 20444 2320
rect 25094 2286 25106 2320
rect 20432 2226 20452 2286
rect 25086 2226 25106 2286
rect 19980 2194 20300 2200
rect 25310 2200 25520 2350
rect 25240 2194 25520 2200
rect 19980 2184 25520 2194
rect 19980 2150 20436 2184
rect 19900 2146 20436 2150
rect 25102 2150 25520 2184
rect 25590 2150 25600 2350
rect 25102 2146 25600 2150
rect 19900 2120 25600 2146
rect 25900 2350 26100 2380
rect 25900 2150 25910 2350
rect 25980 2150 26020 2350
rect 26090 2150 26100 2350
rect 25900 2120 26100 2150
rect 26400 2350 26500 2380
rect 26400 2150 26410 2350
rect 26480 2150 26500 2350
rect 26400 2120 26500 2150
rect 0 2100 120 2120
rect 380 2100 620 2120
rect 880 2100 6620 2120
rect 6880 2100 7120 2120
rect 7380 2100 13120 2120
rect 13380 2100 19620 2120
rect 19880 2100 25620 2120
rect 25880 2100 26120 2120
rect 26380 2100 26500 2120
rect 0 2090 26500 2100
rect 0 2020 150 2090
rect 350 2020 650 2090
rect 850 2020 6650 2090
rect 6850 2020 7150 2090
rect 7350 2020 13150 2090
rect 13350 2020 19650 2090
rect 19850 2020 25650 2090
rect 25850 2020 26150 2090
rect 26350 2020 26500 2090
rect 0 1980 26500 2020
rect 0 1910 150 1980
rect 350 1910 650 1980
rect 850 1910 1150 1980
rect 1350 1910 1650 1980
rect 1850 1910 2150 1980
rect 2350 1910 2650 1980
rect 2850 1910 3150 1980
rect 3350 1910 3650 1980
rect 3850 1910 4150 1980
rect 4350 1910 4650 1980
rect 4850 1910 5150 1980
rect 5350 1910 5650 1980
rect 5850 1910 6150 1980
rect 6350 1910 6650 1980
rect 6850 1910 7150 1980
rect 7350 1910 7650 1980
rect 7850 1910 8150 1980
rect 8350 1910 8650 1980
rect 8850 1910 9150 1980
rect 9350 1910 9650 1980
rect 9850 1910 10150 1980
rect 10350 1910 10650 1980
rect 10850 1910 11150 1980
rect 11350 1910 11650 1980
rect 11850 1910 12150 1980
rect 12350 1910 12650 1980
rect 12850 1910 13150 1980
rect 13350 1910 13650 1980
rect 13850 1910 14150 1980
rect 14350 1910 14650 1980
rect 14850 1910 15150 1980
rect 15350 1910 15650 1980
rect 15850 1910 16150 1980
rect 16350 1910 16650 1980
rect 16850 1910 17150 1980
rect 17350 1910 17650 1980
rect 17850 1910 18150 1980
rect 18350 1910 18650 1980
rect 18850 1910 19150 1980
rect 19350 1910 19650 1980
rect 19850 1910 20150 1980
rect 20350 1910 20650 1980
rect 20850 1910 21150 1980
rect 21350 1910 21650 1980
rect 21850 1910 22150 1980
rect 22350 1910 22650 1980
rect 22850 1910 23150 1980
rect 23350 1910 23650 1980
rect 23850 1910 24150 1980
rect 24350 1910 24650 1980
rect 24850 1910 25150 1980
rect 25350 1910 25650 1980
rect 25850 1910 26150 1980
rect 26350 1910 26500 1980
rect 0 1900 26500 1910
rect 0 1880 120 1900
rect 380 1880 620 1900
rect 880 1880 1120 1900
rect 1380 1880 1620 1900
rect 1880 1880 2120 1900
rect 2380 1880 2620 1900
rect 2880 1880 3120 1900
rect 3380 1880 3620 1900
rect 3880 1880 4120 1900
rect 4380 1880 4620 1900
rect 4880 1880 5120 1900
rect 5380 1880 5620 1900
rect 5880 1880 6120 1900
rect 6380 1880 6620 1900
rect 6880 1880 7120 1900
rect 7380 1880 7620 1900
rect 7880 1880 8120 1900
rect 8380 1880 8620 1900
rect 8880 1880 9120 1900
rect 9380 1880 9620 1900
rect 9880 1880 10120 1900
rect 10380 1880 10620 1900
rect 10880 1880 11120 1900
rect 11380 1880 11620 1900
rect 11880 1880 12120 1900
rect 12380 1880 12620 1900
rect 12880 1880 13120 1900
rect 13380 1880 13620 1900
rect 13880 1880 14120 1900
rect 14380 1880 14620 1900
rect 14880 1880 15120 1900
rect 15380 1880 15620 1900
rect 15880 1880 16120 1900
rect 16380 1880 16620 1900
rect 16880 1880 17120 1900
rect 17380 1880 17620 1900
rect 17880 1880 18120 1900
rect 18380 1880 18620 1900
rect 18880 1880 19120 1900
rect 19380 1880 19620 1900
rect 19880 1880 20120 1900
rect 20380 1880 20620 1900
rect 20880 1880 21120 1900
rect 21380 1880 21620 1900
rect 21880 1880 22120 1900
rect 22380 1880 22620 1900
rect 22880 1880 23120 1900
rect 23380 1880 23620 1900
rect 23880 1880 24120 1900
rect 24380 1880 24620 1900
rect 24880 1880 25120 1900
rect 25380 1880 25620 1900
rect 25880 1880 26120 1900
rect 26380 1880 26500 1900
rect 0 1850 100 1880
rect 0 1650 20 1850
rect 90 1650 100 1850
rect 0 1620 100 1650
rect 400 1850 600 1880
rect 400 1650 410 1850
rect 480 1650 520 1850
rect 590 1650 600 1850
rect 400 1620 600 1650
rect 900 1850 1100 1880
rect 900 1650 910 1850
rect 980 1650 1020 1850
rect 1090 1650 1100 1850
rect 900 1620 1100 1650
rect 1400 1850 1600 1880
rect 1400 1650 1410 1850
rect 1480 1650 1520 1850
rect 1590 1650 1600 1850
rect 1400 1620 1600 1650
rect 1900 1850 2100 1880
rect 1900 1650 1910 1850
rect 1980 1650 2020 1850
rect 2090 1650 2100 1850
rect 1900 1620 2100 1650
rect 2400 1850 2600 1880
rect 2400 1650 2410 1850
rect 2480 1650 2520 1850
rect 2590 1650 2600 1850
rect 2400 1620 2600 1650
rect 2900 1850 3100 1880
rect 2900 1650 2910 1850
rect 2980 1650 3020 1850
rect 3090 1650 3100 1850
rect 2900 1620 3100 1650
rect 3400 1850 3600 1880
rect 3400 1650 3410 1850
rect 3480 1650 3520 1850
rect 3590 1650 3600 1850
rect 3400 1620 3600 1650
rect 3900 1850 4100 1880
rect 3900 1650 3910 1850
rect 3980 1650 4020 1850
rect 4090 1650 4100 1850
rect 3900 1620 4100 1650
rect 4400 1850 4600 1880
rect 4400 1650 4410 1850
rect 4480 1650 4520 1850
rect 4590 1650 4600 1850
rect 4400 1620 4600 1650
rect 4900 1850 5100 1880
rect 4900 1650 4910 1850
rect 4980 1650 5020 1850
rect 5090 1650 5100 1850
rect 4900 1620 5100 1650
rect 5400 1850 5600 1880
rect 5400 1650 5410 1850
rect 5480 1650 5520 1850
rect 5590 1650 5600 1850
rect 5400 1620 5600 1650
rect 5900 1850 6100 1880
rect 5900 1650 5910 1850
rect 5980 1650 6020 1850
rect 6090 1650 6100 1850
rect 5900 1620 6100 1650
rect 6400 1850 6600 1880
rect 6400 1650 6410 1850
rect 6480 1650 6520 1850
rect 6590 1650 6600 1850
rect 6400 1620 6600 1650
rect 6900 1850 7100 1880
rect 6900 1650 6910 1850
rect 6980 1650 7020 1850
rect 7090 1650 7100 1850
rect 6900 1620 7100 1650
rect 7400 1850 7600 1880
rect 7400 1650 7410 1850
rect 7480 1650 7520 1850
rect 7590 1650 7600 1850
rect 7400 1620 7600 1650
rect 7900 1850 8100 1880
rect 7900 1650 7910 1850
rect 7980 1650 8020 1850
rect 8090 1650 8100 1850
rect 7900 1620 8100 1650
rect 8400 1850 8600 1880
rect 8400 1650 8410 1850
rect 8480 1650 8520 1850
rect 8590 1650 8600 1850
rect 8400 1620 8600 1650
rect 8900 1850 9100 1880
rect 8900 1650 8910 1850
rect 8980 1650 9020 1850
rect 9090 1650 9100 1850
rect 8900 1620 9100 1650
rect 9400 1850 9600 1880
rect 9400 1650 9410 1850
rect 9480 1650 9520 1850
rect 9590 1650 9600 1850
rect 9400 1620 9600 1650
rect 9900 1850 10100 1880
rect 9900 1650 9910 1850
rect 9980 1650 10020 1850
rect 10090 1650 10100 1850
rect 9900 1620 10100 1650
rect 10400 1850 10600 1880
rect 10400 1650 10410 1850
rect 10480 1650 10520 1850
rect 10590 1650 10600 1850
rect 10400 1620 10600 1650
rect 10900 1850 11100 1880
rect 10900 1650 10910 1850
rect 10980 1650 11020 1850
rect 11090 1650 11100 1850
rect 10900 1620 11100 1650
rect 11400 1850 11600 1880
rect 11400 1650 11410 1850
rect 11480 1650 11520 1850
rect 11590 1650 11600 1850
rect 11400 1620 11600 1650
rect 11900 1850 12100 1880
rect 11900 1650 11910 1850
rect 11980 1650 12020 1850
rect 12090 1650 12100 1850
rect 11900 1620 12100 1650
rect 12400 1850 12600 1880
rect 12400 1650 12410 1850
rect 12480 1650 12520 1850
rect 12590 1650 12600 1850
rect 12400 1620 12600 1650
rect 12900 1850 13100 1880
rect 12900 1650 12910 1850
rect 12980 1650 13020 1850
rect 13090 1650 13100 1850
rect 12900 1620 13100 1650
rect 13400 1850 13600 1880
rect 13400 1650 13410 1850
rect 13480 1650 13520 1850
rect 13590 1650 13600 1850
rect 13400 1620 13600 1650
rect 13900 1850 14100 1880
rect 13900 1650 13910 1850
rect 13980 1650 14020 1850
rect 14090 1650 14100 1850
rect 13900 1620 14100 1650
rect 14400 1850 14600 1880
rect 14400 1650 14410 1850
rect 14480 1650 14520 1850
rect 14590 1650 14600 1850
rect 14400 1620 14600 1650
rect 14900 1850 15100 1880
rect 14900 1650 14910 1850
rect 14980 1650 15020 1850
rect 15090 1650 15100 1850
rect 14900 1620 15100 1650
rect 15400 1850 15600 1880
rect 15400 1650 15410 1850
rect 15480 1650 15520 1850
rect 15590 1650 15600 1850
rect 15400 1620 15600 1650
rect 15900 1850 16100 1880
rect 15900 1650 15910 1850
rect 15980 1650 16020 1850
rect 16090 1650 16100 1850
rect 15900 1620 16100 1650
rect 16400 1850 16600 1880
rect 16400 1650 16410 1850
rect 16480 1650 16520 1850
rect 16590 1650 16600 1850
rect 16400 1620 16600 1650
rect 16900 1850 17100 1880
rect 16900 1650 16910 1850
rect 16980 1650 17020 1850
rect 17090 1650 17100 1850
rect 16900 1620 17100 1650
rect 17400 1850 17600 1880
rect 17400 1650 17410 1850
rect 17480 1650 17520 1850
rect 17590 1650 17600 1850
rect 17400 1620 17600 1650
rect 17900 1850 18100 1880
rect 17900 1650 17910 1850
rect 17980 1650 18020 1850
rect 18090 1650 18100 1850
rect 17900 1620 18100 1650
rect 18400 1850 18600 1880
rect 18400 1650 18410 1850
rect 18480 1650 18520 1850
rect 18590 1650 18600 1850
rect 18400 1620 18600 1650
rect 18900 1850 19100 1880
rect 18900 1650 18910 1850
rect 18980 1650 19020 1850
rect 19090 1650 19100 1850
rect 18900 1620 19100 1650
rect 19400 1850 19600 1880
rect 19400 1650 19410 1850
rect 19480 1650 19520 1850
rect 19590 1650 19600 1850
rect 19400 1620 19600 1650
rect 19900 1850 20100 1880
rect 19900 1650 19910 1850
rect 19980 1650 20020 1850
rect 20090 1650 20100 1850
rect 19900 1620 20100 1650
rect 20400 1850 20600 1880
rect 20400 1650 20410 1850
rect 20480 1650 20520 1850
rect 20590 1650 20600 1850
rect 20400 1620 20600 1650
rect 20900 1850 21100 1880
rect 20900 1650 20910 1850
rect 20980 1650 21020 1850
rect 21090 1650 21100 1850
rect 20900 1620 21100 1650
rect 21400 1850 21600 1880
rect 21400 1650 21410 1850
rect 21480 1650 21520 1850
rect 21590 1650 21600 1850
rect 21400 1620 21600 1650
rect 21900 1850 22100 1880
rect 21900 1650 21910 1850
rect 21980 1650 22020 1850
rect 22090 1650 22100 1850
rect 21900 1620 22100 1650
rect 22400 1850 22600 1880
rect 22400 1650 22410 1850
rect 22480 1650 22520 1850
rect 22590 1650 22600 1850
rect 22400 1620 22600 1650
rect 22900 1850 23100 1880
rect 22900 1650 22910 1850
rect 22980 1650 23020 1850
rect 23090 1650 23100 1850
rect 22900 1620 23100 1650
rect 23400 1850 23600 1880
rect 23400 1650 23410 1850
rect 23480 1650 23520 1850
rect 23590 1650 23600 1850
rect 23400 1620 23600 1650
rect 23900 1850 24100 1880
rect 23900 1650 23910 1850
rect 23980 1650 24020 1850
rect 24090 1650 24100 1850
rect 23900 1620 24100 1650
rect 24400 1850 24600 1880
rect 24400 1650 24410 1850
rect 24480 1650 24520 1850
rect 24590 1650 24600 1850
rect 24400 1620 24600 1650
rect 24900 1850 25100 1880
rect 24900 1650 24910 1850
rect 24980 1650 25020 1850
rect 25090 1650 25100 1850
rect 24900 1620 25100 1650
rect 25400 1850 25600 1880
rect 25400 1650 25410 1850
rect 25480 1650 25520 1850
rect 25590 1650 25600 1850
rect 25400 1620 25600 1650
rect 25900 1850 26100 1880
rect 25900 1650 25910 1850
rect 25980 1650 26020 1850
rect 26090 1650 26100 1850
rect 25900 1620 26100 1650
rect 26400 1850 26500 1880
rect 26400 1650 26410 1850
rect 26480 1650 26500 1850
rect 26400 1620 26500 1650
rect 0 1600 120 1620
rect 380 1600 620 1620
rect 880 1600 1120 1620
rect 1380 1600 1620 1620
rect 1880 1600 2120 1620
rect 2380 1600 2620 1620
rect 2880 1600 3120 1620
rect 3380 1600 3620 1620
rect 3880 1600 4120 1620
rect 4380 1600 4620 1620
rect 4880 1600 5120 1620
rect 5380 1600 5620 1620
rect 5880 1600 6120 1620
rect 6380 1600 6620 1620
rect 6880 1600 7120 1620
rect 7380 1600 7620 1620
rect 7880 1600 8120 1620
rect 8380 1600 8620 1620
rect 8880 1600 9120 1620
rect 9380 1600 9620 1620
rect 9880 1600 10120 1620
rect 10380 1600 10620 1620
rect 10880 1600 11120 1620
rect 11380 1600 11620 1620
rect 11880 1600 12120 1620
rect 12380 1600 12620 1620
rect 12880 1600 13120 1620
rect 13380 1600 13620 1620
rect 13880 1600 14120 1620
rect 14380 1600 14620 1620
rect 14880 1600 15120 1620
rect 15380 1600 15620 1620
rect 15880 1600 16120 1620
rect 16380 1600 16620 1620
rect 16880 1600 17120 1620
rect 17380 1600 17620 1620
rect 17880 1600 18120 1620
rect 18380 1600 18620 1620
rect 18880 1600 19120 1620
rect 19380 1600 19620 1620
rect 19880 1600 20120 1620
rect 20380 1600 20620 1620
rect 20880 1600 21120 1620
rect 21380 1600 21620 1620
rect 21880 1600 22120 1620
rect 22380 1600 22620 1620
rect 22880 1600 23120 1620
rect 23380 1600 23620 1620
rect 23880 1600 24120 1620
rect 24380 1600 24620 1620
rect 24880 1600 25120 1620
rect 25380 1600 25620 1620
rect 25880 1600 26120 1620
rect 26380 1600 26500 1620
rect 0 1590 26500 1600
rect 0 1520 150 1590
rect 350 1520 650 1590
rect 850 1520 1150 1590
rect 1350 1520 1650 1590
rect 1850 1520 2150 1590
rect 2350 1520 2650 1590
rect 2850 1520 3150 1590
rect 3350 1520 3650 1590
rect 3850 1520 4150 1590
rect 4350 1520 4650 1590
rect 4850 1520 5150 1590
rect 5350 1520 5650 1590
rect 5850 1520 6150 1590
rect 6350 1520 6650 1590
rect 6850 1520 7150 1590
rect 7350 1520 7650 1590
rect 7850 1520 8150 1590
rect 8350 1520 8650 1590
rect 8850 1520 9150 1590
rect 9350 1520 9650 1590
rect 9850 1520 10150 1590
rect 10350 1520 10650 1590
rect 10850 1520 11150 1590
rect 11350 1520 11650 1590
rect 11850 1520 12150 1590
rect 12350 1520 12650 1590
rect 12850 1520 13150 1590
rect 13350 1520 13650 1590
rect 13850 1520 14150 1590
rect 14350 1520 14650 1590
rect 14850 1520 15150 1590
rect 15350 1520 15650 1590
rect 15850 1520 16150 1590
rect 16350 1520 16650 1590
rect 16850 1520 17150 1590
rect 17350 1520 17650 1590
rect 17850 1520 18150 1590
rect 18350 1520 18650 1590
rect 18850 1520 19150 1590
rect 19350 1520 19650 1590
rect 19850 1520 20150 1590
rect 20350 1520 20650 1590
rect 20850 1520 21150 1590
rect 21350 1520 21650 1590
rect 21850 1520 22150 1590
rect 22350 1520 22650 1590
rect 22850 1520 23150 1590
rect 23350 1520 23650 1590
rect 23850 1520 24150 1590
rect 24350 1520 24650 1590
rect 24850 1520 25150 1590
rect 25350 1520 25650 1590
rect 25850 1520 26150 1590
rect 26350 1520 26500 1590
rect 0 1480 26500 1520
rect 0 1410 150 1480
rect 350 1410 650 1480
rect 850 1410 1150 1480
rect 1350 1410 1650 1480
rect 1850 1410 2150 1480
rect 2350 1410 2650 1480
rect 2850 1410 3150 1480
rect 3350 1410 3650 1480
rect 3850 1410 4150 1480
rect 4350 1410 4650 1480
rect 4850 1410 5150 1480
rect 5350 1410 5650 1480
rect 5850 1410 6150 1480
rect 6350 1410 6650 1480
rect 6850 1410 7150 1480
rect 7350 1410 7650 1480
rect 7850 1410 8150 1480
rect 8350 1410 8650 1480
rect 8850 1410 9150 1480
rect 9350 1410 9650 1480
rect 9850 1410 10150 1480
rect 10350 1410 10650 1480
rect 10850 1410 11150 1480
rect 11350 1410 11650 1480
rect 11850 1410 12150 1480
rect 12350 1410 12650 1480
rect 12850 1410 13150 1480
rect 13350 1410 13650 1480
rect 13850 1410 14150 1480
rect 14350 1410 14650 1480
rect 14850 1410 15150 1480
rect 15350 1410 15650 1480
rect 15850 1410 16150 1480
rect 16350 1410 16650 1480
rect 16850 1410 17150 1480
rect 17350 1410 17650 1480
rect 17850 1410 18150 1480
rect 18350 1410 18650 1480
rect 18850 1410 19150 1480
rect 19350 1410 19650 1480
rect 19850 1410 20150 1480
rect 20350 1410 20650 1480
rect 20850 1410 21150 1480
rect 21350 1410 21650 1480
rect 21850 1410 22150 1480
rect 22350 1410 22650 1480
rect 22850 1410 23150 1480
rect 23350 1410 23650 1480
rect 23850 1410 24150 1480
rect 24350 1410 24650 1480
rect 24850 1410 25150 1480
rect 25350 1410 25650 1480
rect 25850 1410 26150 1480
rect 26350 1410 26500 1480
rect 0 1400 26500 1410
rect 0 1380 120 1400
rect 380 1380 620 1400
rect 880 1380 1120 1400
rect 1380 1380 1620 1400
rect 1880 1380 2120 1400
rect 2380 1380 2620 1400
rect 2880 1380 3120 1400
rect 3380 1380 3620 1400
rect 3880 1380 4120 1400
rect 4380 1380 4620 1400
rect 4880 1380 5120 1400
rect 5380 1380 5620 1400
rect 5880 1380 6120 1400
rect 6380 1380 6620 1400
rect 6880 1380 7120 1400
rect 7380 1380 7620 1400
rect 7880 1380 8120 1400
rect 8380 1380 8620 1400
rect 8880 1380 9120 1400
rect 9380 1380 9620 1400
rect 9880 1380 10120 1400
rect 10380 1380 10620 1400
rect 10880 1380 11120 1400
rect 11380 1380 11620 1400
rect 11880 1380 12120 1400
rect 12380 1380 12620 1400
rect 12880 1380 13120 1400
rect 13380 1380 13620 1400
rect 13880 1380 14120 1400
rect 14380 1380 14620 1400
rect 14880 1380 15120 1400
rect 15380 1380 15620 1400
rect 15880 1380 16120 1400
rect 16380 1380 16620 1400
rect 16880 1380 17120 1400
rect 17380 1380 17620 1400
rect 17880 1380 18120 1400
rect 18380 1380 18620 1400
rect 18880 1380 19120 1400
rect 19380 1380 19620 1400
rect 19880 1380 20120 1400
rect 20380 1380 20620 1400
rect 20880 1380 21120 1400
rect 21380 1380 21620 1400
rect 21880 1380 22120 1400
rect 22380 1380 22620 1400
rect 22880 1380 23120 1400
rect 23380 1380 23620 1400
rect 23880 1380 24120 1400
rect 24380 1380 24620 1400
rect 24880 1380 25120 1400
rect 25380 1380 25620 1400
rect 25880 1380 26120 1400
rect 26380 1380 26500 1400
rect 0 1350 100 1380
rect 0 1150 20 1350
rect 90 1150 100 1350
rect 0 1120 100 1150
rect 400 1350 600 1380
rect 400 1150 410 1350
rect 480 1150 520 1350
rect 590 1150 600 1350
rect 400 1120 600 1150
rect 900 1350 1100 1380
rect 900 1150 910 1350
rect 980 1150 1020 1350
rect 1090 1150 1100 1350
rect 900 1120 1100 1150
rect 1400 1350 1600 1380
rect 1400 1150 1410 1350
rect 1480 1150 1520 1350
rect 1590 1150 1600 1350
rect 1400 1120 1600 1150
rect 1900 1350 2100 1380
rect 1900 1150 1910 1350
rect 1980 1150 2020 1350
rect 2090 1150 2100 1350
rect 1900 1120 2100 1150
rect 2400 1350 2600 1380
rect 2400 1150 2410 1350
rect 2480 1150 2520 1350
rect 2590 1150 2600 1350
rect 2400 1120 2600 1150
rect 2900 1350 3100 1380
rect 2900 1150 2910 1350
rect 2980 1150 3020 1350
rect 3090 1150 3100 1350
rect 2900 1120 3100 1150
rect 3400 1350 3600 1380
rect 3400 1150 3410 1350
rect 3480 1150 3520 1350
rect 3590 1150 3600 1350
rect 3400 1120 3600 1150
rect 3900 1350 4100 1380
rect 3900 1150 3910 1350
rect 3980 1150 4020 1350
rect 4090 1150 4100 1350
rect 3900 1120 4100 1150
rect 4400 1350 4600 1380
rect 4400 1150 4410 1350
rect 4480 1150 4520 1350
rect 4590 1150 4600 1350
rect 4400 1120 4600 1150
rect 4900 1350 5100 1380
rect 4900 1150 4910 1350
rect 4980 1150 5020 1350
rect 5090 1150 5100 1350
rect 4900 1120 5100 1150
rect 5400 1350 5600 1380
rect 5400 1150 5410 1350
rect 5480 1150 5520 1350
rect 5590 1150 5600 1350
rect 5400 1120 5600 1150
rect 5900 1350 6100 1380
rect 5900 1150 5910 1350
rect 5980 1150 6020 1350
rect 6090 1150 6100 1350
rect 5900 1120 6100 1150
rect 6400 1350 6600 1380
rect 6400 1150 6410 1350
rect 6480 1150 6520 1350
rect 6590 1150 6600 1350
rect 6400 1120 6600 1150
rect 6900 1350 7100 1380
rect 6900 1150 6910 1350
rect 6980 1150 7020 1350
rect 7090 1150 7100 1350
rect 6900 1120 7100 1150
rect 7400 1350 7600 1380
rect 7400 1150 7410 1350
rect 7480 1150 7520 1350
rect 7590 1150 7600 1350
rect 7400 1120 7600 1150
rect 7900 1350 8100 1380
rect 7900 1150 7910 1350
rect 7980 1150 8020 1350
rect 8090 1150 8100 1350
rect 7900 1120 8100 1150
rect 8400 1350 8600 1380
rect 8400 1150 8410 1350
rect 8480 1150 8520 1350
rect 8590 1150 8600 1350
rect 8400 1120 8600 1150
rect 8900 1350 9100 1380
rect 8900 1150 8910 1350
rect 8980 1150 9020 1350
rect 9090 1150 9100 1350
rect 8900 1120 9100 1150
rect 9400 1350 9600 1380
rect 9400 1150 9410 1350
rect 9480 1150 9520 1350
rect 9590 1150 9600 1350
rect 9400 1120 9600 1150
rect 9900 1350 10100 1380
rect 9900 1150 9910 1350
rect 9980 1150 10020 1350
rect 10090 1150 10100 1350
rect 9900 1120 10100 1150
rect 10400 1350 10600 1380
rect 10400 1150 10410 1350
rect 10480 1150 10520 1350
rect 10590 1150 10600 1350
rect 10400 1120 10600 1150
rect 10900 1350 11100 1380
rect 10900 1150 10910 1350
rect 10980 1150 11020 1350
rect 11090 1150 11100 1350
rect 10900 1120 11100 1150
rect 11400 1350 11600 1380
rect 11400 1150 11410 1350
rect 11480 1150 11520 1350
rect 11590 1150 11600 1350
rect 11400 1120 11600 1150
rect 11900 1350 12100 1380
rect 11900 1150 11910 1350
rect 11980 1150 12020 1350
rect 12090 1150 12100 1350
rect 11900 1120 12100 1150
rect 12400 1350 12600 1380
rect 12400 1150 12410 1350
rect 12480 1150 12520 1350
rect 12590 1150 12600 1350
rect 12400 1120 12600 1150
rect 12900 1350 13100 1380
rect 12900 1150 12910 1350
rect 12980 1150 13020 1350
rect 13090 1150 13100 1350
rect 12900 1120 13100 1150
rect 13400 1350 13600 1380
rect 13400 1150 13410 1350
rect 13480 1150 13520 1350
rect 13590 1150 13600 1350
rect 13400 1120 13600 1150
rect 13900 1350 14100 1380
rect 13900 1150 13910 1350
rect 13980 1150 14020 1350
rect 14090 1150 14100 1350
rect 13900 1120 14100 1150
rect 14400 1350 14600 1380
rect 14400 1150 14410 1350
rect 14480 1150 14520 1350
rect 14590 1150 14600 1350
rect 14400 1120 14600 1150
rect 14900 1350 15100 1380
rect 14900 1150 14910 1350
rect 14980 1150 15020 1350
rect 15090 1150 15100 1350
rect 14900 1120 15100 1150
rect 15400 1350 15600 1380
rect 15400 1150 15410 1350
rect 15480 1150 15520 1350
rect 15590 1150 15600 1350
rect 15400 1120 15600 1150
rect 15900 1350 16100 1380
rect 15900 1150 15910 1350
rect 15980 1150 16020 1350
rect 16090 1150 16100 1350
rect 15900 1120 16100 1150
rect 16400 1350 16600 1380
rect 16400 1150 16410 1350
rect 16480 1150 16520 1350
rect 16590 1150 16600 1350
rect 16400 1120 16600 1150
rect 16900 1350 17100 1380
rect 16900 1150 16910 1350
rect 16980 1150 17020 1350
rect 17090 1150 17100 1350
rect 16900 1120 17100 1150
rect 17400 1350 17600 1380
rect 17400 1150 17410 1350
rect 17480 1150 17520 1350
rect 17590 1150 17600 1350
rect 17400 1120 17600 1150
rect 17900 1350 18100 1380
rect 17900 1150 17910 1350
rect 17980 1150 18020 1350
rect 18090 1150 18100 1350
rect 17900 1120 18100 1150
rect 18400 1350 18600 1380
rect 18400 1150 18410 1350
rect 18480 1150 18520 1350
rect 18590 1150 18600 1350
rect 18400 1120 18600 1150
rect 18900 1350 19100 1380
rect 18900 1150 18910 1350
rect 18980 1150 19020 1350
rect 19090 1150 19100 1350
rect 18900 1120 19100 1150
rect 19400 1350 19600 1380
rect 19400 1150 19410 1350
rect 19480 1150 19520 1350
rect 19590 1150 19600 1350
rect 19400 1120 19600 1150
rect 19900 1350 20100 1380
rect 19900 1150 19910 1350
rect 19980 1150 20020 1350
rect 20090 1150 20100 1350
rect 19900 1120 20100 1150
rect 20400 1350 20600 1380
rect 20400 1150 20410 1350
rect 20480 1150 20520 1350
rect 20590 1150 20600 1350
rect 20400 1120 20600 1150
rect 20900 1350 21100 1380
rect 20900 1150 20910 1350
rect 20980 1150 21020 1350
rect 21090 1150 21100 1350
rect 20900 1120 21100 1150
rect 21400 1350 21600 1380
rect 21400 1150 21410 1350
rect 21480 1150 21520 1350
rect 21590 1150 21600 1350
rect 21400 1120 21600 1150
rect 21900 1350 22100 1380
rect 21900 1150 21910 1350
rect 21980 1150 22020 1350
rect 22090 1150 22100 1350
rect 21900 1120 22100 1150
rect 22400 1350 22600 1380
rect 22400 1150 22410 1350
rect 22480 1150 22520 1350
rect 22590 1150 22600 1350
rect 22400 1120 22600 1150
rect 22900 1350 23100 1380
rect 22900 1150 22910 1350
rect 22980 1150 23020 1350
rect 23090 1150 23100 1350
rect 22900 1120 23100 1150
rect 23400 1350 23600 1380
rect 23400 1150 23410 1350
rect 23480 1150 23520 1350
rect 23590 1150 23600 1350
rect 23400 1120 23600 1150
rect 23900 1350 24100 1380
rect 23900 1150 23910 1350
rect 23980 1150 24020 1350
rect 24090 1150 24100 1350
rect 23900 1120 24100 1150
rect 24400 1350 24600 1380
rect 24400 1150 24410 1350
rect 24480 1150 24520 1350
rect 24590 1150 24600 1350
rect 24400 1120 24600 1150
rect 24900 1350 25100 1380
rect 24900 1150 24910 1350
rect 24980 1150 25020 1350
rect 25090 1150 25100 1350
rect 24900 1120 25100 1150
rect 25400 1350 25600 1380
rect 25400 1150 25410 1350
rect 25480 1150 25520 1350
rect 25590 1150 25600 1350
rect 25400 1120 25600 1150
rect 25900 1350 26100 1380
rect 25900 1150 25910 1350
rect 25980 1150 26020 1350
rect 26090 1150 26100 1350
rect 25900 1120 26100 1150
rect 26400 1350 26500 1380
rect 26400 1150 26410 1350
rect 26480 1150 26500 1350
rect 26400 1120 26500 1150
rect 0 1100 120 1120
rect 380 1100 620 1120
rect 880 1100 1120 1120
rect 1380 1100 1620 1120
rect 1880 1100 2120 1120
rect 2380 1100 2620 1120
rect 2880 1100 3120 1120
rect 3380 1100 3620 1120
rect 3880 1100 4120 1120
rect 4380 1100 4620 1120
rect 4880 1100 5120 1120
rect 5380 1100 5620 1120
rect 5880 1100 6120 1120
rect 6380 1100 6620 1120
rect 6880 1100 7120 1120
rect 7380 1100 7620 1120
rect 7880 1100 8120 1120
rect 8380 1100 8620 1120
rect 8880 1100 9120 1120
rect 9380 1100 9620 1120
rect 9880 1100 10120 1120
rect 10380 1100 10620 1120
rect 10880 1100 11120 1120
rect 11380 1100 11620 1120
rect 11880 1100 12120 1120
rect 12380 1100 12620 1120
rect 12880 1100 13120 1120
rect 13380 1100 13620 1120
rect 13880 1100 14120 1120
rect 14380 1100 14620 1120
rect 14880 1100 15120 1120
rect 15380 1100 15620 1120
rect 15880 1100 16120 1120
rect 16380 1100 16620 1120
rect 16880 1100 17120 1120
rect 17380 1100 17620 1120
rect 17880 1100 18120 1120
rect 18380 1100 18620 1120
rect 18880 1100 19120 1120
rect 19380 1100 19620 1120
rect 19880 1100 20120 1120
rect 20380 1100 20620 1120
rect 20880 1100 21120 1120
rect 21380 1100 21620 1120
rect 21880 1100 22120 1120
rect 22380 1100 22620 1120
rect 22880 1100 23120 1120
rect 23380 1100 23620 1120
rect 23880 1100 24120 1120
rect 24380 1100 24620 1120
rect 24880 1100 25120 1120
rect 25380 1100 25620 1120
rect 25880 1100 26120 1120
rect 26380 1100 26500 1120
rect 0 1090 26500 1100
rect 0 1020 150 1090
rect 350 1020 650 1090
rect 850 1020 1150 1090
rect 1350 1020 1650 1090
rect 1850 1020 2150 1090
rect 2350 1020 2650 1090
rect 2850 1020 3150 1090
rect 3350 1020 3650 1090
rect 3850 1020 4150 1090
rect 4350 1020 4650 1090
rect 4850 1020 5150 1090
rect 5350 1020 5650 1090
rect 5850 1020 6150 1090
rect 6350 1020 6650 1090
rect 6850 1020 7150 1090
rect 7350 1020 7650 1090
rect 7850 1020 8150 1090
rect 8350 1020 8650 1090
rect 8850 1020 9150 1090
rect 9350 1020 9650 1090
rect 9850 1020 10150 1090
rect 10350 1020 10650 1090
rect 10850 1020 11150 1090
rect 11350 1020 11650 1090
rect 11850 1020 12150 1090
rect 12350 1020 12650 1090
rect 12850 1020 13150 1090
rect 13350 1020 13650 1090
rect 13850 1020 14150 1090
rect 14350 1020 14650 1090
rect 14850 1020 15150 1090
rect 15350 1020 15650 1090
rect 15850 1020 16150 1090
rect 16350 1020 16650 1090
rect 16850 1020 17150 1090
rect 17350 1020 17650 1090
rect 17850 1020 18150 1090
rect 18350 1020 18650 1090
rect 18850 1020 19150 1090
rect 19350 1020 19650 1090
rect 19850 1020 20150 1090
rect 20350 1020 20650 1090
rect 20850 1020 21150 1090
rect 21350 1020 21650 1090
rect 21850 1020 22150 1090
rect 22350 1020 22650 1090
rect 22850 1020 23150 1090
rect 23350 1020 23650 1090
rect 23850 1020 24150 1090
rect 24350 1020 24650 1090
rect 24850 1020 25150 1090
rect 25350 1020 25650 1090
rect 25850 1020 26150 1090
rect 26350 1020 26500 1090
rect 0 1000 26500 1020
<< via1 >>
rect 150 47410 350 47480
rect 650 47410 850 47480
rect 1150 47410 1350 47480
rect 1650 47410 1850 47480
rect 2150 47410 2350 47480
rect 2650 47410 2850 47480
rect 3150 47410 3350 47480
rect 3650 47410 3850 47480
rect 4150 47410 4350 47480
rect 4650 47410 4850 47480
rect 5150 47410 5350 47480
rect 5650 47410 5850 47480
rect 6150 47410 6350 47480
rect 6650 47410 6850 47480
rect 7150 47410 7350 47480
rect 7650 47410 7850 47480
rect 8150 47410 8350 47480
rect 8650 47410 8850 47480
rect 9150 47410 9350 47480
rect 9650 47410 9850 47480
rect 10150 47410 10350 47480
rect 10650 47410 10850 47480
rect 11150 47410 11350 47480
rect 11650 47410 11850 47480
rect 12150 47410 12350 47480
rect 12650 47410 12850 47480
rect 13150 47410 13350 47480
rect 13650 47410 13850 47480
rect 14150 47410 14350 47480
rect 14650 47410 14850 47480
rect 15150 47410 15350 47480
rect 15650 47410 15850 47480
rect 16150 47410 16350 47480
rect 16650 47410 16850 47480
rect 17150 47410 17350 47480
rect 17650 47410 17850 47480
rect 18150 47410 18350 47480
rect 18650 47410 18850 47480
rect 19150 47410 19350 47480
rect 19650 47410 19850 47480
rect 20150 47410 20350 47480
rect 20650 47410 20850 47480
rect 21150 47410 21350 47480
rect 21650 47410 21850 47480
rect 22150 47410 22350 47480
rect 22650 47410 22850 47480
rect 23150 47410 23350 47480
rect 23650 47410 23850 47480
rect 24150 47410 24350 47480
rect 24650 47410 24850 47480
rect 25150 47410 25350 47480
rect 25650 47410 25850 47480
rect 26150 47410 26350 47480
rect 20 47150 90 47350
rect 410 47150 480 47350
rect 520 47150 590 47350
rect 910 47150 980 47350
rect 1020 47150 1090 47350
rect 1410 47150 1480 47350
rect 1520 47150 1590 47350
rect 1910 47150 1980 47350
rect 2020 47150 2090 47350
rect 2410 47150 2480 47350
rect 2520 47150 2590 47350
rect 2910 47150 2980 47350
rect 3020 47150 3090 47350
rect 3410 47150 3480 47350
rect 3520 47150 3590 47350
rect 3910 47150 3980 47350
rect 4020 47150 4090 47350
rect 4410 47150 4480 47350
rect 4520 47150 4590 47350
rect 4910 47150 4980 47350
rect 5020 47150 5090 47350
rect 5410 47150 5480 47350
rect 5520 47150 5590 47350
rect 5910 47150 5980 47350
rect 6020 47150 6090 47350
rect 6410 47150 6480 47350
rect 6520 47150 6590 47350
rect 6910 47150 6980 47350
rect 7020 47150 7090 47350
rect 7410 47150 7480 47350
rect 7520 47150 7590 47350
rect 7910 47150 7980 47350
rect 8020 47150 8090 47350
rect 8410 47150 8480 47350
rect 8520 47150 8590 47350
rect 8910 47150 8980 47350
rect 9020 47150 9090 47350
rect 9410 47150 9480 47350
rect 9520 47150 9590 47350
rect 9910 47150 9980 47350
rect 10020 47150 10090 47350
rect 10410 47150 10480 47350
rect 10520 47150 10590 47350
rect 10910 47150 10980 47350
rect 11020 47150 11090 47350
rect 11410 47150 11480 47350
rect 11520 47150 11590 47350
rect 11910 47150 11980 47350
rect 12020 47150 12090 47350
rect 12410 47150 12480 47350
rect 12520 47150 12590 47350
rect 12910 47150 12980 47350
rect 13020 47150 13090 47350
rect 13410 47150 13480 47350
rect 13520 47150 13590 47350
rect 13910 47150 13980 47350
rect 14020 47150 14090 47350
rect 14410 47150 14480 47350
rect 14520 47150 14590 47350
rect 14910 47150 14980 47350
rect 15020 47150 15090 47350
rect 15410 47150 15480 47350
rect 15520 47150 15590 47350
rect 15910 47150 15980 47350
rect 16020 47150 16090 47350
rect 16410 47150 16480 47350
rect 16520 47150 16590 47350
rect 16910 47150 16980 47350
rect 17020 47150 17090 47350
rect 17410 47150 17480 47350
rect 17520 47150 17590 47350
rect 17910 47150 17980 47350
rect 18020 47150 18090 47350
rect 18410 47150 18480 47350
rect 18520 47150 18590 47350
rect 18910 47150 18980 47350
rect 19020 47150 19090 47350
rect 19410 47150 19480 47350
rect 19520 47150 19590 47350
rect 19910 47150 19980 47350
rect 20020 47150 20090 47350
rect 20410 47150 20480 47350
rect 20520 47150 20590 47350
rect 20910 47150 20980 47350
rect 21020 47150 21090 47350
rect 21410 47150 21480 47350
rect 21520 47150 21590 47350
rect 21910 47150 21980 47350
rect 22020 47150 22090 47350
rect 22410 47150 22480 47350
rect 22520 47150 22590 47350
rect 22910 47150 22980 47350
rect 23020 47150 23090 47350
rect 23410 47150 23480 47350
rect 23520 47150 23590 47350
rect 23910 47150 23980 47350
rect 24020 47150 24090 47350
rect 24410 47150 24480 47350
rect 24520 47150 24590 47350
rect 24910 47150 24980 47350
rect 25020 47150 25090 47350
rect 25410 47150 25480 47350
rect 25520 47150 25590 47350
rect 25910 47150 25980 47350
rect 26020 47150 26090 47350
rect 26410 47150 26480 47350
rect 150 47020 350 47090
rect 650 47020 850 47090
rect 1150 47020 1350 47090
rect 1650 47020 1850 47090
rect 2150 47020 2350 47090
rect 2650 47020 2850 47090
rect 3150 47020 3350 47090
rect 3650 47020 3850 47090
rect 4150 47020 4350 47090
rect 4650 47020 4850 47090
rect 5150 47020 5350 47090
rect 5650 47020 5850 47090
rect 6150 47020 6350 47090
rect 6650 47020 6850 47090
rect 7150 47020 7350 47090
rect 7650 47020 7850 47090
rect 8150 47020 8350 47090
rect 8650 47020 8850 47090
rect 9150 47020 9350 47090
rect 9650 47020 9850 47090
rect 10150 47020 10350 47090
rect 10650 47020 10850 47090
rect 11150 47020 11350 47090
rect 11650 47020 11850 47090
rect 12150 47020 12350 47090
rect 12650 47020 12850 47090
rect 13150 47020 13350 47090
rect 13650 47020 13850 47090
rect 14150 47020 14350 47090
rect 14650 47020 14850 47090
rect 15150 47020 15350 47090
rect 15650 47020 15850 47090
rect 16150 47020 16350 47090
rect 16650 47020 16850 47090
rect 17150 47020 17350 47090
rect 17650 47020 17850 47090
rect 18150 47020 18350 47090
rect 18650 47020 18850 47090
rect 19150 47020 19350 47090
rect 19650 47020 19850 47090
rect 20150 47020 20350 47090
rect 20650 47020 20850 47090
rect 21150 47020 21350 47090
rect 21650 47020 21850 47090
rect 22150 47020 22350 47090
rect 22650 47020 22850 47090
rect 23150 47020 23350 47090
rect 23650 47020 23850 47090
rect 24150 47020 24350 47090
rect 24650 47020 24850 47090
rect 25150 47020 25350 47090
rect 25650 47020 25850 47090
rect 26150 47020 26350 47090
rect 150 46910 350 46980
rect 650 46910 850 46980
rect 1150 46910 1350 46980
rect 1650 46910 1850 46980
rect 2150 46910 2350 46980
rect 2650 46910 2850 46980
rect 3150 46910 3350 46980
rect 3650 46910 3850 46980
rect 4150 46910 4350 46980
rect 4650 46910 4850 46980
rect 5150 46910 5350 46980
rect 5650 46910 5850 46980
rect 6150 46910 6350 46980
rect 6650 46910 6850 46980
rect 7150 46910 7350 46980
rect 7650 46910 7850 46980
rect 8150 46910 8350 46980
rect 8650 46910 8850 46980
rect 9150 46910 9350 46980
rect 9650 46910 9850 46980
rect 10150 46910 10350 46980
rect 10650 46910 10850 46980
rect 11150 46910 11350 46980
rect 11650 46910 11850 46980
rect 12150 46910 12350 46980
rect 12650 46910 12850 46980
rect 13150 46910 13350 46980
rect 13650 46910 13850 46980
rect 14150 46910 14350 46980
rect 14650 46910 14850 46980
rect 15150 46910 15350 46980
rect 15650 46910 15850 46980
rect 16150 46910 16350 46980
rect 16650 46910 16850 46980
rect 17150 46910 17350 46980
rect 17650 46910 17850 46980
rect 18150 46910 18350 46980
rect 18650 46910 18850 46980
rect 19150 46910 19350 46980
rect 19650 46910 19850 46980
rect 20150 46910 20350 46980
rect 20650 46910 20850 46980
rect 21150 46910 21350 46980
rect 21650 46910 21850 46980
rect 22150 46910 22350 46980
rect 22650 46910 22850 46980
rect 23150 46910 23350 46980
rect 23650 46910 23850 46980
rect 24150 46910 24350 46980
rect 24650 46910 24850 46980
rect 25150 46910 25350 46980
rect 25650 46910 25850 46980
rect 26150 46910 26350 46980
rect 20 46650 90 46850
rect 410 46650 480 46850
rect 520 46650 590 46850
rect 910 46650 980 46850
rect 1020 46650 1090 46850
rect 1410 46650 1480 46850
rect 1520 46650 1590 46850
rect 1910 46650 1980 46850
rect 2020 46650 2090 46850
rect 2410 46650 2480 46850
rect 2520 46650 2590 46850
rect 2910 46650 2980 46850
rect 3020 46650 3090 46850
rect 3410 46650 3480 46850
rect 3520 46650 3590 46850
rect 3910 46650 3980 46850
rect 4020 46650 4090 46850
rect 4410 46650 4480 46850
rect 4520 46650 4590 46850
rect 4910 46650 4980 46850
rect 5020 46650 5090 46850
rect 5410 46650 5480 46850
rect 5520 46650 5590 46850
rect 5910 46650 5980 46850
rect 6020 46650 6090 46850
rect 6410 46650 6480 46850
rect 6520 46650 6590 46850
rect 6910 46650 6980 46850
rect 7020 46650 7090 46850
rect 7410 46650 7480 46850
rect 7520 46650 7590 46850
rect 7910 46650 7980 46850
rect 8020 46650 8090 46850
rect 8410 46650 8480 46850
rect 8520 46650 8590 46850
rect 8910 46650 8980 46850
rect 9020 46650 9090 46850
rect 9410 46650 9480 46850
rect 9520 46650 9590 46850
rect 9910 46650 9980 46850
rect 10020 46650 10090 46850
rect 10410 46650 10480 46850
rect 10520 46650 10590 46850
rect 10910 46650 10980 46850
rect 11020 46650 11090 46850
rect 11410 46650 11480 46850
rect 11520 46650 11590 46850
rect 11910 46650 11980 46850
rect 12020 46650 12090 46850
rect 12410 46650 12480 46850
rect 12520 46650 12590 46850
rect 12910 46650 12980 46850
rect 13020 46650 13090 46850
rect 13410 46650 13480 46850
rect 13520 46650 13590 46850
rect 13910 46650 13980 46850
rect 14020 46650 14090 46850
rect 14410 46650 14480 46850
rect 14520 46650 14590 46850
rect 14910 46650 14980 46850
rect 15020 46650 15090 46850
rect 15410 46650 15480 46850
rect 15520 46650 15590 46850
rect 15910 46650 15980 46850
rect 16020 46650 16090 46850
rect 16410 46650 16480 46850
rect 16520 46650 16590 46850
rect 16910 46650 16980 46850
rect 17020 46650 17090 46850
rect 17410 46650 17480 46850
rect 17520 46650 17590 46850
rect 17910 46650 17980 46850
rect 18020 46650 18090 46850
rect 18410 46650 18480 46850
rect 18520 46650 18590 46850
rect 18910 46650 18980 46850
rect 19020 46650 19090 46850
rect 19410 46650 19480 46850
rect 19520 46650 19590 46850
rect 19910 46650 19980 46850
rect 20020 46650 20090 46850
rect 20410 46650 20480 46850
rect 20520 46650 20590 46850
rect 20910 46650 20980 46850
rect 21020 46650 21090 46850
rect 21410 46650 21480 46850
rect 21520 46650 21590 46850
rect 21910 46650 21980 46850
rect 22020 46650 22090 46850
rect 22410 46650 22480 46850
rect 22520 46650 22590 46850
rect 22910 46650 22980 46850
rect 23020 46650 23090 46850
rect 23410 46650 23480 46850
rect 23520 46650 23590 46850
rect 23910 46650 23980 46850
rect 24020 46650 24090 46850
rect 24410 46650 24480 46850
rect 24520 46650 24590 46850
rect 24910 46650 24980 46850
rect 25020 46650 25090 46850
rect 25410 46650 25480 46850
rect 25520 46650 25590 46850
rect 25910 46650 25980 46850
rect 26020 46650 26090 46850
rect 26410 46650 26480 46850
rect 150 46520 350 46590
rect 650 46520 850 46590
rect 1150 46520 1350 46590
rect 1650 46520 1850 46590
rect 2150 46520 2350 46590
rect 2650 46520 2850 46590
rect 3150 46520 3350 46590
rect 3650 46520 3850 46590
rect 4150 46520 4350 46590
rect 4650 46520 4850 46590
rect 5150 46520 5350 46590
rect 5650 46520 5850 46590
rect 6150 46520 6350 46590
rect 6650 46520 6850 46590
rect 7150 46520 7350 46590
rect 7650 46520 7850 46590
rect 8150 46520 8350 46590
rect 8650 46520 8850 46590
rect 9150 46520 9350 46590
rect 9650 46520 9850 46590
rect 10150 46520 10350 46590
rect 10650 46520 10850 46590
rect 11150 46520 11350 46590
rect 11650 46520 11850 46590
rect 12150 46520 12350 46590
rect 12650 46520 12850 46590
rect 13150 46520 13350 46590
rect 13650 46520 13850 46590
rect 14150 46520 14350 46590
rect 14650 46520 14850 46590
rect 15150 46520 15350 46590
rect 15650 46520 15850 46590
rect 16150 46520 16350 46590
rect 16650 46520 16850 46590
rect 17150 46520 17350 46590
rect 17650 46520 17850 46590
rect 18150 46520 18350 46590
rect 18650 46520 18850 46590
rect 19150 46520 19350 46590
rect 19650 46520 19850 46590
rect 20150 46520 20350 46590
rect 20650 46520 20850 46590
rect 21150 46520 21350 46590
rect 21650 46520 21850 46590
rect 22150 46520 22350 46590
rect 22650 46520 22850 46590
rect 23150 46520 23350 46590
rect 23650 46520 23850 46590
rect 24150 46520 24350 46590
rect 24650 46520 24850 46590
rect 25150 46520 25350 46590
rect 25650 46520 25850 46590
rect 26150 46520 26350 46590
rect 150 46410 350 46480
rect 650 46410 850 46480
rect 20 46150 90 46350
rect 410 46150 480 46350
rect 520 46150 590 46350
rect 910 46150 980 46350
rect 6650 46410 6850 46480
rect 7150 46410 7350 46480
rect 150 46020 350 46090
rect 650 46020 850 46090
rect 1330 45980 1400 46120
rect 1552 46030 6186 46090
rect 1552 45996 1612 46030
rect 1612 45996 1702 46030
rect 1702 45996 1770 46030
rect 1770 45996 1860 46030
rect 1860 45996 1928 46030
rect 1928 45996 2018 46030
rect 2018 45996 2086 46030
rect 2086 45996 2176 46030
rect 2176 45996 2244 46030
rect 2244 45996 2334 46030
rect 2334 45996 2402 46030
rect 2402 45996 2492 46030
rect 2492 45996 2560 46030
rect 2560 45996 2650 46030
rect 2650 45996 2718 46030
rect 2718 45996 2808 46030
rect 2808 45996 2876 46030
rect 2876 45996 2966 46030
rect 2966 45996 3034 46030
rect 3034 45996 3124 46030
rect 3124 45996 3192 46030
rect 3192 45996 3282 46030
rect 3282 45996 3350 46030
rect 3350 45996 3440 46030
rect 3440 45996 3508 46030
rect 3508 45996 3598 46030
rect 3598 45996 3666 46030
rect 3666 45996 3756 46030
rect 3756 45996 3824 46030
rect 3824 45996 3914 46030
rect 3914 45996 3982 46030
rect 3982 45996 4072 46030
rect 4072 45996 4140 46030
rect 4140 45996 4230 46030
rect 4230 45996 4298 46030
rect 4298 45996 4388 46030
rect 4388 45996 4456 46030
rect 4456 45996 4546 46030
rect 4546 45996 4614 46030
rect 4614 45996 4704 46030
rect 4704 45996 4772 46030
rect 4772 45996 4862 46030
rect 4862 45996 4930 46030
rect 4930 45996 5020 46030
rect 5020 45996 5088 46030
rect 5088 45996 5178 46030
rect 5178 45996 5246 46030
rect 5246 45996 5336 46030
rect 5336 45996 5404 46030
rect 5404 45996 5494 46030
rect 5494 45996 5562 46030
rect 5562 45996 5652 46030
rect 5652 45996 5720 46030
rect 5720 45996 5810 46030
rect 5810 45996 5878 46030
rect 5878 45996 5968 46030
rect 5968 45996 6036 46030
rect 6036 45996 6126 46030
rect 6126 45996 6186 46030
rect 1552 45990 6186 45996
rect 150 45910 350 45980
rect 650 45910 850 45980
rect 20 45650 90 45850
rect 410 45650 480 45850
rect 520 45650 590 45850
rect 910 45650 980 45850
rect 150 45520 350 45590
rect 650 45520 850 45590
rect 150 45410 350 45480
rect 650 45410 850 45480
rect 20 45150 90 45350
rect 410 45150 480 45350
rect 520 45150 590 45350
rect 910 45150 980 45350
rect 150 45020 350 45090
rect 650 45020 850 45090
rect 150 44910 350 44980
rect 650 44910 850 44980
rect 20 44650 90 44850
rect 410 44650 480 44850
rect 520 44650 590 44850
rect 910 44650 980 44850
rect 150 44520 350 44590
rect 650 44520 850 44590
rect 150 44410 350 44480
rect 650 44410 850 44480
rect 20 44150 90 44350
rect 410 44150 480 44350
rect 520 44150 590 44350
rect 910 44150 980 44350
rect 150 44020 350 44090
rect 650 44020 850 44090
rect 150 43910 350 43980
rect 650 43910 850 43980
rect 20 43650 90 43850
rect 410 43650 480 43850
rect 520 43650 590 43850
rect 910 43650 980 43850
rect 150 43520 350 43590
rect 650 43520 850 43590
rect 150 43410 350 43480
rect 650 43410 850 43480
rect 20 43150 90 43350
rect 410 43150 480 43350
rect 520 43150 590 43350
rect 910 43150 980 43350
rect 150 43020 350 43090
rect 650 43020 850 43090
rect 150 42910 350 42980
rect 650 42910 850 42980
rect 20 42650 90 42850
rect 410 42650 480 42850
rect 520 42650 590 42850
rect 910 42650 980 42850
rect 150 42520 350 42590
rect 650 42520 850 42590
rect 150 42410 350 42480
rect 650 42410 850 42480
rect 20 42150 90 42350
rect 410 42150 480 42350
rect 520 42150 590 42350
rect 910 42150 980 42350
rect 150 42020 350 42090
rect 650 42020 850 42090
rect 150 41910 350 41980
rect 650 41910 850 41980
rect 20 41650 90 41850
rect 410 41650 480 41850
rect 520 41650 590 41850
rect 910 41650 980 41850
rect 150 41520 350 41590
rect 650 41520 850 41590
rect 150 41410 350 41480
rect 650 41410 850 41480
rect 20 41150 90 41350
rect 410 41150 480 41350
rect 520 41150 590 41350
rect 910 41150 980 41350
rect 150 41020 350 41090
rect 650 41020 850 41090
rect 150 40910 350 40980
rect 650 40910 850 40980
rect 20 40650 90 40850
rect 410 40650 480 40850
rect 520 40650 590 40850
rect 910 40650 980 40850
rect 150 40520 350 40590
rect 650 40520 850 40590
rect -3290 40276 -3110 40450
rect -3290 40236 -3218 40276
rect -3218 40236 -3184 40276
rect -3184 40236 -3110 40276
rect -3290 40190 -3110 40236
rect -3290 38902 -3110 38910
rect -3290 38862 -3218 38902
rect -3218 38862 -3184 38902
rect -3184 38862 -3110 38902
rect -3290 38690 -3110 38862
rect 150 40410 350 40480
rect 650 40410 850 40480
rect 20 40150 90 40350
rect 410 40150 480 40350
rect 520 40150 590 40350
rect 910 40150 980 40350
rect 150 40020 350 40090
rect 650 40020 850 40090
rect -2850 39910 -2650 39980
rect -2350 39910 -2150 39980
rect -1850 39910 -1650 39980
rect -1350 39910 -1150 39980
rect -850 39910 -650 39980
rect -350 39910 -150 39980
rect 150 39910 350 39980
rect 650 39910 850 39980
rect 1330 39936 1346 45980
rect 1346 39936 1384 45980
rect 1384 39936 1400 45980
rect 6340 45980 6410 46120
rect 6520 46150 6590 46350
rect 6910 46150 6980 46350
rect 7020 46150 7090 46350
rect 7410 46150 7480 46350
rect 13150 46410 13350 46480
rect 13650 46410 13850 46480
rect 6650 46020 6850 46090
rect 7150 46020 7350 46090
rect 1465 39978 1482 45938
rect 1482 39978 1516 45938
rect 1516 39978 1531 45938
rect 1623 39978 1640 45938
rect 1640 39978 1674 45938
rect 1674 39978 1689 45938
rect 1781 39978 1798 45938
rect 1798 39978 1832 45938
rect 1832 39978 1847 45938
rect 1939 39978 1956 45938
rect 1956 39978 1990 45938
rect 1990 39978 2005 45938
rect 2097 39978 2114 45938
rect 2114 39978 2148 45938
rect 2148 39978 2163 45938
rect 2255 39978 2272 45938
rect 2272 39978 2306 45938
rect 2306 39978 2321 45938
rect 2413 39978 2430 45938
rect 2430 39978 2464 45938
rect 2464 39978 2479 45938
rect 2571 39978 2588 45938
rect 2588 39978 2622 45938
rect 2622 39978 2637 45938
rect 2729 39978 2746 45938
rect 2746 39978 2780 45938
rect 2780 39978 2795 45938
rect 2887 39978 2904 45938
rect 2904 39978 2938 45938
rect 2938 39978 2953 45938
rect 3045 39978 3062 45938
rect 3062 39978 3096 45938
rect 3096 39978 3111 45938
rect 3203 39978 3220 45938
rect 3220 39978 3254 45938
rect 3254 39978 3269 45938
rect 3361 39978 3378 45938
rect 3378 39978 3412 45938
rect 3412 39978 3427 45938
rect 3519 39978 3536 45938
rect 3536 39978 3570 45938
rect 3570 39978 3585 45938
rect 3677 39978 3694 45938
rect 3694 39978 3728 45938
rect 3728 39978 3743 45938
rect 3835 39978 3852 45938
rect 3852 39978 3886 45938
rect 3886 39978 3901 45938
rect 3993 39978 4010 45938
rect 4010 39978 4044 45938
rect 4044 39978 4059 45938
rect 4151 39978 4168 45938
rect 4168 39978 4202 45938
rect 4202 39978 4217 45938
rect 4309 39978 4326 45938
rect 4326 39978 4360 45938
rect 4360 39978 4375 45938
rect 4467 39978 4484 45938
rect 4484 39978 4518 45938
rect 4518 39978 4533 45938
rect 4625 39978 4642 45938
rect 4642 39978 4676 45938
rect 4676 39978 4691 45938
rect 4783 39978 4800 45938
rect 4800 39978 4834 45938
rect 4834 39978 4849 45938
rect 4941 39978 4958 45938
rect 4958 39978 4992 45938
rect 4992 39978 5007 45938
rect 5099 39978 5116 45938
rect 5116 39978 5150 45938
rect 5150 39978 5165 45938
rect 5257 39978 5274 45938
rect 5274 39978 5308 45938
rect 5308 39978 5323 45938
rect 5415 39978 5432 45938
rect 5432 39978 5466 45938
rect 5466 39978 5481 45938
rect 5573 39978 5590 45938
rect 5590 39978 5624 45938
rect 5624 39978 5639 45938
rect 5731 39978 5748 45938
rect 5748 39978 5782 45938
rect 5782 39978 5797 45938
rect 5889 39978 5906 45938
rect 5906 39978 5940 45938
rect 5940 39978 5955 45938
rect 6047 39978 6064 45938
rect 6064 39978 6098 45938
rect 6098 39978 6113 45938
rect 6205 39978 6222 45938
rect 6222 39978 6256 45938
rect 6256 39978 6271 45938
rect -2980 39650 -2910 39850
rect -2590 39650 -2520 39850
rect -2480 39650 -2410 39850
rect -2090 39650 -2020 39850
rect -1980 39650 -1910 39850
rect -1590 39650 -1520 39850
rect -1480 39650 -1410 39850
rect -1090 39650 -1020 39850
rect -980 39650 -910 39850
rect -590 39650 -520 39850
rect -480 39650 -410 39850
rect -90 39650 -20 39850
rect 20 39650 90 39850
rect 410 39650 480 39850
rect 520 39650 590 39850
rect 910 39650 980 39850
rect 1330 39800 1400 39936
rect 6340 39936 6354 45980
rect 6354 39936 6392 45980
rect 6392 39936 6410 45980
rect 1552 39920 6186 39926
rect 1552 39886 1612 39920
rect 1612 39886 1702 39920
rect 1702 39886 1770 39920
rect 1770 39886 1860 39920
rect 1860 39886 1928 39920
rect 1928 39886 2018 39920
rect 2018 39886 2086 39920
rect 2086 39886 2176 39920
rect 2176 39886 2244 39920
rect 2244 39886 2334 39920
rect 2334 39886 2402 39920
rect 2402 39886 2492 39920
rect 2492 39886 2560 39920
rect 2560 39886 2650 39920
rect 2650 39886 2718 39920
rect 2718 39886 2808 39920
rect 2808 39886 2876 39920
rect 2876 39886 2966 39920
rect 2966 39886 3034 39920
rect 3034 39886 3124 39920
rect 3124 39886 3192 39920
rect 3192 39886 3282 39920
rect 3282 39886 3350 39920
rect 3350 39886 3440 39920
rect 3440 39886 3508 39920
rect 3508 39886 3598 39920
rect 3598 39886 3666 39920
rect 3666 39886 3756 39920
rect 3756 39886 3824 39920
rect 3824 39886 3914 39920
rect 3914 39886 3982 39920
rect 3982 39886 4072 39920
rect 4072 39886 4140 39920
rect 4140 39886 4230 39920
rect 4230 39886 4298 39920
rect 4298 39886 4388 39920
rect 4388 39886 4456 39920
rect 4456 39886 4546 39920
rect 4546 39886 4614 39920
rect 4614 39886 4704 39920
rect 4704 39886 4772 39920
rect 4772 39886 4862 39920
rect 4862 39886 4930 39920
rect 4930 39886 5020 39920
rect 5020 39886 5088 39920
rect 5088 39886 5178 39920
rect 5178 39886 5246 39920
rect 5246 39886 5336 39920
rect 5336 39886 5404 39920
rect 5404 39886 5494 39920
rect 5494 39886 5562 39920
rect 5562 39886 5652 39920
rect 5652 39886 5720 39920
rect 5720 39886 5810 39920
rect 5810 39886 5878 39920
rect 5878 39886 5968 39920
rect 5968 39886 6036 39920
rect 6036 39886 6126 39920
rect 6126 39886 6186 39920
rect 1552 39826 6186 39886
rect 6340 39800 6410 39936
rect 7630 45980 7700 46120
rect 7852 46030 12486 46090
rect 7852 45996 7912 46030
rect 7912 45996 8002 46030
rect 8002 45996 8070 46030
rect 8070 45996 8160 46030
rect 8160 45996 8228 46030
rect 8228 45996 8318 46030
rect 8318 45996 8386 46030
rect 8386 45996 8476 46030
rect 8476 45996 8544 46030
rect 8544 45996 8634 46030
rect 8634 45996 8702 46030
rect 8702 45996 8792 46030
rect 8792 45996 8860 46030
rect 8860 45996 8950 46030
rect 8950 45996 9018 46030
rect 9018 45996 9108 46030
rect 9108 45996 9176 46030
rect 9176 45996 9266 46030
rect 9266 45996 9334 46030
rect 9334 45996 9424 46030
rect 9424 45996 9492 46030
rect 9492 45996 9582 46030
rect 9582 45996 9650 46030
rect 9650 45996 9740 46030
rect 9740 45996 9808 46030
rect 9808 45996 9898 46030
rect 9898 45996 9966 46030
rect 9966 45996 10056 46030
rect 10056 45996 10124 46030
rect 10124 45996 10214 46030
rect 10214 45996 10282 46030
rect 10282 45996 10372 46030
rect 10372 45996 10440 46030
rect 10440 45996 10530 46030
rect 10530 45996 10598 46030
rect 10598 45996 10688 46030
rect 10688 45996 10756 46030
rect 10756 45996 10846 46030
rect 10846 45996 10914 46030
rect 10914 45996 11004 46030
rect 11004 45996 11072 46030
rect 11072 45996 11162 46030
rect 11162 45996 11230 46030
rect 11230 45996 11320 46030
rect 11320 45996 11388 46030
rect 11388 45996 11478 46030
rect 11478 45996 11546 46030
rect 11546 45996 11636 46030
rect 11636 45996 11704 46030
rect 11704 45996 11794 46030
rect 11794 45996 11862 46030
rect 11862 45996 11952 46030
rect 11952 45996 12020 46030
rect 12020 45996 12110 46030
rect 12110 45996 12178 46030
rect 12178 45996 12268 46030
rect 12268 45996 12336 46030
rect 12336 45996 12426 46030
rect 12426 45996 12486 46030
rect 7852 45990 12486 45996
rect 7630 39936 7646 45980
rect 7646 39936 7684 45980
rect 7684 39936 7700 45980
rect 12640 45980 12710 46120
rect 13020 46150 13090 46350
rect 13410 46150 13480 46350
rect 13520 46150 13590 46350
rect 13910 46150 13980 46350
rect 19150 46410 19350 46480
rect 19650 46410 19850 46480
rect 19020 46150 19090 46350
rect 13150 46020 13350 46090
rect 13650 46020 13850 46090
rect 7765 39978 7782 45938
rect 7782 39978 7816 45938
rect 7816 39978 7831 45938
rect 7923 39978 7940 45938
rect 7940 39978 7974 45938
rect 7974 39978 7989 45938
rect 8081 39978 8098 45938
rect 8098 39978 8132 45938
rect 8132 39978 8147 45938
rect 8239 39978 8256 45938
rect 8256 39978 8290 45938
rect 8290 39978 8305 45938
rect 8397 39978 8414 45938
rect 8414 39978 8448 45938
rect 8448 39978 8463 45938
rect 8555 39978 8572 45938
rect 8572 39978 8606 45938
rect 8606 39978 8621 45938
rect 8713 39978 8730 45938
rect 8730 39978 8764 45938
rect 8764 39978 8779 45938
rect 8871 39978 8888 45938
rect 8888 39978 8922 45938
rect 8922 39978 8937 45938
rect 9029 39978 9046 45938
rect 9046 39978 9080 45938
rect 9080 39978 9095 45938
rect 9187 39978 9204 45938
rect 9204 39978 9238 45938
rect 9238 39978 9253 45938
rect 9345 39978 9362 45938
rect 9362 39978 9396 45938
rect 9396 39978 9411 45938
rect 9503 39978 9520 45938
rect 9520 39978 9554 45938
rect 9554 39978 9569 45938
rect 9661 39978 9678 45938
rect 9678 39978 9712 45938
rect 9712 39978 9727 45938
rect 9819 39978 9836 45938
rect 9836 39978 9870 45938
rect 9870 39978 9885 45938
rect 9977 39978 9994 45938
rect 9994 39978 10028 45938
rect 10028 39978 10043 45938
rect 10135 39978 10152 45938
rect 10152 39978 10186 45938
rect 10186 39978 10201 45938
rect 10293 39978 10310 45938
rect 10310 39978 10344 45938
rect 10344 39978 10359 45938
rect 10451 39978 10468 45938
rect 10468 39978 10502 45938
rect 10502 39978 10517 45938
rect 10609 39978 10626 45938
rect 10626 39978 10660 45938
rect 10660 39978 10675 45938
rect 10767 39978 10784 45938
rect 10784 39978 10818 45938
rect 10818 39978 10833 45938
rect 10925 39978 10942 45938
rect 10942 39978 10976 45938
rect 10976 39978 10991 45938
rect 11083 39978 11100 45938
rect 11100 39978 11134 45938
rect 11134 39978 11149 45938
rect 11241 39978 11258 45938
rect 11258 39978 11292 45938
rect 11292 39978 11307 45938
rect 11399 39978 11416 45938
rect 11416 39978 11450 45938
rect 11450 39978 11465 45938
rect 11557 39978 11574 45938
rect 11574 39978 11608 45938
rect 11608 39978 11623 45938
rect 11715 39978 11732 45938
rect 11732 39978 11766 45938
rect 11766 39978 11781 45938
rect 11873 39978 11890 45938
rect 11890 39978 11924 45938
rect 11924 39978 11939 45938
rect 12031 39978 12048 45938
rect 12048 39978 12082 45938
rect 12082 39978 12097 45938
rect 12189 39978 12206 45938
rect 12206 39978 12240 45938
rect 12240 39978 12255 45938
rect 12347 39978 12364 45938
rect 12364 39978 12398 45938
rect 12398 39978 12413 45938
rect 12505 39978 12522 45938
rect 12522 39978 12556 45938
rect 12556 39978 12571 45938
rect 7630 39800 7700 39936
rect 12640 39936 12654 45980
rect 12654 39936 12692 45980
rect 12692 39936 12710 45980
rect 7852 39920 12486 39926
rect 7852 39886 7912 39920
rect 7912 39886 8002 39920
rect 8002 39886 8070 39920
rect 8070 39886 8160 39920
rect 8160 39886 8228 39920
rect 8228 39886 8318 39920
rect 8318 39886 8386 39920
rect 8386 39886 8476 39920
rect 8476 39886 8544 39920
rect 8544 39886 8634 39920
rect 8634 39886 8702 39920
rect 8702 39886 8792 39920
rect 8792 39886 8860 39920
rect 8860 39886 8950 39920
rect 8950 39886 9018 39920
rect 9018 39886 9108 39920
rect 9108 39886 9176 39920
rect 9176 39886 9266 39920
rect 9266 39886 9334 39920
rect 9334 39886 9424 39920
rect 9424 39886 9492 39920
rect 9492 39886 9582 39920
rect 9582 39886 9650 39920
rect 9650 39886 9740 39920
rect 9740 39886 9808 39920
rect 9808 39886 9898 39920
rect 9898 39886 9966 39920
rect 9966 39886 10056 39920
rect 10056 39886 10124 39920
rect 10124 39886 10214 39920
rect 10214 39886 10282 39920
rect 10282 39886 10372 39920
rect 10372 39886 10440 39920
rect 10440 39886 10530 39920
rect 10530 39886 10598 39920
rect 10598 39886 10688 39920
rect 10688 39886 10756 39920
rect 10756 39886 10846 39920
rect 10846 39886 10914 39920
rect 10914 39886 11004 39920
rect 11004 39886 11072 39920
rect 11072 39886 11162 39920
rect 11162 39886 11230 39920
rect 11230 39886 11320 39920
rect 11320 39886 11388 39920
rect 11388 39886 11478 39920
rect 11478 39886 11546 39920
rect 11546 39886 11636 39920
rect 11636 39886 11704 39920
rect 11704 39886 11794 39920
rect 11794 39886 11862 39920
rect 11862 39886 11952 39920
rect 11952 39886 12020 39920
rect 12020 39886 12110 39920
rect 12110 39886 12178 39920
rect 12178 39886 12268 39920
rect 12268 39886 12336 39920
rect 12336 39886 12426 39920
rect 12426 39886 12486 39920
rect 7852 39826 12486 39886
rect 12640 39800 12710 39936
rect 13930 45980 14000 46120
rect 19410 46150 19480 46350
rect 19520 46150 19590 46350
rect 19910 46150 19980 46350
rect 25650 46410 25850 46480
rect 26150 46410 26350 46480
rect 14152 46030 18786 46090
rect 14152 45996 14212 46030
rect 14212 45996 14302 46030
rect 14302 45996 14370 46030
rect 14370 45996 14460 46030
rect 14460 45996 14528 46030
rect 14528 45996 14618 46030
rect 14618 45996 14686 46030
rect 14686 45996 14776 46030
rect 14776 45996 14844 46030
rect 14844 45996 14934 46030
rect 14934 45996 15002 46030
rect 15002 45996 15092 46030
rect 15092 45996 15160 46030
rect 15160 45996 15250 46030
rect 15250 45996 15318 46030
rect 15318 45996 15408 46030
rect 15408 45996 15476 46030
rect 15476 45996 15566 46030
rect 15566 45996 15634 46030
rect 15634 45996 15724 46030
rect 15724 45996 15792 46030
rect 15792 45996 15882 46030
rect 15882 45996 15950 46030
rect 15950 45996 16040 46030
rect 16040 45996 16108 46030
rect 16108 45996 16198 46030
rect 16198 45996 16266 46030
rect 16266 45996 16356 46030
rect 16356 45996 16424 46030
rect 16424 45996 16514 46030
rect 16514 45996 16582 46030
rect 16582 45996 16672 46030
rect 16672 45996 16740 46030
rect 16740 45996 16830 46030
rect 16830 45996 16898 46030
rect 16898 45996 16988 46030
rect 16988 45996 17056 46030
rect 17056 45996 17146 46030
rect 17146 45996 17214 46030
rect 17214 45996 17304 46030
rect 17304 45996 17372 46030
rect 17372 45996 17462 46030
rect 17462 45996 17530 46030
rect 17530 45996 17620 46030
rect 17620 45996 17688 46030
rect 17688 45996 17778 46030
rect 17778 45996 17846 46030
rect 17846 45996 17936 46030
rect 17936 45996 18004 46030
rect 18004 45996 18094 46030
rect 18094 45996 18162 46030
rect 18162 45996 18252 46030
rect 18252 45996 18320 46030
rect 18320 45996 18410 46030
rect 18410 45996 18478 46030
rect 18478 45996 18568 46030
rect 18568 45996 18636 46030
rect 18636 45996 18726 46030
rect 18726 45996 18786 46030
rect 14152 45990 18786 45996
rect 13930 39936 13946 45980
rect 13946 39936 13984 45980
rect 13984 39936 14000 45980
rect 18940 45980 19010 46120
rect 19150 46020 19350 46090
rect 19650 46020 19850 46090
rect 25520 46150 25590 46350
rect 14065 39978 14082 45938
rect 14082 39978 14116 45938
rect 14116 39978 14131 45938
rect 14223 39978 14240 45938
rect 14240 39978 14274 45938
rect 14274 39978 14289 45938
rect 14381 39978 14398 45938
rect 14398 39978 14432 45938
rect 14432 39978 14447 45938
rect 14539 39978 14556 45938
rect 14556 39978 14590 45938
rect 14590 39978 14605 45938
rect 14697 39978 14714 45938
rect 14714 39978 14748 45938
rect 14748 39978 14763 45938
rect 14855 39978 14872 45938
rect 14872 39978 14906 45938
rect 14906 39978 14921 45938
rect 15013 39978 15030 45938
rect 15030 39978 15064 45938
rect 15064 39978 15079 45938
rect 15171 39978 15188 45938
rect 15188 39978 15222 45938
rect 15222 39978 15237 45938
rect 15329 39978 15346 45938
rect 15346 39978 15380 45938
rect 15380 39978 15395 45938
rect 15487 39978 15504 45938
rect 15504 39978 15538 45938
rect 15538 39978 15553 45938
rect 15645 39978 15662 45938
rect 15662 39978 15696 45938
rect 15696 39978 15711 45938
rect 15803 39978 15820 45938
rect 15820 39978 15854 45938
rect 15854 39978 15869 45938
rect 15961 39978 15978 45938
rect 15978 39978 16012 45938
rect 16012 39978 16027 45938
rect 16119 39978 16136 45938
rect 16136 39978 16170 45938
rect 16170 39978 16185 45938
rect 16277 39978 16294 45938
rect 16294 39978 16328 45938
rect 16328 39978 16343 45938
rect 16435 39978 16452 45938
rect 16452 39978 16486 45938
rect 16486 39978 16501 45938
rect 16593 39978 16610 45938
rect 16610 39978 16644 45938
rect 16644 39978 16659 45938
rect 16751 39978 16768 45938
rect 16768 39978 16802 45938
rect 16802 39978 16817 45938
rect 16909 39978 16926 45938
rect 16926 39978 16960 45938
rect 16960 39978 16975 45938
rect 17067 39978 17084 45938
rect 17084 39978 17118 45938
rect 17118 39978 17133 45938
rect 17225 39978 17242 45938
rect 17242 39978 17276 45938
rect 17276 39978 17291 45938
rect 17383 39978 17400 45938
rect 17400 39978 17434 45938
rect 17434 39978 17449 45938
rect 17541 39978 17558 45938
rect 17558 39978 17592 45938
rect 17592 39978 17607 45938
rect 17699 39978 17716 45938
rect 17716 39978 17750 45938
rect 17750 39978 17765 45938
rect 17857 39978 17874 45938
rect 17874 39978 17908 45938
rect 17908 39978 17923 45938
rect 18015 39978 18032 45938
rect 18032 39978 18066 45938
rect 18066 39978 18081 45938
rect 18173 39978 18190 45938
rect 18190 39978 18224 45938
rect 18224 39978 18239 45938
rect 18331 39978 18348 45938
rect 18348 39978 18382 45938
rect 18382 39978 18397 45938
rect 18489 39978 18506 45938
rect 18506 39978 18540 45938
rect 18540 39978 18555 45938
rect 18647 39978 18664 45938
rect 18664 39978 18698 45938
rect 18698 39978 18713 45938
rect 18805 39978 18822 45938
rect 18822 39978 18856 45938
rect 18856 39978 18871 45938
rect 13930 39800 14000 39936
rect 18940 39936 18954 45980
rect 18954 39936 18992 45980
rect 18992 39936 19010 45980
rect 14152 39920 18786 39926
rect 14152 39886 14212 39920
rect 14212 39886 14302 39920
rect 14302 39886 14370 39920
rect 14370 39886 14460 39920
rect 14460 39886 14528 39920
rect 14528 39886 14618 39920
rect 14618 39886 14686 39920
rect 14686 39886 14776 39920
rect 14776 39886 14844 39920
rect 14844 39886 14934 39920
rect 14934 39886 15002 39920
rect 15002 39886 15092 39920
rect 15092 39886 15160 39920
rect 15160 39886 15250 39920
rect 15250 39886 15318 39920
rect 15318 39886 15408 39920
rect 15408 39886 15476 39920
rect 15476 39886 15566 39920
rect 15566 39886 15634 39920
rect 15634 39886 15724 39920
rect 15724 39886 15792 39920
rect 15792 39886 15882 39920
rect 15882 39886 15950 39920
rect 15950 39886 16040 39920
rect 16040 39886 16108 39920
rect 16108 39886 16198 39920
rect 16198 39886 16266 39920
rect 16266 39886 16356 39920
rect 16356 39886 16424 39920
rect 16424 39886 16514 39920
rect 16514 39886 16582 39920
rect 16582 39886 16672 39920
rect 16672 39886 16740 39920
rect 16740 39886 16830 39920
rect 16830 39886 16898 39920
rect 16898 39886 16988 39920
rect 16988 39886 17056 39920
rect 17056 39886 17146 39920
rect 17146 39886 17214 39920
rect 17214 39886 17304 39920
rect 17304 39886 17372 39920
rect 17372 39886 17462 39920
rect 17462 39886 17530 39920
rect 17530 39886 17620 39920
rect 17620 39886 17688 39920
rect 17688 39886 17778 39920
rect 17778 39886 17846 39920
rect 17846 39886 17936 39920
rect 17936 39886 18004 39920
rect 18004 39886 18094 39920
rect 18094 39886 18162 39920
rect 18162 39886 18252 39920
rect 18252 39886 18320 39920
rect 18320 39886 18410 39920
rect 18410 39886 18478 39920
rect 18478 39886 18568 39920
rect 18568 39886 18636 39920
rect 18636 39886 18726 39920
rect 18726 39886 18786 39920
rect 14152 39826 18786 39886
rect 18940 39800 19010 39936
rect 20230 45980 20300 46120
rect 25910 46150 25980 46350
rect 26020 46150 26090 46350
rect 26410 46150 26480 46350
rect 20452 46030 25086 46090
rect 20452 45996 20512 46030
rect 20512 45996 20602 46030
rect 20602 45996 20670 46030
rect 20670 45996 20760 46030
rect 20760 45996 20828 46030
rect 20828 45996 20918 46030
rect 20918 45996 20986 46030
rect 20986 45996 21076 46030
rect 21076 45996 21144 46030
rect 21144 45996 21234 46030
rect 21234 45996 21302 46030
rect 21302 45996 21392 46030
rect 21392 45996 21460 46030
rect 21460 45996 21550 46030
rect 21550 45996 21618 46030
rect 21618 45996 21708 46030
rect 21708 45996 21776 46030
rect 21776 45996 21866 46030
rect 21866 45996 21934 46030
rect 21934 45996 22024 46030
rect 22024 45996 22092 46030
rect 22092 45996 22182 46030
rect 22182 45996 22250 46030
rect 22250 45996 22340 46030
rect 22340 45996 22408 46030
rect 22408 45996 22498 46030
rect 22498 45996 22566 46030
rect 22566 45996 22656 46030
rect 22656 45996 22724 46030
rect 22724 45996 22814 46030
rect 22814 45996 22882 46030
rect 22882 45996 22972 46030
rect 22972 45996 23040 46030
rect 23040 45996 23130 46030
rect 23130 45996 23198 46030
rect 23198 45996 23288 46030
rect 23288 45996 23356 46030
rect 23356 45996 23446 46030
rect 23446 45996 23514 46030
rect 23514 45996 23604 46030
rect 23604 45996 23672 46030
rect 23672 45996 23762 46030
rect 23762 45996 23830 46030
rect 23830 45996 23920 46030
rect 23920 45996 23988 46030
rect 23988 45996 24078 46030
rect 24078 45996 24146 46030
rect 24146 45996 24236 46030
rect 24236 45996 24304 46030
rect 24304 45996 24394 46030
rect 24394 45996 24462 46030
rect 24462 45996 24552 46030
rect 24552 45996 24620 46030
rect 24620 45996 24710 46030
rect 24710 45996 24778 46030
rect 24778 45996 24868 46030
rect 24868 45996 24936 46030
rect 24936 45996 25026 46030
rect 25026 45996 25086 46030
rect 20452 45990 25086 45996
rect 20230 39936 20246 45980
rect 20246 39936 20284 45980
rect 20284 39936 20300 45980
rect 25240 45980 25310 46120
rect 25650 46020 25850 46090
rect 26150 46020 26350 46090
rect 20365 39978 20382 45938
rect 20382 39978 20416 45938
rect 20416 39978 20431 45938
rect 20523 39978 20540 45938
rect 20540 39978 20574 45938
rect 20574 39978 20589 45938
rect 20681 39978 20698 45938
rect 20698 39978 20732 45938
rect 20732 39978 20747 45938
rect 20839 39978 20856 45938
rect 20856 39978 20890 45938
rect 20890 39978 20905 45938
rect 20997 39978 21014 45938
rect 21014 39978 21048 45938
rect 21048 39978 21063 45938
rect 21155 39978 21172 45938
rect 21172 39978 21206 45938
rect 21206 39978 21221 45938
rect 21313 39978 21330 45938
rect 21330 39978 21364 45938
rect 21364 39978 21379 45938
rect 21471 39978 21488 45938
rect 21488 39978 21522 45938
rect 21522 39978 21537 45938
rect 21629 39978 21646 45938
rect 21646 39978 21680 45938
rect 21680 39978 21695 45938
rect 21787 39978 21804 45938
rect 21804 39978 21838 45938
rect 21838 39978 21853 45938
rect 21945 39978 21962 45938
rect 21962 39978 21996 45938
rect 21996 39978 22011 45938
rect 22103 39978 22120 45938
rect 22120 39978 22154 45938
rect 22154 39978 22169 45938
rect 22261 39978 22278 45938
rect 22278 39978 22312 45938
rect 22312 39978 22327 45938
rect 22419 39978 22436 45938
rect 22436 39978 22470 45938
rect 22470 39978 22485 45938
rect 22577 39978 22594 45938
rect 22594 39978 22628 45938
rect 22628 39978 22643 45938
rect 22735 39978 22752 45938
rect 22752 39978 22786 45938
rect 22786 39978 22801 45938
rect 22893 39978 22910 45938
rect 22910 39978 22944 45938
rect 22944 39978 22959 45938
rect 23051 39978 23068 45938
rect 23068 39978 23102 45938
rect 23102 39978 23117 45938
rect 23209 39978 23226 45938
rect 23226 39978 23260 45938
rect 23260 39978 23275 45938
rect 23367 39978 23384 45938
rect 23384 39978 23418 45938
rect 23418 39978 23433 45938
rect 23525 39978 23542 45938
rect 23542 39978 23576 45938
rect 23576 39978 23591 45938
rect 23683 39978 23700 45938
rect 23700 39978 23734 45938
rect 23734 39978 23749 45938
rect 23841 39978 23858 45938
rect 23858 39978 23892 45938
rect 23892 39978 23907 45938
rect 23999 39978 24016 45938
rect 24016 39978 24050 45938
rect 24050 39978 24065 45938
rect 24157 39978 24174 45938
rect 24174 39978 24208 45938
rect 24208 39978 24223 45938
rect 24315 39978 24332 45938
rect 24332 39978 24366 45938
rect 24366 39978 24381 45938
rect 24473 39978 24490 45938
rect 24490 39978 24524 45938
rect 24524 39978 24539 45938
rect 24631 39978 24648 45938
rect 24648 39978 24682 45938
rect 24682 39978 24697 45938
rect 24789 39978 24806 45938
rect 24806 39978 24840 45938
rect 24840 39978 24855 45938
rect 24947 39978 24964 45938
rect 24964 39978 24998 45938
rect 24998 39978 25013 45938
rect 25105 39978 25122 45938
rect 25122 39978 25156 45938
rect 25156 39978 25171 45938
rect 20230 39800 20300 39936
rect 25240 39936 25254 45980
rect 25254 39936 25292 45980
rect 25292 39936 25310 45980
rect 25650 45910 25850 45980
rect 26150 45910 26350 45980
rect 25520 45650 25590 45850
rect 25910 45650 25980 45850
rect 26020 45650 26090 45850
rect 26410 45650 26480 45850
rect 25650 45520 25850 45590
rect 26150 45520 26350 45590
rect 25650 45410 25850 45480
rect 26150 45410 26350 45480
rect 25520 45150 25590 45350
rect 25910 45150 25980 45350
rect 26020 45150 26090 45350
rect 26410 45150 26480 45350
rect 25650 45020 25850 45090
rect 26150 45020 26350 45090
rect 25650 44910 25850 44980
rect 26150 44910 26350 44980
rect 25520 44650 25590 44850
rect 25910 44650 25980 44850
rect 26020 44650 26090 44850
rect 26410 44650 26480 44850
rect 25650 44520 25850 44590
rect 26150 44520 26350 44590
rect 25650 44410 25850 44480
rect 26150 44410 26350 44480
rect 25520 44150 25590 44350
rect 25910 44150 25980 44350
rect 26020 44150 26090 44350
rect 26410 44150 26480 44350
rect 25650 44020 25850 44090
rect 26150 44020 26350 44090
rect 25650 43910 25850 43980
rect 26150 43910 26350 43980
rect 25520 43650 25590 43850
rect 25910 43650 25980 43850
rect 26020 43650 26090 43850
rect 26410 43650 26480 43850
rect 25650 43520 25850 43590
rect 26150 43520 26350 43590
rect 25650 43410 25850 43480
rect 26150 43410 26350 43480
rect 25520 43150 25590 43350
rect 25910 43150 25980 43350
rect 26020 43150 26090 43350
rect 26410 43150 26480 43350
rect 25650 43020 25850 43090
rect 26150 43020 26350 43090
rect 25650 42910 25850 42980
rect 26150 42910 26350 42980
rect 25520 42650 25590 42850
rect 25910 42650 25980 42850
rect 26020 42650 26090 42850
rect 26410 42650 26480 42850
rect 25650 42520 25850 42590
rect 26150 42520 26350 42590
rect 25650 42410 25850 42480
rect 26150 42410 26350 42480
rect 25520 42150 25590 42350
rect 25910 42150 25980 42350
rect 26020 42150 26090 42350
rect 26410 42150 26480 42350
rect 25650 42020 25850 42090
rect 26150 42020 26350 42090
rect 25650 41910 25850 41980
rect 26150 41910 26350 41980
rect 25520 41650 25590 41850
rect 25910 41650 25980 41850
rect 26020 41650 26090 41850
rect 26410 41650 26480 41850
rect 25650 41520 25850 41590
rect 26150 41520 26350 41590
rect 25650 41410 25850 41480
rect 26150 41410 26350 41480
rect 25520 41150 25590 41350
rect 25910 41150 25980 41350
rect 26020 41150 26090 41350
rect 26410 41150 26480 41350
rect 25650 41020 25850 41090
rect 26150 41020 26350 41090
rect 25650 40910 25850 40980
rect 26150 40910 26350 40980
rect 25520 40650 25590 40850
rect 25910 40650 25980 40850
rect 26020 40650 26090 40850
rect 26410 40650 26480 40850
rect 25650 40520 25850 40590
rect 26150 40520 26350 40590
rect 25650 40410 25850 40480
rect 26150 40410 26350 40480
rect 25520 40150 25590 40350
rect 25910 40150 25980 40350
rect 26020 40150 26090 40350
rect 26410 40150 26480 40350
rect 25650 40020 25850 40090
rect 26150 40020 26350 40090
rect 20452 39920 25086 39926
rect 20452 39886 20512 39920
rect 20512 39886 20602 39920
rect 20602 39886 20670 39920
rect 20670 39886 20760 39920
rect 20760 39886 20828 39920
rect 20828 39886 20918 39920
rect 20918 39886 20986 39920
rect 20986 39886 21076 39920
rect 21076 39886 21144 39920
rect 21144 39886 21234 39920
rect 21234 39886 21302 39920
rect 21302 39886 21392 39920
rect 21392 39886 21460 39920
rect 21460 39886 21550 39920
rect 21550 39886 21618 39920
rect 21618 39886 21708 39920
rect 21708 39886 21776 39920
rect 21776 39886 21866 39920
rect 21866 39886 21934 39920
rect 21934 39886 22024 39920
rect 22024 39886 22092 39920
rect 22092 39886 22182 39920
rect 22182 39886 22250 39920
rect 22250 39886 22340 39920
rect 22340 39886 22408 39920
rect 22408 39886 22498 39920
rect 22498 39886 22566 39920
rect 22566 39886 22656 39920
rect 22656 39886 22724 39920
rect 22724 39886 22814 39920
rect 22814 39886 22882 39920
rect 22882 39886 22972 39920
rect 22972 39886 23040 39920
rect 23040 39886 23130 39920
rect 23130 39886 23198 39920
rect 23198 39886 23288 39920
rect 23288 39886 23356 39920
rect 23356 39886 23446 39920
rect 23446 39886 23514 39920
rect 23514 39886 23604 39920
rect 23604 39886 23672 39920
rect 23672 39886 23762 39920
rect 23762 39886 23830 39920
rect 23830 39886 23920 39920
rect 23920 39886 23988 39920
rect 23988 39886 24078 39920
rect 24078 39886 24146 39920
rect 24146 39886 24236 39920
rect 24236 39886 24304 39920
rect 24304 39886 24394 39920
rect 24394 39886 24462 39920
rect 24462 39886 24552 39920
rect 24552 39886 24620 39920
rect 24620 39886 24710 39920
rect 24710 39886 24778 39920
rect 24778 39886 24868 39920
rect 24868 39886 24936 39920
rect 24936 39886 25026 39920
rect 25026 39886 25086 39920
rect 20452 39826 25086 39886
rect 25240 39800 25310 39936
rect 25650 39910 25850 39980
rect 26150 39910 26350 39980
rect 26650 39910 26850 39980
rect 27150 39910 27350 39980
rect 27650 39910 27850 39980
rect 28150 39910 28350 39980
rect 28650 39910 28850 39980
rect 29150 39910 29350 39980
rect -2850 39520 -2650 39590
rect -2350 39520 -2150 39590
rect -1850 39520 -1650 39590
rect -1350 39520 -1150 39590
rect -850 39520 -650 39590
rect -350 39520 -150 39590
rect 150 39520 350 39590
rect 650 39520 850 39590
rect -2850 39410 -2650 39480
rect -2350 39410 -2150 39480
rect -1850 39410 -1650 39480
rect -1350 39410 -1150 39480
rect -850 39410 -650 39480
rect -350 39410 -150 39480
rect 150 39410 350 39480
rect 650 39410 850 39480
rect -2980 39150 -2910 39350
rect -2590 39150 -2520 39350
rect -2480 39150 -2410 39350
rect -2090 39150 -2020 39350
rect -1980 39150 -1910 39350
rect -1590 39150 -1520 39350
rect -1480 39150 -1410 39350
rect -1090 39150 -1020 39350
rect -980 39150 -910 39350
rect -590 39150 -520 39350
rect -480 39150 -410 39350
rect -90 39150 -20 39350
rect 20 39150 90 39350
rect 410 39150 480 39350
rect 520 39150 590 39350
rect 910 39150 980 39350
rect 25520 39650 25590 39850
rect 25910 39650 25980 39850
rect 26020 39650 26090 39850
rect 26410 39650 26480 39850
rect 26520 39650 26590 39850
rect 26910 39650 26980 39850
rect 27020 39650 27090 39850
rect 27410 39650 27480 39850
rect 27520 39650 27590 39850
rect 27910 39650 27980 39850
rect 28020 39650 28090 39850
rect 28410 39650 28480 39850
rect 28520 39650 28590 39850
rect 28910 39650 28980 39850
rect 29020 39650 29090 39850
rect 29410 39650 29480 39850
rect 25650 39520 25850 39590
rect 26150 39520 26350 39590
rect 26650 39520 26850 39590
rect 27150 39520 27350 39590
rect 27650 39520 27850 39590
rect 28150 39520 28350 39590
rect 28650 39520 28850 39590
rect 29150 39520 29350 39590
rect 25650 39410 25850 39480
rect 26150 39410 26350 39480
rect 26650 39410 26850 39480
rect 27150 39410 27350 39480
rect 27650 39410 27850 39480
rect 28150 39410 28350 39480
rect 28650 39410 28850 39480
rect 29150 39410 29350 39480
rect -2850 39020 -2650 39090
rect -2350 39020 -2150 39090
rect -1850 39020 -1650 39090
rect -1350 39020 -1150 39090
rect -850 39020 -650 39090
rect -350 39020 -150 39090
rect 150 39020 350 39090
rect 650 39020 850 39090
rect 1330 38980 1400 39120
rect 1552 39030 6186 39090
rect 1552 38996 1612 39030
rect 1612 38996 1702 39030
rect 1702 38996 1770 39030
rect 1770 38996 1860 39030
rect 1860 38996 1928 39030
rect 1928 38996 2018 39030
rect 2018 38996 2086 39030
rect 2086 38996 2176 39030
rect 2176 38996 2244 39030
rect 2244 38996 2334 39030
rect 2334 38996 2402 39030
rect 2402 38996 2492 39030
rect 2492 38996 2560 39030
rect 2560 38996 2650 39030
rect 2650 38996 2718 39030
rect 2718 38996 2808 39030
rect 2808 38996 2876 39030
rect 2876 38996 2966 39030
rect 2966 38996 3034 39030
rect 3034 38996 3124 39030
rect 3124 38996 3192 39030
rect 3192 38996 3282 39030
rect 3282 38996 3350 39030
rect 3350 38996 3440 39030
rect 3440 38996 3508 39030
rect 3508 38996 3598 39030
rect 3598 38996 3666 39030
rect 3666 38996 3756 39030
rect 3756 38996 3824 39030
rect 3824 38996 3914 39030
rect 3914 38996 3982 39030
rect 3982 38996 4072 39030
rect 4072 38996 4140 39030
rect 4140 38996 4230 39030
rect 4230 38996 4298 39030
rect 4298 38996 4388 39030
rect 4388 38996 4456 39030
rect 4456 38996 4546 39030
rect 4546 38996 4614 39030
rect 4614 38996 4704 39030
rect 4704 38996 4772 39030
rect 4772 38996 4862 39030
rect 4862 38996 4930 39030
rect 4930 38996 5020 39030
rect 5020 38996 5088 39030
rect 5088 38996 5178 39030
rect 5178 38996 5246 39030
rect 5246 38996 5336 39030
rect 5336 38996 5404 39030
rect 5404 38996 5494 39030
rect 5494 38996 5562 39030
rect 5562 38996 5652 39030
rect 5652 38996 5720 39030
rect 5720 38996 5810 39030
rect 5810 38996 5878 39030
rect 5878 38996 5968 39030
rect 5968 38996 6036 39030
rect 6036 38996 6126 39030
rect 6126 38996 6186 39030
rect 1552 38990 6186 38996
rect 150 38910 350 38980
rect 650 38910 850 38980
rect 20 38650 90 38850
rect 410 38650 480 38850
rect 520 38650 590 38850
rect 910 38650 980 38850
rect 150 38520 350 38590
rect 650 38520 850 38590
rect 150 38410 350 38480
rect 650 38410 850 38480
rect 20 38150 90 38350
rect 410 38150 480 38350
rect 520 38150 590 38350
rect 910 38150 980 38350
rect 150 38020 350 38090
rect 650 38020 850 38090
rect 150 37910 350 37980
rect 650 37910 850 37980
rect 20 37650 90 37850
rect 410 37650 480 37850
rect 520 37650 590 37850
rect 910 37650 980 37850
rect 150 37520 350 37590
rect 650 37520 850 37590
rect 150 37410 350 37480
rect 650 37410 850 37480
rect 20 37150 90 37350
rect 410 37150 480 37350
rect 520 37150 590 37350
rect 910 37150 980 37350
rect 150 37020 350 37090
rect 650 37020 850 37090
rect 150 36910 350 36980
rect 650 36910 850 36980
rect 20 36650 90 36850
rect 410 36650 480 36850
rect 520 36650 590 36850
rect 910 36650 980 36850
rect 150 36520 350 36590
rect 650 36520 850 36590
rect 150 36410 350 36480
rect 650 36410 850 36480
rect 20 36150 90 36350
rect 410 36150 480 36350
rect 520 36150 590 36350
rect 910 36150 980 36350
rect 150 36020 350 36090
rect 650 36020 850 36090
rect 150 35910 350 35980
rect 650 35910 850 35980
rect 20 35650 90 35850
rect 410 35650 480 35850
rect 520 35650 590 35850
rect 910 35650 980 35850
rect 150 35520 350 35590
rect 650 35520 850 35590
rect 150 35410 350 35480
rect 650 35410 850 35480
rect 20 35150 90 35350
rect 410 35150 480 35350
rect 520 35150 590 35350
rect 910 35150 980 35350
rect 150 35020 350 35090
rect 650 35020 850 35090
rect 150 34910 350 34980
rect 650 34910 850 34980
rect 20 34650 90 34850
rect 410 34650 480 34850
rect 520 34650 590 34850
rect 910 34650 980 34850
rect 150 34520 350 34590
rect 650 34520 850 34590
rect 150 34410 350 34480
rect 650 34410 850 34480
rect 20 34150 90 34350
rect 410 34150 480 34350
rect 520 34150 590 34350
rect 910 34150 980 34350
rect 150 34020 350 34090
rect 650 34020 850 34090
rect 150 33910 350 33980
rect 650 33910 850 33980
rect 20 33650 90 33850
rect 410 33650 480 33850
rect 520 33650 590 33850
rect 910 33650 980 33850
rect 150 33520 350 33590
rect 650 33520 850 33590
rect 150 33410 350 33480
rect 650 33410 850 33480
rect 20 33150 90 33350
rect 410 33150 480 33350
rect 520 33150 590 33350
rect 910 33150 980 33350
rect 150 33020 350 33090
rect 650 33020 850 33090
rect 150 32910 350 32980
rect 650 32910 850 32980
rect 1330 32936 1346 38980
rect 1346 32936 1384 38980
rect 1384 32936 1400 38980
rect 6340 38980 6410 39120
rect 1465 32978 1482 38938
rect 1482 32978 1516 38938
rect 1516 32978 1531 38938
rect 1623 32978 1640 38938
rect 1640 32978 1674 38938
rect 1674 32978 1689 38938
rect 1781 32978 1798 38938
rect 1798 32978 1832 38938
rect 1832 32978 1847 38938
rect 1939 32978 1956 38938
rect 1956 32978 1990 38938
rect 1990 32978 2005 38938
rect 2097 32978 2114 38938
rect 2114 32978 2148 38938
rect 2148 32978 2163 38938
rect 2255 32978 2272 38938
rect 2272 32978 2306 38938
rect 2306 32978 2321 38938
rect 2413 32978 2430 38938
rect 2430 32978 2464 38938
rect 2464 32978 2479 38938
rect 2571 32978 2588 38938
rect 2588 32978 2622 38938
rect 2622 32978 2637 38938
rect 2729 32978 2746 38938
rect 2746 32978 2780 38938
rect 2780 32978 2795 38938
rect 2887 32978 2904 38938
rect 2904 32978 2938 38938
rect 2938 32978 2953 38938
rect 3045 32978 3062 38938
rect 3062 32978 3096 38938
rect 3096 32978 3111 38938
rect 3203 32978 3220 38938
rect 3220 32978 3254 38938
rect 3254 32978 3269 38938
rect 3361 32978 3378 38938
rect 3378 32978 3412 38938
rect 3412 32978 3427 38938
rect 3519 32978 3536 38938
rect 3536 32978 3570 38938
rect 3570 32978 3585 38938
rect 3677 32978 3694 38938
rect 3694 32978 3728 38938
rect 3728 32978 3743 38938
rect 3835 32978 3852 38938
rect 3852 32978 3886 38938
rect 3886 32978 3901 38938
rect 3993 32978 4010 38938
rect 4010 32978 4044 38938
rect 4044 32978 4059 38938
rect 4151 32978 4168 38938
rect 4168 32978 4202 38938
rect 4202 32978 4217 38938
rect 4309 32978 4326 38938
rect 4326 32978 4360 38938
rect 4360 32978 4375 38938
rect 4467 32978 4484 38938
rect 4484 32978 4518 38938
rect 4518 32978 4533 38938
rect 4625 32978 4642 38938
rect 4642 32978 4676 38938
rect 4676 32978 4691 38938
rect 4783 32978 4800 38938
rect 4800 32978 4834 38938
rect 4834 32978 4849 38938
rect 4941 32978 4958 38938
rect 4958 32978 4992 38938
rect 4992 32978 5007 38938
rect 5099 32978 5116 38938
rect 5116 32978 5150 38938
rect 5150 32978 5165 38938
rect 5257 32978 5274 38938
rect 5274 32978 5308 38938
rect 5308 32978 5323 38938
rect 5415 32978 5432 38938
rect 5432 32978 5466 38938
rect 5466 32978 5481 38938
rect 5573 32978 5590 38938
rect 5590 32978 5624 38938
rect 5624 32978 5639 38938
rect 5731 32978 5748 38938
rect 5748 32978 5782 38938
rect 5782 32978 5797 38938
rect 5889 32978 5906 38938
rect 5906 32978 5940 38938
rect 5940 32978 5955 38938
rect 6047 32978 6064 38938
rect 6064 32978 6098 38938
rect 6098 32978 6113 38938
rect 6205 32978 6222 38938
rect 6222 32978 6256 38938
rect 6256 32978 6271 38938
rect 20 32650 90 32850
rect 410 32650 480 32850
rect 520 32650 590 32850
rect 910 32650 980 32850
rect 1330 32800 1400 32936
rect 6340 32936 6354 38980
rect 6354 32936 6392 38980
rect 6392 32936 6410 38980
rect 7630 38980 7700 39120
rect 7852 39030 12486 39090
rect 7852 38996 7912 39030
rect 7912 38996 8002 39030
rect 8002 38996 8070 39030
rect 8070 38996 8160 39030
rect 8160 38996 8228 39030
rect 8228 38996 8318 39030
rect 8318 38996 8386 39030
rect 8386 38996 8476 39030
rect 8476 38996 8544 39030
rect 8544 38996 8634 39030
rect 8634 38996 8702 39030
rect 8702 38996 8792 39030
rect 8792 38996 8860 39030
rect 8860 38996 8950 39030
rect 8950 38996 9018 39030
rect 9018 38996 9108 39030
rect 9108 38996 9176 39030
rect 9176 38996 9266 39030
rect 9266 38996 9334 39030
rect 9334 38996 9424 39030
rect 9424 38996 9492 39030
rect 9492 38996 9582 39030
rect 9582 38996 9650 39030
rect 9650 38996 9740 39030
rect 9740 38996 9808 39030
rect 9808 38996 9898 39030
rect 9898 38996 9966 39030
rect 9966 38996 10056 39030
rect 10056 38996 10124 39030
rect 10124 38996 10214 39030
rect 10214 38996 10282 39030
rect 10282 38996 10372 39030
rect 10372 38996 10440 39030
rect 10440 38996 10530 39030
rect 10530 38996 10598 39030
rect 10598 38996 10688 39030
rect 10688 38996 10756 39030
rect 10756 38996 10846 39030
rect 10846 38996 10914 39030
rect 10914 38996 11004 39030
rect 11004 38996 11072 39030
rect 11072 38996 11162 39030
rect 11162 38996 11230 39030
rect 11230 38996 11320 39030
rect 11320 38996 11388 39030
rect 11388 38996 11478 39030
rect 11478 38996 11546 39030
rect 11546 38996 11636 39030
rect 11636 38996 11704 39030
rect 11704 38996 11794 39030
rect 11794 38996 11862 39030
rect 11862 38996 11952 39030
rect 11952 38996 12020 39030
rect 12020 38996 12110 39030
rect 12110 38996 12178 39030
rect 12178 38996 12268 39030
rect 12268 38996 12336 39030
rect 12336 38996 12426 39030
rect 12426 38996 12486 39030
rect 7852 38990 12486 38996
rect 1552 32920 6186 32926
rect 1552 32886 1612 32920
rect 1612 32886 1702 32920
rect 1702 32886 1770 32920
rect 1770 32886 1860 32920
rect 1860 32886 1928 32920
rect 1928 32886 2018 32920
rect 2018 32886 2086 32920
rect 2086 32886 2176 32920
rect 2176 32886 2244 32920
rect 2244 32886 2334 32920
rect 2334 32886 2402 32920
rect 2402 32886 2492 32920
rect 2492 32886 2560 32920
rect 2560 32886 2650 32920
rect 2650 32886 2718 32920
rect 2718 32886 2808 32920
rect 2808 32886 2876 32920
rect 2876 32886 2966 32920
rect 2966 32886 3034 32920
rect 3034 32886 3124 32920
rect 3124 32886 3192 32920
rect 3192 32886 3282 32920
rect 3282 32886 3350 32920
rect 3350 32886 3440 32920
rect 3440 32886 3508 32920
rect 3508 32886 3598 32920
rect 3598 32886 3666 32920
rect 3666 32886 3756 32920
rect 3756 32886 3824 32920
rect 3824 32886 3914 32920
rect 3914 32886 3982 32920
rect 3982 32886 4072 32920
rect 4072 32886 4140 32920
rect 4140 32886 4230 32920
rect 4230 32886 4298 32920
rect 4298 32886 4388 32920
rect 4388 32886 4456 32920
rect 4456 32886 4546 32920
rect 4546 32886 4614 32920
rect 4614 32886 4704 32920
rect 4704 32886 4772 32920
rect 4772 32886 4862 32920
rect 4862 32886 4930 32920
rect 4930 32886 5020 32920
rect 5020 32886 5088 32920
rect 5088 32886 5178 32920
rect 5178 32886 5246 32920
rect 5246 32886 5336 32920
rect 5336 32886 5404 32920
rect 5404 32886 5494 32920
rect 5494 32886 5562 32920
rect 5562 32886 5652 32920
rect 5652 32886 5720 32920
rect 5720 32886 5810 32920
rect 5810 32886 5878 32920
rect 5878 32886 5968 32920
rect 5968 32886 6036 32920
rect 6036 32886 6126 32920
rect 6126 32886 6186 32920
rect 1552 32826 6186 32886
rect 6340 32800 6410 32936
rect 6650 32910 6850 32980
rect 7150 32910 7350 32980
rect 150 32520 350 32590
rect 650 32520 850 32590
rect 6520 32650 6590 32850
rect 6910 32650 6980 32850
rect 7020 32650 7090 32850
rect 7410 32650 7480 32850
rect 7630 32936 7646 38980
rect 7646 32936 7684 38980
rect 7684 32936 7700 38980
rect 12640 38980 12710 39120
rect 7765 32978 7782 38938
rect 7782 32978 7816 38938
rect 7816 32978 7831 38938
rect 7923 32978 7940 38938
rect 7940 32978 7974 38938
rect 7974 32978 7989 38938
rect 8081 32978 8098 38938
rect 8098 32978 8132 38938
rect 8132 32978 8147 38938
rect 8239 32978 8256 38938
rect 8256 32978 8290 38938
rect 8290 32978 8305 38938
rect 8397 32978 8414 38938
rect 8414 32978 8448 38938
rect 8448 32978 8463 38938
rect 8555 32978 8572 38938
rect 8572 32978 8606 38938
rect 8606 32978 8621 38938
rect 8713 32978 8730 38938
rect 8730 32978 8764 38938
rect 8764 32978 8779 38938
rect 8871 32978 8888 38938
rect 8888 32978 8922 38938
rect 8922 32978 8937 38938
rect 9029 32978 9046 38938
rect 9046 32978 9080 38938
rect 9080 32978 9095 38938
rect 9187 32978 9204 38938
rect 9204 32978 9238 38938
rect 9238 32978 9253 38938
rect 9345 32978 9362 38938
rect 9362 32978 9396 38938
rect 9396 32978 9411 38938
rect 9503 32978 9520 38938
rect 9520 32978 9554 38938
rect 9554 32978 9569 38938
rect 9661 32978 9678 38938
rect 9678 32978 9712 38938
rect 9712 32978 9727 38938
rect 9819 32978 9836 38938
rect 9836 32978 9870 38938
rect 9870 32978 9885 38938
rect 9977 32978 9994 38938
rect 9994 32978 10028 38938
rect 10028 32978 10043 38938
rect 10135 32978 10152 38938
rect 10152 32978 10186 38938
rect 10186 32978 10201 38938
rect 10293 32978 10310 38938
rect 10310 32978 10344 38938
rect 10344 32978 10359 38938
rect 10451 32978 10468 38938
rect 10468 32978 10502 38938
rect 10502 32978 10517 38938
rect 10609 32978 10626 38938
rect 10626 32978 10660 38938
rect 10660 32978 10675 38938
rect 10767 32978 10784 38938
rect 10784 32978 10818 38938
rect 10818 32978 10833 38938
rect 10925 32978 10942 38938
rect 10942 32978 10976 38938
rect 10976 32978 10991 38938
rect 11083 32978 11100 38938
rect 11100 32978 11134 38938
rect 11134 32978 11149 38938
rect 11241 32978 11258 38938
rect 11258 32978 11292 38938
rect 11292 32978 11307 38938
rect 11399 32978 11416 38938
rect 11416 32978 11450 38938
rect 11450 32978 11465 38938
rect 11557 32978 11574 38938
rect 11574 32978 11608 38938
rect 11608 32978 11623 38938
rect 11715 32978 11732 38938
rect 11732 32978 11766 38938
rect 11766 32978 11781 38938
rect 11873 32978 11890 38938
rect 11890 32978 11924 38938
rect 11924 32978 11939 38938
rect 12031 32978 12048 38938
rect 12048 32978 12082 38938
rect 12082 32978 12097 38938
rect 12189 32978 12206 38938
rect 12206 32978 12240 38938
rect 12240 32978 12255 38938
rect 12347 32978 12364 38938
rect 12364 32978 12398 38938
rect 12398 32978 12413 38938
rect 12505 32978 12522 38938
rect 12522 32978 12556 38938
rect 12556 32978 12571 38938
rect 7630 32800 7700 32936
rect 12640 32936 12654 38980
rect 12654 32936 12692 38980
rect 12692 32936 12710 38980
rect 13930 38980 14000 39120
rect 14152 39030 18786 39090
rect 14152 38996 14212 39030
rect 14212 38996 14302 39030
rect 14302 38996 14370 39030
rect 14370 38996 14460 39030
rect 14460 38996 14528 39030
rect 14528 38996 14618 39030
rect 14618 38996 14686 39030
rect 14686 38996 14776 39030
rect 14776 38996 14844 39030
rect 14844 38996 14934 39030
rect 14934 38996 15002 39030
rect 15002 38996 15092 39030
rect 15092 38996 15160 39030
rect 15160 38996 15250 39030
rect 15250 38996 15318 39030
rect 15318 38996 15408 39030
rect 15408 38996 15476 39030
rect 15476 38996 15566 39030
rect 15566 38996 15634 39030
rect 15634 38996 15724 39030
rect 15724 38996 15792 39030
rect 15792 38996 15882 39030
rect 15882 38996 15950 39030
rect 15950 38996 16040 39030
rect 16040 38996 16108 39030
rect 16108 38996 16198 39030
rect 16198 38996 16266 39030
rect 16266 38996 16356 39030
rect 16356 38996 16424 39030
rect 16424 38996 16514 39030
rect 16514 38996 16582 39030
rect 16582 38996 16672 39030
rect 16672 38996 16740 39030
rect 16740 38996 16830 39030
rect 16830 38996 16898 39030
rect 16898 38996 16988 39030
rect 16988 38996 17056 39030
rect 17056 38996 17146 39030
rect 17146 38996 17214 39030
rect 17214 38996 17304 39030
rect 17304 38996 17372 39030
rect 17372 38996 17462 39030
rect 17462 38996 17530 39030
rect 17530 38996 17620 39030
rect 17620 38996 17688 39030
rect 17688 38996 17778 39030
rect 17778 38996 17846 39030
rect 17846 38996 17936 39030
rect 17936 38996 18004 39030
rect 18004 38996 18094 39030
rect 18094 38996 18162 39030
rect 18162 38996 18252 39030
rect 18252 38996 18320 39030
rect 18320 38996 18410 39030
rect 18410 38996 18478 39030
rect 18478 38996 18568 39030
rect 18568 38996 18636 39030
rect 18636 38996 18726 39030
rect 18726 38996 18786 39030
rect 14152 38990 18786 38996
rect 7852 32920 12486 32926
rect 7852 32886 7912 32920
rect 7912 32886 8002 32920
rect 8002 32886 8070 32920
rect 8070 32886 8160 32920
rect 8160 32886 8228 32920
rect 8228 32886 8318 32920
rect 8318 32886 8386 32920
rect 8386 32886 8476 32920
rect 8476 32886 8544 32920
rect 8544 32886 8634 32920
rect 8634 32886 8702 32920
rect 8702 32886 8792 32920
rect 8792 32886 8860 32920
rect 8860 32886 8950 32920
rect 8950 32886 9018 32920
rect 9018 32886 9108 32920
rect 9108 32886 9176 32920
rect 9176 32886 9266 32920
rect 9266 32886 9334 32920
rect 9334 32886 9424 32920
rect 9424 32886 9492 32920
rect 9492 32886 9582 32920
rect 9582 32886 9650 32920
rect 9650 32886 9740 32920
rect 9740 32886 9808 32920
rect 9808 32886 9898 32920
rect 9898 32886 9966 32920
rect 9966 32886 10056 32920
rect 10056 32886 10124 32920
rect 10124 32886 10214 32920
rect 10214 32886 10282 32920
rect 10282 32886 10372 32920
rect 10372 32886 10440 32920
rect 10440 32886 10530 32920
rect 10530 32886 10598 32920
rect 10598 32886 10688 32920
rect 10688 32886 10756 32920
rect 10756 32886 10846 32920
rect 10846 32886 10914 32920
rect 10914 32886 11004 32920
rect 11004 32886 11072 32920
rect 11072 32886 11162 32920
rect 11162 32886 11230 32920
rect 11230 32886 11320 32920
rect 11320 32886 11388 32920
rect 11388 32886 11478 32920
rect 11478 32886 11546 32920
rect 11546 32886 11636 32920
rect 11636 32886 11704 32920
rect 11704 32886 11794 32920
rect 11794 32886 11862 32920
rect 11862 32886 11952 32920
rect 11952 32886 12020 32920
rect 12020 32886 12110 32920
rect 12110 32886 12178 32920
rect 12178 32886 12268 32920
rect 12268 32886 12336 32920
rect 12336 32886 12426 32920
rect 12426 32886 12486 32920
rect 7852 32826 12486 32886
rect 12640 32800 12710 32936
rect 13150 32910 13350 32980
rect 6650 32520 6850 32590
rect 7150 32520 7350 32590
rect 13020 32650 13090 32850
rect 13410 32650 13480 32850
rect 13930 32936 13946 38980
rect 13946 32936 13984 38980
rect 13984 32936 14000 38980
rect 18940 38980 19010 39120
rect 14065 32978 14082 38938
rect 14082 32978 14116 38938
rect 14116 32978 14131 38938
rect 14223 32978 14240 38938
rect 14240 32978 14274 38938
rect 14274 32978 14289 38938
rect 14381 32978 14398 38938
rect 14398 32978 14432 38938
rect 14432 32978 14447 38938
rect 14539 32978 14556 38938
rect 14556 32978 14590 38938
rect 14590 32978 14605 38938
rect 14697 32978 14714 38938
rect 14714 32978 14748 38938
rect 14748 32978 14763 38938
rect 14855 32978 14872 38938
rect 14872 32978 14906 38938
rect 14906 32978 14921 38938
rect 15013 32978 15030 38938
rect 15030 32978 15064 38938
rect 15064 32978 15079 38938
rect 15171 32978 15188 38938
rect 15188 32978 15222 38938
rect 15222 32978 15237 38938
rect 15329 32978 15346 38938
rect 15346 32978 15380 38938
rect 15380 32978 15395 38938
rect 15487 32978 15504 38938
rect 15504 32978 15538 38938
rect 15538 32978 15553 38938
rect 15645 32978 15662 38938
rect 15662 32978 15696 38938
rect 15696 32978 15711 38938
rect 15803 32978 15820 38938
rect 15820 32978 15854 38938
rect 15854 32978 15869 38938
rect 15961 32978 15978 38938
rect 15978 32978 16012 38938
rect 16012 32978 16027 38938
rect 16119 32978 16136 38938
rect 16136 32978 16170 38938
rect 16170 32978 16185 38938
rect 16277 32978 16294 38938
rect 16294 32978 16328 38938
rect 16328 32978 16343 38938
rect 16435 32978 16452 38938
rect 16452 32978 16486 38938
rect 16486 32978 16501 38938
rect 16593 32978 16610 38938
rect 16610 32978 16644 38938
rect 16644 32978 16659 38938
rect 16751 32978 16768 38938
rect 16768 32978 16802 38938
rect 16802 32978 16817 38938
rect 16909 32978 16926 38938
rect 16926 32978 16960 38938
rect 16960 32978 16975 38938
rect 17067 32978 17084 38938
rect 17084 32978 17118 38938
rect 17118 32978 17133 38938
rect 17225 32978 17242 38938
rect 17242 32978 17276 38938
rect 17276 32978 17291 38938
rect 17383 32978 17400 38938
rect 17400 32978 17434 38938
rect 17434 32978 17449 38938
rect 17541 32978 17558 38938
rect 17558 32978 17592 38938
rect 17592 32978 17607 38938
rect 17699 32978 17716 38938
rect 17716 32978 17750 38938
rect 17750 32978 17765 38938
rect 17857 32978 17874 38938
rect 17874 32978 17908 38938
rect 17908 32978 17923 38938
rect 18015 32978 18032 38938
rect 18032 32978 18066 38938
rect 18066 32978 18081 38938
rect 18173 32978 18190 38938
rect 18190 32978 18224 38938
rect 18224 32978 18239 38938
rect 18331 32978 18348 38938
rect 18348 32978 18382 38938
rect 18382 32978 18397 38938
rect 18489 32978 18506 38938
rect 18506 32978 18540 38938
rect 18540 32978 18555 38938
rect 18647 32978 18664 38938
rect 18664 32978 18698 38938
rect 18698 32978 18713 38938
rect 18805 32978 18822 38938
rect 18822 32978 18856 38938
rect 18856 32978 18871 38938
rect 13930 32800 14000 32936
rect 18940 32936 18954 38980
rect 18954 32936 18992 38980
rect 18992 32936 19010 38980
rect 25520 39150 25590 39350
rect 20230 38980 20300 39120
rect 25910 39150 25980 39350
rect 26020 39150 26090 39350
rect 26410 39150 26480 39350
rect 26520 39150 26590 39350
rect 26910 39150 26980 39350
rect 27020 39150 27090 39350
rect 27410 39150 27480 39350
rect 27520 39150 27590 39350
rect 27910 39150 27980 39350
rect 28020 39150 28090 39350
rect 28410 39150 28480 39350
rect 28520 39150 28590 39350
rect 28910 39150 28980 39350
rect 29020 39150 29090 39350
rect 29410 39150 29480 39350
rect 20452 39030 25086 39090
rect 20452 38996 20512 39030
rect 20512 38996 20602 39030
rect 20602 38996 20670 39030
rect 20670 38996 20760 39030
rect 20760 38996 20828 39030
rect 20828 38996 20918 39030
rect 20918 38996 20986 39030
rect 20986 38996 21076 39030
rect 21076 38996 21144 39030
rect 21144 38996 21234 39030
rect 21234 38996 21302 39030
rect 21302 38996 21392 39030
rect 21392 38996 21460 39030
rect 21460 38996 21550 39030
rect 21550 38996 21618 39030
rect 21618 38996 21708 39030
rect 21708 38996 21776 39030
rect 21776 38996 21866 39030
rect 21866 38996 21934 39030
rect 21934 38996 22024 39030
rect 22024 38996 22092 39030
rect 22092 38996 22182 39030
rect 22182 38996 22250 39030
rect 22250 38996 22340 39030
rect 22340 38996 22408 39030
rect 22408 38996 22498 39030
rect 22498 38996 22566 39030
rect 22566 38996 22656 39030
rect 22656 38996 22724 39030
rect 22724 38996 22814 39030
rect 22814 38996 22882 39030
rect 22882 38996 22972 39030
rect 22972 38996 23040 39030
rect 23040 38996 23130 39030
rect 23130 38996 23198 39030
rect 23198 38996 23288 39030
rect 23288 38996 23356 39030
rect 23356 38996 23446 39030
rect 23446 38996 23514 39030
rect 23514 38996 23604 39030
rect 23604 38996 23672 39030
rect 23672 38996 23762 39030
rect 23762 38996 23830 39030
rect 23830 38996 23920 39030
rect 23920 38996 23988 39030
rect 23988 38996 24078 39030
rect 24078 38996 24146 39030
rect 24146 38996 24236 39030
rect 24236 38996 24304 39030
rect 24304 38996 24394 39030
rect 24394 38996 24462 39030
rect 24462 38996 24552 39030
rect 24552 38996 24620 39030
rect 24620 38996 24710 39030
rect 24710 38996 24778 39030
rect 24778 38996 24868 39030
rect 24868 38996 24936 39030
rect 24936 38996 25026 39030
rect 25026 38996 25086 39030
rect 20452 38990 25086 38996
rect 14152 32920 18786 32926
rect 14152 32886 14212 32920
rect 14212 32886 14302 32920
rect 14302 32886 14370 32920
rect 14370 32886 14460 32920
rect 14460 32886 14528 32920
rect 14528 32886 14618 32920
rect 14618 32886 14686 32920
rect 14686 32886 14776 32920
rect 14776 32886 14844 32920
rect 14844 32886 14934 32920
rect 14934 32886 15002 32920
rect 15002 32886 15092 32920
rect 15092 32886 15160 32920
rect 15160 32886 15250 32920
rect 15250 32886 15318 32920
rect 15318 32886 15408 32920
rect 15408 32886 15476 32920
rect 15476 32886 15566 32920
rect 15566 32886 15634 32920
rect 15634 32886 15724 32920
rect 15724 32886 15792 32920
rect 15792 32886 15882 32920
rect 15882 32886 15950 32920
rect 15950 32886 16040 32920
rect 16040 32886 16108 32920
rect 16108 32886 16198 32920
rect 16198 32886 16266 32920
rect 16266 32886 16356 32920
rect 16356 32886 16424 32920
rect 16424 32886 16514 32920
rect 16514 32886 16582 32920
rect 16582 32886 16672 32920
rect 16672 32886 16740 32920
rect 16740 32886 16830 32920
rect 16830 32886 16898 32920
rect 16898 32886 16988 32920
rect 16988 32886 17056 32920
rect 17056 32886 17146 32920
rect 17146 32886 17214 32920
rect 17214 32886 17304 32920
rect 17304 32886 17372 32920
rect 17372 32886 17462 32920
rect 17462 32886 17530 32920
rect 17530 32886 17620 32920
rect 17620 32886 17688 32920
rect 17688 32886 17778 32920
rect 17778 32886 17846 32920
rect 17846 32886 17936 32920
rect 17936 32886 18004 32920
rect 18004 32886 18094 32920
rect 18094 32886 18162 32920
rect 18162 32886 18252 32920
rect 18252 32886 18320 32920
rect 18320 32886 18410 32920
rect 18410 32886 18478 32920
rect 18478 32886 18568 32920
rect 18568 32886 18636 32920
rect 18636 32886 18726 32920
rect 18726 32886 18786 32920
rect 14152 32826 18786 32886
rect 18940 32800 19010 32936
rect 19650 32910 19850 32980
rect 13150 32520 13350 32590
rect 19520 32650 19590 32850
rect 19910 32650 19980 32850
rect 20230 32936 20246 38980
rect 20246 32936 20284 38980
rect 20284 32936 20300 38980
rect 25240 38980 25310 39120
rect 25650 39020 25850 39090
rect 26150 39020 26350 39090
rect 26650 39020 26850 39090
rect 27150 39020 27350 39090
rect 27650 39020 27850 39090
rect 28150 39020 28350 39090
rect 28650 39020 28850 39090
rect 29150 39020 29350 39090
rect 20365 32978 20382 38938
rect 20382 32978 20416 38938
rect 20416 32978 20431 38938
rect 20523 32978 20540 38938
rect 20540 32978 20574 38938
rect 20574 32978 20589 38938
rect 20681 32978 20698 38938
rect 20698 32978 20732 38938
rect 20732 32978 20747 38938
rect 20839 32978 20856 38938
rect 20856 32978 20890 38938
rect 20890 32978 20905 38938
rect 20997 32978 21014 38938
rect 21014 32978 21048 38938
rect 21048 32978 21063 38938
rect 21155 32978 21172 38938
rect 21172 32978 21206 38938
rect 21206 32978 21221 38938
rect 21313 32978 21330 38938
rect 21330 32978 21364 38938
rect 21364 32978 21379 38938
rect 21471 32978 21488 38938
rect 21488 32978 21522 38938
rect 21522 32978 21537 38938
rect 21629 32978 21646 38938
rect 21646 32978 21680 38938
rect 21680 32978 21695 38938
rect 21787 32978 21804 38938
rect 21804 32978 21838 38938
rect 21838 32978 21853 38938
rect 21945 32978 21962 38938
rect 21962 32978 21996 38938
rect 21996 32978 22011 38938
rect 22103 32978 22120 38938
rect 22120 32978 22154 38938
rect 22154 32978 22169 38938
rect 22261 32978 22278 38938
rect 22278 32978 22312 38938
rect 22312 32978 22327 38938
rect 22419 32978 22436 38938
rect 22436 32978 22470 38938
rect 22470 32978 22485 38938
rect 22577 32978 22594 38938
rect 22594 32978 22628 38938
rect 22628 32978 22643 38938
rect 22735 32978 22752 38938
rect 22752 32978 22786 38938
rect 22786 32978 22801 38938
rect 22893 32978 22910 38938
rect 22910 32978 22944 38938
rect 22944 32978 22959 38938
rect 23051 32978 23068 38938
rect 23068 32978 23102 38938
rect 23102 32978 23117 38938
rect 23209 32978 23226 38938
rect 23226 32978 23260 38938
rect 23260 32978 23275 38938
rect 23367 32978 23384 38938
rect 23384 32978 23418 38938
rect 23418 32978 23433 38938
rect 23525 32978 23542 38938
rect 23542 32978 23576 38938
rect 23576 32978 23591 38938
rect 23683 32978 23700 38938
rect 23700 32978 23734 38938
rect 23734 32978 23749 38938
rect 23841 32978 23858 38938
rect 23858 32978 23892 38938
rect 23892 32978 23907 38938
rect 23999 32978 24016 38938
rect 24016 32978 24050 38938
rect 24050 32978 24065 38938
rect 24157 32978 24174 38938
rect 24174 32978 24208 38938
rect 24208 32978 24223 38938
rect 24315 32978 24332 38938
rect 24332 32978 24366 38938
rect 24366 32978 24381 38938
rect 24473 32978 24490 38938
rect 24490 32978 24524 38938
rect 24524 32978 24539 38938
rect 24631 32978 24648 38938
rect 24648 32978 24682 38938
rect 24682 32978 24697 38938
rect 24789 32978 24806 38938
rect 24806 32978 24840 38938
rect 24840 32978 24855 38938
rect 24947 32978 24964 38938
rect 24964 32978 24998 38938
rect 24998 32978 25013 38938
rect 25105 32978 25122 38938
rect 25122 32978 25156 38938
rect 25156 32978 25171 38938
rect 20230 32800 20300 32936
rect 25240 32936 25254 38980
rect 25254 32936 25292 38980
rect 25292 32936 25310 38980
rect 25650 38910 25850 38980
rect 26150 38910 26350 38980
rect 25520 38650 25590 38850
rect 25910 38650 25980 38850
rect 26020 38650 26090 38850
rect 26410 38650 26480 38850
rect 29910 40276 30090 40450
rect 29910 40236 29984 40276
rect 29984 40236 30018 40276
rect 30018 40236 30090 40276
rect 29910 40190 30090 40236
rect 29910 38902 30090 38910
rect 29910 38862 29984 38902
rect 29984 38862 30018 38902
rect 30018 38862 30090 38902
rect 29910 38690 30090 38862
rect 25650 38520 25850 38590
rect 26150 38520 26350 38590
rect 25650 38410 25850 38480
rect 26150 38410 26350 38480
rect 25520 38150 25590 38350
rect 25910 38150 25980 38350
rect 26020 38150 26090 38350
rect 26410 38150 26480 38350
rect 25650 38020 25850 38090
rect 26150 38020 26350 38090
rect 25650 37910 25850 37980
rect 26150 37910 26350 37980
rect 25520 37650 25590 37850
rect 25910 37650 25980 37850
rect 26020 37650 26090 37850
rect 26410 37650 26480 37850
rect 25650 37520 25850 37590
rect 26150 37520 26350 37590
rect 25650 37410 25850 37480
rect 26150 37410 26350 37480
rect 25520 37150 25590 37350
rect 25910 37150 25980 37350
rect 26020 37150 26090 37350
rect 26410 37150 26480 37350
rect 25650 37020 25850 37090
rect 26150 37020 26350 37090
rect 25650 36910 25850 36980
rect 26150 36910 26350 36980
rect 25520 36650 25590 36850
rect 25910 36650 25980 36850
rect 26020 36650 26090 36850
rect 26410 36650 26480 36850
rect 25650 36520 25850 36590
rect 26150 36520 26350 36590
rect 25650 36410 25850 36480
rect 26150 36410 26350 36480
rect 25520 36150 25590 36350
rect 25910 36150 25980 36350
rect 26020 36150 26090 36350
rect 26410 36150 26480 36350
rect 25650 36020 25850 36090
rect 26150 36020 26350 36090
rect 25650 35910 25850 35980
rect 26150 35910 26350 35980
rect 25520 35650 25590 35850
rect 25910 35650 25980 35850
rect 26020 35650 26090 35850
rect 26410 35650 26480 35850
rect 25650 35520 25850 35590
rect 26150 35520 26350 35590
rect 25650 35410 25850 35480
rect 26150 35410 26350 35480
rect 25520 35150 25590 35350
rect 25910 35150 25980 35350
rect 26020 35150 26090 35350
rect 26410 35150 26480 35350
rect 25650 35020 25850 35090
rect 26150 35020 26350 35090
rect 25650 34910 25850 34980
rect 26150 34910 26350 34980
rect 25520 34650 25590 34850
rect 25910 34650 25980 34850
rect 26020 34650 26090 34850
rect 26410 34650 26480 34850
rect 25650 34520 25850 34590
rect 26150 34520 26350 34590
rect 25650 34410 25850 34480
rect 26150 34410 26350 34480
rect 25520 34150 25590 34350
rect 25910 34150 25980 34350
rect 26020 34150 26090 34350
rect 26410 34150 26480 34350
rect 25650 34020 25850 34090
rect 26150 34020 26350 34090
rect 25650 33910 25850 33980
rect 26150 33910 26350 33980
rect 25520 33650 25590 33850
rect 25910 33650 25980 33850
rect 26020 33650 26090 33850
rect 26410 33650 26480 33850
rect 25650 33520 25850 33590
rect 26150 33520 26350 33590
rect 25650 33410 25850 33480
rect 26150 33410 26350 33480
rect 25520 33150 25590 33350
rect 25910 33150 25980 33350
rect 26020 33150 26090 33350
rect 26410 33150 26480 33350
rect 25650 33020 25850 33090
rect 26150 33020 26350 33090
rect 20452 32920 25086 32926
rect 20452 32886 20512 32920
rect 20512 32886 20602 32920
rect 20602 32886 20670 32920
rect 20670 32886 20760 32920
rect 20760 32886 20828 32920
rect 20828 32886 20918 32920
rect 20918 32886 20986 32920
rect 20986 32886 21076 32920
rect 21076 32886 21144 32920
rect 21144 32886 21234 32920
rect 21234 32886 21302 32920
rect 21302 32886 21392 32920
rect 21392 32886 21460 32920
rect 21460 32886 21550 32920
rect 21550 32886 21618 32920
rect 21618 32886 21708 32920
rect 21708 32886 21776 32920
rect 21776 32886 21866 32920
rect 21866 32886 21934 32920
rect 21934 32886 22024 32920
rect 22024 32886 22092 32920
rect 22092 32886 22182 32920
rect 22182 32886 22250 32920
rect 22250 32886 22340 32920
rect 22340 32886 22408 32920
rect 22408 32886 22498 32920
rect 22498 32886 22566 32920
rect 22566 32886 22656 32920
rect 22656 32886 22724 32920
rect 22724 32886 22814 32920
rect 22814 32886 22882 32920
rect 22882 32886 22972 32920
rect 22972 32886 23040 32920
rect 23040 32886 23130 32920
rect 23130 32886 23198 32920
rect 23198 32886 23288 32920
rect 23288 32886 23356 32920
rect 23356 32886 23446 32920
rect 23446 32886 23514 32920
rect 23514 32886 23604 32920
rect 23604 32886 23672 32920
rect 23672 32886 23762 32920
rect 23762 32886 23830 32920
rect 23830 32886 23920 32920
rect 23920 32886 23988 32920
rect 23988 32886 24078 32920
rect 24078 32886 24146 32920
rect 24146 32886 24236 32920
rect 24236 32886 24304 32920
rect 24304 32886 24394 32920
rect 24394 32886 24462 32920
rect 24462 32886 24552 32920
rect 24552 32886 24620 32920
rect 24620 32886 24710 32920
rect 24710 32886 24778 32920
rect 24778 32886 24868 32920
rect 24868 32886 24936 32920
rect 24936 32886 25026 32920
rect 25026 32886 25086 32920
rect 20452 32826 25086 32886
rect 25240 32800 25310 32936
rect 25650 32910 25850 32980
rect 26150 32910 26350 32980
rect 19650 32520 19850 32590
rect 25520 32650 25590 32850
rect 25910 32650 25980 32850
rect 26020 32650 26090 32850
rect 26410 32650 26480 32850
rect 25650 32520 25850 32590
rect 26150 32520 26350 32590
rect 150 32410 350 32480
rect 650 32410 850 32480
rect 1150 32410 1350 32480
rect 1650 32410 1850 32480
rect 2150 32410 2350 32480
rect 2650 32410 2850 32480
rect 3150 32410 3350 32480
rect 3650 32410 3850 32480
rect 4150 32410 4350 32480
rect 4650 32410 4850 32480
rect 5150 32410 5350 32480
rect 5650 32410 5850 32480
rect 6150 32410 6350 32480
rect 6650 32410 6850 32480
rect 7150 32410 7350 32480
rect 7650 32410 7850 32480
rect 8150 32410 8350 32480
rect 8650 32410 8850 32480
rect 9150 32410 9350 32480
rect 9650 32410 9850 32480
rect 10150 32410 10350 32480
rect 10650 32410 10850 32480
rect 11150 32410 11350 32480
rect 11650 32410 11850 32480
rect 12150 32410 12350 32480
rect 12650 32410 12850 32480
rect 13150 32410 13350 32480
rect 13650 32410 13850 32480
rect 14150 32410 14350 32480
rect 14650 32410 14850 32480
rect 15150 32410 15350 32480
rect 15650 32410 15850 32480
rect 16150 32410 16350 32480
rect 16650 32410 16850 32480
rect 17150 32410 17350 32480
rect 17650 32410 17850 32480
rect 18150 32410 18350 32480
rect 18650 32410 18850 32480
rect 19150 32410 19350 32480
rect 19650 32410 19850 32480
rect 20150 32410 20350 32480
rect 20650 32410 20850 32480
rect 21150 32410 21350 32480
rect 21650 32410 21850 32480
rect 22150 32410 22350 32480
rect 22650 32410 22850 32480
rect 23150 32410 23350 32480
rect 23650 32410 23850 32480
rect 24150 32410 24350 32480
rect 24650 32410 24850 32480
rect 25150 32410 25350 32480
rect 25650 32410 25850 32480
rect 26150 32410 26350 32480
rect 20 32150 90 32350
rect 410 32150 480 32350
rect 520 32150 590 32350
rect 910 32150 980 32350
rect 1020 32150 1090 32350
rect 1410 32150 1480 32350
rect 1520 32150 1590 32350
rect 1910 32150 1980 32350
rect 2020 32150 2090 32350
rect 2410 32150 2480 32350
rect 2520 32150 2590 32350
rect 2910 32150 2980 32350
rect 3020 32150 3090 32350
rect 3410 32150 3480 32350
rect 3520 32150 3590 32350
rect 3910 32150 3980 32350
rect 4020 32150 4090 32350
rect 4410 32150 4480 32350
rect 4520 32150 4590 32350
rect 4910 32150 4980 32350
rect 5020 32150 5090 32350
rect 5410 32150 5480 32350
rect 5520 32150 5590 32350
rect 5910 32150 5980 32350
rect 6020 32150 6090 32350
rect 6410 32150 6480 32350
rect 6520 32150 6590 32350
rect 6910 32150 6980 32350
rect 7020 32150 7090 32350
rect 7410 32150 7480 32350
rect 7520 32150 7590 32350
rect 7910 32150 7980 32350
rect 8020 32150 8090 32350
rect 8410 32150 8480 32350
rect 8520 32150 8590 32350
rect 8910 32150 8980 32350
rect 9020 32150 9090 32350
rect 9410 32150 9480 32350
rect 9520 32150 9590 32350
rect 9910 32150 9980 32350
rect 10020 32150 10090 32350
rect 10410 32150 10480 32350
rect 10520 32150 10590 32350
rect 10910 32150 10980 32350
rect 11020 32150 11090 32350
rect 11410 32150 11480 32350
rect 11520 32150 11590 32350
rect 11910 32150 11980 32350
rect 12020 32150 12090 32350
rect 12410 32150 12480 32350
rect 12520 32150 12590 32350
rect 12910 32150 12980 32350
rect 13020 32150 13090 32350
rect 13410 32150 13480 32350
rect 13520 32150 13590 32350
rect 13910 32150 13980 32350
rect 14020 32150 14090 32350
rect 14410 32150 14480 32350
rect 14520 32150 14590 32350
rect 14910 32150 14980 32350
rect 15020 32150 15090 32350
rect 15410 32150 15480 32350
rect 15520 32150 15590 32350
rect 15910 32150 15980 32350
rect 16020 32150 16090 32350
rect 16410 32150 16480 32350
rect 16520 32150 16590 32350
rect 16910 32150 16980 32350
rect 17020 32150 17090 32350
rect 17410 32150 17480 32350
rect 17520 32150 17590 32350
rect 17910 32150 17980 32350
rect 18020 32150 18090 32350
rect 18410 32150 18480 32350
rect 18520 32150 18590 32350
rect 18910 32150 18980 32350
rect 19020 32150 19090 32350
rect 19410 32150 19480 32350
rect 19520 32150 19590 32350
rect 19910 32150 19980 32350
rect 20020 32150 20090 32350
rect 20410 32150 20480 32350
rect 20520 32150 20590 32350
rect 20910 32150 20980 32350
rect 21020 32150 21090 32350
rect 21410 32150 21480 32350
rect 21520 32150 21590 32350
rect 21910 32150 21980 32350
rect 22020 32150 22090 32350
rect 22410 32150 22480 32350
rect 22520 32150 22590 32350
rect 22910 32150 22980 32350
rect 23020 32150 23090 32350
rect 23410 32150 23480 32350
rect 23520 32150 23590 32350
rect 23910 32150 23980 32350
rect 24020 32150 24090 32350
rect 24410 32150 24480 32350
rect 24520 32150 24590 32350
rect 24910 32150 24980 32350
rect 25020 32150 25090 32350
rect 25410 32150 25480 32350
rect 25520 32150 25590 32350
rect 25910 32150 25980 32350
rect 26020 32150 26090 32350
rect 26410 32150 26480 32350
rect 150 32020 350 32090
rect 650 32020 850 32090
rect 1150 32020 1350 32090
rect 1650 32020 1850 32090
rect 2150 32020 2350 32090
rect 2650 32020 2850 32090
rect 3150 32020 3350 32090
rect 3650 32020 3850 32090
rect 4150 32020 4350 32090
rect 4650 32020 4850 32090
rect 5150 32020 5350 32090
rect 5650 32020 5850 32090
rect 6150 32020 6350 32090
rect 6650 32020 6850 32090
rect 7150 32020 7350 32090
rect 7650 32020 7850 32090
rect 8150 32020 8350 32090
rect 8650 32020 8850 32090
rect 9150 32020 9350 32090
rect 9650 32020 9850 32090
rect 10150 32020 10350 32090
rect 10650 32020 10850 32090
rect 11150 32020 11350 32090
rect 11650 32020 11850 32090
rect 12150 32020 12350 32090
rect 12650 32020 12850 32090
rect 13150 32020 13350 32090
rect 13650 32020 13850 32090
rect 14150 32020 14350 32090
rect 14650 32020 14850 32090
rect 15150 32020 15350 32090
rect 15650 32020 15850 32090
rect 16150 32020 16350 32090
rect 16650 32020 16850 32090
rect 17150 32020 17350 32090
rect 17650 32020 17850 32090
rect 18150 32020 18350 32090
rect 18650 32020 18850 32090
rect 19150 32020 19350 32090
rect 19650 32020 19850 32090
rect 20150 32020 20350 32090
rect 20650 32020 20850 32090
rect 21150 32020 21350 32090
rect 21650 32020 21850 32090
rect 22150 32020 22350 32090
rect 22650 32020 22850 32090
rect 23150 32020 23350 32090
rect 23650 32020 23850 32090
rect 24150 32020 24350 32090
rect 24650 32020 24850 32090
rect 25150 32020 25350 32090
rect 25650 32020 25850 32090
rect 26150 32020 26350 32090
rect 150 31910 350 31980
rect 650 31910 850 31980
rect 1150 31910 1350 31980
rect 1650 31910 1850 31980
rect 2150 31910 2350 31980
rect 2650 31910 2850 31980
rect 3150 31910 3350 31980
rect 3650 31910 3850 31980
rect 4150 31910 4350 31980
rect 4650 31910 4850 31980
rect 5150 31910 5350 31980
rect 5650 31910 5850 31980
rect 6150 31910 6350 31980
rect 6650 31910 6850 31980
rect 7150 31910 7350 31980
rect 7650 31910 7850 31980
rect 8150 31910 8350 31980
rect 8650 31910 8850 31980
rect 9150 31910 9350 31980
rect 9650 31910 9850 31980
rect 10150 31910 10350 31980
rect 10650 31910 10850 31980
rect 11150 31910 11350 31980
rect 11650 31910 11850 31980
rect 12150 31910 12350 31980
rect 12650 31910 12850 31980
rect 13150 31910 13350 31980
rect 13650 31910 13850 31980
rect 14150 31910 14350 31980
rect 14650 31910 14850 31980
rect 15150 31910 15350 31980
rect 15650 31910 15850 31980
rect 16150 31910 16350 31980
rect 16650 31910 16850 31980
rect 17150 31910 17350 31980
rect 17650 31910 17850 31980
rect 18150 31910 18350 31980
rect 18650 31910 18850 31980
rect 19150 31910 19350 31980
rect 19650 31910 19850 31980
rect 20150 31910 20350 31980
rect 20650 31910 20850 31980
rect 21150 31910 21350 31980
rect 21650 31910 21850 31980
rect 22150 31910 22350 31980
rect 22650 31910 22850 31980
rect 23150 31910 23350 31980
rect 23650 31910 23850 31980
rect 24150 31910 24350 31980
rect 24650 31910 24850 31980
rect 25150 31910 25350 31980
rect 25650 31910 25850 31980
rect 26150 31910 26350 31980
rect 20 31650 90 31850
rect 410 31650 480 31850
rect 520 31650 590 31850
rect 910 31650 980 31850
rect 1020 31650 1090 31850
rect 1410 31650 1480 31850
rect 1520 31650 1590 31850
rect 1910 31650 1980 31850
rect 2020 31650 2090 31850
rect 2410 31650 2480 31850
rect 2520 31650 2590 31850
rect 2910 31650 2980 31850
rect 3020 31650 3090 31850
rect 3410 31650 3480 31850
rect 3520 31650 3590 31850
rect 3910 31650 3980 31850
rect 4020 31650 4090 31850
rect 4410 31650 4480 31850
rect 4520 31650 4590 31850
rect 4910 31650 4980 31850
rect 5020 31650 5090 31850
rect 5410 31650 5480 31850
rect 5520 31650 5590 31850
rect 5910 31650 5980 31850
rect 6020 31650 6090 31850
rect 6410 31650 6480 31850
rect 6520 31650 6590 31850
rect 6910 31650 6980 31850
rect 7020 31650 7090 31850
rect 7410 31650 7480 31850
rect 7520 31650 7590 31850
rect 7910 31650 7980 31850
rect 8020 31650 8090 31850
rect 8410 31650 8480 31850
rect 8520 31650 8590 31850
rect 8910 31650 8980 31850
rect 9020 31650 9090 31850
rect 9410 31650 9480 31850
rect 9520 31650 9590 31850
rect 9910 31650 9980 31850
rect 10020 31650 10090 31850
rect 10410 31650 10480 31850
rect 10520 31650 10590 31850
rect 10910 31650 10980 31850
rect 11020 31650 11090 31850
rect 11410 31650 11480 31850
rect 11520 31650 11590 31850
rect 11910 31650 11980 31850
rect 12020 31650 12090 31850
rect 12410 31650 12480 31850
rect 12520 31650 12590 31850
rect 12910 31650 12980 31850
rect 13020 31650 13090 31850
rect 13410 31650 13480 31850
rect 13520 31650 13590 31850
rect 13910 31650 13980 31850
rect 14020 31650 14090 31850
rect 14410 31650 14480 31850
rect 14520 31650 14590 31850
rect 14910 31650 14980 31850
rect 15020 31650 15090 31850
rect 15410 31650 15480 31850
rect 15520 31650 15590 31850
rect 15910 31650 15980 31850
rect 16020 31650 16090 31850
rect 16410 31650 16480 31850
rect 16520 31650 16590 31850
rect 16910 31650 16980 31850
rect 17020 31650 17090 31850
rect 17410 31650 17480 31850
rect 17520 31650 17590 31850
rect 17910 31650 17980 31850
rect 18020 31650 18090 31850
rect 18410 31650 18480 31850
rect 18520 31650 18590 31850
rect 18910 31650 18980 31850
rect 19020 31650 19090 31850
rect 19410 31650 19480 31850
rect 19520 31650 19590 31850
rect 19910 31650 19980 31850
rect 20020 31650 20090 31850
rect 20410 31650 20480 31850
rect 20520 31650 20590 31850
rect 20910 31650 20980 31850
rect 21020 31650 21090 31850
rect 21410 31650 21480 31850
rect 21520 31650 21590 31850
rect 21910 31650 21980 31850
rect 22020 31650 22090 31850
rect 22410 31650 22480 31850
rect 22520 31650 22590 31850
rect 22910 31650 22980 31850
rect 23020 31650 23090 31850
rect 23410 31650 23480 31850
rect 23520 31650 23590 31850
rect 23910 31650 23980 31850
rect 24020 31650 24090 31850
rect 24410 31650 24480 31850
rect 24520 31650 24590 31850
rect 24910 31650 24980 31850
rect 25020 31650 25090 31850
rect 25410 31650 25480 31850
rect 25520 31650 25590 31850
rect 25910 31650 25980 31850
rect 26020 31650 26090 31850
rect 26410 31650 26480 31850
rect 150 31520 350 31590
rect 650 31520 850 31590
rect 1150 31520 1350 31590
rect 1650 31520 1850 31590
rect 2150 31520 2350 31590
rect 2650 31520 2850 31590
rect 3150 31520 3350 31590
rect 3650 31520 3850 31590
rect 4150 31520 4350 31590
rect 4650 31520 4850 31590
rect 5150 31520 5350 31590
rect 5650 31520 5850 31590
rect 6150 31520 6350 31590
rect 6650 31520 6850 31590
rect 7150 31520 7350 31590
rect 7650 31520 7850 31590
rect 8150 31520 8350 31590
rect 8650 31520 8850 31590
rect 9150 31520 9350 31590
rect 9650 31520 9850 31590
rect 10150 31520 10350 31590
rect 10650 31520 10850 31590
rect 11150 31520 11350 31590
rect 11650 31520 11850 31590
rect 12150 31520 12350 31590
rect 12650 31520 12850 31590
rect 13150 31520 13350 31590
rect 13650 31520 13850 31590
rect 14150 31520 14350 31590
rect 14650 31520 14850 31590
rect 15150 31520 15350 31590
rect 15650 31520 15850 31590
rect 16150 31520 16350 31590
rect 16650 31520 16850 31590
rect 17150 31520 17350 31590
rect 17650 31520 17850 31590
rect 18150 31520 18350 31590
rect 18650 31520 18850 31590
rect 19150 31520 19350 31590
rect 19650 31520 19850 31590
rect 20150 31520 20350 31590
rect 20650 31520 20850 31590
rect 21150 31520 21350 31590
rect 21650 31520 21850 31590
rect 22150 31520 22350 31590
rect 22650 31520 22850 31590
rect 23150 31520 23350 31590
rect 23650 31520 23850 31590
rect 24150 31520 24350 31590
rect 24650 31520 24850 31590
rect 25150 31520 25350 31590
rect 25650 31520 25850 31590
rect 26150 31520 26350 31590
rect 150 31410 350 31480
rect 650 31410 850 31480
rect 20 31150 90 31350
rect 410 31150 480 31350
rect 520 31150 590 31350
rect 910 31150 980 31350
rect 150 31020 350 31090
rect 650 31020 850 31090
rect 150 30910 350 30980
rect 650 30910 850 30980
rect 6650 31410 6850 31480
rect 7150 31410 7350 31480
rect 6520 31150 6590 31350
rect 6910 31150 6980 31350
rect 7020 31150 7090 31350
rect 7410 31150 7480 31350
rect 6650 31020 6850 31090
rect 7150 31020 7350 31090
rect 13150 31410 13350 31480
rect 13020 31150 13090 31350
rect 13410 31150 13480 31350
rect 13150 31020 13350 31090
rect 19650 31410 19850 31480
rect 19520 31150 19590 31350
rect 19910 31150 19980 31350
rect 19650 31020 19850 31090
rect 6650 30910 6850 30980
rect 7150 30910 7350 30980
rect 19650 30910 19850 30980
rect 25650 31410 25850 31480
rect 26150 31410 26350 31480
rect 25520 31150 25590 31350
rect 25910 31150 25980 31350
rect 26020 31150 26090 31350
rect 26410 31150 26480 31350
rect 25650 31020 25850 31090
rect 26150 31020 26350 31090
rect 25650 30910 25850 30980
rect 26150 30910 26350 30980
rect 20 30650 90 30850
rect 410 30650 480 30850
rect 520 30650 590 30850
rect 910 30650 980 30850
rect 1330 30680 1400 30820
rect 1552 30730 6186 30790
rect 1552 30696 1612 30730
rect 1612 30696 1702 30730
rect 1702 30696 1770 30730
rect 1770 30696 1860 30730
rect 1860 30696 1928 30730
rect 1928 30696 2018 30730
rect 2018 30696 2086 30730
rect 2086 30696 2176 30730
rect 2176 30696 2244 30730
rect 2244 30696 2334 30730
rect 2334 30696 2402 30730
rect 2402 30696 2492 30730
rect 2492 30696 2560 30730
rect 2560 30696 2650 30730
rect 2650 30696 2718 30730
rect 2718 30696 2808 30730
rect 2808 30696 2876 30730
rect 2876 30696 2966 30730
rect 2966 30696 3034 30730
rect 3034 30696 3124 30730
rect 3124 30696 3192 30730
rect 3192 30696 3282 30730
rect 3282 30696 3350 30730
rect 3350 30696 3440 30730
rect 3440 30696 3508 30730
rect 3508 30696 3598 30730
rect 3598 30696 3666 30730
rect 3666 30696 3756 30730
rect 3756 30696 3824 30730
rect 3824 30696 3914 30730
rect 3914 30696 3982 30730
rect 3982 30696 4072 30730
rect 4072 30696 4140 30730
rect 4140 30696 4230 30730
rect 4230 30696 4298 30730
rect 4298 30696 4388 30730
rect 4388 30696 4456 30730
rect 4456 30696 4546 30730
rect 4546 30696 4614 30730
rect 4614 30696 4704 30730
rect 4704 30696 4772 30730
rect 4772 30696 4862 30730
rect 4862 30696 4930 30730
rect 4930 30696 5020 30730
rect 5020 30696 5088 30730
rect 5088 30696 5178 30730
rect 5178 30696 5246 30730
rect 5246 30696 5336 30730
rect 5336 30696 5404 30730
rect 5404 30696 5494 30730
rect 5494 30696 5562 30730
rect 5562 30696 5652 30730
rect 5652 30696 5720 30730
rect 5720 30696 5810 30730
rect 5810 30696 5878 30730
rect 5878 30696 5968 30730
rect 5968 30696 6036 30730
rect 6036 30696 6126 30730
rect 6126 30696 6186 30730
rect 1552 30690 6186 30696
rect 150 30520 350 30590
rect 650 30520 850 30590
rect 150 30410 350 30480
rect 650 30410 850 30480
rect 20 30150 90 30350
rect 410 30150 480 30350
rect 520 30150 590 30350
rect 910 30150 980 30350
rect 150 30020 350 30090
rect 650 30020 850 30090
rect 150 29910 350 29980
rect 650 29910 850 29980
rect 20 29650 90 29850
rect 410 29650 480 29850
rect 520 29650 590 29850
rect 910 29650 980 29850
rect 150 29520 350 29590
rect 650 29520 850 29590
rect 150 29410 350 29480
rect 650 29410 850 29480
rect 20 29150 90 29350
rect 410 29150 480 29350
rect 520 29150 590 29350
rect 910 29150 980 29350
rect 150 29020 350 29090
rect 650 29020 850 29090
rect 150 28910 350 28980
rect 650 28910 850 28980
rect 20 28650 90 28850
rect 410 28650 480 28850
rect 520 28650 590 28850
rect 910 28650 980 28850
rect 150 28520 350 28590
rect 650 28520 850 28590
rect 150 28410 350 28480
rect 650 28410 850 28480
rect 20 28150 90 28350
rect 410 28150 480 28350
rect 520 28150 590 28350
rect 910 28150 980 28350
rect 150 28020 350 28090
rect 650 28020 850 28090
rect 150 27910 350 27980
rect 650 27910 850 27980
rect 20 27650 90 27850
rect 410 27650 480 27850
rect 520 27650 590 27850
rect 910 27650 980 27850
rect 150 27520 350 27590
rect 650 27520 850 27590
rect 150 27410 350 27480
rect 650 27410 850 27480
rect -4290 27076 -4110 27250
rect -4290 27036 -4218 27076
rect -4218 27036 -4184 27076
rect -4184 27036 -4110 27076
rect -4290 27030 -4110 27036
rect -4290 25702 -4110 25710
rect -4290 25662 -4218 25702
rect -4218 25662 -4184 25702
rect -4184 25662 -4110 25702
rect -4290 25490 -4110 25662
rect 20 27150 90 27350
rect 410 27150 480 27350
rect 520 27150 590 27350
rect 910 27150 980 27350
rect 150 27020 350 27090
rect 650 27020 850 27090
rect -3850 26910 -3650 26980
rect -3350 26910 -3150 26980
rect -2850 26910 -2650 26980
rect -2350 26910 -2150 26980
rect -1850 26910 -1650 26980
rect -1350 26910 -1150 26980
rect -850 26910 -650 26980
rect -350 26910 -150 26980
rect 150 26910 350 26980
rect 650 26910 850 26980
rect -3980 26650 -3910 26850
rect -3590 26650 -3520 26850
rect -3480 26650 -3410 26850
rect -3090 26650 -3020 26850
rect -2980 26650 -2910 26850
rect -2590 26650 -2520 26850
rect -2480 26650 -2410 26850
rect -2090 26650 -2020 26850
rect -1980 26650 -1910 26850
rect -1590 26650 -1520 26850
rect -1480 26650 -1410 26850
rect -1090 26650 -1020 26850
rect -980 26650 -910 26850
rect -590 26650 -520 26850
rect -480 26650 -410 26850
rect -90 26650 -20 26850
rect 20 26650 90 26850
rect 410 26650 480 26850
rect 520 26650 590 26850
rect 910 26650 980 26850
rect -3850 26520 -3650 26590
rect -3350 26520 -3150 26590
rect -2850 26520 -2650 26590
rect -2350 26520 -2150 26590
rect -1850 26520 -1650 26590
rect -1350 26520 -1150 26590
rect -850 26520 -650 26590
rect -350 26520 -150 26590
rect 150 26520 350 26590
rect 650 26520 850 26590
rect -3850 26410 -3650 26480
rect -3350 26410 -3150 26480
rect -2850 26410 -2650 26480
rect -2350 26410 -2150 26480
rect -1850 26410 -1650 26480
rect -1350 26410 -1150 26480
rect -850 26410 -650 26480
rect -350 26410 -150 26480
rect 150 26410 350 26480
rect 650 26410 850 26480
rect -3980 26150 -3910 26350
rect -3590 26150 -3520 26350
rect -3480 26150 -3410 26350
rect -3090 26150 -3020 26350
rect -2980 26150 -2910 26350
rect -2590 26150 -2520 26350
rect -2480 26150 -2410 26350
rect -2090 26150 -2020 26350
rect -1980 26150 -1910 26350
rect -1590 26150 -1520 26350
rect -1480 26150 -1410 26350
rect -1090 26150 -1020 26350
rect -980 26150 -910 26350
rect -590 26150 -520 26350
rect -480 26150 -410 26350
rect -90 26150 -20 26350
rect 20 26150 90 26350
rect 410 26150 480 26350
rect 520 26150 590 26350
rect 910 26150 980 26350
rect -3850 26020 -3650 26090
rect -3350 26020 -3150 26090
rect -2850 26020 -2650 26090
rect -2350 26020 -2150 26090
rect -1850 26020 -1650 26090
rect -1350 26020 -1150 26090
rect -850 26020 -650 26090
rect -350 26020 -150 26090
rect 150 26020 350 26090
rect 650 26020 850 26090
rect 150 25910 350 25980
rect 650 25910 850 25980
rect 20 25650 90 25850
rect 410 25650 480 25850
rect 520 25650 590 25850
rect 910 25650 980 25850
rect 150 25520 350 25590
rect 650 25520 850 25590
rect 150 25410 350 25480
rect 650 25410 850 25480
rect 20 25150 90 25350
rect 410 25150 480 25350
rect 520 25150 590 25350
rect 910 25150 980 25350
rect 150 25020 350 25090
rect 650 25020 850 25090
rect 150 24910 350 24980
rect 650 24910 850 24980
rect 20 24650 90 24850
rect 410 24650 480 24850
rect 520 24650 590 24850
rect 910 24650 980 24850
rect 1330 24636 1346 30680
rect 1346 24636 1384 30680
rect 1384 24636 1400 30680
rect 6340 30680 6410 30820
rect 1465 24678 1482 30638
rect 1482 24678 1516 30638
rect 1516 24678 1531 30638
rect 1623 24678 1640 30638
rect 1640 24678 1674 30638
rect 1674 24678 1689 30638
rect 1781 24678 1798 30638
rect 1798 24678 1832 30638
rect 1832 24678 1847 30638
rect 1939 24678 1956 30638
rect 1956 24678 1990 30638
rect 1990 24678 2005 30638
rect 2097 24678 2114 30638
rect 2114 24678 2148 30638
rect 2148 24678 2163 30638
rect 2255 24678 2272 30638
rect 2272 24678 2306 30638
rect 2306 24678 2321 30638
rect 2413 24678 2430 30638
rect 2430 24678 2464 30638
rect 2464 24678 2479 30638
rect 2571 24678 2588 30638
rect 2588 24678 2622 30638
rect 2622 24678 2637 30638
rect 2729 24678 2746 30638
rect 2746 24678 2780 30638
rect 2780 24678 2795 30638
rect 2887 24678 2904 30638
rect 2904 24678 2938 30638
rect 2938 24678 2953 30638
rect 3045 24678 3062 30638
rect 3062 24678 3096 30638
rect 3096 24678 3111 30638
rect 3203 24678 3220 30638
rect 3220 24678 3254 30638
rect 3254 24678 3269 30638
rect 3361 24678 3378 30638
rect 3378 24678 3412 30638
rect 3412 24678 3427 30638
rect 3519 24678 3536 30638
rect 3536 24678 3570 30638
rect 3570 24678 3585 30638
rect 3677 24678 3694 30638
rect 3694 24678 3728 30638
rect 3728 24678 3743 30638
rect 3835 24678 3852 30638
rect 3852 24678 3886 30638
rect 3886 24678 3901 30638
rect 3993 24678 4010 30638
rect 4010 24678 4044 30638
rect 4044 24678 4059 30638
rect 4151 24678 4168 30638
rect 4168 24678 4202 30638
rect 4202 24678 4217 30638
rect 4309 24678 4326 30638
rect 4326 24678 4360 30638
rect 4360 24678 4375 30638
rect 4467 24678 4484 30638
rect 4484 24678 4518 30638
rect 4518 24678 4533 30638
rect 4625 24678 4642 30638
rect 4642 24678 4676 30638
rect 4676 24678 4691 30638
rect 4783 24678 4800 30638
rect 4800 24678 4834 30638
rect 4834 24678 4849 30638
rect 4941 24678 4958 30638
rect 4958 24678 4992 30638
rect 4992 24678 5007 30638
rect 5099 24678 5116 30638
rect 5116 24678 5150 30638
rect 5150 24678 5165 30638
rect 5257 24678 5274 30638
rect 5274 24678 5308 30638
rect 5308 24678 5323 30638
rect 5415 24678 5432 30638
rect 5432 24678 5466 30638
rect 5466 24678 5481 30638
rect 5573 24678 5590 30638
rect 5590 24678 5624 30638
rect 5624 24678 5639 30638
rect 5731 24678 5748 30638
rect 5748 24678 5782 30638
rect 5782 24678 5797 30638
rect 5889 24678 5906 30638
rect 5906 24678 5940 30638
rect 5940 24678 5955 30638
rect 6047 24678 6064 30638
rect 6064 24678 6098 30638
rect 6098 24678 6113 30638
rect 6205 24678 6222 30638
rect 6222 24678 6256 30638
rect 6256 24678 6271 30638
rect 150 24520 350 24590
rect 650 24520 850 24590
rect 1330 24500 1400 24636
rect 6340 24636 6354 30680
rect 6354 24636 6392 30680
rect 6392 24636 6410 30680
rect 6520 30650 6590 30850
rect 6910 30650 6980 30850
rect 7020 30650 7090 30850
rect 7410 30650 7480 30850
rect 6650 30520 6850 30590
rect 7150 30520 7350 30590
rect 7630 30680 7700 30820
rect 7852 30730 12486 30790
rect 7852 30696 7912 30730
rect 7912 30696 8002 30730
rect 8002 30696 8070 30730
rect 8070 30696 8160 30730
rect 8160 30696 8228 30730
rect 8228 30696 8318 30730
rect 8318 30696 8386 30730
rect 8386 30696 8476 30730
rect 8476 30696 8544 30730
rect 8544 30696 8634 30730
rect 8634 30696 8702 30730
rect 8702 30696 8792 30730
rect 8792 30696 8860 30730
rect 8860 30696 8950 30730
rect 8950 30696 9018 30730
rect 9018 30696 9108 30730
rect 9108 30696 9176 30730
rect 9176 30696 9266 30730
rect 9266 30696 9334 30730
rect 9334 30696 9424 30730
rect 9424 30696 9492 30730
rect 9492 30696 9582 30730
rect 9582 30696 9650 30730
rect 9650 30696 9740 30730
rect 9740 30696 9808 30730
rect 9808 30696 9898 30730
rect 9898 30696 9966 30730
rect 9966 30696 10056 30730
rect 10056 30696 10124 30730
rect 10124 30696 10214 30730
rect 10214 30696 10282 30730
rect 10282 30696 10372 30730
rect 10372 30696 10440 30730
rect 10440 30696 10530 30730
rect 10530 30696 10598 30730
rect 10598 30696 10688 30730
rect 10688 30696 10756 30730
rect 10756 30696 10846 30730
rect 10846 30696 10914 30730
rect 10914 30696 11004 30730
rect 11004 30696 11072 30730
rect 11072 30696 11162 30730
rect 11162 30696 11230 30730
rect 11230 30696 11320 30730
rect 11320 30696 11388 30730
rect 11388 30696 11478 30730
rect 11478 30696 11546 30730
rect 11546 30696 11636 30730
rect 11636 30696 11704 30730
rect 11704 30696 11794 30730
rect 11794 30696 11862 30730
rect 11862 30696 11952 30730
rect 11952 30696 12020 30730
rect 12020 30696 12110 30730
rect 12110 30696 12178 30730
rect 12178 30696 12268 30730
rect 12268 30696 12336 30730
rect 12336 30696 12426 30730
rect 12426 30696 12486 30730
rect 7852 30690 12486 30696
rect 1552 24620 6186 24626
rect 1552 24586 1612 24620
rect 1612 24586 1702 24620
rect 1702 24586 1770 24620
rect 1770 24586 1860 24620
rect 1860 24586 1928 24620
rect 1928 24586 2018 24620
rect 2018 24586 2086 24620
rect 2086 24586 2176 24620
rect 2176 24586 2244 24620
rect 2244 24586 2334 24620
rect 2334 24586 2402 24620
rect 2402 24586 2492 24620
rect 2492 24586 2560 24620
rect 2560 24586 2650 24620
rect 2650 24586 2718 24620
rect 2718 24586 2808 24620
rect 2808 24586 2876 24620
rect 2876 24586 2966 24620
rect 2966 24586 3034 24620
rect 3034 24586 3124 24620
rect 3124 24586 3192 24620
rect 3192 24586 3282 24620
rect 3282 24586 3350 24620
rect 3350 24586 3440 24620
rect 3440 24586 3508 24620
rect 3508 24586 3598 24620
rect 3598 24586 3666 24620
rect 3666 24586 3756 24620
rect 3756 24586 3824 24620
rect 3824 24586 3914 24620
rect 3914 24586 3982 24620
rect 3982 24586 4072 24620
rect 4072 24586 4140 24620
rect 4140 24586 4230 24620
rect 4230 24586 4298 24620
rect 4298 24586 4388 24620
rect 4388 24586 4456 24620
rect 4456 24586 4546 24620
rect 4546 24586 4614 24620
rect 4614 24586 4704 24620
rect 4704 24586 4772 24620
rect 4772 24586 4862 24620
rect 4862 24586 4930 24620
rect 4930 24586 5020 24620
rect 5020 24586 5088 24620
rect 5088 24586 5178 24620
rect 5178 24586 5246 24620
rect 5246 24586 5336 24620
rect 5336 24586 5404 24620
rect 5404 24586 5494 24620
rect 5494 24586 5562 24620
rect 5562 24586 5652 24620
rect 5652 24586 5720 24620
rect 5720 24586 5810 24620
rect 5810 24586 5878 24620
rect 5878 24586 5968 24620
rect 5968 24586 6036 24620
rect 6036 24586 6126 24620
rect 6126 24586 6186 24620
rect 1552 24526 6186 24586
rect 6340 24500 6410 24636
rect 150 24410 350 24480
rect 650 24410 850 24480
rect 7630 24636 7646 30680
rect 7646 24636 7684 30680
rect 7684 24636 7700 30680
rect 12640 30680 12710 30820
rect 7765 24678 7782 30638
rect 7782 24678 7816 30638
rect 7816 24678 7831 30638
rect 7923 24678 7940 30638
rect 7940 24678 7974 30638
rect 7974 24678 7989 30638
rect 8081 24678 8098 30638
rect 8098 24678 8132 30638
rect 8132 24678 8147 30638
rect 8239 24678 8256 30638
rect 8256 24678 8290 30638
rect 8290 24678 8305 30638
rect 8397 24678 8414 30638
rect 8414 24678 8448 30638
rect 8448 24678 8463 30638
rect 8555 24678 8572 30638
rect 8572 24678 8606 30638
rect 8606 24678 8621 30638
rect 8713 24678 8730 30638
rect 8730 24678 8764 30638
rect 8764 24678 8779 30638
rect 8871 24678 8888 30638
rect 8888 24678 8922 30638
rect 8922 24678 8937 30638
rect 9029 24678 9046 30638
rect 9046 24678 9080 30638
rect 9080 24678 9095 30638
rect 9187 24678 9204 30638
rect 9204 24678 9238 30638
rect 9238 24678 9253 30638
rect 9345 24678 9362 30638
rect 9362 24678 9396 30638
rect 9396 24678 9411 30638
rect 9503 24678 9520 30638
rect 9520 24678 9554 30638
rect 9554 24678 9569 30638
rect 9661 24678 9678 30638
rect 9678 24678 9712 30638
rect 9712 24678 9727 30638
rect 9819 24678 9836 30638
rect 9836 24678 9870 30638
rect 9870 24678 9885 30638
rect 9977 24678 9994 30638
rect 9994 24678 10028 30638
rect 10028 24678 10043 30638
rect 10135 24678 10152 30638
rect 10152 24678 10186 30638
rect 10186 24678 10201 30638
rect 10293 24678 10310 30638
rect 10310 24678 10344 30638
rect 10344 24678 10359 30638
rect 10451 24678 10468 30638
rect 10468 24678 10502 30638
rect 10502 24678 10517 30638
rect 10609 24678 10626 30638
rect 10626 24678 10660 30638
rect 10660 24678 10675 30638
rect 10767 24678 10784 30638
rect 10784 24678 10818 30638
rect 10818 24678 10833 30638
rect 10925 24678 10942 30638
rect 10942 24678 10976 30638
rect 10976 24678 10991 30638
rect 11083 24678 11100 30638
rect 11100 24678 11134 30638
rect 11134 24678 11149 30638
rect 11241 24678 11258 30638
rect 11258 24678 11292 30638
rect 11292 24678 11307 30638
rect 11399 24678 11416 30638
rect 11416 24678 11450 30638
rect 11450 24678 11465 30638
rect 11557 24678 11574 30638
rect 11574 24678 11608 30638
rect 11608 24678 11623 30638
rect 11715 24678 11732 30638
rect 11732 24678 11766 30638
rect 11766 24678 11781 30638
rect 11873 24678 11890 30638
rect 11890 24678 11924 30638
rect 11924 24678 11939 30638
rect 12031 24678 12048 30638
rect 12048 24678 12082 30638
rect 12082 24678 12097 30638
rect 12189 24678 12206 30638
rect 12206 24678 12240 30638
rect 12240 24678 12255 30638
rect 12347 24678 12364 30638
rect 12364 24678 12398 30638
rect 12398 24678 12413 30638
rect 12505 24678 12522 30638
rect 12522 24678 12556 30638
rect 12556 24678 12571 30638
rect 7630 24500 7700 24636
rect 12640 24636 12654 30680
rect 12654 24636 12692 30680
rect 12692 24636 12710 30680
rect 7852 24620 12486 24626
rect 7852 24586 7912 24620
rect 7912 24586 8002 24620
rect 8002 24586 8070 24620
rect 8070 24586 8160 24620
rect 8160 24586 8228 24620
rect 8228 24586 8318 24620
rect 8318 24586 8386 24620
rect 8386 24586 8476 24620
rect 8476 24586 8544 24620
rect 8544 24586 8634 24620
rect 8634 24586 8702 24620
rect 8702 24586 8792 24620
rect 8792 24586 8860 24620
rect 8860 24586 8950 24620
rect 8950 24586 9018 24620
rect 9018 24586 9108 24620
rect 9108 24586 9176 24620
rect 9176 24586 9266 24620
rect 9266 24586 9334 24620
rect 9334 24586 9424 24620
rect 9424 24586 9492 24620
rect 9492 24586 9582 24620
rect 9582 24586 9650 24620
rect 9650 24586 9740 24620
rect 9740 24586 9808 24620
rect 9808 24586 9898 24620
rect 9898 24586 9966 24620
rect 9966 24586 10056 24620
rect 10056 24586 10124 24620
rect 10124 24586 10214 24620
rect 10214 24586 10282 24620
rect 10282 24586 10372 24620
rect 10372 24586 10440 24620
rect 10440 24586 10530 24620
rect 10530 24586 10598 24620
rect 10598 24586 10688 24620
rect 10688 24586 10756 24620
rect 10756 24586 10846 24620
rect 10846 24586 10914 24620
rect 10914 24586 11004 24620
rect 11004 24586 11072 24620
rect 11072 24586 11162 24620
rect 11162 24586 11230 24620
rect 11230 24586 11320 24620
rect 11320 24586 11388 24620
rect 11388 24586 11478 24620
rect 11478 24586 11546 24620
rect 11546 24586 11636 24620
rect 11636 24586 11704 24620
rect 11704 24586 11794 24620
rect 11794 24586 11862 24620
rect 11862 24586 11952 24620
rect 11952 24586 12020 24620
rect 12020 24586 12110 24620
rect 12110 24586 12178 24620
rect 12178 24586 12268 24620
rect 12268 24586 12336 24620
rect 12336 24586 12426 24620
rect 12426 24586 12486 24620
rect 7852 24526 12486 24586
rect 12640 24500 12710 24636
rect 13930 30680 14000 30820
rect 14152 30730 18786 30790
rect 14152 30696 14212 30730
rect 14212 30696 14302 30730
rect 14302 30696 14370 30730
rect 14370 30696 14460 30730
rect 14460 30696 14528 30730
rect 14528 30696 14618 30730
rect 14618 30696 14686 30730
rect 14686 30696 14776 30730
rect 14776 30696 14844 30730
rect 14844 30696 14934 30730
rect 14934 30696 15002 30730
rect 15002 30696 15092 30730
rect 15092 30696 15160 30730
rect 15160 30696 15250 30730
rect 15250 30696 15318 30730
rect 15318 30696 15408 30730
rect 15408 30696 15476 30730
rect 15476 30696 15566 30730
rect 15566 30696 15634 30730
rect 15634 30696 15724 30730
rect 15724 30696 15792 30730
rect 15792 30696 15882 30730
rect 15882 30696 15950 30730
rect 15950 30696 16040 30730
rect 16040 30696 16108 30730
rect 16108 30696 16198 30730
rect 16198 30696 16266 30730
rect 16266 30696 16356 30730
rect 16356 30696 16424 30730
rect 16424 30696 16514 30730
rect 16514 30696 16582 30730
rect 16582 30696 16672 30730
rect 16672 30696 16740 30730
rect 16740 30696 16830 30730
rect 16830 30696 16898 30730
rect 16898 30696 16988 30730
rect 16988 30696 17056 30730
rect 17056 30696 17146 30730
rect 17146 30696 17214 30730
rect 17214 30696 17304 30730
rect 17304 30696 17372 30730
rect 17372 30696 17462 30730
rect 17462 30696 17530 30730
rect 17530 30696 17620 30730
rect 17620 30696 17688 30730
rect 17688 30696 17778 30730
rect 17778 30696 17846 30730
rect 17846 30696 17936 30730
rect 17936 30696 18004 30730
rect 18004 30696 18094 30730
rect 18094 30696 18162 30730
rect 18162 30696 18252 30730
rect 18252 30696 18320 30730
rect 18320 30696 18410 30730
rect 18410 30696 18478 30730
rect 18478 30696 18568 30730
rect 18568 30696 18636 30730
rect 18636 30696 18726 30730
rect 18726 30696 18786 30730
rect 14152 30690 18786 30696
rect 13930 24636 13946 30680
rect 13946 24636 13984 30680
rect 13984 24636 14000 30680
rect 18940 30680 19010 30820
rect 14065 24678 14082 30638
rect 14082 24678 14116 30638
rect 14116 24678 14131 30638
rect 14223 24678 14240 30638
rect 14240 24678 14274 30638
rect 14274 24678 14289 30638
rect 14381 24678 14398 30638
rect 14398 24678 14432 30638
rect 14432 24678 14447 30638
rect 14539 24678 14556 30638
rect 14556 24678 14590 30638
rect 14590 24678 14605 30638
rect 14697 24678 14714 30638
rect 14714 24678 14748 30638
rect 14748 24678 14763 30638
rect 14855 24678 14872 30638
rect 14872 24678 14906 30638
rect 14906 24678 14921 30638
rect 15013 24678 15030 30638
rect 15030 24678 15064 30638
rect 15064 24678 15079 30638
rect 15171 24678 15188 30638
rect 15188 24678 15222 30638
rect 15222 24678 15237 30638
rect 15329 24678 15346 30638
rect 15346 24678 15380 30638
rect 15380 24678 15395 30638
rect 15487 24678 15504 30638
rect 15504 24678 15538 30638
rect 15538 24678 15553 30638
rect 15645 24678 15662 30638
rect 15662 24678 15696 30638
rect 15696 24678 15711 30638
rect 15803 24678 15820 30638
rect 15820 24678 15854 30638
rect 15854 24678 15869 30638
rect 15961 24678 15978 30638
rect 15978 24678 16012 30638
rect 16012 24678 16027 30638
rect 16119 24678 16136 30638
rect 16136 24678 16170 30638
rect 16170 24678 16185 30638
rect 16277 24678 16294 30638
rect 16294 24678 16328 30638
rect 16328 24678 16343 30638
rect 16435 24678 16452 30638
rect 16452 24678 16486 30638
rect 16486 24678 16501 30638
rect 16593 24678 16610 30638
rect 16610 24678 16644 30638
rect 16644 24678 16659 30638
rect 16751 24678 16768 30638
rect 16768 24678 16802 30638
rect 16802 24678 16817 30638
rect 16909 24678 16926 30638
rect 16926 24678 16960 30638
rect 16960 24678 16975 30638
rect 17067 24678 17084 30638
rect 17084 24678 17118 30638
rect 17118 24678 17133 30638
rect 17225 24678 17242 30638
rect 17242 24678 17276 30638
rect 17276 24678 17291 30638
rect 17383 24678 17400 30638
rect 17400 24678 17434 30638
rect 17434 24678 17449 30638
rect 17541 24678 17558 30638
rect 17558 24678 17592 30638
rect 17592 24678 17607 30638
rect 17699 24678 17716 30638
rect 17716 24678 17750 30638
rect 17750 24678 17765 30638
rect 17857 24678 17874 30638
rect 17874 24678 17908 30638
rect 17908 24678 17923 30638
rect 18015 24678 18032 30638
rect 18032 24678 18066 30638
rect 18066 24678 18081 30638
rect 18173 24678 18190 30638
rect 18190 24678 18224 30638
rect 18224 24678 18239 30638
rect 18331 24678 18348 30638
rect 18348 24678 18382 30638
rect 18382 24678 18397 30638
rect 18489 24678 18506 30638
rect 18506 24678 18540 30638
rect 18540 24678 18555 30638
rect 18647 24678 18664 30638
rect 18664 24678 18698 30638
rect 18698 24678 18713 30638
rect 18805 24678 18822 30638
rect 18822 24678 18856 30638
rect 18856 24678 18871 30638
rect 13930 24500 14000 24636
rect 18940 24636 18954 30680
rect 18954 24636 18992 30680
rect 18992 24636 19010 30680
rect 19520 30650 19590 30850
rect 19910 30650 19980 30850
rect 19650 30520 19850 30590
rect 20230 30680 20300 30820
rect 20452 30730 25086 30790
rect 20452 30696 20512 30730
rect 20512 30696 20602 30730
rect 20602 30696 20670 30730
rect 20670 30696 20760 30730
rect 20760 30696 20828 30730
rect 20828 30696 20918 30730
rect 20918 30696 20986 30730
rect 20986 30696 21076 30730
rect 21076 30696 21144 30730
rect 21144 30696 21234 30730
rect 21234 30696 21302 30730
rect 21302 30696 21392 30730
rect 21392 30696 21460 30730
rect 21460 30696 21550 30730
rect 21550 30696 21618 30730
rect 21618 30696 21708 30730
rect 21708 30696 21776 30730
rect 21776 30696 21866 30730
rect 21866 30696 21934 30730
rect 21934 30696 22024 30730
rect 22024 30696 22092 30730
rect 22092 30696 22182 30730
rect 22182 30696 22250 30730
rect 22250 30696 22340 30730
rect 22340 30696 22408 30730
rect 22408 30696 22498 30730
rect 22498 30696 22566 30730
rect 22566 30696 22656 30730
rect 22656 30696 22724 30730
rect 22724 30696 22814 30730
rect 22814 30696 22882 30730
rect 22882 30696 22972 30730
rect 22972 30696 23040 30730
rect 23040 30696 23130 30730
rect 23130 30696 23198 30730
rect 23198 30696 23288 30730
rect 23288 30696 23356 30730
rect 23356 30696 23446 30730
rect 23446 30696 23514 30730
rect 23514 30696 23604 30730
rect 23604 30696 23672 30730
rect 23672 30696 23762 30730
rect 23762 30696 23830 30730
rect 23830 30696 23920 30730
rect 23920 30696 23988 30730
rect 23988 30696 24078 30730
rect 24078 30696 24146 30730
rect 24146 30696 24236 30730
rect 24236 30696 24304 30730
rect 24304 30696 24394 30730
rect 24394 30696 24462 30730
rect 24462 30696 24552 30730
rect 24552 30696 24620 30730
rect 24620 30696 24710 30730
rect 24710 30696 24778 30730
rect 24778 30696 24868 30730
rect 24868 30696 24936 30730
rect 24936 30696 25026 30730
rect 25026 30696 25086 30730
rect 20452 30690 25086 30696
rect 14152 24620 18786 24626
rect 14152 24586 14212 24620
rect 14212 24586 14302 24620
rect 14302 24586 14370 24620
rect 14370 24586 14460 24620
rect 14460 24586 14528 24620
rect 14528 24586 14618 24620
rect 14618 24586 14686 24620
rect 14686 24586 14776 24620
rect 14776 24586 14844 24620
rect 14844 24586 14934 24620
rect 14934 24586 15002 24620
rect 15002 24586 15092 24620
rect 15092 24586 15160 24620
rect 15160 24586 15250 24620
rect 15250 24586 15318 24620
rect 15318 24586 15408 24620
rect 15408 24586 15476 24620
rect 15476 24586 15566 24620
rect 15566 24586 15634 24620
rect 15634 24586 15724 24620
rect 15724 24586 15792 24620
rect 15792 24586 15882 24620
rect 15882 24586 15950 24620
rect 15950 24586 16040 24620
rect 16040 24586 16108 24620
rect 16108 24586 16198 24620
rect 16198 24586 16266 24620
rect 16266 24586 16356 24620
rect 16356 24586 16424 24620
rect 16424 24586 16514 24620
rect 16514 24586 16582 24620
rect 16582 24586 16672 24620
rect 16672 24586 16740 24620
rect 16740 24586 16830 24620
rect 16830 24586 16898 24620
rect 16898 24586 16988 24620
rect 16988 24586 17056 24620
rect 17056 24586 17146 24620
rect 17146 24586 17214 24620
rect 17214 24586 17304 24620
rect 17304 24586 17372 24620
rect 17372 24586 17462 24620
rect 17462 24586 17530 24620
rect 17530 24586 17620 24620
rect 17620 24586 17688 24620
rect 17688 24586 17778 24620
rect 17778 24586 17846 24620
rect 17846 24586 17936 24620
rect 17936 24586 18004 24620
rect 18004 24586 18094 24620
rect 18094 24586 18162 24620
rect 18162 24586 18252 24620
rect 18252 24586 18320 24620
rect 18320 24586 18410 24620
rect 18410 24586 18478 24620
rect 18478 24586 18568 24620
rect 18568 24586 18636 24620
rect 18636 24586 18726 24620
rect 18726 24586 18786 24620
rect 14152 24526 18786 24586
rect 18940 24500 19010 24636
rect 20230 24636 20246 30680
rect 20246 24636 20284 30680
rect 20284 24636 20300 30680
rect 25240 30680 25310 30820
rect 20365 24678 20382 30638
rect 20382 24678 20416 30638
rect 20416 24678 20431 30638
rect 20523 24678 20540 30638
rect 20540 24678 20574 30638
rect 20574 24678 20589 30638
rect 20681 24678 20698 30638
rect 20698 24678 20732 30638
rect 20732 24678 20747 30638
rect 20839 24678 20856 30638
rect 20856 24678 20890 30638
rect 20890 24678 20905 30638
rect 20997 24678 21014 30638
rect 21014 24678 21048 30638
rect 21048 24678 21063 30638
rect 21155 24678 21172 30638
rect 21172 24678 21206 30638
rect 21206 24678 21221 30638
rect 21313 24678 21330 30638
rect 21330 24678 21364 30638
rect 21364 24678 21379 30638
rect 21471 24678 21488 30638
rect 21488 24678 21522 30638
rect 21522 24678 21537 30638
rect 21629 24678 21646 30638
rect 21646 24678 21680 30638
rect 21680 24678 21695 30638
rect 21787 24678 21804 30638
rect 21804 24678 21838 30638
rect 21838 24678 21853 30638
rect 21945 24678 21962 30638
rect 21962 24678 21996 30638
rect 21996 24678 22011 30638
rect 22103 24678 22120 30638
rect 22120 24678 22154 30638
rect 22154 24678 22169 30638
rect 22261 24678 22278 30638
rect 22278 24678 22312 30638
rect 22312 24678 22327 30638
rect 22419 24678 22436 30638
rect 22436 24678 22470 30638
rect 22470 24678 22485 30638
rect 22577 24678 22594 30638
rect 22594 24678 22628 30638
rect 22628 24678 22643 30638
rect 22735 24678 22752 30638
rect 22752 24678 22786 30638
rect 22786 24678 22801 30638
rect 22893 24678 22910 30638
rect 22910 24678 22944 30638
rect 22944 24678 22959 30638
rect 23051 24678 23068 30638
rect 23068 24678 23102 30638
rect 23102 24678 23117 30638
rect 23209 24678 23226 30638
rect 23226 24678 23260 30638
rect 23260 24678 23275 30638
rect 23367 24678 23384 30638
rect 23384 24678 23418 30638
rect 23418 24678 23433 30638
rect 23525 24678 23542 30638
rect 23542 24678 23576 30638
rect 23576 24678 23591 30638
rect 23683 24678 23700 30638
rect 23700 24678 23734 30638
rect 23734 24678 23749 30638
rect 23841 24678 23858 30638
rect 23858 24678 23892 30638
rect 23892 24678 23907 30638
rect 23999 24678 24016 30638
rect 24016 24678 24050 30638
rect 24050 24678 24065 30638
rect 24157 24678 24174 30638
rect 24174 24678 24208 30638
rect 24208 24678 24223 30638
rect 24315 24678 24332 30638
rect 24332 24678 24366 30638
rect 24366 24678 24381 30638
rect 24473 24678 24490 30638
rect 24490 24678 24524 30638
rect 24524 24678 24539 30638
rect 24631 24678 24648 30638
rect 24648 24678 24682 30638
rect 24682 24678 24697 30638
rect 24789 24678 24806 30638
rect 24806 24678 24840 30638
rect 24840 24678 24855 30638
rect 24947 24678 24964 30638
rect 24964 24678 24998 30638
rect 24998 24678 25013 30638
rect 25105 24678 25122 30638
rect 25122 24678 25156 30638
rect 25156 24678 25171 30638
rect 20230 24500 20300 24636
rect 25240 24636 25254 30680
rect 25254 24636 25292 30680
rect 25292 24636 25310 30680
rect 25520 30650 25590 30850
rect 25910 30650 25980 30850
rect 26020 30650 26090 30850
rect 26410 30650 26480 30850
rect 25650 30520 25850 30590
rect 26150 30520 26350 30590
rect 25650 30410 25850 30480
rect 26150 30410 26350 30480
rect 25520 30150 25590 30350
rect 25910 30150 25980 30350
rect 26020 30150 26090 30350
rect 26410 30150 26480 30350
rect 25650 30020 25850 30090
rect 26150 30020 26350 30090
rect 25650 29910 25850 29980
rect 26150 29910 26350 29980
rect 25520 29650 25590 29850
rect 25910 29650 25980 29850
rect 26020 29650 26090 29850
rect 26410 29650 26480 29850
rect 25650 29520 25850 29590
rect 26150 29520 26350 29590
rect 25650 29410 25850 29480
rect 26150 29410 26350 29480
rect 25520 29150 25590 29350
rect 25910 29150 25980 29350
rect 26020 29150 26090 29350
rect 26410 29150 26480 29350
rect 25650 29020 25850 29090
rect 26150 29020 26350 29090
rect 25650 28910 25850 28980
rect 26150 28910 26350 28980
rect 25520 28650 25590 28850
rect 25910 28650 25980 28850
rect 26020 28650 26090 28850
rect 26410 28650 26480 28850
rect 25650 28520 25850 28590
rect 26150 28520 26350 28590
rect 25650 28410 25850 28480
rect 26150 28410 26350 28480
rect 25520 28150 25590 28350
rect 25910 28150 25980 28350
rect 26020 28150 26090 28350
rect 26410 28150 26480 28350
rect 25650 28020 25850 28090
rect 26150 28020 26350 28090
rect 25650 27910 25850 27980
rect 26150 27910 26350 27980
rect 25520 27650 25590 27850
rect 25910 27650 25980 27850
rect 26020 27650 26090 27850
rect 26410 27650 26480 27850
rect 25650 27520 25850 27590
rect 26150 27520 26350 27590
rect 25650 27410 25850 27480
rect 26150 27410 26350 27480
rect 25520 27150 25590 27350
rect 25910 27150 25980 27350
rect 26020 27150 26090 27350
rect 26410 27150 26480 27350
rect 25650 27020 25850 27090
rect 26150 27020 26350 27090
rect 30910 27076 31090 27250
rect 30910 27036 30984 27076
rect 30984 27036 31018 27076
rect 31018 27036 31090 27076
rect 30910 27030 31090 27036
rect 25650 26910 25850 26980
rect 26150 26910 26350 26980
rect 26650 26910 26850 26980
rect 27150 26910 27350 26980
rect 27650 26910 27850 26980
rect 28150 26910 28350 26980
rect 28650 26910 28850 26980
rect 29150 26910 29350 26980
rect 29650 26910 29850 26980
rect 30150 26910 30350 26980
rect 25520 26650 25590 26850
rect 25910 26650 25980 26850
rect 26020 26650 26090 26850
rect 26410 26650 26480 26850
rect 26520 26650 26590 26850
rect 26910 26650 26980 26850
rect 27020 26650 27090 26850
rect 27410 26650 27480 26850
rect 27520 26650 27590 26850
rect 27910 26650 27980 26850
rect 28020 26650 28090 26850
rect 28410 26650 28480 26850
rect 28520 26650 28590 26850
rect 28910 26650 28980 26850
rect 29020 26650 29090 26850
rect 29410 26650 29480 26850
rect 29520 26650 29590 26850
rect 29910 26650 29980 26850
rect 30020 26650 30090 26850
rect 30410 26650 30480 26850
rect 25650 26520 25850 26590
rect 26150 26520 26350 26590
rect 26650 26520 26850 26590
rect 27150 26520 27350 26590
rect 27650 26520 27850 26590
rect 28150 26520 28350 26590
rect 28650 26520 28850 26590
rect 29150 26520 29350 26590
rect 29650 26520 29850 26590
rect 30150 26520 30350 26590
rect 25650 26410 25850 26480
rect 26150 26410 26350 26480
rect 26650 26410 26850 26480
rect 27150 26410 27350 26480
rect 27650 26410 27850 26480
rect 28150 26410 28350 26480
rect 28650 26410 28850 26480
rect 29150 26410 29350 26480
rect 29650 26410 29850 26480
rect 30150 26410 30350 26480
rect 25520 26150 25590 26350
rect 25910 26150 25980 26350
rect 26020 26150 26090 26350
rect 26410 26150 26480 26350
rect 26520 26150 26590 26350
rect 26910 26150 26980 26350
rect 27020 26150 27090 26350
rect 27410 26150 27480 26350
rect 27520 26150 27590 26350
rect 27910 26150 27980 26350
rect 28020 26150 28090 26350
rect 28410 26150 28480 26350
rect 28520 26150 28590 26350
rect 28910 26150 28980 26350
rect 29020 26150 29090 26350
rect 29410 26150 29480 26350
rect 29520 26150 29590 26350
rect 29910 26150 29980 26350
rect 30020 26150 30090 26350
rect 30410 26150 30480 26350
rect 25650 26020 25850 26090
rect 26150 26020 26350 26090
rect 26650 26020 26850 26090
rect 27150 26020 27350 26090
rect 27650 26020 27850 26090
rect 28150 26020 28350 26090
rect 28650 26020 28850 26090
rect 29150 26020 29350 26090
rect 29650 26020 29850 26090
rect 30150 26020 30350 26090
rect 25650 25910 25850 25980
rect 26150 25910 26350 25980
rect 25520 25650 25590 25850
rect 25910 25650 25980 25850
rect 26020 25650 26090 25850
rect 26410 25650 26480 25850
rect 25650 25520 25850 25590
rect 26150 25520 26350 25590
rect 30910 25702 31090 25710
rect 30910 25662 30984 25702
rect 30984 25662 31018 25702
rect 31018 25662 31090 25702
rect 30910 25490 31090 25662
rect 25650 25410 25850 25480
rect 26150 25410 26350 25480
rect 25520 25150 25590 25350
rect 25910 25150 25980 25350
rect 26020 25150 26090 25350
rect 26410 25150 26480 25350
rect 25650 25020 25850 25090
rect 26150 25020 26350 25090
rect 25650 24910 25850 24980
rect 26150 24910 26350 24980
rect 25520 24650 25590 24850
rect 20452 24620 25086 24626
rect 20452 24586 20512 24620
rect 20512 24586 20602 24620
rect 20602 24586 20670 24620
rect 20670 24586 20760 24620
rect 20760 24586 20828 24620
rect 20828 24586 20918 24620
rect 20918 24586 20986 24620
rect 20986 24586 21076 24620
rect 21076 24586 21144 24620
rect 21144 24586 21234 24620
rect 21234 24586 21302 24620
rect 21302 24586 21392 24620
rect 21392 24586 21460 24620
rect 21460 24586 21550 24620
rect 21550 24586 21618 24620
rect 21618 24586 21708 24620
rect 21708 24586 21776 24620
rect 21776 24586 21866 24620
rect 21866 24586 21934 24620
rect 21934 24586 22024 24620
rect 22024 24586 22092 24620
rect 22092 24586 22182 24620
rect 22182 24586 22250 24620
rect 22250 24586 22340 24620
rect 22340 24586 22408 24620
rect 22408 24586 22498 24620
rect 22498 24586 22566 24620
rect 22566 24586 22656 24620
rect 22656 24586 22724 24620
rect 22724 24586 22814 24620
rect 22814 24586 22882 24620
rect 22882 24586 22972 24620
rect 22972 24586 23040 24620
rect 23040 24586 23130 24620
rect 23130 24586 23198 24620
rect 23198 24586 23288 24620
rect 23288 24586 23356 24620
rect 23356 24586 23446 24620
rect 23446 24586 23514 24620
rect 23514 24586 23604 24620
rect 23604 24586 23672 24620
rect 23672 24586 23762 24620
rect 23762 24586 23830 24620
rect 23830 24586 23920 24620
rect 23920 24586 23988 24620
rect 23988 24586 24078 24620
rect 24078 24586 24146 24620
rect 24146 24586 24236 24620
rect 24236 24586 24304 24620
rect 24304 24586 24394 24620
rect 24394 24586 24462 24620
rect 24462 24586 24552 24620
rect 24552 24586 24620 24620
rect 24620 24586 24710 24620
rect 24710 24586 24778 24620
rect 24778 24586 24868 24620
rect 24868 24586 24936 24620
rect 24936 24586 25026 24620
rect 25026 24586 25086 24620
rect 20452 24526 25086 24586
rect 25240 24500 25310 24636
rect 25910 24650 25980 24850
rect 26020 24650 26090 24850
rect 26410 24650 26480 24850
rect 25650 24520 25850 24590
rect 26150 24520 26350 24590
rect 20 24150 90 24350
rect 410 24150 480 24350
rect 520 24150 590 24350
rect 910 24150 980 24350
rect 150 24020 350 24090
rect 650 24020 850 24090
rect 150 23910 350 23980
rect 650 23910 850 23980
rect 25650 24410 25850 24480
rect 26150 24410 26350 24480
rect 25520 24150 25590 24350
rect 25910 24150 25980 24350
rect 26020 24150 26090 24350
rect 26410 24150 26480 24350
rect 25650 24020 25850 24090
rect 26150 24020 26350 24090
rect 25650 23910 25850 23980
rect 26150 23910 26350 23980
rect 20 23650 90 23850
rect 410 23650 480 23850
rect 520 23650 590 23850
rect 910 23650 980 23850
rect 1330 23680 1400 23820
rect 1552 23730 6186 23790
rect 1552 23696 1612 23730
rect 1612 23696 1702 23730
rect 1702 23696 1770 23730
rect 1770 23696 1860 23730
rect 1860 23696 1928 23730
rect 1928 23696 2018 23730
rect 2018 23696 2086 23730
rect 2086 23696 2176 23730
rect 2176 23696 2244 23730
rect 2244 23696 2334 23730
rect 2334 23696 2402 23730
rect 2402 23696 2492 23730
rect 2492 23696 2560 23730
rect 2560 23696 2650 23730
rect 2650 23696 2718 23730
rect 2718 23696 2808 23730
rect 2808 23696 2876 23730
rect 2876 23696 2966 23730
rect 2966 23696 3034 23730
rect 3034 23696 3124 23730
rect 3124 23696 3192 23730
rect 3192 23696 3282 23730
rect 3282 23696 3350 23730
rect 3350 23696 3440 23730
rect 3440 23696 3508 23730
rect 3508 23696 3598 23730
rect 3598 23696 3666 23730
rect 3666 23696 3756 23730
rect 3756 23696 3824 23730
rect 3824 23696 3914 23730
rect 3914 23696 3982 23730
rect 3982 23696 4072 23730
rect 4072 23696 4140 23730
rect 4140 23696 4230 23730
rect 4230 23696 4298 23730
rect 4298 23696 4388 23730
rect 4388 23696 4456 23730
rect 4456 23696 4546 23730
rect 4546 23696 4614 23730
rect 4614 23696 4704 23730
rect 4704 23696 4772 23730
rect 4772 23696 4862 23730
rect 4862 23696 4930 23730
rect 4930 23696 5020 23730
rect 5020 23696 5088 23730
rect 5088 23696 5178 23730
rect 5178 23696 5246 23730
rect 5246 23696 5336 23730
rect 5336 23696 5404 23730
rect 5404 23696 5494 23730
rect 5494 23696 5562 23730
rect 5562 23696 5652 23730
rect 5652 23696 5720 23730
rect 5720 23696 5810 23730
rect 5810 23696 5878 23730
rect 5878 23696 5968 23730
rect 5968 23696 6036 23730
rect 6036 23696 6126 23730
rect 6126 23696 6186 23730
rect 1552 23690 6186 23696
rect 150 23520 350 23590
rect 650 23520 850 23590
rect 150 23410 350 23480
rect 650 23410 850 23480
rect 20 23150 90 23350
rect 410 23150 480 23350
rect 520 23150 590 23350
rect 910 23150 980 23350
rect 150 23020 350 23090
rect 650 23020 850 23090
rect 150 22910 350 22980
rect 650 22910 850 22980
rect 20 22650 90 22850
rect 410 22650 480 22850
rect 520 22650 590 22850
rect 910 22650 980 22850
rect 150 22520 350 22590
rect 650 22520 850 22590
rect 150 22410 350 22480
rect 650 22410 850 22480
rect 20 22150 90 22350
rect 410 22150 480 22350
rect 520 22150 590 22350
rect 910 22150 980 22350
rect 150 22020 350 22090
rect 650 22020 850 22090
rect 150 21910 350 21980
rect 650 21910 850 21980
rect 20 21650 90 21850
rect 410 21650 480 21850
rect 520 21650 590 21850
rect 910 21650 980 21850
rect 150 21520 350 21590
rect 650 21520 850 21590
rect 150 21410 350 21480
rect 650 21410 850 21480
rect 20 21150 90 21350
rect 410 21150 480 21350
rect 520 21150 590 21350
rect 910 21150 980 21350
rect 150 21020 350 21090
rect 650 21020 850 21090
rect 150 20910 350 20980
rect 650 20910 850 20980
rect 20 20650 90 20850
rect 410 20650 480 20850
rect 520 20650 590 20850
rect 910 20650 980 20850
rect 150 20520 350 20590
rect 650 20520 850 20590
rect 150 20410 350 20480
rect 650 20410 850 20480
rect 20 20150 90 20350
rect 410 20150 480 20350
rect 520 20150 590 20350
rect 910 20150 980 20350
rect 150 20020 350 20090
rect 650 20020 850 20090
rect 150 19910 350 19980
rect 650 19910 850 19980
rect 20 19650 90 19850
rect 410 19650 480 19850
rect 520 19650 590 19850
rect 910 19650 980 19850
rect 150 19520 350 19590
rect 650 19520 850 19590
rect 150 19410 350 19480
rect 650 19410 850 19480
rect 20 19150 90 19350
rect 410 19150 480 19350
rect 520 19150 590 19350
rect 910 19150 980 19350
rect 150 19020 350 19090
rect 650 19020 850 19090
rect 150 18910 350 18980
rect 650 18910 850 18980
rect 20 18650 90 18850
rect 410 18650 480 18850
rect 520 18650 590 18850
rect 910 18650 980 18850
rect 150 18520 350 18590
rect 650 18520 850 18590
rect 150 18410 350 18480
rect 650 18410 850 18480
rect 20 18150 90 18350
rect 410 18150 480 18350
rect 520 18150 590 18350
rect 910 18150 980 18350
rect 150 18020 350 18090
rect 650 18020 850 18090
rect 150 17910 350 17980
rect 650 17910 850 17980
rect 20 17650 90 17850
rect 410 17650 480 17850
rect 520 17650 590 17850
rect 910 17650 980 17850
rect 1330 17636 1346 23680
rect 1346 17636 1384 23680
rect 1384 17636 1400 23680
rect 6340 23680 6410 23820
rect 1465 17678 1482 23638
rect 1482 17678 1516 23638
rect 1516 17678 1531 23638
rect 1623 17678 1640 23638
rect 1640 17678 1674 23638
rect 1674 17678 1689 23638
rect 1781 17678 1798 23638
rect 1798 17678 1832 23638
rect 1832 17678 1847 23638
rect 1939 17678 1956 23638
rect 1956 17678 1990 23638
rect 1990 17678 2005 23638
rect 2097 17678 2114 23638
rect 2114 17678 2148 23638
rect 2148 17678 2163 23638
rect 2255 17678 2272 23638
rect 2272 17678 2306 23638
rect 2306 17678 2321 23638
rect 2413 17678 2430 23638
rect 2430 17678 2464 23638
rect 2464 17678 2479 23638
rect 2571 17678 2588 23638
rect 2588 17678 2622 23638
rect 2622 17678 2637 23638
rect 2729 17678 2746 23638
rect 2746 17678 2780 23638
rect 2780 17678 2795 23638
rect 2887 17678 2904 23638
rect 2904 17678 2938 23638
rect 2938 17678 2953 23638
rect 3045 17678 3062 23638
rect 3062 17678 3096 23638
rect 3096 17678 3111 23638
rect 3203 17678 3220 23638
rect 3220 17678 3254 23638
rect 3254 17678 3269 23638
rect 3361 17678 3378 23638
rect 3378 17678 3412 23638
rect 3412 17678 3427 23638
rect 3519 17678 3536 23638
rect 3536 17678 3570 23638
rect 3570 17678 3585 23638
rect 3677 17678 3694 23638
rect 3694 17678 3728 23638
rect 3728 17678 3743 23638
rect 3835 17678 3852 23638
rect 3852 17678 3886 23638
rect 3886 17678 3901 23638
rect 3993 17678 4010 23638
rect 4010 17678 4044 23638
rect 4044 17678 4059 23638
rect 4151 17678 4168 23638
rect 4168 17678 4202 23638
rect 4202 17678 4217 23638
rect 4309 17678 4326 23638
rect 4326 17678 4360 23638
rect 4360 17678 4375 23638
rect 4467 17678 4484 23638
rect 4484 17678 4518 23638
rect 4518 17678 4533 23638
rect 4625 17678 4642 23638
rect 4642 17678 4676 23638
rect 4676 17678 4691 23638
rect 4783 17678 4800 23638
rect 4800 17678 4834 23638
rect 4834 17678 4849 23638
rect 4941 17678 4958 23638
rect 4958 17678 4992 23638
rect 4992 17678 5007 23638
rect 5099 17678 5116 23638
rect 5116 17678 5150 23638
rect 5150 17678 5165 23638
rect 5257 17678 5274 23638
rect 5274 17678 5308 23638
rect 5308 17678 5323 23638
rect 5415 17678 5432 23638
rect 5432 17678 5466 23638
rect 5466 17678 5481 23638
rect 5573 17678 5590 23638
rect 5590 17678 5624 23638
rect 5624 17678 5639 23638
rect 5731 17678 5748 23638
rect 5748 17678 5782 23638
rect 5782 17678 5797 23638
rect 5889 17678 5906 23638
rect 5906 17678 5940 23638
rect 5940 17678 5955 23638
rect 6047 17678 6064 23638
rect 6064 17678 6098 23638
rect 6098 17678 6113 23638
rect 6205 17678 6222 23638
rect 6222 17678 6256 23638
rect 6256 17678 6271 23638
rect 150 17520 350 17590
rect 650 17520 850 17590
rect 1330 17500 1400 17636
rect 6340 17636 6354 23680
rect 6354 17636 6392 23680
rect 6392 17636 6410 23680
rect 1552 17620 6186 17626
rect 1552 17586 1612 17620
rect 1612 17586 1702 17620
rect 1702 17586 1770 17620
rect 1770 17586 1860 17620
rect 1860 17586 1928 17620
rect 1928 17586 2018 17620
rect 2018 17586 2086 17620
rect 2086 17586 2176 17620
rect 2176 17586 2244 17620
rect 2244 17586 2334 17620
rect 2334 17586 2402 17620
rect 2402 17586 2492 17620
rect 2492 17586 2560 17620
rect 2560 17586 2650 17620
rect 2650 17586 2718 17620
rect 2718 17586 2808 17620
rect 2808 17586 2876 17620
rect 2876 17586 2966 17620
rect 2966 17586 3034 17620
rect 3034 17586 3124 17620
rect 3124 17586 3192 17620
rect 3192 17586 3282 17620
rect 3282 17586 3350 17620
rect 3350 17586 3440 17620
rect 3440 17586 3508 17620
rect 3508 17586 3598 17620
rect 3598 17586 3666 17620
rect 3666 17586 3756 17620
rect 3756 17586 3824 17620
rect 3824 17586 3914 17620
rect 3914 17586 3982 17620
rect 3982 17586 4072 17620
rect 4072 17586 4140 17620
rect 4140 17586 4230 17620
rect 4230 17586 4298 17620
rect 4298 17586 4388 17620
rect 4388 17586 4456 17620
rect 4456 17586 4546 17620
rect 4546 17586 4614 17620
rect 4614 17586 4704 17620
rect 4704 17586 4772 17620
rect 4772 17586 4862 17620
rect 4862 17586 4930 17620
rect 4930 17586 5020 17620
rect 5020 17586 5088 17620
rect 5088 17586 5178 17620
rect 5178 17586 5246 17620
rect 5246 17586 5336 17620
rect 5336 17586 5404 17620
rect 5404 17586 5494 17620
rect 5494 17586 5562 17620
rect 5562 17586 5652 17620
rect 5652 17586 5720 17620
rect 5720 17586 5810 17620
rect 5810 17586 5878 17620
rect 5878 17586 5968 17620
rect 5968 17586 6036 17620
rect 6036 17586 6126 17620
rect 6126 17586 6186 17620
rect 1552 17526 6186 17586
rect 6340 17500 6410 17636
rect 7630 23680 7700 23820
rect 7852 23730 12486 23790
rect 7852 23696 7912 23730
rect 7912 23696 8002 23730
rect 8002 23696 8070 23730
rect 8070 23696 8160 23730
rect 8160 23696 8228 23730
rect 8228 23696 8318 23730
rect 8318 23696 8386 23730
rect 8386 23696 8476 23730
rect 8476 23696 8544 23730
rect 8544 23696 8634 23730
rect 8634 23696 8702 23730
rect 8702 23696 8792 23730
rect 8792 23696 8860 23730
rect 8860 23696 8950 23730
rect 8950 23696 9018 23730
rect 9018 23696 9108 23730
rect 9108 23696 9176 23730
rect 9176 23696 9266 23730
rect 9266 23696 9334 23730
rect 9334 23696 9424 23730
rect 9424 23696 9492 23730
rect 9492 23696 9582 23730
rect 9582 23696 9650 23730
rect 9650 23696 9740 23730
rect 9740 23696 9808 23730
rect 9808 23696 9898 23730
rect 9898 23696 9966 23730
rect 9966 23696 10056 23730
rect 10056 23696 10124 23730
rect 10124 23696 10214 23730
rect 10214 23696 10282 23730
rect 10282 23696 10372 23730
rect 10372 23696 10440 23730
rect 10440 23696 10530 23730
rect 10530 23696 10598 23730
rect 10598 23696 10688 23730
rect 10688 23696 10756 23730
rect 10756 23696 10846 23730
rect 10846 23696 10914 23730
rect 10914 23696 11004 23730
rect 11004 23696 11072 23730
rect 11072 23696 11162 23730
rect 11162 23696 11230 23730
rect 11230 23696 11320 23730
rect 11320 23696 11388 23730
rect 11388 23696 11478 23730
rect 11478 23696 11546 23730
rect 11546 23696 11636 23730
rect 11636 23696 11704 23730
rect 11704 23696 11794 23730
rect 11794 23696 11862 23730
rect 11862 23696 11952 23730
rect 11952 23696 12020 23730
rect 12020 23696 12110 23730
rect 12110 23696 12178 23730
rect 12178 23696 12268 23730
rect 12268 23696 12336 23730
rect 12336 23696 12426 23730
rect 12426 23696 12486 23730
rect 7852 23690 12486 23696
rect 7630 17636 7646 23680
rect 7646 17636 7684 23680
rect 7684 17636 7700 23680
rect 12640 23680 12710 23820
rect 7765 17678 7782 23638
rect 7782 17678 7816 23638
rect 7816 17678 7831 23638
rect 7923 17678 7940 23638
rect 7940 17678 7974 23638
rect 7974 17678 7989 23638
rect 8081 17678 8098 23638
rect 8098 17678 8132 23638
rect 8132 17678 8147 23638
rect 8239 17678 8256 23638
rect 8256 17678 8290 23638
rect 8290 17678 8305 23638
rect 8397 17678 8414 23638
rect 8414 17678 8448 23638
rect 8448 17678 8463 23638
rect 8555 17678 8572 23638
rect 8572 17678 8606 23638
rect 8606 17678 8621 23638
rect 8713 17678 8730 23638
rect 8730 17678 8764 23638
rect 8764 17678 8779 23638
rect 8871 17678 8888 23638
rect 8888 17678 8922 23638
rect 8922 17678 8937 23638
rect 9029 17678 9046 23638
rect 9046 17678 9080 23638
rect 9080 17678 9095 23638
rect 9187 17678 9204 23638
rect 9204 17678 9238 23638
rect 9238 17678 9253 23638
rect 9345 17678 9362 23638
rect 9362 17678 9396 23638
rect 9396 17678 9411 23638
rect 9503 17678 9520 23638
rect 9520 17678 9554 23638
rect 9554 17678 9569 23638
rect 9661 17678 9678 23638
rect 9678 17678 9712 23638
rect 9712 17678 9727 23638
rect 9819 17678 9836 23638
rect 9836 17678 9870 23638
rect 9870 17678 9885 23638
rect 9977 17678 9994 23638
rect 9994 17678 10028 23638
rect 10028 17678 10043 23638
rect 10135 17678 10152 23638
rect 10152 17678 10186 23638
rect 10186 17678 10201 23638
rect 10293 17678 10310 23638
rect 10310 17678 10344 23638
rect 10344 17678 10359 23638
rect 10451 17678 10468 23638
rect 10468 17678 10502 23638
rect 10502 17678 10517 23638
rect 10609 17678 10626 23638
rect 10626 17678 10660 23638
rect 10660 17678 10675 23638
rect 10767 17678 10784 23638
rect 10784 17678 10818 23638
rect 10818 17678 10833 23638
rect 10925 17678 10942 23638
rect 10942 17678 10976 23638
rect 10976 17678 10991 23638
rect 11083 17678 11100 23638
rect 11100 17678 11134 23638
rect 11134 17678 11149 23638
rect 11241 17678 11258 23638
rect 11258 17678 11292 23638
rect 11292 17678 11307 23638
rect 11399 17678 11416 23638
rect 11416 17678 11450 23638
rect 11450 17678 11465 23638
rect 11557 17678 11574 23638
rect 11574 17678 11608 23638
rect 11608 17678 11623 23638
rect 11715 17678 11732 23638
rect 11732 17678 11766 23638
rect 11766 17678 11781 23638
rect 11873 17678 11890 23638
rect 11890 17678 11924 23638
rect 11924 17678 11939 23638
rect 12031 17678 12048 23638
rect 12048 17678 12082 23638
rect 12082 17678 12097 23638
rect 12189 17678 12206 23638
rect 12206 17678 12240 23638
rect 12240 17678 12255 23638
rect 12347 17678 12364 23638
rect 12364 17678 12398 23638
rect 12398 17678 12413 23638
rect 12505 17678 12522 23638
rect 12522 17678 12556 23638
rect 12556 17678 12571 23638
rect 7630 17500 7700 17636
rect 12640 17636 12654 23680
rect 12654 17636 12692 23680
rect 12692 17636 12710 23680
rect 7852 17620 12486 17626
rect 7852 17586 7912 17620
rect 7912 17586 8002 17620
rect 8002 17586 8070 17620
rect 8070 17586 8160 17620
rect 8160 17586 8228 17620
rect 8228 17586 8318 17620
rect 8318 17586 8386 17620
rect 8386 17586 8476 17620
rect 8476 17586 8544 17620
rect 8544 17586 8634 17620
rect 8634 17586 8702 17620
rect 8702 17586 8792 17620
rect 8792 17586 8860 17620
rect 8860 17586 8950 17620
rect 8950 17586 9018 17620
rect 9018 17586 9108 17620
rect 9108 17586 9176 17620
rect 9176 17586 9266 17620
rect 9266 17586 9334 17620
rect 9334 17586 9424 17620
rect 9424 17586 9492 17620
rect 9492 17586 9582 17620
rect 9582 17586 9650 17620
rect 9650 17586 9740 17620
rect 9740 17586 9808 17620
rect 9808 17586 9898 17620
rect 9898 17586 9966 17620
rect 9966 17586 10056 17620
rect 10056 17586 10124 17620
rect 10124 17586 10214 17620
rect 10214 17586 10282 17620
rect 10282 17586 10372 17620
rect 10372 17586 10440 17620
rect 10440 17586 10530 17620
rect 10530 17586 10598 17620
rect 10598 17586 10688 17620
rect 10688 17586 10756 17620
rect 10756 17586 10846 17620
rect 10846 17586 10914 17620
rect 10914 17586 11004 17620
rect 11004 17586 11072 17620
rect 11072 17586 11162 17620
rect 11162 17586 11230 17620
rect 11230 17586 11320 17620
rect 11320 17586 11388 17620
rect 11388 17586 11478 17620
rect 11478 17586 11546 17620
rect 11546 17586 11636 17620
rect 11636 17586 11704 17620
rect 11704 17586 11794 17620
rect 11794 17586 11862 17620
rect 11862 17586 11952 17620
rect 11952 17586 12020 17620
rect 12020 17586 12110 17620
rect 12110 17586 12178 17620
rect 12178 17586 12268 17620
rect 12268 17586 12336 17620
rect 12336 17586 12426 17620
rect 12426 17586 12486 17620
rect 7852 17526 12486 17586
rect 150 17410 350 17480
rect 650 17410 850 17480
rect 20 17150 90 17350
rect 410 17150 480 17350
rect 520 17150 590 17350
rect 910 17150 980 17350
rect 150 17020 350 17090
rect 650 17020 850 17090
rect 6650 17410 6850 17480
rect 7150 17410 7350 17480
rect 12640 17500 12710 17636
rect 13930 23680 14000 23820
rect 14152 23730 18786 23790
rect 14152 23696 14212 23730
rect 14212 23696 14302 23730
rect 14302 23696 14370 23730
rect 14370 23696 14460 23730
rect 14460 23696 14528 23730
rect 14528 23696 14618 23730
rect 14618 23696 14686 23730
rect 14686 23696 14776 23730
rect 14776 23696 14844 23730
rect 14844 23696 14934 23730
rect 14934 23696 15002 23730
rect 15002 23696 15092 23730
rect 15092 23696 15160 23730
rect 15160 23696 15250 23730
rect 15250 23696 15318 23730
rect 15318 23696 15408 23730
rect 15408 23696 15476 23730
rect 15476 23696 15566 23730
rect 15566 23696 15634 23730
rect 15634 23696 15724 23730
rect 15724 23696 15792 23730
rect 15792 23696 15882 23730
rect 15882 23696 15950 23730
rect 15950 23696 16040 23730
rect 16040 23696 16108 23730
rect 16108 23696 16198 23730
rect 16198 23696 16266 23730
rect 16266 23696 16356 23730
rect 16356 23696 16424 23730
rect 16424 23696 16514 23730
rect 16514 23696 16582 23730
rect 16582 23696 16672 23730
rect 16672 23696 16740 23730
rect 16740 23696 16830 23730
rect 16830 23696 16898 23730
rect 16898 23696 16988 23730
rect 16988 23696 17056 23730
rect 17056 23696 17146 23730
rect 17146 23696 17214 23730
rect 17214 23696 17304 23730
rect 17304 23696 17372 23730
rect 17372 23696 17462 23730
rect 17462 23696 17530 23730
rect 17530 23696 17620 23730
rect 17620 23696 17688 23730
rect 17688 23696 17778 23730
rect 17778 23696 17846 23730
rect 17846 23696 17936 23730
rect 17936 23696 18004 23730
rect 18004 23696 18094 23730
rect 18094 23696 18162 23730
rect 18162 23696 18252 23730
rect 18252 23696 18320 23730
rect 18320 23696 18410 23730
rect 18410 23696 18478 23730
rect 18478 23696 18568 23730
rect 18568 23696 18636 23730
rect 18636 23696 18726 23730
rect 18726 23696 18786 23730
rect 14152 23690 18786 23696
rect 13930 17636 13946 23680
rect 13946 17636 13984 23680
rect 13984 17636 14000 23680
rect 18940 23680 19010 23820
rect 14065 17678 14082 23638
rect 14082 17678 14116 23638
rect 14116 17678 14131 23638
rect 14223 17678 14240 23638
rect 14240 17678 14274 23638
rect 14274 17678 14289 23638
rect 14381 17678 14398 23638
rect 14398 17678 14432 23638
rect 14432 17678 14447 23638
rect 14539 17678 14556 23638
rect 14556 17678 14590 23638
rect 14590 17678 14605 23638
rect 14697 17678 14714 23638
rect 14714 17678 14748 23638
rect 14748 17678 14763 23638
rect 14855 17678 14872 23638
rect 14872 17678 14906 23638
rect 14906 17678 14921 23638
rect 15013 17678 15030 23638
rect 15030 17678 15064 23638
rect 15064 17678 15079 23638
rect 15171 17678 15188 23638
rect 15188 17678 15222 23638
rect 15222 17678 15237 23638
rect 15329 17678 15346 23638
rect 15346 17678 15380 23638
rect 15380 17678 15395 23638
rect 15487 17678 15504 23638
rect 15504 17678 15538 23638
rect 15538 17678 15553 23638
rect 15645 17678 15662 23638
rect 15662 17678 15696 23638
rect 15696 17678 15711 23638
rect 15803 17678 15820 23638
rect 15820 17678 15854 23638
rect 15854 17678 15869 23638
rect 15961 17678 15978 23638
rect 15978 17678 16012 23638
rect 16012 17678 16027 23638
rect 16119 17678 16136 23638
rect 16136 17678 16170 23638
rect 16170 17678 16185 23638
rect 16277 17678 16294 23638
rect 16294 17678 16328 23638
rect 16328 17678 16343 23638
rect 16435 17678 16452 23638
rect 16452 17678 16486 23638
rect 16486 17678 16501 23638
rect 16593 17678 16610 23638
rect 16610 17678 16644 23638
rect 16644 17678 16659 23638
rect 16751 17678 16768 23638
rect 16768 17678 16802 23638
rect 16802 17678 16817 23638
rect 16909 17678 16926 23638
rect 16926 17678 16960 23638
rect 16960 17678 16975 23638
rect 17067 17678 17084 23638
rect 17084 17678 17118 23638
rect 17118 17678 17133 23638
rect 17225 17678 17242 23638
rect 17242 17678 17276 23638
rect 17276 17678 17291 23638
rect 17383 17678 17400 23638
rect 17400 17678 17434 23638
rect 17434 17678 17449 23638
rect 17541 17678 17558 23638
rect 17558 17678 17592 23638
rect 17592 17678 17607 23638
rect 17699 17678 17716 23638
rect 17716 17678 17750 23638
rect 17750 17678 17765 23638
rect 17857 17678 17874 23638
rect 17874 17678 17908 23638
rect 17908 17678 17923 23638
rect 18015 17678 18032 23638
rect 18032 17678 18066 23638
rect 18066 17678 18081 23638
rect 18173 17678 18190 23638
rect 18190 17678 18224 23638
rect 18224 17678 18239 23638
rect 18331 17678 18348 23638
rect 18348 17678 18382 23638
rect 18382 17678 18397 23638
rect 18489 17678 18506 23638
rect 18506 17678 18540 23638
rect 18540 17678 18555 23638
rect 18647 17678 18664 23638
rect 18664 17678 18698 23638
rect 18698 17678 18713 23638
rect 18805 17678 18822 23638
rect 18822 17678 18856 23638
rect 18856 17678 18871 23638
rect 13930 17500 14000 17636
rect 18940 17636 18954 23680
rect 18954 17636 18992 23680
rect 18992 17636 19010 23680
rect 14152 17620 18786 17626
rect 14152 17586 14212 17620
rect 14212 17586 14302 17620
rect 14302 17586 14370 17620
rect 14370 17586 14460 17620
rect 14460 17586 14528 17620
rect 14528 17586 14618 17620
rect 14618 17586 14686 17620
rect 14686 17586 14776 17620
rect 14776 17586 14844 17620
rect 14844 17586 14934 17620
rect 14934 17586 15002 17620
rect 15002 17586 15092 17620
rect 15092 17586 15160 17620
rect 15160 17586 15250 17620
rect 15250 17586 15318 17620
rect 15318 17586 15408 17620
rect 15408 17586 15476 17620
rect 15476 17586 15566 17620
rect 15566 17586 15634 17620
rect 15634 17586 15724 17620
rect 15724 17586 15792 17620
rect 15792 17586 15882 17620
rect 15882 17586 15950 17620
rect 15950 17586 16040 17620
rect 16040 17586 16108 17620
rect 16108 17586 16198 17620
rect 16198 17586 16266 17620
rect 16266 17586 16356 17620
rect 16356 17586 16424 17620
rect 16424 17586 16514 17620
rect 16514 17586 16582 17620
rect 16582 17586 16672 17620
rect 16672 17586 16740 17620
rect 16740 17586 16830 17620
rect 16830 17586 16898 17620
rect 16898 17586 16988 17620
rect 16988 17586 17056 17620
rect 17056 17586 17146 17620
rect 17146 17586 17214 17620
rect 17214 17586 17304 17620
rect 17304 17586 17372 17620
rect 17372 17586 17462 17620
rect 17462 17586 17530 17620
rect 17530 17586 17620 17620
rect 17620 17586 17688 17620
rect 17688 17586 17778 17620
rect 17778 17586 17846 17620
rect 17846 17586 17936 17620
rect 17936 17586 18004 17620
rect 18004 17586 18094 17620
rect 18094 17586 18162 17620
rect 18162 17586 18252 17620
rect 18252 17586 18320 17620
rect 18320 17586 18410 17620
rect 18410 17586 18478 17620
rect 18478 17586 18568 17620
rect 18568 17586 18636 17620
rect 18636 17586 18726 17620
rect 18726 17586 18786 17620
rect 14152 17526 18786 17586
rect 18940 17500 19010 17636
rect 20230 23680 20300 23820
rect 20452 23730 25086 23790
rect 20452 23696 20512 23730
rect 20512 23696 20602 23730
rect 20602 23696 20670 23730
rect 20670 23696 20760 23730
rect 20760 23696 20828 23730
rect 20828 23696 20918 23730
rect 20918 23696 20986 23730
rect 20986 23696 21076 23730
rect 21076 23696 21144 23730
rect 21144 23696 21234 23730
rect 21234 23696 21302 23730
rect 21302 23696 21392 23730
rect 21392 23696 21460 23730
rect 21460 23696 21550 23730
rect 21550 23696 21618 23730
rect 21618 23696 21708 23730
rect 21708 23696 21776 23730
rect 21776 23696 21866 23730
rect 21866 23696 21934 23730
rect 21934 23696 22024 23730
rect 22024 23696 22092 23730
rect 22092 23696 22182 23730
rect 22182 23696 22250 23730
rect 22250 23696 22340 23730
rect 22340 23696 22408 23730
rect 22408 23696 22498 23730
rect 22498 23696 22566 23730
rect 22566 23696 22656 23730
rect 22656 23696 22724 23730
rect 22724 23696 22814 23730
rect 22814 23696 22882 23730
rect 22882 23696 22972 23730
rect 22972 23696 23040 23730
rect 23040 23696 23130 23730
rect 23130 23696 23198 23730
rect 23198 23696 23288 23730
rect 23288 23696 23356 23730
rect 23356 23696 23446 23730
rect 23446 23696 23514 23730
rect 23514 23696 23604 23730
rect 23604 23696 23672 23730
rect 23672 23696 23762 23730
rect 23762 23696 23830 23730
rect 23830 23696 23920 23730
rect 23920 23696 23988 23730
rect 23988 23696 24078 23730
rect 24078 23696 24146 23730
rect 24146 23696 24236 23730
rect 24236 23696 24304 23730
rect 24304 23696 24394 23730
rect 24394 23696 24462 23730
rect 24462 23696 24552 23730
rect 24552 23696 24620 23730
rect 24620 23696 24710 23730
rect 24710 23696 24778 23730
rect 24778 23696 24868 23730
rect 24868 23696 24936 23730
rect 24936 23696 25026 23730
rect 25026 23696 25086 23730
rect 20452 23690 25086 23696
rect 20230 17636 20246 23680
rect 20246 17636 20284 23680
rect 20284 17636 20300 23680
rect 25240 23680 25310 23820
rect 20365 17678 20382 23638
rect 20382 17678 20416 23638
rect 20416 17678 20431 23638
rect 20523 17678 20540 23638
rect 20540 17678 20574 23638
rect 20574 17678 20589 23638
rect 20681 17678 20698 23638
rect 20698 17678 20732 23638
rect 20732 17678 20747 23638
rect 20839 17678 20856 23638
rect 20856 17678 20890 23638
rect 20890 17678 20905 23638
rect 20997 17678 21014 23638
rect 21014 17678 21048 23638
rect 21048 17678 21063 23638
rect 21155 17678 21172 23638
rect 21172 17678 21206 23638
rect 21206 17678 21221 23638
rect 21313 17678 21330 23638
rect 21330 17678 21364 23638
rect 21364 17678 21379 23638
rect 21471 17678 21488 23638
rect 21488 17678 21522 23638
rect 21522 17678 21537 23638
rect 21629 17678 21646 23638
rect 21646 17678 21680 23638
rect 21680 17678 21695 23638
rect 21787 17678 21804 23638
rect 21804 17678 21838 23638
rect 21838 17678 21853 23638
rect 21945 17678 21962 23638
rect 21962 17678 21996 23638
rect 21996 17678 22011 23638
rect 22103 17678 22120 23638
rect 22120 17678 22154 23638
rect 22154 17678 22169 23638
rect 22261 17678 22278 23638
rect 22278 17678 22312 23638
rect 22312 17678 22327 23638
rect 22419 17678 22436 23638
rect 22436 17678 22470 23638
rect 22470 17678 22485 23638
rect 22577 17678 22594 23638
rect 22594 17678 22628 23638
rect 22628 17678 22643 23638
rect 22735 17678 22752 23638
rect 22752 17678 22786 23638
rect 22786 17678 22801 23638
rect 22893 17678 22910 23638
rect 22910 17678 22944 23638
rect 22944 17678 22959 23638
rect 23051 17678 23068 23638
rect 23068 17678 23102 23638
rect 23102 17678 23117 23638
rect 23209 17678 23226 23638
rect 23226 17678 23260 23638
rect 23260 17678 23275 23638
rect 23367 17678 23384 23638
rect 23384 17678 23418 23638
rect 23418 17678 23433 23638
rect 23525 17678 23542 23638
rect 23542 17678 23576 23638
rect 23576 17678 23591 23638
rect 23683 17678 23700 23638
rect 23700 17678 23734 23638
rect 23734 17678 23749 23638
rect 23841 17678 23858 23638
rect 23858 17678 23892 23638
rect 23892 17678 23907 23638
rect 23999 17678 24016 23638
rect 24016 17678 24050 23638
rect 24050 17678 24065 23638
rect 24157 17678 24174 23638
rect 24174 17678 24208 23638
rect 24208 17678 24223 23638
rect 24315 17678 24332 23638
rect 24332 17678 24366 23638
rect 24366 17678 24381 23638
rect 24473 17678 24490 23638
rect 24490 17678 24524 23638
rect 24524 17678 24539 23638
rect 24631 17678 24648 23638
rect 24648 17678 24682 23638
rect 24682 17678 24697 23638
rect 24789 17678 24806 23638
rect 24806 17678 24840 23638
rect 24840 17678 24855 23638
rect 24947 17678 24964 23638
rect 24964 17678 24998 23638
rect 24998 17678 25013 23638
rect 25105 17678 25122 23638
rect 25122 17678 25156 23638
rect 25156 17678 25171 23638
rect 20230 17500 20300 17636
rect 25240 17636 25254 23680
rect 25254 17636 25292 23680
rect 25292 17636 25310 23680
rect 25520 23650 25590 23850
rect 25910 23650 25980 23850
rect 26020 23650 26090 23850
rect 26410 23650 26480 23850
rect 25650 23520 25850 23590
rect 26150 23520 26350 23590
rect 25650 23410 25850 23480
rect 26150 23410 26350 23480
rect 25520 23150 25590 23350
rect 25910 23150 25980 23350
rect 26020 23150 26090 23350
rect 26410 23150 26480 23350
rect 25650 23020 25850 23090
rect 26150 23020 26350 23090
rect 25650 22910 25850 22980
rect 26150 22910 26350 22980
rect 25520 22650 25590 22850
rect 25910 22650 25980 22850
rect 26020 22650 26090 22850
rect 26410 22650 26480 22850
rect 25650 22520 25850 22590
rect 26150 22520 26350 22590
rect 25650 22410 25850 22480
rect 26150 22410 26350 22480
rect 25520 22150 25590 22350
rect 25910 22150 25980 22350
rect 26020 22150 26090 22350
rect 26410 22150 26480 22350
rect 25650 22020 25850 22090
rect 26150 22020 26350 22090
rect 25650 21910 25850 21980
rect 26150 21910 26350 21980
rect 25520 21650 25590 21850
rect 25910 21650 25980 21850
rect 26020 21650 26090 21850
rect 26410 21650 26480 21850
rect 25650 21520 25850 21590
rect 26150 21520 26350 21590
rect 25650 21410 25850 21480
rect 26150 21410 26350 21480
rect 25520 21150 25590 21350
rect 25910 21150 25980 21350
rect 26020 21150 26090 21350
rect 26410 21150 26480 21350
rect 25650 21020 25850 21090
rect 26150 21020 26350 21090
rect 25650 20910 25850 20980
rect 26150 20910 26350 20980
rect 25520 20650 25590 20850
rect 25910 20650 25980 20850
rect 26020 20650 26090 20850
rect 26410 20650 26480 20850
rect 25650 20520 25850 20590
rect 26150 20520 26350 20590
rect 25650 20410 25850 20480
rect 26150 20410 26350 20480
rect 25520 20150 25590 20350
rect 25910 20150 25980 20350
rect 26020 20150 26090 20350
rect 26410 20150 26480 20350
rect 25650 20020 25850 20090
rect 26150 20020 26350 20090
rect 25650 19910 25850 19980
rect 26150 19910 26350 19980
rect 25520 19650 25590 19850
rect 25910 19650 25980 19850
rect 26020 19650 26090 19850
rect 26410 19650 26480 19850
rect 25650 19520 25850 19590
rect 26150 19520 26350 19590
rect 25650 19410 25850 19480
rect 26150 19410 26350 19480
rect 25520 19150 25590 19350
rect 25910 19150 25980 19350
rect 26020 19150 26090 19350
rect 26410 19150 26480 19350
rect 25650 19020 25850 19090
rect 26150 19020 26350 19090
rect 25650 18910 25850 18980
rect 26150 18910 26350 18980
rect 25520 18650 25590 18850
rect 25910 18650 25980 18850
rect 26020 18650 26090 18850
rect 26410 18650 26480 18850
rect 25650 18520 25850 18590
rect 26150 18520 26350 18590
rect 25650 18410 25850 18480
rect 26150 18410 26350 18480
rect 25520 18150 25590 18350
rect 25910 18150 25980 18350
rect 26020 18150 26090 18350
rect 26410 18150 26480 18350
rect 25650 18020 25850 18090
rect 26150 18020 26350 18090
rect 25650 17910 25850 17980
rect 26150 17910 26350 17980
rect 25520 17650 25590 17850
rect 20452 17620 25086 17626
rect 20452 17586 20512 17620
rect 20512 17586 20602 17620
rect 20602 17586 20670 17620
rect 20670 17586 20760 17620
rect 20760 17586 20828 17620
rect 20828 17586 20918 17620
rect 20918 17586 20986 17620
rect 20986 17586 21076 17620
rect 21076 17586 21144 17620
rect 21144 17586 21234 17620
rect 21234 17586 21302 17620
rect 21302 17586 21392 17620
rect 21392 17586 21460 17620
rect 21460 17586 21550 17620
rect 21550 17586 21618 17620
rect 21618 17586 21708 17620
rect 21708 17586 21776 17620
rect 21776 17586 21866 17620
rect 21866 17586 21934 17620
rect 21934 17586 22024 17620
rect 22024 17586 22092 17620
rect 22092 17586 22182 17620
rect 22182 17586 22250 17620
rect 22250 17586 22340 17620
rect 22340 17586 22408 17620
rect 22408 17586 22498 17620
rect 22498 17586 22566 17620
rect 22566 17586 22656 17620
rect 22656 17586 22724 17620
rect 22724 17586 22814 17620
rect 22814 17586 22882 17620
rect 22882 17586 22972 17620
rect 22972 17586 23040 17620
rect 23040 17586 23130 17620
rect 23130 17586 23198 17620
rect 23198 17586 23288 17620
rect 23288 17586 23356 17620
rect 23356 17586 23446 17620
rect 23446 17586 23514 17620
rect 23514 17586 23604 17620
rect 23604 17586 23672 17620
rect 23672 17586 23762 17620
rect 23762 17586 23830 17620
rect 23830 17586 23920 17620
rect 23920 17586 23988 17620
rect 23988 17586 24078 17620
rect 24078 17586 24146 17620
rect 24146 17586 24236 17620
rect 24236 17586 24304 17620
rect 24304 17586 24394 17620
rect 24394 17586 24462 17620
rect 24462 17586 24552 17620
rect 24552 17586 24620 17620
rect 24620 17586 24710 17620
rect 24710 17586 24778 17620
rect 24778 17586 24868 17620
rect 24868 17586 24936 17620
rect 24936 17586 25026 17620
rect 25026 17586 25086 17620
rect 20452 17526 25086 17586
rect 6520 17150 6590 17350
rect 6910 17150 6980 17350
rect 7020 17150 7090 17350
rect 7410 17150 7480 17350
rect 6650 17020 6850 17090
rect 7150 17020 7350 17090
rect 13150 17410 13350 17480
rect 13650 17410 13850 17480
rect 13020 17150 13090 17350
rect 13410 17150 13480 17350
rect 13520 17150 13590 17350
rect 13910 17150 13980 17350
rect 13150 17020 13350 17090
rect 13650 17020 13850 17090
rect 19150 17410 19350 17480
rect 19650 17410 19850 17480
rect 25240 17500 25310 17636
rect 25910 17650 25980 17850
rect 26020 17650 26090 17850
rect 26410 17650 26480 17850
rect 25650 17520 25850 17590
rect 26150 17520 26350 17590
rect 19020 17150 19090 17350
rect 19410 17150 19480 17350
rect 19520 17150 19590 17350
rect 19910 17150 19980 17350
rect 19150 17020 19350 17090
rect 19650 17020 19850 17090
rect 25650 17410 25850 17480
rect 26150 17410 26350 17480
rect 25520 17150 25590 17350
rect 25910 17150 25980 17350
rect 26020 17150 26090 17350
rect 26410 17150 26480 17350
rect 25650 17020 25850 17090
rect 26150 17020 26350 17090
rect 150 16910 350 16980
rect 650 16910 850 16980
rect 1150 16910 1350 16980
rect 1650 16910 1850 16980
rect 2150 16910 2350 16980
rect 2650 16910 2850 16980
rect 3150 16910 3350 16980
rect 3650 16910 3850 16980
rect 4150 16910 4350 16980
rect 4650 16910 4850 16980
rect 5150 16910 5350 16980
rect 5650 16910 5850 16980
rect 6150 16910 6350 16980
rect 6650 16910 6850 16980
rect 7150 16910 7350 16980
rect 7650 16910 7850 16980
rect 8150 16910 8350 16980
rect 8650 16910 8850 16980
rect 9150 16910 9350 16980
rect 9650 16910 9850 16980
rect 10150 16910 10350 16980
rect 10650 16910 10850 16980
rect 11150 16910 11350 16980
rect 11650 16910 11850 16980
rect 12150 16910 12350 16980
rect 12650 16910 12850 16980
rect 13150 16910 13350 16980
rect 13650 16910 13850 16980
rect 14150 16910 14350 16980
rect 14650 16910 14850 16980
rect 15150 16910 15350 16980
rect 15650 16910 15850 16980
rect 16150 16910 16350 16980
rect 16650 16910 16850 16980
rect 17150 16910 17350 16980
rect 17650 16910 17850 16980
rect 18150 16910 18350 16980
rect 18650 16910 18850 16980
rect 19150 16910 19350 16980
rect 19650 16910 19850 16980
rect 20150 16910 20350 16980
rect 20650 16910 20850 16980
rect 21150 16910 21350 16980
rect 21650 16910 21850 16980
rect 22150 16910 22350 16980
rect 22650 16910 22850 16980
rect 23150 16910 23350 16980
rect 23650 16910 23850 16980
rect 24150 16910 24350 16980
rect 24650 16910 24850 16980
rect 25150 16910 25350 16980
rect 25650 16910 25850 16980
rect 26150 16910 26350 16980
rect 20 16650 90 16850
rect 410 16650 480 16850
rect 520 16650 590 16850
rect 910 16650 980 16850
rect 1020 16650 1090 16850
rect 1410 16650 1480 16850
rect 1520 16650 1590 16850
rect 1910 16650 1980 16850
rect 2020 16650 2090 16850
rect 2410 16650 2480 16850
rect 2520 16650 2590 16850
rect 2910 16650 2980 16850
rect 3020 16650 3090 16850
rect 3410 16650 3480 16850
rect 3520 16650 3590 16850
rect 3910 16650 3980 16850
rect 4020 16650 4090 16850
rect 4410 16650 4480 16850
rect 4520 16650 4590 16850
rect 4910 16650 4980 16850
rect 5020 16650 5090 16850
rect 5410 16650 5480 16850
rect 5520 16650 5590 16850
rect 5910 16650 5980 16850
rect 6020 16650 6090 16850
rect 6410 16650 6480 16850
rect 6520 16650 6590 16850
rect 6910 16650 6980 16850
rect 7020 16650 7090 16850
rect 7410 16650 7480 16850
rect 7520 16650 7590 16850
rect 7910 16650 7980 16850
rect 8020 16650 8090 16850
rect 8410 16650 8480 16850
rect 8520 16650 8590 16850
rect 8910 16650 8980 16850
rect 9020 16650 9090 16850
rect 9410 16650 9480 16850
rect 9520 16650 9590 16850
rect 9910 16650 9980 16850
rect 10020 16650 10090 16850
rect 10410 16650 10480 16850
rect 10520 16650 10590 16850
rect 10910 16650 10980 16850
rect 11020 16650 11090 16850
rect 11410 16650 11480 16850
rect 11520 16650 11590 16850
rect 11910 16650 11980 16850
rect 12020 16650 12090 16850
rect 12410 16650 12480 16850
rect 12520 16650 12590 16850
rect 12910 16650 12980 16850
rect 13020 16650 13090 16850
rect 13410 16650 13480 16850
rect 13520 16650 13590 16850
rect 13910 16650 13980 16850
rect 14020 16650 14090 16850
rect 14410 16650 14480 16850
rect 14520 16650 14590 16850
rect 14910 16650 14980 16850
rect 15020 16650 15090 16850
rect 15410 16650 15480 16850
rect 15520 16650 15590 16850
rect 15910 16650 15980 16850
rect 16020 16650 16090 16850
rect 16410 16650 16480 16850
rect 16520 16650 16590 16850
rect 16910 16650 16980 16850
rect 17020 16650 17090 16850
rect 17410 16650 17480 16850
rect 17520 16650 17590 16850
rect 17910 16650 17980 16850
rect 18020 16650 18090 16850
rect 18410 16650 18480 16850
rect 18520 16650 18590 16850
rect 18910 16650 18980 16850
rect 19020 16650 19090 16850
rect 19410 16650 19480 16850
rect 19520 16650 19590 16850
rect 19910 16650 19980 16850
rect 20020 16650 20090 16850
rect 20410 16650 20480 16850
rect 20520 16650 20590 16850
rect 20910 16650 20980 16850
rect 21020 16650 21090 16850
rect 21410 16650 21480 16850
rect 21520 16650 21590 16850
rect 21910 16650 21980 16850
rect 22020 16650 22090 16850
rect 22410 16650 22480 16850
rect 22520 16650 22590 16850
rect 22910 16650 22980 16850
rect 23020 16650 23090 16850
rect 23410 16650 23480 16850
rect 23520 16650 23590 16850
rect 23910 16650 23980 16850
rect 24020 16650 24090 16850
rect 24410 16650 24480 16850
rect 24520 16650 24590 16850
rect 24910 16650 24980 16850
rect 25020 16650 25090 16850
rect 25410 16650 25480 16850
rect 25520 16650 25590 16850
rect 25910 16650 25980 16850
rect 26020 16650 26090 16850
rect 26410 16650 26480 16850
rect 150 16520 350 16590
rect 650 16520 850 16590
rect 1150 16520 1350 16590
rect 1650 16520 1850 16590
rect 2150 16520 2350 16590
rect 2650 16520 2850 16590
rect 3150 16520 3350 16590
rect 3650 16520 3850 16590
rect 4150 16520 4350 16590
rect 4650 16520 4850 16590
rect 5150 16520 5350 16590
rect 5650 16520 5850 16590
rect 6150 16520 6350 16590
rect 6650 16520 6850 16590
rect 7150 16520 7350 16590
rect 7650 16520 7850 16590
rect 8150 16520 8350 16590
rect 8650 16520 8850 16590
rect 9150 16520 9350 16590
rect 9650 16520 9850 16590
rect 10150 16520 10350 16590
rect 10650 16520 10850 16590
rect 11150 16520 11350 16590
rect 11650 16520 11850 16590
rect 12150 16520 12350 16590
rect 12650 16520 12850 16590
rect 13150 16520 13350 16590
rect 13650 16520 13850 16590
rect 14150 16520 14350 16590
rect 14650 16520 14850 16590
rect 15150 16520 15350 16590
rect 15650 16520 15850 16590
rect 16150 16520 16350 16590
rect 16650 16520 16850 16590
rect 17150 16520 17350 16590
rect 17650 16520 17850 16590
rect 18150 16520 18350 16590
rect 18650 16520 18850 16590
rect 19150 16520 19350 16590
rect 19650 16520 19850 16590
rect 20150 16520 20350 16590
rect 20650 16520 20850 16590
rect 21150 16520 21350 16590
rect 21650 16520 21850 16590
rect 22150 16520 22350 16590
rect 22650 16520 22850 16590
rect 23150 16520 23350 16590
rect 23650 16520 23850 16590
rect 24150 16520 24350 16590
rect 24650 16520 24850 16590
rect 25150 16520 25350 16590
rect 25650 16520 25850 16590
rect 26150 16520 26350 16590
rect 150 16410 350 16480
rect 650 16410 850 16480
rect 1150 16410 1350 16480
rect 1650 16410 1850 16480
rect 2150 16410 2350 16480
rect 2650 16410 2850 16480
rect 3150 16410 3350 16480
rect 3650 16410 3850 16480
rect 4150 16410 4350 16480
rect 4650 16410 4850 16480
rect 5150 16410 5350 16480
rect 5650 16410 5850 16480
rect 6150 16410 6350 16480
rect 6650 16410 6850 16480
rect 7150 16410 7350 16480
rect 7650 16410 7850 16480
rect 8150 16410 8350 16480
rect 8650 16410 8850 16480
rect 9150 16410 9350 16480
rect 9650 16410 9850 16480
rect 10150 16410 10350 16480
rect 10650 16410 10850 16480
rect 11150 16410 11350 16480
rect 11650 16410 11850 16480
rect 12150 16410 12350 16480
rect 12650 16410 12850 16480
rect 13150 16410 13350 16480
rect 13650 16410 13850 16480
rect 14150 16410 14350 16480
rect 14650 16410 14850 16480
rect 15150 16410 15350 16480
rect 15650 16410 15850 16480
rect 16150 16410 16350 16480
rect 16650 16410 16850 16480
rect 17150 16410 17350 16480
rect 17650 16410 17850 16480
rect 18150 16410 18350 16480
rect 18650 16410 18850 16480
rect 19150 16410 19350 16480
rect 19650 16410 19850 16480
rect 20150 16410 20350 16480
rect 20650 16410 20850 16480
rect 21150 16410 21350 16480
rect 21650 16410 21850 16480
rect 22150 16410 22350 16480
rect 22650 16410 22850 16480
rect 23150 16410 23350 16480
rect 23650 16410 23850 16480
rect 24150 16410 24350 16480
rect 24650 16410 24850 16480
rect 25150 16410 25350 16480
rect 25650 16410 25850 16480
rect 26150 16410 26350 16480
rect 20 16150 90 16350
rect 410 16150 480 16350
rect 520 16150 590 16350
rect 910 16150 980 16350
rect 1020 16150 1090 16350
rect 1410 16150 1480 16350
rect 1520 16150 1590 16350
rect 1910 16150 1980 16350
rect 2020 16150 2090 16350
rect 2410 16150 2480 16350
rect 2520 16150 2590 16350
rect 2910 16150 2980 16350
rect 3020 16150 3090 16350
rect 3410 16150 3480 16350
rect 3520 16150 3590 16350
rect 3910 16150 3980 16350
rect 4020 16150 4090 16350
rect 4410 16150 4480 16350
rect 4520 16150 4590 16350
rect 4910 16150 4980 16350
rect 5020 16150 5090 16350
rect 5410 16150 5480 16350
rect 5520 16150 5590 16350
rect 5910 16150 5980 16350
rect 6020 16150 6090 16350
rect 6410 16150 6480 16350
rect 6520 16150 6590 16350
rect 6910 16150 6980 16350
rect 7020 16150 7090 16350
rect 7410 16150 7480 16350
rect 7520 16150 7590 16350
rect 7910 16150 7980 16350
rect 8020 16150 8090 16350
rect 8410 16150 8480 16350
rect 8520 16150 8590 16350
rect 8910 16150 8980 16350
rect 9020 16150 9090 16350
rect 9410 16150 9480 16350
rect 9520 16150 9590 16350
rect 9910 16150 9980 16350
rect 10020 16150 10090 16350
rect 10410 16150 10480 16350
rect 10520 16150 10590 16350
rect 10910 16150 10980 16350
rect 11020 16150 11090 16350
rect 11410 16150 11480 16350
rect 11520 16150 11590 16350
rect 11910 16150 11980 16350
rect 12020 16150 12090 16350
rect 12410 16150 12480 16350
rect 12520 16150 12590 16350
rect 12910 16150 12980 16350
rect 13020 16150 13090 16350
rect 13410 16150 13480 16350
rect 13520 16150 13590 16350
rect 13910 16150 13980 16350
rect 14020 16150 14090 16350
rect 14410 16150 14480 16350
rect 14520 16150 14590 16350
rect 14910 16150 14980 16350
rect 15020 16150 15090 16350
rect 15410 16150 15480 16350
rect 15520 16150 15590 16350
rect 15910 16150 15980 16350
rect 16020 16150 16090 16350
rect 16410 16150 16480 16350
rect 16520 16150 16590 16350
rect 16910 16150 16980 16350
rect 17020 16150 17090 16350
rect 17410 16150 17480 16350
rect 17520 16150 17590 16350
rect 17910 16150 17980 16350
rect 18020 16150 18090 16350
rect 18410 16150 18480 16350
rect 18520 16150 18590 16350
rect 18910 16150 18980 16350
rect 19020 16150 19090 16350
rect 19410 16150 19480 16350
rect 19520 16150 19590 16350
rect 19910 16150 19980 16350
rect 20020 16150 20090 16350
rect 20410 16150 20480 16350
rect 20520 16150 20590 16350
rect 20910 16150 20980 16350
rect 21020 16150 21090 16350
rect 21410 16150 21480 16350
rect 21520 16150 21590 16350
rect 21910 16150 21980 16350
rect 22020 16150 22090 16350
rect 22410 16150 22480 16350
rect 22520 16150 22590 16350
rect 22910 16150 22980 16350
rect 23020 16150 23090 16350
rect 23410 16150 23480 16350
rect 23520 16150 23590 16350
rect 23910 16150 23980 16350
rect 24020 16150 24090 16350
rect 24410 16150 24480 16350
rect 24520 16150 24590 16350
rect 24910 16150 24980 16350
rect 25020 16150 25090 16350
rect 25410 16150 25480 16350
rect 25520 16150 25590 16350
rect 25910 16150 25980 16350
rect 26020 16150 26090 16350
rect 26410 16150 26480 16350
rect 150 16020 350 16090
rect 650 16020 850 16090
rect 1150 16020 1350 16090
rect 1650 16020 1850 16090
rect 2150 16020 2350 16090
rect 2650 16020 2850 16090
rect 3150 16020 3350 16090
rect 3650 16020 3850 16090
rect 4150 16020 4350 16090
rect 4650 16020 4850 16090
rect 5150 16020 5350 16090
rect 5650 16020 5850 16090
rect 6150 16020 6350 16090
rect 6650 16020 6850 16090
rect 7150 16020 7350 16090
rect 7650 16020 7850 16090
rect 8150 16020 8350 16090
rect 8650 16020 8850 16090
rect 9150 16020 9350 16090
rect 9650 16020 9850 16090
rect 10150 16020 10350 16090
rect 10650 16020 10850 16090
rect 11150 16020 11350 16090
rect 11650 16020 11850 16090
rect 12150 16020 12350 16090
rect 12650 16020 12850 16090
rect 13150 16020 13350 16090
rect 13650 16020 13850 16090
rect 14150 16020 14350 16090
rect 14650 16020 14850 16090
rect 15150 16020 15350 16090
rect 15650 16020 15850 16090
rect 16150 16020 16350 16090
rect 16650 16020 16850 16090
rect 17150 16020 17350 16090
rect 17650 16020 17850 16090
rect 18150 16020 18350 16090
rect 18650 16020 18850 16090
rect 19150 16020 19350 16090
rect 19650 16020 19850 16090
rect 20150 16020 20350 16090
rect 20650 16020 20850 16090
rect 21150 16020 21350 16090
rect 21650 16020 21850 16090
rect 22150 16020 22350 16090
rect 22650 16020 22850 16090
rect 23150 16020 23350 16090
rect 23650 16020 23850 16090
rect 24150 16020 24350 16090
rect 24650 16020 24850 16090
rect 25150 16020 25350 16090
rect 25650 16020 25850 16090
rect 26150 16020 26350 16090
rect 150 15910 350 15980
rect 650 15910 850 15980
rect 20 15650 90 15850
rect 410 15650 480 15850
rect 520 15650 590 15850
rect 910 15650 980 15850
rect 150 15520 350 15590
rect 650 15520 850 15590
rect 6650 15910 6850 15980
rect 7150 15910 7350 15980
rect 6520 15650 6590 15850
rect 6910 15650 6980 15850
rect 7020 15650 7090 15850
rect 7410 15650 7480 15850
rect 150 15410 350 15480
rect 650 15410 850 15480
rect 1330 15380 1400 15520
rect 1552 15430 6186 15490
rect 1552 15396 1612 15430
rect 1612 15396 1702 15430
rect 1702 15396 1770 15430
rect 1770 15396 1860 15430
rect 1860 15396 1928 15430
rect 1928 15396 2018 15430
rect 2018 15396 2086 15430
rect 2086 15396 2176 15430
rect 2176 15396 2244 15430
rect 2244 15396 2334 15430
rect 2334 15396 2402 15430
rect 2402 15396 2492 15430
rect 2492 15396 2560 15430
rect 2560 15396 2650 15430
rect 2650 15396 2718 15430
rect 2718 15396 2808 15430
rect 2808 15396 2876 15430
rect 2876 15396 2966 15430
rect 2966 15396 3034 15430
rect 3034 15396 3124 15430
rect 3124 15396 3192 15430
rect 3192 15396 3282 15430
rect 3282 15396 3350 15430
rect 3350 15396 3440 15430
rect 3440 15396 3508 15430
rect 3508 15396 3598 15430
rect 3598 15396 3666 15430
rect 3666 15396 3756 15430
rect 3756 15396 3824 15430
rect 3824 15396 3914 15430
rect 3914 15396 3982 15430
rect 3982 15396 4072 15430
rect 4072 15396 4140 15430
rect 4140 15396 4230 15430
rect 4230 15396 4298 15430
rect 4298 15396 4388 15430
rect 4388 15396 4456 15430
rect 4456 15396 4546 15430
rect 4546 15396 4614 15430
rect 4614 15396 4704 15430
rect 4704 15396 4772 15430
rect 4772 15396 4862 15430
rect 4862 15396 4930 15430
rect 4930 15396 5020 15430
rect 5020 15396 5088 15430
rect 5088 15396 5178 15430
rect 5178 15396 5246 15430
rect 5246 15396 5336 15430
rect 5336 15396 5404 15430
rect 5404 15396 5494 15430
rect 5494 15396 5562 15430
rect 5562 15396 5652 15430
rect 5652 15396 5720 15430
rect 5720 15396 5810 15430
rect 5810 15396 5878 15430
rect 5878 15396 5968 15430
rect 5968 15396 6036 15430
rect 6036 15396 6126 15430
rect 6126 15396 6186 15430
rect 1552 15390 6186 15396
rect 20 15150 90 15350
rect 410 15150 480 15350
rect 520 15150 590 15350
rect 910 15150 980 15350
rect 150 15020 350 15090
rect 650 15020 850 15090
rect 150 14910 350 14980
rect 650 14910 850 14980
rect 20 14650 90 14850
rect 410 14650 480 14850
rect 520 14650 590 14850
rect 910 14650 980 14850
rect 150 14520 350 14590
rect 650 14520 850 14590
rect 150 14410 350 14480
rect 650 14410 850 14480
rect 20 14150 90 14350
rect 410 14150 480 14350
rect 520 14150 590 14350
rect 910 14150 980 14350
rect 150 14020 350 14090
rect 650 14020 850 14090
rect -4290 13832 -4110 13900
rect -4290 13435 -4218 13832
rect -4218 13435 -4180 13832
rect -4180 13435 -4110 13832
rect -4290 13420 -4110 13435
rect -4290 13081 -4110 13090
rect -4290 12684 -4218 13081
rect -4218 12684 -4180 13081
rect -4180 12684 -4110 13081
rect -4290 12610 -4110 12684
rect -3850 13910 -3650 13980
rect -3350 13910 -3150 13980
rect -2850 13910 -2650 13980
rect -2350 13910 -2150 13980
rect -1850 13910 -1650 13980
rect -1350 13910 -1150 13980
rect -850 13910 -650 13980
rect -350 13910 -150 13980
rect 150 13910 350 13980
rect 650 13910 850 13980
rect -3980 13650 -3910 13850
rect -3590 13650 -3520 13850
rect -3480 13650 -3410 13850
rect -3090 13650 -3020 13850
rect -2980 13650 -2910 13850
rect -2590 13650 -2520 13850
rect -2480 13650 -2410 13850
rect -2090 13650 -2020 13850
rect -1980 13650 -1910 13850
rect -1590 13650 -1520 13850
rect -1480 13650 -1410 13850
rect -1090 13650 -1020 13850
rect -980 13650 -910 13850
rect -590 13650 -520 13850
rect -480 13650 -410 13850
rect -90 13650 -20 13850
rect 20 13650 90 13850
rect 410 13650 480 13850
rect 520 13650 590 13850
rect 910 13650 980 13850
rect -3850 13520 -3650 13590
rect -3350 13520 -3150 13590
rect -2850 13520 -2650 13590
rect -2350 13520 -2150 13590
rect -1850 13520 -1650 13590
rect -1350 13520 -1150 13590
rect -850 13520 -650 13590
rect -350 13520 -150 13590
rect 150 13520 350 13590
rect 650 13520 850 13590
rect -3850 13410 -3650 13480
rect -3350 13410 -3150 13480
rect -2850 13410 -2650 13480
rect -2350 13410 -2150 13480
rect -1850 13410 -1650 13480
rect -1350 13410 -1150 13480
rect -850 13410 -650 13480
rect -350 13410 -150 13480
rect 150 13410 350 13480
rect 650 13410 850 13480
rect -3980 13150 -3910 13350
rect -3590 13150 -3520 13350
rect -3480 13150 -3410 13350
rect -3090 13150 -3020 13350
rect -2980 13150 -2910 13350
rect -2590 13150 -2520 13350
rect -2480 13150 -2410 13350
rect -2090 13150 -2020 13350
rect -1980 13150 -1910 13350
rect -1590 13150 -1520 13350
rect -1480 13150 -1410 13350
rect -1090 13150 -1020 13350
rect -980 13150 -910 13350
rect -590 13150 -520 13350
rect -480 13150 -410 13350
rect -90 13150 -20 13350
rect 20 13150 90 13350
rect 410 13150 480 13350
rect 520 13150 590 13350
rect 910 13150 980 13350
rect -3850 13020 -3650 13090
rect -3350 13020 -3150 13090
rect -2850 13020 -2650 13090
rect -2350 13020 -2150 13090
rect -1850 13020 -1650 13090
rect -1350 13020 -1150 13090
rect -850 13020 -650 13090
rect -350 13020 -150 13090
rect 150 13020 350 13090
rect 650 13020 850 13090
rect 150 12910 350 12980
rect 650 12910 850 12980
rect 20 12650 90 12850
rect 410 12650 480 12850
rect 520 12650 590 12850
rect 910 12650 980 12850
rect 150 12520 350 12590
rect 650 12520 850 12590
rect 150 12410 350 12480
rect 650 12410 850 12480
rect 20 12150 90 12350
rect 410 12150 480 12350
rect 520 12150 590 12350
rect 910 12150 980 12350
rect 150 12020 350 12090
rect 650 12020 850 12090
rect 150 11910 350 11980
rect 650 11910 850 11980
rect 20 11650 90 11850
rect 410 11650 480 11850
rect 520 11650 590 11850
rect 910 11650 980 11850
rect 150 11520 350 11590
rect 650 11520 850 11590
rect 150 11410 350 11480
rect 650 11410 850 11480
rect 20 11150 90 11350
rect 410 11150 480 11350
rect 520 11150 590 11350
rect 910 11150 980 11350
rect 150 11020 350 11090
rect 650 11020 850 11090
rect 150 10910 350 10980
rect 650 10910 850 10980
rect 20 10650 90 10850
rect 410 10650 480 10850
rect 520 10650 590 10850
rect 910 10650 980 10850
rect 150 10520 350 10590
rect 650 10520 850 10590
rect 150 10410 350 10480
rect 650 10410 850 10480
rect 20 10150 90 10350
rect 410 10150 480 10350
rect 520 10150 590 10350
rect 910 10150 980 10350
rect 150 10020 350 10090
rect 650 10020 850 10090
rect 150 9910 350 9980
rect 650 9910 850 9980
rect 20 9650 90 9850
rect 410 9650 480 9850
rect 520 9650 590 9850
rect 910 9650 980 9850
rect 150 9520 350 9590
rect 650 9520 850 9590
rect 150 9410 350 9480
rect 650 9410 850 9480
rect 20 9150 90 9350
rect 410 9150 480 9350
rect 520 9150 590 9350
rect 910 9150 980 9350
rect 1330 9336 1346 15380
rect 1346 9336 1384 15380
rect 1384 9336 1400 15380
rect 6340 15380 6410 15520
rect 6650 15520 6850 15590
rect 7150 15520 7350 15590
rect 13150 15910 13350 15980
rect 13650 15910 13850 15980
rect 13020 15650 13090 15850
rect 13410 15650 13480 15850
rect 13520 15650 13590 15850
rect 13910 15650 13980 15850
rect 1465 9378 1482 15338
rect 1482 9378 1516 15338
rect 1516 9378 1531 15338
rect 1623 9378 1640 15338
rect 1640 9378 1674 15338
rect 1674 9378 1689 15338
rect 1781 9378 1798 15338
rect 1798 9378 1832 15338
rect 1832 9378 1847 15338
rect 1939 9378 1956 15338
rect 1956 9378 1990 15338
rect 1990 9378 2005 15338
rect 2097 9378 2114 15338
rect 2114 9378 2148 15338
rect 2148 9378 2163 15338
rect 2255 9378 2272 15338
rect 2272 9378 2306 15338
rect 2306 9378 2321 15338
rect 2413 9378 2430 15338
rect 2430 9378 2464 15338
rect 2464 9378 2479 15338
rect 2571 9378 2588 15338
rect 2588 9378 2622 15338
rect 2622 9378 2637 15338
rect 2729 9378 2746 15338
rect 2746 9378 2780 15338
rect 2780 9378 2795 15338
rect 2887 9378 2904 15338
rect 2904 9378 2938 15338
rect 2938 9378 2953 15338
rect 3045 9378 3062 15338
rect 3062 9378 3096 15338
rect 3096 9378 3111 15338
rect 3203 9378 3220 15338
rect 3220 9378 3254 15338
rect 3254 9378 3269 15338
rect 3361 9378 3378 15338
rect 3378 9378 3412 15338
rect 3412 9378 3427 15338
rect 3519 9378 3536 15338
rect 3536 9378 3570 15338
rect 3570 9378 3585 15338
rect 3677 9378 3694 15338
rect 3694 9378 3728 15338
rect 3728 9378 3743 15338
rect 3835 9378 3852 15338
rect 3852 9378 3886 15338
rect 3886 9378 3901 15338
rect 3993 9378 4010 15338
rect 4010 9378 4044 15338
rect 4044 9378 4059 15338
rect 4151 9378 4168 15338
rect 4168 9378 4202 15338
rect 4202 9378 4217 15338
rect 4309 9378 4326 15338
rect 4326 9378 4360 15338
rect 4360 9378 4375 15338
rect 4467 9378 4484 15338
rect 4484 9378 4518 15338
rect 4518 9378 4533 15338
rect 4625 9378 4642 15338
rect 4642 9378 4676 15338
rect 4676 9378 4691 15338
rect 4783 9378 4800 15338
rect 4800 9378 4834 15338
rect 4834 9378 4849 15338
rect 4941 9378 4958 15338
rect 4958 9378 4992 15338
rect 4992 9378 5007 15338
rect 5099 9378 5116 15338
rect 5116 9378 5150 15338
rect 5150 9378 5165 15338
rect 5257 9378 5274 15338
rect 5274 9378 5308 15338
rect 5308 9378 5323 15338
rect 5415 9378 5432 15338
rect 5432 9378 5466 15338
rect 5466 9378 5481 15338
rect 5573 9378 5590 15338
rect 5590 9378 5624 15338
rect 5624 9378 5639 15338
rect 5731 9378 5748 15338
rect 5748 9378 5782 15338
rect 5782 9378 5797 15338
rect 5889 9378 5906 15338
rect 5906 9378 5940 15338
rect 5940 9378 5955 15338
rect 6047 9378 6064 15338
rect 6064 9378 6098 15338
rect 6098 9378 6113 15338
rect 6205 9378 6222 15338
rect 6222 9378 6256 15338
rect 6256 9378 6271 15338
rect 1330 9200 1400 9336
rect 6340 9336 6354 15380
rect 6354 9336 6392 15380
rect 6392 9336 6410 15380
rect 1552 9320 6186 9326
rect 1552 9286 1612 9320
rect 1612 9286 1702 9320
rect 1702 9286 1770 9320
rect 1770 9286 1860 9320
rect 1860 9286 1928 9320
rect 1928 9286 2018 9320
rect 2018 9286 2086 9320
rect 2086 9286 2176 9320
rect 2176 9286 2244 9320
rect 2244 9286 2334 9320
rect 2334 9286 2402 9320
rect 2402 9286 2492 9320
rect 2492 9286 2560 9320
rect 2560 9286 2650 9320
rect 2650 9286 2718 9320
rect 2718 9286 2808 9320
rect 2808 9286 2876 9320
rect 2876 9286 2966 9320
rect 2966 9286 3034 9320
rect 3034 9286 3124 9320
rect 3124 9286 3192 9320
rect 3192 9286 3282 9320
rect 3282 9286 3350 9320
rect 3350 9286 3440 9320
rect 3440 9286 3508 9320
rect 3508 9286 3598 9320
rect 3598 9286 3666 9320
rect 3666 9286 3756 9320
rect 3756 9286 3824 9320
rect 3824 9286 3914 9320
rect 3914 9286 3982 9320
rect 3982 9286 4072 9320
rect 4072 9286 4140 9320
rect 4140 9286 4230 9320
rect 4230 9286 4298 9320
rect 4298 9286 4388 9320
rect 4388 9286 4456 9320
rect 4456 9286 4546 9320
rect 4546 9286 4614 9320
rect 4614 9286 4704 9320
rect 4704 9286 4772 9320
rect 4772 9286 4862 9320
rect 4862 9286 4930 9320
rect 4930 9286 5020 9320
rect 5020 9286 5088 9320
rect 5088 9286 5178 9320
rect 5178 9286 5246 9320
rect 5246 9286 5336 9320
rect 5336 9286 5404 9320
rect 5404 9286 5494 9320
rect 5494 9286 5562 9320
rect 5562 9286 5652 9320
rect 5652 9286 5720 9320
rect 5720 9286 5810 9320
rect 5810 9286 5878 9320
rect 5878 9286 5968 9320
rect 5968 9286 6036 9320
rect 6036 9286 6126 9320
rect 6126 9286 6186 9320
rect 1552 9226 6186 9286
rect 6340 9200 6410 9336
rect 7630 15380 7700 15520
rect 7852 15430 12486 15490
rect 7852 15396 7912 15430
rect 7912 15396 8002 15430
rect 8002 15396 8070 15430
rect 8070 15396 8160 15430
rect 8160 15396 8228 15430
rect 8228 15396 8318 15430
rect 8318 15396 8386 15430
rect 8386 15396 8476 15430
rect 8476 15396 8544 15430
rect 8544 15396 8634 15430
rect 8634 15396 8702 15430
rect 8702 15396 8792 15430
rect 8792 15396 8860 15430
rect 8860 15396 8950 15430
rect 8950 15396 9018 15430
rect 9018 15396 9108 15430
rect 9108 15396 9176 15430
rect 9176 15396 9266 15430
rect 9266 15396 9334 15430
rect 9334 15396 9424 15430
rect 9424 15396 9492 15430
rect 9492 15396 9582 15430
rect 9582 15396 9650 15430
rect 9650 15396 9740 15430
rect 9740 15396 9808 15430
rect 9808 15396 9898 15430
rect 9898 15396 9966 15430
rect 9966 15396 10056 15430
rect 10056 15396 10124 15430
rect 10124 15396 10214 15430
rect 10214 15396 10282 15430
rect 10282 15396 10372 15430
rect 10372 15396 10440 15430
rect 10440 15396 10530 15430
rect 10530 15396 10598 15430
rect 10598 15396 10688 15430
rect 10688 15396 10756 15430
rect 10756 15396 10846 15430
rect 10846 15396 10914 15430
rect 10914 15396 11004 15430
rect 11004 15396 11072 15430
rect 11072 15396 11162 15430
rect 11162 15396 11230 15430
rect 11230 15396 11320 15430
rect 11320 15396 11388 15430
rect 11388 15396 11478 15430
rect 11478 15396 11546 15430
rect 11546 15396 11636 15430
rect 11636 15396 11704 15430
rect 11704 15396 11794 15430
rect 11794 15396 11862 15430
rect 11862 15396 11952 15430
rect 11952 15396 12020 15430
rect 12020 15396 12110 15430
rect 12110 15396 12178 15430
rect 12178 15396 12268 15430
rect 12268 15396 12336 15430
rect 12336 15396 12426 15430
rect 12426 15396 12486 15430
rect 7852 15390 12486 15396
rect 7630 9336 7646 15380
rect 7646 9336 7684 15380
rect 7684 9336 7700 15380
rect 12640 15380 12710 15520
rect 13150 15520 13350 15590
rect 13650 15520 13850 15590
rect 19150 15910 19350 15980
rect 19650 15910 19850 15980
rect 19020 15650 19090 15850
rect 19410 15650 19480 15850
rect 19520 15650 19590 15850
rect 19910 15650 19980 15850
rect 7765 9378 7782 15338
rect 7782 9378 7816 15338
rect 7816 9378 7831 15338
rect 7923 9378 7940 15338
rect 7940 9378 7974 15338
rect 7974 9378 7989 15338
rect 8081 9378 8098 15338
rect 8098 9378 8132 15338
rect 8132 9378 8147 15338
rect 8239 9378 8256 15338
rect 8256 9378 8290 15338
rect 8290 9378 8305 15338
rect 8397 9378 8414 15338
rect 8414 9378 8448 15338
rect 8448 9378 8463 15338
rect 8555 9378 8572 15338
rect 8572 9378 8606 15338
rect 8606 9378 8621 15338
rect 8713 9378 8730 15338
rect 8730 9378 8764 15338
rect 8764 9378 8779 15338
rect 8871 9378 8888 15338
rect 8888 9378 8922 15338
rect 8922 9378 8937 15338
rect 9029 9378 9046 15338
rect 9046 9378 9080 15338
rect 9080 9378 9095 15338
rect 9187 9378 9204 15338
rect 9204 9378 9238 15338
rect 9238 9378 9253 15338
rect 9345 9378 9362 15338
rect 9362 9378 9396 15338
rect 9396 9378 9411 15338
rect 9503 9378 9520 15338
rect 9520 9378 9554 15338
rect 9554 9378 9569 15338
rect 9661 9378 9678 15338
rect 9678 9378 9712 15338
rect 9712 9378 9727 15338
rect 9819 9378 9836 15338
rect 9836 9378 9870 15338
rect 9870 9378 9885 15338
rect 9977 9378 9994 15338
rect 9994 9378 10028 15338
rect 10028 9378 10043 15338
rect 10135 9378 10152 15338
rect 10152 9378 10186 15338
rect 10186 9378 10201 15338
rect 10293 9378 10310 15338
rect 10310 9378 10344 15338
rect 10344 9378 10359 15338
rect 10451 9378 10468 15338
rect 10468 9378 10502 15338
rect 10502 9378 10517 15338
rect 10609 9378 10626 15338
rect 10626 9378 10660 15338
rect 10660 9378 10675 15338
rect 10767 9378 10784 15338
rect 10784 9378 10818 15338
rect 10818 9378 10833 15338
rect 10925 9378 10942 15338
rect 10942 9378 10976 15338
rect 10976 9378 10991 15338
rect 11083 9378 11100 15338
rect 11100 9378 11134 15338
rect 11134 9378 11149 15338
rect 11241 9378 11258 15338
rect 11258 9378 11292 15338
rect 11292 9378 11307 15338
rect 11399 9378 11416 15338
rect 11416 9378 11450 15338
rect 11450 9378 11465 15338
rect 11557 9378 11574 15338
rect 11574 9378 11608 15338
rect 11608 9378 11623 15338
rect 11715 9378 11732 15338
rect 11732 9378 11766 15338
rect 11766 9378 11781 15338
rect 11873 9378 11890 15338
rect 11890 9378 11924 15338
rect 11924 9378 11939 15338
rect 12031 9378 12048 15338
rect 12048 9378 12082 15338
rect 12082 9378 12097 15338
rect 12189 9378 12206 15338
rect 12206 9378 12240 15338
rect 12240 9378 12255 15338
rect 12347 9378 12364 15338
rect 12364 9378 12398 15338
rect 12398 9378 12413 15338
rect 12505 9378 12522 15338
rect 12522 9378 12556 15338
rect 12556 9378 12571 15338
rect 7630 9200 7700 9336
rect 12640 9336 12654 15380
rect 12654 9336 12692 15380
rect 12692 9336 12710 15380
rect 7852 9320 12486 9326
rect 7852 9286 7912 9320
rect 7912 9286 8002 9320
rect 8002 9286 8070 9320
rect 8070 9286 8160 9320
rect 8160 9286 8228 9320
rect 8228 9286 8318 9320
rect 8318 9286 8386 9320
rect 8386 9286 8476 9320
rect 8476 9286 8544 9320
rect 8544 9286 8634 9320
rect 8634 9286 8702 9320
rect 8702 9286 8792 9320
rect 8792 9286 8860 9320
rect 8860 9286 8950 9320
rect 8950 9286 9018 9320
rect 9018 9286 9108 9320
rect 9108 9286 9176 9320
rect 9176 9286 9266 9320
rect 9266 9286 9334 9320
rect 9334 9286 9424 9320
rect 9424 9286 9492 9320
rect 9492 9286 9582 9320
rect 9582 9286 9650 9320
rect 9650 9286 9740 9320
rect 9740 9286 9808 9320
rect 9808 9286 9898 9320
rect 9898 9286 9966 9320
rect 9966 9286 10056 9320
rect 10056 9286 10124 9320
rect 10124 9286 10214 9320
rect 10214 9286 10282 9320
rect 10282 9286 10372 9320
rect 10372 9286 10440 9320
rect 10440 9286 10530 9320
rect 10530 9286 10598 9320
rect 10598 9286 10688 9320
rect 10688 9286 10756 9320
rect 10756 9286 10846 9320
rect 10846 9286 10914 9320
rect 10914 9286 11004 9320
rect 11004 9286 11072 9320
rect 11072 9286 11162 9320
rect 11162 9286 11230 9320
rect 11230 9286 11320 9320
rect 11320 9286 11388 9320
rect 11388 9286 11478 9320
rect 11478 9286 11546 9320
rect 11546 9286 11636 9320
rect 11636 9286 11704 9320
rect 11704 9286 11794 9320
rect 11794 9286 11862 9320
rect 11862 9286 11952 9320
rect 11952 9286 12020 9320
rect 12020 9286 12110 9320
rect 12110 9286 12178 9320
rect 12178 9286 12268 9320
rect 12268 9286 12336 9320
rect 12336 9286 12426 9320
rect 12426 9286 12486 9320
rect 7852 9226 12486 9286
rect 12640 9200 12710 9336
rect 13930 15380 14000 15520
rect 19150 15520 19350 15590
rect 19650 15520 19850 15590
rect 25650 15910 25850 15980
rect 26150 15910 26350 15980
rect 25520 15650 25590 15850
rect 25910 15650 25980 15850
rect 26020 15650 26090 15850
rect 26410 15650 26480 15850
rect 14152 15430 18786 15490
rect 14152 15396 14212 15430
rect 14212 15396 14302 15430
rect 14302 15396 14370 15430
rect 14370 15396 14460 15430
rect 14460 15396 14528 15430
rect 14528 15396 14618 15430
rect 14618 15396 14686 15430
rect 14686 15396 14776 15430
rect 14776 15396 14844 15430
rect 14844 15396 14934 15430
rect 14934 15396 15002 15430
rect 15002 15396 15092 15430
rect 15092 15396 15160 15430
rect 15160 15396 15250 15430
rect 15250 15396 15318 15430
rect 15318 15396 15408 15430
rect 15408 15396 15476 15430
rect 15476 15396 15566 15430
rect 15566 15396 15634 15430
rect 15634 15396 15724 15430
rect 15724 15396 15792 15430
rect 15792 15396 15882 15430
rect 15882 15396 15950 15430
rect 15950 15396 16040 15430
rect 16040 15396 16108 15430
rect 16108 15396 16198 15430
rect 16198 15396 16266 15430
rect 16266 15396 16356 15430
rect 16356 15396 16424 15430
rect 16424 15396 16514 15430
rect 16514 15396 16582 15430
rect 16582 15396 16672 15430
rect 16672 15396 16740 15430
rect 16740 15396 16830 15430
rect 16830 15396 16898 15430
rect 16898 15396 16988 15430
rect 16988 15396 17056 15430
rect 17056 15396 17146 15430
rect 17146 15396 17214 15430
rect 17214 15396 17304 15430
rect 17304 15396 17372 15430
rect 17372 15396 17462 15430
rect 17462 15396 17530 15430
rect 17530 15396 17620 15430
rect 17620 15396 17688 15430
rect 17688 15396 17778 15430
rect 17778 15396 17846 15430
rect 17846 15396 17936 15430
rect 17936 15396 18004 15430
rect 18004 15396 18094 15430
rect 18094 15396 18162 15430
rect 18162 15396 18252 15430
rect 18252 15396 18320 15430
rect 18320 15396 18410 15430
rect 18410 15396 18478 15430
rect 18478 15396 18568 15430
rect 18568 15396 18636 15430
rect 18636 15396 18726 15430
rect 18726 15396 18786 15430
rect 14152 15390 18786 15396
rect 13930 9336 13946 15380
rect 13946 9336 13984 15380
rect 13984 9336 14000 15380
rect 18940 15380 19010 15520
rect 14065 9378 14082 15338
rect 14082 9378 14116 15338
rect 14116 9378 14131 15338
rect 14223 9378 14240 15338
rect 14240 9378 14274 15338
rect 14274 9378 14289 15338
rect 14381 9378 14398 15338
rect 14398 9378 14432 15338
rect 14432 9378 14447 15338
rect 14539 9378 14556 15338
rect 14556 9378 14590 15338
rect 14590 9378 14605 15338
rect 14697 9378 14714 15338
rect 14714 9378 14748 15338
rect 14748 9378 14763 15338
rect 14855 9378 14872 15338
rect 14872 9378 14906 15338
rect 14906 9378 14921 15338
rect 15013 9378 15030 15338
rect 15030 9378 15064 15338
rect 15064 9378 15079 15338
rect 15171 9378 15188 15338
rect 15188 9378 15222 15338
rect 15222 9378 15237 15338
rect 15329 9378 15346 15338
rect 15346 9378 15380 15338
rect 15380 9378 15395 15338
rect 15487 9378 15504 15338
rect 15504 9378 15538 15338
rect 15538 9378 15553 15338
rect 15645 9378 15662 15338
rect 15662 9378 15696 15338
rect 15696 9378 15711 15338
rect 15803 9378 15820 15338
rect 15820 9378 15854 15338
rect 15854 9378 15869 15338
rect 15961 9378 15978 15338
rect 15978 9378 16012 15338
rect 16012 9378 16027 15338
rect 16119 9378 16136 15338
rect 16136 9378 16170 15338
rect 16170 9378 16185 15338
rect 16277 9378 16294 15338
rect 16294 9378 16328 15338
rect 16328 9378 16343 15338
rect 16435 9378 16452 15338
rect 16452 9378 16486 15338
rect 16486 9378 16501 15338
rect 16593 9378 16610 15338
rect 16610 9378 16644 15338
rect 16644 9378 16659 15338
rect 16751 9378 16768 15338
rect 16768 9378 16802 15338
rect 16802 9378 16817 15338
rect 16909 9378 16926 15338
rect 16926 9378 16960 15338
rect 16960 9378 16975 15338
rect 17067 9378 17084 15338
rect 17084 9378 17118 15338
rect 17118 9378 17133 15338
rect 17225 9378 17242 15338
rect 17242 9378 17276 15338
rect 17276 9378 17291 15338
rect 17383 9378 17400 15338
rect 17400 9378 17434 15338
rect 17434 9378 17449 15338
rect 17541 9378 17558 15338
rect 17558 9378 17592 15338
rect 17592 9378 17607 15338
rect 17699 9378 17716 15338
rect 17716 9378 17750 15338
rect 17750 9378 17765 15338
rect 17857 9378 17874 15338
rect 17874 9378 17908 15338
rect 17908 9378 17923 15338
rect 18015 9378 18032 15338
rect 18032 9378 18066 15338
rect 18066 9378 18081 15338
rect 18173 9378 18190 15338
rect 18190 9378 18224 15338
rect 18224 9378 18239 15338
rect 18331 9378 18348 15338
rect 18348 9378 18382 15338
rect 18382 9378 18397 15338
rect 18489 9378 18506 15338
rect 18506 9378 18540 15338
rect 18540 9378 18555 15338
rect 18647 9378 18664 15338
rect 18664 9378 18698 15338
rect 18698 9378 18713 15338
rect 18805 9378 18822 15338
rect 18822 9378 18856 15338
rect 18856 9378 18871 15338
rect 13930 9200 14000 9336
rect 18940 9336 18954 15380
rect 18954 9336 18992 15380
rect 18992 9336 19010 15380
rect 14152 9320 18786 9326
rect 14152 9286 14212 9320
rect 14212 9286 14302 9320
rect 14302 9286 14370 9320
rect 14370 9286 14460 9320
rect 14460 9286 14528 9320
rect 14528 9286 14618 9320
rect 14618 9286 14686 9320
rect 14686 9286 14776 9320
rect 14776 9286 14844 9320
rect 14844 9286 14934 9320
rect 14934 9286 15002 9320
rect 15002 9286 15092 9320
rect 15092 9286 15160 9320
rect 15160 9286 15250 9320
rect 15250 9286 15318 9320
rect 15318 9286 15408 9320
rect 15408 9286 15476 9320
rect 15476 9286 15566 9320
rect 15566 9286 15634 9320
rect 15634 9286 15724 9320
rect 15724 9286 15792 9320
rect 15792 9286 15882 9320
rect 15882 9286 15950 9320
rect 15950 9286 16040 9320
rect 16040 9286 16108 9320
rect 16108 9286 16198 9320
rect 16198 9286 16266 9320
rect 16266 9286 16356 9320
rect 16356 9286 16424 9320
rect 16424 9286 16514 9320
rect 16514 9286 16582 9320
rect 16582 9286 16672 9320
rect 16672 9286 16740 9320
rect 16740 9286 16830 9320
rect 16830 9286 16898 9320
rect 16898 9286 16988 9320
rect 16988 9286 17056 9320
rect 17056 9286 17146 9320
rect 17146 9286 17214 9320
rect 17214 9286 17304 9320
rect 17304 9286 17372 9320
rect 17372 9286 17462 9320
rect 17462 9286 17530 9320
rect 17530 9286 17620 9320
rect 17620 9286 17688 9320
rect 17688 9286 17778 9320
rect 17778 9286 17846 9320
rect 17846 9286 17936 9320
rect 17936 9286 18004 9320
rect 18004 9286 18094 9320
rect 18094 9286 18162 9320
rect 18162 9286 18252 9320
rect 18252 9286 18320 9320
rect 18320 9286 18410 9320
rect 18410 9286 18478 9320
rect 18478 9286 18568 9320
rect 18568 9286 18636 9320
rect 18636 9286 18726 9320
rect 18726 9286 18786 9320
rect 14152 9226 18786 9286
rect 18940 9200 19010 9336
rect 20230 15380 20300 15520
rect 25650 15520 25850 15590
rect 26150 15520 26350 15590
rect 20452 15430 25086 15490
rect 20452 15396 20512 15430
rect 20512 15396 20602 15430
rect 20602 15396 20670 15430
rect 20670 15396 20760 15430
rect 20760 15396 20828 15430
rect 20828 15396 20918 15430
rect 20918 15396 20986 15430
rect 20986 15396 21076 15430
rect 21076 15396 21144 15430
rect 21144 15396 21234 15430
rect 21234 15396 21302 15430
rect 21302 15396 21392 15430
rect 21392 15396 21460 15430
rect 21460 15396 21550 15430
rect 21550 15396 21618 15430
rect 21618 15396 21708 15430
rect 21708 15396 21776 15430
rect 21776 15396 21866 15430
rect 21866 15396 21934 15430
rect 21934 15396 22024 15430
rect 22024 15396 22092 15430
rect 22092 15396 22182 15430
rect 22182 15396 22250 15430
rect 22250 15396 22340 15430
rect 22340 15396 22408 15430
rect 22408 15396 22498 15430
rect 22498 15396 22566 15430
rect 22566 15396 22656 15430
rect 22656 15396 22724 15430
rect 22724 15396 22814 15430
rect 22814 15396 22882 15430
rect 22882 15396 22972 15430
rect 22972 15396 23040 15430
rect 23040 15396 23130 15430
rect 23130 15396 23198 15430
rect 23198 15396 23288 15430
rect 23288 15396 23356 15430
rect 23356 15396 23446 15430
rect 23446 15396 23514 15430
rect 23514 15396 23604 15430
rect 23604 15396 23672 15430
rect 23672 15396 23762 15430
rect 23762 15396 23830 15430
rect 23830 15396 23920 15430
rect 23920 15396 23988 15430
rect 23988 15396 24078 15430
rect 24078 15396 24146 15430
rect 24146 15396 24236 15430
rect 24236 15396 24304 15430
rect 24304 15396 24394 15430
rect 24394 15396 24462 15430
rect 24462 15396 24552 15430
rect 24552 15396 24620 15430
rect 24620 15396 24710 15430
rect 24710 15396 24778 15430
rect 24778 15396 24868 15430
rect 24868 15396 24936 15430
rect 24936 15396 25026 15430
rect 25026 15396 25086 15430
rect 20452 15390 25086 15396
rect 20230 9336 20246 15380
rect 20246 9336 20284 15380
rect 20284 9336 20300 15380
rect 25240 15380 25310 15520
rect 25650 15410 25850 15480
rect 26150 15410 26350 15480
rect 20365 9378 20382 15338
rect 20382 9378 20416 15338
rect 20416 9378 20431 15338
rect 20523 9378 20540 15338
rect 20540 9378 20574 15338
rect 20574 9378 20589 15338
rect 20681 9378 20698 15338
rect 20698 9378 20732 15338
rect 20732 9378 20747 15338
rect 20839 9378 20856 15338
rect 20856 9378 20890 15338
rect 20890 9378 20905 15338
rect 20997 9378 21014 15338
rect 21014 9378 21048 15338
rect 21048 9378 21063 15338
rect 21155 9378 21172 15338
rect 21172 9378 21206 15338
rect 21206 9378 21221 15338
rect 21313 9378 21330 15338
rect 21330 9378 21364 15338
rect 21364 9378 21379 15338
rect 21471 9378 21488 15338
rect 21488 9378 21522 15338
rect 21522 9378 21537 15338
rect 21629 9378 21646 15338
rect 21646 9378 21680 15338
rect 21680 9378 21695 15338
rect 21787 9378 21804 15338
rect 21804 9378 21838 15338
rect 21838 9378 21853 15338
rect 21945 9378 21962 15338
rect 21962 9378 21996 15338
rect 21996 9378 22011 15338
rect 22103 9378 22120 15338
rect 22120 9378 22154 15338
rect 22154 9378 22169 15338
rect 22261 9378 22278 15338
rect 22278 9378 22312 15338
rect 22312 9378 22327 15338
rect 22419 9378 22436 15338
rect 22436 9378 22470 15338
rect 22470 9378 22485 15338
rect 22577 9378 22594 15338
rect 22594 9378 22628 15338
rect 22628 9378 22643 15338
rect 22735 9378 22752 15338
rect 22752 9378 22786 15338
rect 22786 9378 22801 15338
rect 22893 9378 22910 15338
rect 22910 9378 22944 15338
rect 22944 9378 22959 15338
rect 23051 9378 23068 15338
rect 23068 9378 23102 15338
rect 23102 9378 23117 15338
rect 23209 9378 23226 15338
rect 23226 9378 23260 15338
rect 23260 9378 23275 15338
rect 23367 9378 23384 15338
rect 23384 9378 23418 15338
rect 23418 9378 23433 15338
rect 23525 9378 23542 15338
rect 23542 9378 23576 15338
rect 23576 9378 23591 15338
rect 23683 9378 23700 15338
rect 23700 9378 23734 15338
rect 23734 9378 23749 15338
rect 23841 9378 23858 15338
rect 23858 9378 23892 15338
rect 23892 9378 23907 15338
rect 23999 9378 24016 15338
rect 24016 9378 24050 15338
rect 24050 9378 24065 15338
rect 24157 9378 24174 15338
rect 24174 9378 24208 15338
rect 24208 9378 24223 15338
rect 24315 9378 24332 15338
rect 24332 9378 24366 15338
rect 24366 9378 24381 15338
rect 24473 9378 24490 15338
rect 24490 9378 24524 15338
rect 24524 9378 24539 15338
rect 24631 9378 24648 15338
rect 24648 9378 24682 15338
rect 24682 9378 24697 15338
rect 24789 9378 24806 15338
rect 24806 9378 24840 15338
rect 24840 9378 24855 15338
rect 24947 9378 24964 15338
rect 24964 9378 24998 15338
rect 24998 9378 25013 15338
rect 25105 9378 25122 15338
rect 25122 9378 25156 15338
rect 25156 9378 25171 15338
rect 20230 9200 20300 9336
rect 25240 9336 25254 15380
rect 25254 9336 25292 15380
rect 25292 9336 25310 15380
rect 25520 15150 25590 15350
rect 25910 15150 25980 15350
rect 26020 15150 26090 15350
rect 26410 15150 26480 15350
rect 25650 15020 25850 15090
rect 26150 15020 26350 15090
rect 25650 14910 25850 14980
rect 26150 14910 26350 14980
rect 25520 14650 25590 14850
rect 25910 14650 25980 14850
rect 26020 14650 26090 14850
rect 26410 14650 26480 14850
rect 25650 14520 25850 14590
rect 26150 14520 26350 14590
rect 25650 14410 25850 14480
rect 26150 14410 26350 14480
rect 25520 14150 25590 14350
rect 25910 14150 25980 14350
rect 26020 14150 26090 14350
rect 26410 14150 26480 14350
rect 25650 14020 25850 14090
rect 26150 14020 26350 14090
rect 25650 13910 25850 13980
rect 26150 13910 26350 13980
rect 26650 13910 26850 13980
rect 27150 13910 27350 13980
rect 27650 13910 27850 13980
rect 28150 13910 28350 13980
rect 28650 13910 28850 13980
rect 29150 13910 29350 13980
rect 29650 13910 29850 13980
rect 30150 13910 30350 13980
rect 25520 13650 25590 13850
rect 25910 13650 25980 13850
rect 26020 13650 26090 13850
rect 26410 13650 26480 13850
rect 26520 13650 26590 13850
rect 26910 13650 26980 13850
rect 27020 13650 27090 13850
rect 27410 13650 27480 13850
rect 27520 13650 27590 13850
rect 27910 13650 27980 13850
rect 28020 13650 28090 13850
rect 28410 13650 28480 13850
rect 28520 13650 28590 13850
rect 28910 13650 28980 13850
rect 29020 13650 29090 13850
rect 29410 13650 29480 13850
rect 29520 13650 29590 13850
rect 29910 13650 29980 13850
rect 30020 13650 30090 13850
rect 30410 13650 30480 13850
rect 25650 13520 25850 13590
rect 26150 13520 26350 13590
rect 26650 13520 26850 13590
rect 27150 13520 27350 13590
rect 27650 13520 27850 13590
rect 28150 13520 28350 13590
rect 28650 13520 28850 13590
rect 29150 13520 29350 13590
rect 29650 13520 29850 13590
rect 30150 13520 30350 13590
rect 25650 13410 25850 13480
rect 26150 13410 26350 13480
rect 26650 13410 26850 13480
rect 27150 13410 27350 13480
rect 27650 13410 27850 13480
rect 28150 13410 28350 13480
rect 28650 13410 28850 13480
rect 29150 13410 29350 13480
rect 29650 13410 29850 13480
rect 30150 13410 30350 13480
rect 25520 13150 25590 13350
rect 25910 13150 25980 13350
rect 26020 13150 26090 13350
rect 26410 13150 26480 13350
rect 26520 13150 26590 13350
rect 26910 13150 26980 13350
rect 27020 13150 27090 13350
rect 27410 13150 27480 13350
rect 27520 13150 27590 13350
rect 27910 13150 27980 13350
rect 28020 13150 28090 13350
rect 28410 13150 28480 13350
rect 28520 13150 28590 13350
rect 28910 13150 28980 13350
rect 29020 13150 29090 13350
rect 29410 13150 29480 13350
rect 29520 13150 29590 13350
rect 29910 13150 29980 13350
rect 30020 13150 30090 13350
rect 30410 13150 30480 13350
rect 25650 13020 25850 13090
rect 26150 13020 26350 13090
rect 26650 13020 26850 13090
rect 27150 13020 27350 13090
rect 27650 13020 27850 13090
rect 28150 13020 28350 13090
rect 28650 13020 28850 13090
rect 29150 13020 29350 13090
rect 29650 13020 29850 13090
rect 30150 13020 30350 13090
rect 25650 12910 25850 12980
rect 26150 12910 26350 12980
rect 25520 12650 25590 12850
rect 25910 12650 25980 12850
rect 26020 12650 26090 12850
rect 26410 12650 26480 12850
rect 25650 12520 25850 12590
rect 26150 12520 26350 12590
rect 30910 13832 31090 13900
rect 30910 13435 30980 13832
rect 30980 13435 31018 13832
rect 31018 13435 31090 13832
rect 30910 13420 31090 13435
rect 30910 13081 31090 13090
rect 30910 12684 30980 13081
rect 30980 12684 31018 13081
rect 31018 12684 31090 13081
rect 30910 12610 31090 12684
rect 25650 12410 25850 12480
rect 26150 12410 26350 12480
rect 25520 12150 25590 12350
rect 25910 12150 25980 12350
rect 26020 12150 26090 12350
rect 26410 12150 26480 12350
rect 25650 12020 25850 12090
rect 26150 12020 26350 12090
rect 25650 11910 25850 11980
rect 26150 11910 26350 11980
rect 25520 11650 25590 11850
rect 25910 11650 25980 11850
rect 26020 11650 26090 11850
rect 26410 11650 26480 11850
rect 25650 11520 25850 11590
rect 26150 11520 26350 11590
rect 25650 11410 25850 11480
rect 26150 11410 26350 11480
rect 25520 11150 25590 11350
rect 25910 11150 25980 11350
rect 26020 11150 26090 11350
rect 26410 11150 26480 11350
rect 25650 11020 25850 11090
rect 26150 11020 26350 11090
rect 25650 10910 25850 10980
rect 26150 10910 26350 10980
rect 25520 10650 25590 10850
rect 25910 10650 25980 10850
rect 26020 10650 26090 10850
rect 26410 10650 26480 10850
rect 25650 10520 25850 10590
rect 26150 10520 26350 10590
rect 25650 10410 25850 10480
rect 26150 10410 26350 10480
rect 25520 10150 25590 10350
rect 25910 10150 25980 10350
rect 26020 10150 26090 10350
rect 26410 10150 26480 10350
rect 25650 10020 25850 10090
rect 26150 10020 26350 10090
rect 25650 9910 25850 9980
rect 26150 9910 26350 9980
rect 25520 9650 25590 9850
rect 25910 9650 25980 9850
rect 26020 9650 26090 9850
rect 26410 9650 26480 9850
rect 25650 9520 25850 9590
rect 26150 9520 26350 9590
rect 25650 9410 25850 9480
rect 26150 9410 26350 9480
rect 20452 9320 25086 9326
rect 20452 9286 20512 9320
rect 20512 9286 20602 9320
rect 20602 9286 20670 9320
rect 20670 9286 20760 9320
rect 20760 9286 20828 9320
rect 20828 9286 20918 9320
rect 20918 9286 20986 9320
rect 20986 9286 21076 9320
rect 21076 9286 21144 9320
rect 21144 9286 21234 9320
rect 21234 9286 21302 9320
rect 21302 9286 21392 9320
rect 21392 9286 21460 9320
rect 21460 9286 21550 9320
rect 21550 9286 21618 9320
rect 21618 9286 21708 9320
rect 21708 9286 21776 9320
rect 21776 9286 21866 9320
rect 21866 9286 21934 9320
rect 21934 9286 22024 9320
rect 22024 9286 22092 9320
rect 22092 9286 22182 9320
rect 22182 9286 22250 9320
rect 22250 9286 22340 9320
rect 22340 9286 22408 9320
rect 22408 9286 22498 9320
rect 22498 9286 22566 9320
rect 22566 9286 22656 9320
rect 22656 9286 22724 9320
rect 22724 9286 22814 9320
rect 22814 9286 22882 9320
rect 22882 9286 22972 9320
rect 22972 9286 23040 9320
rect 23040 9286 23130 9320
rect 23130 9286 23198 9320
rect 23198 9286 23288 9320
rect 23288 9286 23356 9320
rect 23356 9286 23446 9320
rect 23446 9286 23514 9320
rect 23514 9286 23604 9320
rect 23604 9286 23672 9320
rect 23672 9286 23762 9320
rect 23762 9286 23830 9320
rect 23830 9286 23920 9320
rect 23920 9286 23988 9320
rect 23988 9286 24078 9320
rect 24078 9286 24146 9320
rect 24146 9286 24236 9320
rect 24236 9286 24304 9320
rect 24304 9286 24394 9320
rect 24394 9286 24462 9320
rect 24462 9286 24552 9320
rect 24552 9286 24620 9320
rect 24620 9286 24710 9320
rect 24710 9286 24778 9320
rect 24778 9286 24868 9320
rect 24868 9286 24936 9320
rect 24936 9286 25026 9320
rect 25026 9286 25086 9320
rect 20452 9226 25086 9286
rect 25240 9200 25310 9336
rect 25520 9150 25590 9350
rect 150 9020 350 9090
rect 650 9020 850 9090
rect 150 8910 350 8980
rect 650 8910 850 8980
rect 20 8650 90 8850
rect 410 8650 480 8850
rect 520 8650 590 8850
rect 910 8650 980 8850
rect 150 8520 350 8590
rect 650 8520 850 8590
rect 25910 9150 25980 9350
rect 26020 9150 26090 9350
rect 26410 9150 26480 9350
rect 25650 9020 25850 9090
rect 26150 9020 26350 9090
rect 25650 8910 25850 8980
rect 26150 8910 26350 8980
rect 25520 8650 25590 8850
rect 25910 8650 25980 8850
rect 26020 8650 26090 8850
rect 26410 8650 26480 8850
rect 150 8410 350 8480
rect 650 8410 850 8480
rect 1330 8380 1400 8520
rect 1552 8430 6186 8490
rect 1552 8396 1612 8430
rect 1612 8396 1702 8430
rect 1702 8396 1770 8430
rect 1770 8396 1860 8430
rect 1860 8396 1928 8430
rect 1928 8396 2018 8430
rect 2018 8396 2086 8430
rect 2086 8396 2176 8430
rect 2176 8396 2244 8430
rect 2244 8396 2334 8430
rect 2334 8396 2402 8430
rect 2402 8396 2492 8430
rect 2492 8396 2560 8430
rect 2560 8396 2650 8430
rect 2650 8396 2718 8430
rect 2718 8396 2808 8430
rect 2808 8396 2876 8430
rect 2876 8396 2966 8430
rect 2966 8396 3034 8430
rect 3034 8396 3124 8430
rect 3124 8396 3192 8430
rect 3192 8396 3282 8430
rect 3282 8396 3350 8430
rect 3350 8396 3440 8430
rect 3440 8396 3508 8430
rect 3508 8396 3598 8430
rect 3598 8396 3666 8430
rect 3666 8396 3756 8430
rect 3756 8396 3824 8430
rect 3824 8396 3914 8430
rect 3914 8396 3982 8430
rect 3982 8396 4072 8430
rect 4072 8396 4140 8430
rect 4140 8396 4230 8430
rect 4230 8396 4298 8430
rect 4298 8396 4388 8430
rect 4388 8396 4456 8430
rect 4456 8396 4546 8430
rect 4546 8396 4614 8430
rect 4614 8396 4704 8430
rect 4704 8396 4772 8430
rect 4772 8396 4862 8430
rect 4862 8396 4930 8430
rect 4930 8396 5020 8430
rect 5020 8396 5088 8430
rect 5088 8396 5178 8430
rect 5178 8396 5246 8430
rect 5246 8396 5336 8430
rect 5336 8396 5404 8430
rect 5404 8396 5494 8430
rect 5494 8396 5562 8430
rect 5562 8396 5652 8430
rect 5652 8396 5720 8430
rect 5720 8396 5810 8430
rect 5810 8396 5878 8430
rect 5878 8396 5968 8430
rect 5968 8396 6036 8430
rect 6036 8396 6126 8430
rect 6126 8396 6186 8430
rect 1552 8390 6186 8396
rect 20 8150 90 8350
rect 410 8150 480 8350
rect 520 8150 590 8350
rect 910 8150 980 8350
rect 150 8020 350 8090
rect 650 8020 850 8090
rect 150 7910 350 7980
rect 650 7910 850 7980
rect 20 7650 90 7850
rect 410 7650 480 7850
rect 520 7650 590 7850
rect 910 7650 980 7850
rect 150 7520 350 7590
rect 650 7520 850 7590
rect 150 7410 350 7480
rect 650 7410 850 7480
rect 20 7150 90 7350
rect 410 7150 480 7350
rect 520 7150 590 7350
rect 910 7150 980 7350
rect 150 7020 350 7090
rect 650 7020 850 7090
rect 150 6910 350 6980
rect 650 6910 850 6980
rect 20 6650 90 6850
rect 410 6650 480 6850
rect 520 6650 590 6850
rect 910 6650 980 6850
rect 150 6520 350 6590
rect 650 6520 850 6590
rect 150 6410 350 6480
rect 650 6410 850 6480
rect 20 6150 90 6350
rect 410 6150 480 6350
rect 520 6150 590 6350
rect 910 6150 980 6350
rect 150 6020 350 6090
rect 650 6020 850 6090
rect 150 5910 350 5980
rect 650 5910 850 5980
rect 20 5650 90 5850
rect 410 5650 480 5850
rect 520 5650 590 5850
rect 910 5650 980 5850
rect 150 5520 350 5590
rect 650 5520 850 5590
rect 150 5410 350 5480
rect 650 5410 850 5480
rect 20 5150 90 5350
rect 410 5150 480 5350
rect 520 5150 590 5350
rect 910 5150 980 5350
rect 150 5020 350 5090
rect 650 5020 850 5090
rect 150 4910 350 4980
rect 650 4910 850 4980
rect 20 4650 90 4850
rect 410 4650 480 4850
rect 520 4650 590 4850
rect 910 4650 980 4850
rect 150 4520 350 4590
rect 650 4520 850 4590
rect 150 4410 350 4480
rect 650 4410 850 4480
rect 20 4150 90 4350
rect 410 4150 480 4350
rect 520 4150 590 4350
rect 910 4150 980 4350
rect 150 4020 350 4090
rect 650 4020 850 4090
rect 150 3910 350 3980
rect 650 3910 850 3980
rect 20 3650 90 3850
rect 410 3650 480 3850
rect 520 3650 590 3850
rect 910 3650 980 3850
rect 150 3520 350 3590
rect 650 3520 850 3590
rect 150 3410 350 3480
rect 650 3410 850 3480
rect 20 3150 90 3350
rect 410 3150 480 3350
rect 520 3150 590 3350
rect 910 3150 980 3350
rect 150 3020 350 3090
rect 650 3020 850 3090
rect 150 2910 350 2980
rect 650 2910 850 2980
rect 20 2650 90 2850
rect 410 2650 480 2850
rect 520 2650 590 2850
rect 910 2650 980 2850
rect 150 2520 350 2590
rect 650 2520 850 2590
rect 150 2410 350 2480
rect 650 2410 850 2480
rect 20 2150 90 2350
rect 410 2150 480 2350
rect 520 2150 590 2350
rect 910 2150 980 2350
rect 1330 2336 1346 8380
rect 1346 2336 1384 8380
rect 1384 2336 1400 8380
rect 6340 8380 6410 8520
rect 1465 2378 1482 8338
rect 1482 2378 1516 8338
rect 1516 2378 1531 8338
rect 1623 2378 1640 8338
rect 1640 2378 1674 8338
rect 1674 2378 1689 8338
rect 1781 2378 1798 8338
rect 1798 2378 1832 8338
rect 1832 2378 1847 8338
rect 1939 2378 1956 8338
rect 1956 2378 1990 8338
rect 1990 2378 2005 8338
rect 2097 2378 2114 8338
rect 2114 2378 2148 8338
rect 2148 2378 2163 8338
rect 2255 2378 2272 8338
rect 2272 2378 2306 8338
rect 2306 2378 2321 8338
rect 2413 2378 2430 8338
rect 2430 2378 2464 8338
rect 2464 2378 2479 8338
rect 2571 2378 2588 8338
rect 2588 2378 2622 8338
rect 2622 2378 2637 8338
rect 2729 2378 2746 8338
rect 2746 2378 2780 8338
rect 2780 2378 2795 8338
rect 2887 2378 2904 8338
rect 2904 2378 2938 8338
rect 2938 2378 2953 8338
rect 3045 2378 3062 8338
rect 3062 2378 3096 8338
rect 3096 2378 3111 8338
rect 3203 2378 3220 8338
rect 3220 2378 3254 8338
rect 3254 2378 3269 8338
rect 3361 2378 3378 8338
rect 3378 2378 3412 8338
rect 3412 2378 3427 8338
rect 3519 2378 3536 8338
rect 3536 2378 3570 8338
rect 3570 2378 3585 8338
rect 3677 2378 3694 8338
rect 3694 2378 3728 8338
rect 3728 2378 3743 8338
rect 3835 2378 3852 8338
rect 3852 2378 3886 8338
rect 3886 2378 3901 8338
rect 3993 2378 4010 8338
rect 4010 2378 4044 8338
rect 4044 2378 4059 8338
rect 4151 2378 4168 8338
rect 4168 2378 4202 8338
rect 4202 2378 4217 8338
rect 4309 2378 4326 8338
rect 4326 2378 4360 8338
rect 4360 2378 4375 8338
rect 4467 2378 4484 8338
rect 4484 2378 4518 8338
rect 4518 2378 4533 8338
rect 4625 2378 4642 8338
rect 4642 2378 4676 8338
rect 4676 2378 4691 8338
rect 4783 2378 4800 8338
rect 4800 2378 4834 8338
rect 4834 2378 4849 8338
rect 4941 2378 4958 8338
rect 4958 2378 4992 8338
rect 4992 2378 5007 8338
rect 5099 2378 5116 8338
rect 5116 2378 5150 8338
rect 5150 2378 5165 8338
rect 5257 2378 5274 8338
rect 5274 2378 5308 8338
rect 5308 2378 5323 8338
rect 5415 2378 5432 8338
rect 5432 2378 5466 8338
rect 5466 2378 5481 8338
rect 5573 2378 5590 8338
rect 5590 2378 5624 8338
rect 5624 2378 5639 8338
rect 5731 2378 5748 8338
rect 5748 2378 5782 8338
rect 5782 2378 5797 8338
rect 5889 2378 5906 8338
rect 5906 2378 5940 8338
rect 5940 2378 5955 8338
rect 6047 2378 6064 8338
rect 6064 2378 6098 8338
rect 6098 2378 6113 8338
rect 6205 2378 6222 8338
rect 6222 2378 6256 8338
rect 6256 2378 6271 8338
rect 1330 2200 1400 2336
rect 6340 2336 6354 8380
rect 6354 2336 6392 8380
rect 6392 2336 6410 8380
rect 7630 8380 7700 8520
rect 7852 8430 12486 8490
rect 7852 8396 7912 8430
rect 7912 8396 8002 8430
rect 8002 8396 8070 8430
rect 8070 8396 8160 8430
rect 8160 8396 8228 8430
rect 8228 8396 8318 8430
rect 8318 8396 8386 8430
rect 8386 8396 8476 8430
rect 8476 8396 8544 8430
rect 8544 8396 8634 8430
rect 8634 8396 8702 8430
rect 8702 8396 8792 8430
rect 8792 8396 8860 8430
rect 8860 8396 8950 8430
rect 8950 8396 9018 8430
rect 9018 8396 9108 8430
rect 9108 8396 9176 8430
rect 9176 8396 9266 8430
rect 9266 8396 9334 8430
rect 9334 8396 9424 8430
rect 9424 8396 9492 8430
rect 9492 8396 9582 8430
rect 9582 8396 9650 8430
rect 9650 8396 9740 8430
rect 9740 8396 9808 8430
rect 9808 8396 9898 8430
rect 9898 8396 9966 8430
rect 9966 8396 10056 8430
rect 10056 8396 10124 8430
rect 10124 8396 10214 8430
rect 10214 8396 10282 8430
rect 10282 8396 10372 8430
rect 10372 8396 10440 8430
rect 10440 8396 10530 8430
rect 10530 8396 10598 8430
rect 10598 8396 10688 8430
rect 10688 8396 10756 8430
rect 10756 8396 10846 8430
rect 10846 8396 10914 8430
rect 10914 8396 11004 8430
rect 11004 8396 11072 8430
rect 11072 8396 11162 8430
rect 11162 8396 11230 8430
rect 11230 8396 11320 8430
rect 11320 8396 11388 8430
rect 11388 8396 11478 8430
rect 11478 8396 11546 8430
rect 11546 8396 11636 8430
rect 11636 8396 11704 8430
rect 11704 8396 11794 8430
rect 11794 8396 11862 8430
rect 11862 8396 11952 8430
rect 11952 8396 12020 8430
rect 12020 8396 12110 8430
rect 12110 8396 12178 8430
rect 12178 8396 12268 8430
rect 12268 8396 12336 8430
rect 12336 8396 12426 8430
rect 12426 8396 12486 8430
rect 7852 8390 12486 8396
rect 6650 2410 6850 2480
rect 7150 2410 7350 2480
rect 1552 2320 6186 2326
rect 1552 2286 1612 2320
rect 1612 2286 1702 2320
rect 1702 2286 1770 2320
rect 1770 2286 1860 2320
rect 1860 2286 1928 2320
rect 1928 2286 2018 2320
rect 2018 2286 2086 2320
rect 2086 2286 2176 2320
rect 2176 2286 2244 2320
rect 2244 2286 2334 2320
rect 2334 2286 2402 2320
rect 2402 2286 2492 2320
rect 2492 2286 2560 2320
rect 2560 2286 2650 2320
rect 2650 2286 2718 2320
rect 2718 2286 2808 2320
rect 2808 2286 2876 2320
rect 2876 2286 2966 2320
rect 2966 2286 3034 2320
rect 3034 2286 3124 2320
rect 3124 2286 3192 2320
rect 3192 2286 3282 2320
rect 3282 2286 3350 2320
rect 3350 2286 3440 2320
rect 3440 2286 3508 2320
rect 3508 2286 3598 2320
rect 3598 2286 3666 2320
rect 3666 2286 3756 2320
rect 3756 2286 3824 2320
rect 3824 2286 3914 2320
rect 3914 2286 3982 2320
rect 3982 2286 4072 2320
rect 4072 2286 4140 2320
rect 4140 2286 4230 2320
rect 4230 2286 4298 2320
rect 4298 2286 4388 2320
rect 4388 2286 4456 2320
rect 4456 2286 4546 2320
rect 4546 2286 4614 2320
rect 4614 2286 4704 2320
rect 4704 2286 4772 2320
rect 4772 2286 4862 2320
rect 4862 2286 4930 2320
rect 4930 2286 5020 2320
rect 5020 2286 5088 2320
rect 5088 2286 5178 2320
rect 5178 2286 5246 2320
rect 5246 2286 5336 2320
rect 5336 2286 5404 2320
rect 5404 2286 5494 2320
rect 5494 2286 5562 2320
rect 5562 2286 5652 2320
rect 5652 2286 5720 2320
rect 5720 2286 5810 2320
rect 5810 2286 5878 2320
rect 5878 2286 5968 2320
rect 5968 2286 6036 2320
rect 6036 2286 6126 2320
rect 6126 2286 6186 2320
rect 1552 2226 6186 2286
rect 6340 2200 6410 2336
rect 6520 2150 6590 2350
rect 6910 2150 6980 2350
rect 7020 2150 7090 2350
rect 7410 2150 7480 2350
rect 7630 2336 7646 8380
rect 7646 2336 7684 8380
rect 7684 2336 7700 8380
rect 12640 8380 12710 8520
rect 7765 2378 7782 8338
rect 7782 2378 7816 8338
rect 7816 2378 7831 8338
rect 7923 2378 7940 8338
rect 7940 2378 7974 8338
rect 7974 2378 7989 8338
rect 8081 2378 8098 8338
rect 8098 2378 8132 8338
rect 8132 2378 8147 8338
rect 8239 2378 8256 8338
rect 8256 2378 8290 8338
rect 8290 2378 8305 8338
rect 8397 2378 8414 8338
rect 8414 2378 8448 8338
rect 8448 2378 8463 8338
rect 8555 2378 8572 8338
rect 8572 2378 8606 8338
rect 8606 2378 8621 8338
rect 8713 2378 8730 8338
rect 8730 2378 8764 8338
rect 8764 2378 8779 8338
rect 8871 2378 8888 8338
rect 8888 2378 8922 8338
rect 8922 2378 8937 8338
rect 9029 2378 9046 8338
rect 9046 2378 9080 8338
rect 9080 2378 9095 8338
rect 9187 2378 9204 8338
rect 9204 2378 9238 8338
rect 9238 2378 9253 8338
rect 9345 2378 9362 8338
rect 9362 2378 9396 8338
rect 9396 2378 9411 8338
rect 9503 2378 9520 8338
rect 9520 2378 9554 8338
rect 9554 2378 9569 8338
rect 9661 2378 9678 8338
rect 9678 2378 9712 8338
rect 9712 2378 9727 8338
rect 9819 2378 9836 8338
rect 9836 2378 9870 8338
rect 9870 2378 9885 8338
rect 9977 2378 9994 8338
rect 9994 2378 10028 8338
rect 10028 2378 10043 8338
rect 10135 2378 10152 8338
rect 10152 2378 10186 8338
rect 10186 2378 10201 8338
rect 10293 2378 10310 8338
rect 10310 2378 10344 8338
rect 10344 2378 10359 8338
rect 10451 2378 10468 8338
rect 10468 2378 10502 8338
rect 10502 2378 10517 8338
rect 10609 2378 10626 8338
rect 10626 2378 10660 8338
rect 10660 2378 10675 8338
rect 10767 2378 10784 8338
rect 10784 2378 10818 8338
rect 10818 2378 10833 8338
rect 10925 2378 10942 8338
rect 10942 2378 10976 8338
rect 10976 2378 10991 8338
rect 11083 2378 11100 8338
rect 11100 2378 11134 8338
rect 11134 2378 11149 8338
rect 11241 2378 11258 8338
rect 11258 2378 11292 8338
rect 11292 2378 11307 8338
rect 11399 2378 11416 8338
rect 11416 2378 11450 8338
rect 11450 2378 11465 8338
rect 11557 2378 11574 8338
rect 11574 2378 11608 8338
rect 11608 2378 11623 8338
rect 11715 2378 11732 8338
rect 11732 2378 11766 8338
rect 11766 2378 11781 8338
rect 11873 2378 11890 8338
rect 11890 2378 11924 8338
rect 11924 2378 11939 8338
rect 12031 2378 12048 8338
rect 12048 2378 12082 8338
rect 12082 2378 12097 8338
rect 12189 2378 12206 8338
rect 12206 2378 12240 8338
rect 12240 2378 12255 8338
rect 12347 2378 12364 8338
rect 12364 2378 12398 8338
rect 12398 2378 12413 8338
rect 12505 2378 12522 8338
rect 12522 2378 12556 8338
rect 12556 2378 12571 8338
rect 7630 2200 7700 2336
rect 12640 2336 12654 8380
rect 12654 2336 12692 8380
rect 12692 2336 12710 8380
rect 13930 8380 14000 8520
rect 14152 8430 18786 8490
rect 14152 8396 14212 8430
rect 14212 8396 14302 8430
rect 14302 8396 14370 8430
rect 14370 8396 14460 8430
rect 14460 8396 14528 8430
rect 14528 8396 14618 8430
rect 14618 8396 14686 8430
rect 14686 8396 14776 8430
rect 14776 8396 14844 8430
rect 14844 8396 14934 8430
rect 14934 8396 15002 8430
rect 15002 8396 15092 8430
rect 15092 8396 15160 8430
rect 15160 8396 15250 8430
rect 15250 8396 15318 8430
rect 15318 8396 15408 8430
rect 15408 8396 15476 8430
rect 15476 8396 15566 8430
rect 15566 8396 15634 8430
rect 15634 8396 15724 8430
rect 15724 8396 15792 8430
rect 15792 8396 15882 8430
rect 15882 8396 15950 8430
rect 15950 8396 16040 8430
rect 16040 8396 16108 8430
rect 16108 8396 16198 8430
rect 16198 8396 16266 8430
rect 16266 8396 16356 8430
rect 16356 8396 16424 8430
rect 16424 8396 16514 8430
rect 16514 8396 16582 8430
rect 16582 8396 16672 8430
rect 16672 8396 16740 8430
rect 16740 8396 16830 8430
rect 16830 8396 16898 8430
rect 16898 8396 16988 8430
rect 16988 8396 17056 8430
rect 17056 8396 17146 8430
rect 17146 8396 17214 8430
rect 17214 8396 17304 8430
rect 17304 8396 17372 8430
rect 17372 8396 17462 8430
rect 17462 8396 17530 8430
rect 17530 8396 17620 8430
rect 17620 8396 17688 8430
rect 17688 8396 17778 8430
rect 17778 8396 17846 8430
rect 17846 8396 17936 8430
rect 17936 8396 18004 8430
rect 18004 8396 18094 8430
rect 18094 8396 18162 8430
rect 18162 8396 18252 8430
rect 18252 8396 18320 8430
rect 18320 8396 18410 8430
rect 18410 8396 18478 8430
rect 18478 8396 18568 8430
rect 18568 8396 18636 8430
rect 18636 8396 18726 8430
rect 18726 8396 18786 8430
rect 14152 8390 18786 8396
rect 13150 2410 13350 2480
rect 7852 2320 12486 2326
rect 7852 2286 7912 2320
rect 7912 2286 8002 2320
rect 8002 2286 8070 2320
rect 8070 2286 8160 2320
rect 8160 2286 8228 2320
rect 8228 2286 8318 2320
rect 8318 2286 8386 2320
rect 8386 2286 8476 2320
rect 8476 2286 8544 2320
rect 8544 2286 8634 2320
rect 8634 2286 8702 2320
rect 8702 2286 8792 2320
rect 8792 2286 8860 2320
rect 8860 2286 8950 2320
rect 8950 2286 9018 2320
rect 9018 2286 9108 2320
rect 9108 2286 9176 2320
rect 9176 2286 9266 2320
rect 9266 2286 9334 2320
rect 9334 2286 9424 2320
rect 9424 2286 9492 2320
rect 9492 2286 9582 2320
rect 9582 2286 9650 2320
rect 9650 2286 9740 2320
rect 9740 2286 9808 2320
rect 9808 2286 9898 2320
rect 9898 2286 9966 2320
rect 9966 2286 10056 2320
rect 10056 2286 10124 2320
rect 10124 2286 10214 2320
rect 10214 2286 10282 2320
rect 10282 2286 10372 2320
rect 10372 2286 10440 2320
rect 10440 2286 10530 2320
rect 10530 2286 10598 2320
rect 10598 2286 10688 2320
rect 10688 2286 10756 2320
rect 10756 2286 10846 2320
rect 10846 2286 10914 2320
rect 10914 2286 11004 2320
rect 11004 2286 11072 2320
rect 11072 2286 11162 2320
rect 11162 2286 11230 2320
rect 11230 2286 11320 2320
rect 11320 2286 11388 2320
rect 11388 2286 11478 2320
rect 11478 2286 11546 2320
rect 11546 2286 11636 2320
rect 11636 2286 11704 2320
rect 11704 2286 11794 2320
rect 11794 2286 11862 2320
rect 11862 2286 11952 2320
rect 11952 2286 12020 2320
rect 12020 2286 12110 2320
rect 12110 2286 12178 2320
rect 12178 2286 12268 2320
rect 12268 2286 12336 2320
rect 12336 2286 12426 2320
rect 12426 2286 12486 2320
rect 7852 2226 12486 2286
rect 12640 2200 12710 2336
rect 13020 2150 13090 2350
rect 13410 2150 13480 2350
rect 13930 2336 13946 8380
rect 13946 2336 13984 8380
rect 13984 2336 14000 8380
rect 18940 8380 19010 8520
rect 14065 2378 14082 8338
rect 14082 2378 14116 8338
rect 14116 2378 14131 8338
rect 14223 2378 14240 8338
rect 14240 2378 14274 8338
rect 14274 2378 14289 8338
rect 14381 2378 14398 8338
rect 14398 2378 14432 8338
rect 14432 2378 14447 8338
rect 14539 2378 14556 8338
rect 14556 2378 14590 8338
rect 14590 2378 14605 8338
rect 14697 2378 14714 8338
rect 14714 2378 14748 8338
rect 14748 2378 14763 8338
rect 14855 2378 14872 8338
rect 14872 2378 14906 8338
rect 14906 2378 14921 8338
rect 15013 2378 15030 8338
rect 15030 2378 15064 8338
rect 15064 2378 15079 8338
rect 15171 2378 15188 8338
rect 15188 2378 15222 8338
rect 15222 2378 15237 8338
rect 15329 2378 15346 8338
rect 15346 2378 15380 8338
rect 15380 2378 15395 8338
rect 15487 2378 15504 8338
rect 15504 2378 15538 8338
rect 15538 2378 15553 8338
rect 15645 2378 15662 8338
rect 15662 2378 15696 8338
rect 15696 2378 15711 8338
rect 15803 2378 15820 8338
rect 15820 2378 15854 8338
rect 15854 2378 15869 8338
rect 15961 2378 15978 8338
rect 15978 2378 16012 8338
rect 16012 2378 16027 8338
rect 16119 2378 16136 8338
rect 16136 2378 16170 8338
rect 16170 2378 16185 8338
rect 16277 2378 16294 8338
rect 16294 2378 16328 8338
rect 16328 2378 16343 8338
rect 16435 2378 16452 8338
rect 16452 2378 16486 8338
rect 16486 2378 16501 8338
rect 16593 2378 16610 8338
rect 16610 2378 16644 8338
rect 16644 2378 16659 8338
rect 16751 2378 16768 8338
rect 16768 2378 16802 8338
rect 16802 2378 16817 8338
rect 16909 2378 16926 8338
rect 16926 2378 16960 8338
rect 16960 2378 16975 8338
rect 17067 2378 17084 8338
rect 17084 2378 17118 8338
rect 17118 2378 17133 8338
rect 17225 2378 17242 8338
rect 17242 2378 17276 8338
rect 17276 2378 17291 8338
rect 17383 2378 17400 8338
rect 17400 2378 17434 8338
rect 17434 2378 17449 8338
rect 17541 2378 17558 8338
rect 17558 2378 17592 8338
rect 17592 2378 17607 8338
rect 17699 2378 17716 8338
rect 17716 2378 17750 8338
rect 17750 2378 17765 8338
rect 17857 2378 17874 8338
rect 17874 2378 17908 8338
rect 17908 2378 17923 8338
rect 18015 2378 18032 8338
rect 18032 2378 18066 8338
rect 18066 2378 18081 8338
rect 18173 2378 18190 8338
rect 18190 2378 18224 8338
rect 18224 2378 18239 8338
rect 18331 2378 18348 8338
rect 18348 2378 18382 8338
rect 18382 2378 18397 8338
rect 18489 2378 18506 8338
rect 18506 2378 18540 8338
rect 18540 2378 18555 8338
rect 18647 2378 18664 8338
rect 18664 2378 18698 8338
rect 18698 2378 18713 8338
rect 18805 2378 18822 8338
rect 18822 2378 18856 8338
rect 18856 2378 18871 8338
rect 13930 2200 14000 2336
rect 18940 2336 18954 8380
rect 18954 2336 18992 8380
rect 18992 2336 19010 8380
rect 20230 8380 20300 8520
rect 25650 8520 25850 8590
rect 26150 8520 26350 8590
rect 20452 8430 25086 8490
rect 20452 8396 20512 8430
rect 20512 8396 20602 8430
rect 20602 8396 20670 8430
rect 20670 8396 20760 8430
rect 20760 8396 20828 8430
rect 20828 8396 20918 8430
rect 20918 8396 20986 8430
rect 20986 8396 21076 8430
rect 21076 8396 21144 8430
rect 21144 8396 21234 8430
rect 21234 8396 21302 8430
rect 21302 8396 21392 8430
rect 21392 8396 21460 8430
rect 21460 8396 21550 8430
rect 21550 8396 21618 8430
rect 21618 8396 21708 8430
rect 21708 8396 21776 8430
rect 21776 8396 21866 8430
rect 21866 8396 21934 8430
rect 21934 8396 22024 8430
rect 22024 8396 22092 8430
rect 22092 8396 22182 8430
rect 22182 8396 22250 8430
rect 22250 8396 22340 8430
rect 22340 8396 22408 8430
rect 22408 8396 22498 8430
rect 22498 8396 22566 8430
rect 22566 8396 22656 8430
rect 22656 8396 22724 8430
rect 22724 8396 22814 8430
rect 22814 8396 22882 8430
rect 22882 8396 22972 8430
rect 22972 8396 23040 8430
rect 23040 8396 23130 8430
rect 23130 8396 23198 8430
rect 23198 8396 23288 8430
rect 23288 8396 23356 8430
rect 23356 8396 23446 8430
rect 23446 8396 23514 8430
rect 23514 8396 23604 8430
rect 23604 8396 23672 8430
rect 23672 8396 23762 8430
rect 23762 8396 23830 8430
rect 23830 8396 23920 8430
rect 23920 8396 23988 8430
rect 23988 8396 24078 8430
rect 24078 8396 24146 8430
rect 24146 8396 24236 8430
rect 24236 8396 24304 8430
rect 24304 8396 24394 8430
rect 24394 8396 24462 8430
rect 24462 8396 24552 8430
rect 24552 8396 24620 8430
rect 24620 8396 24710 8430
rect 24710 8396 24778 8430
rect 24778 8396 24868 8430
rect 24868 8396 24936 8430
rect 24936 8396 25026 8430
rect 25026 8396 25086 8430
rect 20452 8390 25086 8396
rect 19650 2410 19850 2480
rect 14152 2320 18786 2326
rect 14152 2286 14212 2320
rect 14212 2286 14302 2320
rect 14302 2286 14370 2320
rect 14370 2286 14460 2320
rect 14460 2286 14528 2320
rect 14528 2286 14618 2320
rect 14618 2286 14686 2320
rect 14686 2286 14776 2320
rect 14776 2286 14844 2320
rect 14844 2286 14934 2320
rect 14934 2286 15002 2320
rect 15002 2286 15092 2320
rect 15092 2286 15160 2320
rect 15160 2286 15250 2320
rect 15250 2286 15318 2320
rect 15318 2286 15408 2320
rect 15408 2286 15476 2320
rect 15476 2286 15566 2320
rect 15566 2286 15634 2320
rect 15634 2286 15724 2320
rect 15724 2286 15792 2320
rect 15792 2286 15882 2320
rect 15882 2286 15950 2320
rect 15950 2286 16040 2320
rect 16040 2286 16108 2320
rect 16108 2286 16198 2320
rect 16198 2286 16266 2320
rect 16266 2286 16356 2320
rect 16356 2286 16424 2320
rect 16424 2286 16514 2320
rect 16514 2286 16582 2320
rect 16582 2286 16672 2320
rect 16672 2286 16740 2320
rect 16740 2286 16830 2320
rect 16830 2286 16898 2320
rect 16898 2286 16988 2320
rect 16988 2286 17056 2320
rect 17056 2286 17146 2320
rect 17146 2286 17214 2320
rect 17214 2286 17304 2320
rect 17304 2286 17372 2320
rect 17372 2286 17462 2320
rect 17462 2286 17530 2320
rect 17530 2286 17620 2320
rect 17620 2286 17688 2320
rect 17688 2286 17778 2320
rect 17778 2286 17846 2320
rect 17846 2286 17936 2320
rect 17936 2286 18004 2320
rect 18004 2286 18094 2320
rect 18094 2286 18162 2320
rect 18162 2286 18252 2320
rect 18252 2286 18320 2320
rect 18320 2286 18410 2320
rect 18410 2286 18478 2320
rect 18478 2286 18568 2320
rect 18568 2286 18636 2320
rect 18636 2286 18726 2320
rect 18726 2286 18786 2320
rect 14152 2226 18786 2286
rect 18940 2200 19010 2336
rect 19520 2150 19590 2350
rect 19910 2150 19980 2350
rect 20230 2336 20246 8380
rect 20246 2336 20284 8380
rect 20284 2336 20300 8380
rect 25240 8380 25310 8520
rect 25650 8410 25850 8480
rect 26150 8410 26350 8480
rect 20365 2378 20382 8338
rect 20382 2378 20416 8338
rect 20416 2378 20431 8338
rect 20523 2378 20540 8338
rect 20540 2378 20574 8338
rect 20574 2378 20589 8338
rect 20681 2378 20698 8338
rect 20698 2378 20732 8338
rect 20732 2378 20747 8338
rect 20839 2378 20856 8338
rect 20856 2378 20890 8338
rect 20890 2378 20905 8338
rect 20997 2378 21014 8338
rect 21014 2378 21048 8338
rect 21048 2378 21063 8338
rect 21155 2378 21172 8338
rect 21172 2378 21206 8338
rect 21206 2378 21221 8338
rect 21313 2378 21330 8338
rect 21330 2378 21364 8338
rect 21364 2378 21379 8338
rect 21471 2378 21488 8338
rect 21488 2378 21522 8338
rect 21522 2378 21537 8338
rect 21629 2378 21646 8338
rect 21646 2378 21680 8338
rect 21680 2378 21695 8338
rect 21787 2378 21804 8338
rect 21804 2378 21838 8338
rect 21838 2378 21853 8338
rect 21945 2378 21962 8338
rect 21962 2378 21996 8338
rect 21996 2378 22011 8338
rect 22103 2378 22120 8338
rect 22120 2378 22154 8338
rect 22154 2378 22169 8338
rect 22261 2378 22278 8338
rect 22278 2378 22312 8338
rect 22312 2378 22327 8338
rect 22419 2378 22436 8338
rect 22436 2378 22470 8338
rect 22470 2378 22485 8338
rect 22577 2378 22594 8338
rect 22594 2378 22628 8338
rect 22628 2378 22643 8338
rect 22735 2378 22752 8338
rect 22752 2378 22786 8338
rect 22786 2378 22801 8338
rect 22893 2378 22910 8338
rect 22910 2378 22944 8338
rect 22944 2378 22959 8338
rect 23051 2378 23068 8338
rect 23068 2378 23102 8338
rect 23102 2378 23117 8338
rect 23209 2378 23226 8338
rect 23226 2378 23260 8338
rect 23260 2378 23275 8338
rect 23367 2378 23384 8338
rect 23384 2378 23418 8338
rect 23418 2378 23433 8338
rect 23525 2378 23542 8338
rect 23542 2378 23576 8338
rect 23576 2378 23591 8338
rect 23683 2378 23700 8338
rect 23700 2378 23734 8338
rect 23734 2378 23749 8338
rect 23841 2378 23858 8338
rect 23858 2378 23892 8338
rect 23892 2378 23907 8338
rect 23999 2378 24016 8338
rect 24016 2378 24050 8338
rect 24050 2378 24065 8338
rect 24157 2378 24174 8338
rect 24174 2378 24208 8338
rect 24208 2378 24223 8338
rect 24315 2378 24332 8338
rect 24332 2378 24366 8338
rect 24366 2378 24381 8338
rect 24473 2378 24490 8338
rect 24490 2378 24524 8338
rect 24524 2378 24539 8338
rect 24631 2378 24648 8338
rect 24648 2378 24682 8338
rect 24682 2378 24697 8338
rect 24789 2378 24806 8338
rect 24806 2378 24840 8338
rect 24840 2378 24855 8338
rect 24947 2378 24964 8338
rect 24964 2378 24998 8338
rect 24998 2378 25013 8338
rect 25105 2378 25122 8338
rect 25122 2378 25156 8338
rect 25156 2378 25171 8338
rect 20230 2200 20300 2336
rect 25240 2336 25254 8380
rect 25254 2336 25292 8380
rect 25292 2336 25310 8380
rect 25520 8150 25590 8350
rect 25910 8150 25980 8350
rect 26020 8150 26090 8350
rect 26410 8150 26480 8350
rect 25650 8020 25850 8090
rect 26150 8020 26350 8090
rect 25650 7910 25850 7980
rect 26150 7910 26350 7980
rect 25520 7650 25590 7850
rect 25910 7650 25980 7850
rect 26020 7650 26090 7850
rect 26410 7650 26480 7850
rect 25650 7520 25850 7590
rect 26150 7520 26350 7590
rect 25650 7410 25850 7480
rect 26150 7410 26350 7480
rect 25520 7150 25590 7350
rect 25910 7150 25980 7350
rect 26020 7150 26090 7350
rect 26410 7150 26480 7350
rect 25650 7020 25850 7090
rect 26150 7020 26350 7090
rect 25650 6910 25850 6980
rect 26150 6910 26350 6980
rect 25520 6650 25590 6850
rect 25910 6650 25980 6850
rect 26020 6650 26090 6850
rect 26410 6650 26480 6850
rect 25650 6520 25850 6590
rect 26150 6520 26350 6590
rect 25650 6410 25850 6480
rect 26150 6410 26350 6480
rect 25520 6150 25590 6350
rect 25910 6150 25980 6350
rect 26020 6150 26090 6350
rect 26410 6150 26480 6350
rect 25650 6020 25850 6090
rect 26150 6020 26350 6090
rect 25650 5910 25850 5980
rect 26150 5910 26350 5980
rect 25520 5650 25590 5850
rect 25910 5650 25980 5850
rect 26020 5650 26090 5850
rect 26410 5650 26480 5850
rect 25650 5520 25850 5590
rect 26150 5520 26350 5590
rect 25650 5410 25850 5480
rect 26150 5410 26350 5480
rect 25520 5150 25590 5350
rect 25910 5150 25980 5350
rect 26020 5150 26090 5350
rect 26410 5150 26480 5350
rect 25650 5020 25850 5090
rect 26150 5020 26350 5090
rect 25650 4910 25850 4980
rect 26150 4910 26350 4980
rect 25520 4650 25590 4850
rect 25910 4650 25980 4850
rect 26020 4650 26090 4850
rect 26410 4650 26480 4850
rect 25650 4520 25850 4590
rect 26150 4520 26350 4590
rect 25650 4410 25850 4480
rect 26150 4410 26350 4480
rect 25520 4150 25590 4350
rect 25910 4150 25980 4350
rect 26020 4150 26090 4350
rect 26410 4150 26480 4350
rect 25650 4020 25850 4090
rect 26150 4020 26350 4090
rect 25650 3910 25850 3980
rect 26150 3910 26350 3980
rect 25520 3650 25590 3850
rect 25910 3650 25980 3850
rect 26020 3650 26090 3850
rect 26410 3650 26480 3850
rect 25650 3520 25850 3590
rect 26150 3520 26350 3590
rect 25650 3410 25850 3480
rect 26150 3410 26350 3480
rect 25520 3150 25590 3350
rect 25910 3150 25980 3350
rect 26020 3150 26090 3350
rect 26410 3150 26480 3350
rect 25650 3020 25850 3090
rect 26150 3020 26350 3090
rect 25650 2910 25850 2980
rect 26150 2910 26350 2980
rect 25520 2650 25590 2850
rect 25910 2650 25980 2850
rect 26020 2650 26090 2850
rect 26410 2650 26480 2850
rect 25650 2520 25850 2590
rect 26150 2520 26350 2590
rect 25650 2410 25850 2480
rect 26150 2410 26350 2480
rect 20452 2320 25086 2326
rect 20452 2286 20512 2320
rect 20512 2286 20602 2320
rect 20602 2286 20670 2320
rect 20670 2286 20760 2320
rect 20760 2286 20828 2320
rect 20828 2286 20918 2320
rect 20918 2286 20986 2320
rect 20986 2286 21076 2320
rect 21076 2286 21144 2320
rect 21144 2286 21234 2320
rect 21234 2286 21302 2320
rect 21302 2286 21392 2320
rect 21392 2286 21460 2320
rect 21460 2286 21550 2320
rect 21550 2286 21618 2320
rect 21618 2286 21708 2320
rect 21708 2286 21776 2320
rect 21776 2286 21866 2320
rect 21866 2286 21934 2320
rect 21934 2286 22024 2320
rect 22024 2286 22092 2320
rect 22092 2286 22182 2320
rect 22182 2286 22250 2320
rect 22250 2286 22340 2320
rect 22340 2286 22408 2320
rect 22408 2286 22498 2320
rect 22498 2286 22566 2320
rect 22566 2286 22656 2320
rect 22656 2286 22724 2320
rect 22724 2286 22814 2320
rect 22814 2286 22882 2320
rect 22882 2286 22972 2320
rect 22972 2286 23040 2320
rect 23040 2286 23130 2320
rect 23130 2286 23198 2320
rect 23198 2286 23288 2320
rect 23288 2286 23356 2320
rect 23356 2286 23446 2320
rect 23446 2286 23514 2320
rect 23514 2286 23604 2320
rect 23604 2286 23672 2320
rect 23672 2286 23762 2320
rect 23762 2286 23830 2320
rect 23830 2286 23920 2320
rect 23920 2286 23988 2320
rect 23988 2286 24078 2320
rect 24078 2286 24146 2320
rect 24146 2286 24236 2320
rect 24236 2286 24304 2320
rect 24304 2286 24394 2320
rect 24394 2286 24462 2320
rect 24462 2286 24552 2320
rect 24552 2286 24620 2320
rect 24620 2286 24710 2320
rect 24710 2286 24778 2320
rect 24778 2286 24868 2320
rect 24868 2286 24936 2320
rect 24936 2286 25026 2320
rect 25026 2286 25086 2320
rect 20452 2226 25086 2286
rect 25240 2200 25310 2336
rect 25520 2150 25590 2350
rect 25910 2150 25980 2350
rect 26020 2150 26090 2350
rect 26410 2150 26480 2350
rect 150 2020 350 2090
rect 650 2020 850 2090
rect 6650 2020 6850 2090
rect 7150 2020 7350 2090
rect 13150 2020 13350 2090
rect 19650 2020 19850 2090
rect 25650 2020 25850 2090
rect 26150 2020 26350 2090
rect 150 1910 350 1980
rect 650 1910 850 1980
rect 1150 1910 1350 1980
rect 1650 1910 1850 1980
rect 2150 1910 2350 1980
rect 2650 1910 2850 1980
rect 3150 1910 3350 1980
rect 3650 1910 3850 1980
rect 4150 1910 4350 1980
rect 4650 1910 4850 1980
rect 5150 1910 5350 1980
rect 5650 1910 5850 1980
rect 6150 1910 6350 1980
rect 6650 1910 6850 1980
rect 7150 1910 7350 1980
rect 7650 1910 7850 1980
rect 8150 1910 8350 1980
rect 8650 1910 8850 1980
rect 9150 1910 9350 1980
rect 9650 1910 9850 1980
rect 10150 1910 10350 1980
rect 10650 1910 10850 1980
rect 11150 1910 11350 1980
rect 11650 1910 11850 1980
rect 12150 1910 12350 1980
rect 12650 1910 12850 1980
rect 13150 1910 13350 1980
rect 13650 1910 13850 1980
rect 14150 1910 14350 1980
rect 14650 1910 14850 1980
rect 15150 1910 15350 1980
rect 15650 1910 15850 1980
rect 16150 1910 16350 1980
rect 16650 1910 16850 1980
rect 17150 1910 17350 1980
rect 17650 1910 17850 1980
rect 18150 1910 18350 1980
rect 18650 1910 18850 1980
rect 19150 1910 19350 1980
rect 19650 1910 19850 1980
rect 20150 1910 20350 1980
rect 20650 1910 20850 1980
rect 21150 1910 21350 1980
rect 21650 1910 21850 1980
rect 22150 1910 22350 1980
rect 22650 1910 22850 1980
rect 23150 1910 23350 1980
rect 23650 1910 23850 1980
rect 24150 1910 24350 1980
rect 24650 1910 24850 1980
rect 25150 1910 25350 1980
rect 25650 1910 25850 1980
rect 26150 1910 26350 1980
rect 20 1650 90 1850
rect 410 1650 480 1850
rect 520 1650 590 1850
rect 910 1650 980 1850
rect 1020 1650 1090 1850
rect 1410 1650 1480 1850
rect 1520 1650 1590 1850
rect 1910 1650 1980 1850
rect 2020 1650 2090 1850
rect 2410 1650 2480 1850
rect 2520 1650 2590 1850
rect 2910 1650 2980 1850
rect 3020 1650 3090 1850
rect 3410 1650 3480 1850
rect 3520 1650 3590 1850
rect 3910 1650 3980 1850
rect 4020 1650 4090 1850
rect 4410 1650 4480 1850
rect 4520 1650 4590 1850
rect 4910 1650 4980 1850
rect 5020 1650 5090 1850
rect 5410 1650 5480 1850
rect 5520 1650 5590 1850
rect 5910 1650 5980 1850
rect 6020 1650 6090 1850
rect 6410 1650 6480 1850
rect 6520 1650 6590 1850
rect 6910 1650 6980 1850
rect 7020 1650 7090 1850
rect 7410 1650 7480 1850
rect 7520 1650 7590 1850
rect 7910 1650 7980 1850
rect 8020 1650 8090 1850
rect 8410 1650 8480 1850
rect 8520 1650 8590 1850
rect 8910 1650 8980 1850
rect 9020 1650 9090 1850
rect 9410 1650 9480 1850
rect 9520 1650 9590 1850
rect 9910 1650 9980 1850
rect 10020 1650 10090 1850
rect 10410 1650 10480 1850
rect 10520 1650 10590 1850
rect 10910 1650 10980 1850
rect 11020 1650 11090 1850
rect 11410 1650 11480 1850
rect 11520 1650 11590 1850
rect 11910 1650 11980 1850
rect 12020 1650 12090 1850
rect 12410 1650 12480 1850
rect 12520 1650 12590 1850
rect 12910 1650 12980 1850
rect 13020 1650 13090 1850
rect 13410 1650 13480 1850
rect 13520 1650 13590 1850
rect 13910 1650 13980 1850
rect 14020 1650 14090 1850
rect 14410 1650 14480 1850
rect 14520 1650 14590 1850
rect 14910 1650 14980 1850
rect 15020 1650 15090 1850
rect 15410 1650 15480 1850
rect 15520 1650 15590 1850
rect 15910 1650 15980 1850
rect 16020 1650 16090 1850
rect 16410 1650 16480 1850
rect 16520 1650 16590 1850
rect 16910 1650 16980 1850
rect 17020 1650 17090 1850
rect 17410 1650 17480 1850
rect 17520 1650 17590 1850
rect 17910 1650 17980 1850
rect 18020 1650 18090 1850
rect 18410 1650 18480 1850
rect 18520 1650 18590 1850
rect 18910 1650 18980 1850
rect 19020 1650 19090 1850
rect 19410 1650 19480 1850
rect 19520 1650 19590 1850
rect 19910 1650 19980 1850
rect 20020 1650 20090 1850
rect 20410 1650 20480 1850
rect 20520 1650 20590 1850
rect 20910 1650 20980 1850
rect 21020 1650 21090 1850
rect 21410 1650 21480 1850
rect 21520 1650 21590 1850
rect 21910 1650 21980 1850
rect 22020 1650 22090 1850
rect 22410 1650 22480 1850
rect 22520 1650 22590 1850
rect 22910 1650 22980 1850
rect 23020 1650 23090 1850
rect 23410 1650 23480 1850
rect 23520 1650 23590 1850
rect 23910 1650 23980 1850
rect 24020 1650 24090 1850
rect 24410 1650 24480 1850
rect 24520 1650 24590 1850
rect 24910 1650 24980 1850
rect 25020 1650 25090 1850
rect 25410 1650 25480 1850
rect 25520 1650 25590 1850
rect 25910 1650 25980 1850
rect 26020 1650 26090 1850
rect 26410 1650 26480 1850
rect 150 1520 350 1590
rect 650 1520 850 1590
rect 1150 1520 1350 1590
rect 1650 1520 1850 1590
rect 2150 1520 2350 1590
rect 2650 1520 2850 1590
rect 3150 1520 3350 1590
rect 3650 1520 3850 1590
rect 4150 1520 4350 1590
rect 4650 1520 4850 1590
rect 5150 1520 5350 1590
rect 5650 1520 5850 1590
rect 6150 1520 6350 1590
rect 6650 1520 6850 1590
rect 7150 1520 7350 1590
rect 7650 1520 7850 1590
rect 8150 1520 8350 1590
rect 8650 1520 8850 1590
rect 9150 1520 9350 1590
rect 9650 1520 9850 1590
rect 10150 1520 10350 1590
rect 10650 1520 10850 1590
rect 11150 1520 11350 1590
rect 11650 1520 11850 1590
rect 12150 1520 12350 1590
rect 12650 1520 12850 1590
rect 13150 1520 13350 1590
rect 13650 1520 13850 1590
rect 14150 1520 14350 1590
rect 14650 1520 14850 1590
rect 15150 1520 15350 1590
rect 15650 1520 15850 1590
rect 16150 1520 16350 1590
rect 16650 1520 16850 1590
rect 17150 1520 17350 1590
rect 17650 1520 17850 1590
rect 18150 1520 18350 1590
rect 18650 1520 18850 1590
rect 19150 1520 19350 1590
rect 19650 1520 19850 1590
rect 20150 1520 20350 1590
rect 20650 1520 20850 1590
rect 21150 1520 21350 1590
rect 21650 1520 21850 1590
rect 22150 1520 22350 1590
rect 22650 1520 22850 1590
rect 23150 1520 23350 1590
rect 23650 1520 23850 1590
rect 24150 1520 24350 1590
rect 24650 1520 24850 1590
rect 25150 1520 25350 1590
rect 25650 1520 25850 1590
rect 26150 1520 26350 1590
rect 150 1410 350 1480
rect 650 1410 850 1480
rect 1150 1410 1350 1480
rect 1650 1410 1850 1480
rect 2150 1410 2350 1480
rect 2650 1410 2850 1480
rect 3150 1410 3350 1480
rect 3650 1410 3850 1480
rect 4150 1410 4350 1480
rect 4650 1410 4850 1480
rect 5150 1410 5350 1480
rect 5650 1410 5850 1480
rect 6150 1410 6350 1480
rect 6650 1410 6850 1480
rect 7150 1410 7350 1480
rect 7650 1410 7850 1480
rect 8150 1410 8350 1480
rect 8650 1410 8850 1480
rect 9150 1410 9350 1480
rect 9650 1410 9850 1480
rect 10150 1410 10350 1480
rect 10650 1410 10850 1480
rect 11150 1410 11350 1480
rect 11650 1410 11850 1480
rect 12150 1410 12350 1480
rect 12650 1410 12850 1480
rect 13150 1410 13350 1480
rect 13650 1410 13850 1480
rect 14150 1410 14350 1480
rect 14650 1410 14850 1480
rect 15150 1410 15350 1480
rect 15650 1410 15850 1480
rect 16150 1410 16350 1480
rect 16650 1410 16850 1480
rect 17150 1410 17350 1480
rect 17650 1410 17850 1480
rect 18150 1410 18350 1480
rect 18650 1410 18850 1480
rect 19150 1410 19350 1480
rect 19650 1410 19850 1480
rect 20150 1410 20350 1480
rect 20650 1410 20850 1480
rect 21150 1410 21350 1480
rect 21650 1410 21850 1480
rect 22150 1410 22350 1480
rect 22650 1410 22850 1480
rect 23150 1410 23350 1480
rect 23650 1410 23850 1480
rect 24150 1410 24350 1480
rect 24650 1410 24850 1480
rect 25150 1410 25350 1480
rect 25650 1410 25850 1480
rect 26150 1410 26350 1480
rect 20 1150 90 1350
rect 410 1150 480 1350
rect 520 1150 590 1350
rect 910 1150 980 1350
rect 1020 1150 1090 1350
rect 1410 1150 1480 1350
rect 1520 1150 1590 1350
rect 1910 1150 1980 1350
rect 2020 1150 2090 1350
rect 2410 1150 2480 1350
rect 2520 1150 2590 1350
rect 2910 1150 2980 1350
rect 3020 1150 3090 1350
rect 3410 1150 3480 1350
rect 3520 1150 3590 1350
rect 3910 1150 3980 1350
rect 4020 1150 4090 1350
rect 4410 1150 4480 1350
rect 4520 1150 4590 1350
rect 4910 1150 4980 1350
rect 5020 1150 5090 1350
rect 5410 1150 5480 1350
rect 5520 1150 5590 1350
rect 5910 1150 5980 1350
rect 6020 1150 6090 1350
rect 6410 1150 6480 1350
rect 6520 1150 6590 1350
rect 6910 1150 6980 1350
rect 7020 1150 7090 1350
rect 7410 1150 7480 1350
rect 7520 1150 7590 1350
rect 7910 1150 7980 1350
rect 8020 1150 8090 1350
rect 8410 1150 8480 1350
rect 8520 1150 8590 1350
rect 8910 1150 8980 1350
rect 9020 1150 9090 1350
rect 9410 1150 9480 1350
rect 9520 1150 9590 1350
rect 9910 1150 9980 1350
rect 10020 1150 10090 1350
rect 10410 1150 10480 1350
rect 10520 1150 10590 1350
rect 10910 1150 10980 1350
rect 11020 1150 11090 1350
rect 11410 1150 11480 1350
rect 11520 1150 11590 1350
rect 11910 1150 11980 1350
rect 12020 1150 12090 1350
rect 12410 1150 12480 1350
rect 12520 1150 12590 1350
rect 12910 1150 12980 1350
rect 13020 1150 13090 1350
rect 13410 1150 13480 1350
rect 13520 1150 13590 1350
rect 13910 1150 13980 1350
rect 14020 1150 14090 1350
rect 14410 1150 14480 1350
rect 14520 1150 14590 1350
rect 14910 1150 14980 1350
rect 15020 1150 15090 1350
rect 15410 1150 15480 1350
rect 15520 1150 15590 1350
rect 15910 1150 15980 1350
rect 16020 1150 16090 1350
rect 16410 1150 16480 1350
rect 16520 1150 16590 1350
rect 16910 1150 16980 1350
rect 17020 1150 17090 1350
rect 17410 1150 17480 1350
rect 17520 1150 17590 1350
rect 17910 1150 17980 1350
rect 18020 1150 18090 1350
rect 18410 1150 18480 1350
rect 18520 1150 18590 1350
rect 18910 1150 18980 1350
rect 19020 1150 19090 1350
rect 19410 1150 19480 1350
rect 19520 1150 19590 1350
rect 19910 1150 19980 1350
rect 20020 1150 20090 1350
rect 20410 1150 20480 1350
rect 20520 1150 20590 1350
rect 20910 1150 20980 1350
rect 21020 1150 21090 1350
rect 21410 1150 21480 1350
rect 21520 1150 21590 1350
rect 21910 1150 21980 1350
rect 22020 1150 22090 1350
rect 22410 1150 22480 1350
rect 22520 1150 22590 1350
rect 22910 1150 22980 1350
rect 23020 1150 23090 1350
rect 23410 1150 23480 1350
rect 23520 1150 23590 1350
rect 23910 1150 23980 1350
rect 24020 1150 24090 1350
rect 24410 1150 24480 1350
rect 24520 1150 24590 1350
rect 24910 1150 24980 1350
rect 25020 1150 25090 1350
rect 25410 1150 25480 1350
rect 25520 1150 25590 1350
rect 25910 1150 25980 1350
rect 26020 1150 26090 1350
rect 26410 1150 26480 1350
rect 150 1020 350 1090
rect 650 1020 850 1090
rect 1150 1020 1350 1090
rect 1650 1020 1850 1090
rect 2150 1020 2350 1090
rect 2650 1020 2850 1090
rect 3150 1020 3350 1090
rect 3650 1020 3850 1090
rect 4150 1020 4350 1090
rect 4650 1020 4850 1090
rect 5150 1020 5350 1090
rect 5650 1020 5850 1090
rect 6150 1020 6350 1090
rect 6650 1020 6850 1090
rect 7150 1020 7350 1090
rect 7650 1020 7850 1090
rect 8150 1020 8350 1090
rect 8650 1020 8850 1090
rect 9150 1020 9350 1090
rect 9650 1020 9850 1090
rect 10150 1020 10350 1090
rect 10650 1020 10850 1090
rect 11150 1020 11350 1090
rect 11650 1020 11850 1090
rect 12150 1020 12350 1090
rect 12650 1020 12850 1090
rect 13150 1020 13350 1090
rect 13650 1020 13850 1090
rect 14150 1020 14350 1090
rect 14650 1020 14850 1090
rect 15150 1020 15350 1090
rect 15650 1020 15850 1090
rect 16150 1020 16350 1090
rect 16650 1020 16850 1090
rect 17150 1020 17350 1090
rect 17650 1020 17850 1090
rect 18150 1020 18350 1090
rect 18650 1020 18850 1090
rect 19150 1020 19350 1090
rect 19650 1020 19850 1090
rect 20150 1020 20350 1090
rect 20650 1020 20850 1090
rect 21150 1020 21350 1090
rect 21650 1020 21850 1090
rect 22150 1020 22350 1090
rect 22650 1020 22850 1090
rect 23150 1020 23350 1090
rect 23650 1020 23850 1090
rect 24150 1020 24350 1090
rect 24650 1020 24850 1090
rect 25150 1020 25350 1090
rect 25650 1020 25850 1090
rect 26150 1020 26350 1090
<< metal2 >>
rect 140 47480 360 47500
rect 140 47410 150 47480
rect 350 47410 360 47480
rect 140 47360 360 47410
rect 640 47480 860 47500
rect 640 47410 650 47480
rect 850 47410 860 47480
rect 640 47360 860 47410
rect 1140 47480 1360 47500
rect 1140 47410 1150 47480
rect 1350 47410 1360 47480
rect 1140 47360 1360 47410
rect 1640 47480 1860 47500
rect 1640 47410 1650 47480
rect 1850 47410 1860 47480
rect 1640 47360 1860 47410
rect 2140 47480 2360 47500
rect 2140 47410 2150 47480
rect 2350 47410 2360 47480
rect 2140 47360 2360 47410
rect 2640 47480 2860 47500
rect 2640 47410 2650 47480
rect 2850 47410 2860 47480
rect 2640 47360 2860 47410
rect 3140 47480 3360 47500
rect 3140 47410 3150 47480
rect 3350 47410 3360 47480
rect 3140 47360 3360 47410
rect 3640 47480 3860 47500
rect 3640 47410 3650 47480
rect 3850 47410 3860 47480
rect 3640 47360 3860 47410
rect 4140 47480 4360 47500
rect 4140 47410 4150 47480
rect 4350 47410 4360 47480
rect 4140 47360 4360 47410
rect 4640 47480 4860 47500
rect 4640 47410 4650 47480
rect 4850 47410 4860 47480
rect 4640 47360 4860 47410
rect 5140 47480 5360 47500
rect 5140 47410 5150 47480
rect 5350 47410 5360 47480
rect 5140 47360 5360 47410
rect 5640 47480 5860 47500
rect 5640 47410 5650 47480
rect 5850 47410 5860 47480
rect 5640 47360 5860 47410
rect 6140 47480 6360 47500
rect 6140 47410 6150 47480
rect 6350 47410 6360 47480
rect 6140 47360 6360 47410
rect 6640 47480 6860 47500
rect 6640 47410 6650 47480
rect 6850 47410 6860 47480
rect 6640 47360 6860 47410
rect 7140 47480 7360 47500
rect 7140 47410 7150 47480
rect 7350 47410 7360 47480
rect 7140 47360 7360 47410
rect 7640 47480 7860 47500
rect 7640 47410 7650 47480
rect 7850 47410 7860 47480
rect 7640 47360 7860 47410
rect 8140 47480 8360 47500
rect 8140 47410 8150 47480
rect 8350 47410 8360 47480
rect 8140 47360 8360 47410
rect 8640 47480 8860 47500
rect 8640 47410 8650 47480
rect 8850 47410 8860 47480
rect 8640 47360 8860 47410
rect 9140 47480 9360 47500
rect 9140 47410 9150 47480
rect 9350 47410 9360 47480
rect 9140 47360 9360 47410
rect 9640 47480 9860 47500
rect 9640 47410 9650 47480
rect 9850 47410 9860 47480
rect 9640 47360 9860 47410
rect 10140 47480 10360 47500
rect 10140 47410 10150 47480
rect 10350 47410 10360 47480
rect 10140 47360 10360 47410
rect 10640 47480 10860 47500
rect 10640 47410 10650 47480
rect 10850 47410 10860 47480
rect 10640 47360 10860 47410
rect 11140 47480 11360 47500
rect 11140 47410 11150 47480
rect 11350 47410 11360 47480
rect 11140 47360 11360 47410
rect 11640 47480 11860 47500
rect 11640 47410 11650 47480
rect 11850 47410 11860 47480
rect 11640 47360 11860 47410
rect 12140 47480 12360 47500
rect 12140 47410 12150 47480
rect 12350 47410 12360 47480
rect 12140 47360 12360 47410
rect 12640 47480 12860 47500
rect 12640 47410 12650 47480
rect 12850 47410 12860 47480
rect 12640 47360 12860 47410
rect 13140 47480 13360 47500
rect 13140 47410 13150 47480
rect 13350 47410 13360 47480
rect 13140 47360 13360 47410
rect 13640 47480 13860 47500
rect 13640 47410 13650 47480
rect 13850 47410 13860 47480
rect 13640 47360 13860 47410
rect 14140 47480 14360 47500
rect 14140 47410 14150 47480
rect 14350 47410 14360 47480
rect 14140 47360 14360 47410
rect 14640 47480 14860 47500
rect 14640 47410 14650 47480
rect 14850 47410 14860 47480
rect 14640 47360 14860 47410
rect 15140 47480 15360 47500
rect 15140 47410 15150 47480
rect 15350 47410 15360 47480
rect 15140 47360 15360 47410
rect 15640 47480 15860 47500
rect 15640 47410 15650 47480
rect 15850 47410 15860 47480
rect 15640 47360 15860 47410
rect 16140 47480 16360 47500
rect 16140 47410 16150 47480
rect 16350 47410 16360 47480
rect 16140 47360 16360 47410
rect 16640 47480 16860 47500
rect 16640 47410 16650 47480
rect 16850 47410 16860 47480
rect 16640 47360 16860 47410
rect 17140 47480 17360 47500
rect 17140 47410 17150 47480
rect 17350 47410 17360 47480
rect 17140 47360 17360 47410
rect 17640 47480 17860 47500
rect 17640 47410 17650 47480
rect 17850 47410 17860 47480
rect 17640 47360 17860 47410
rect 18140 47480 18360 47500
rect 18140 47410 18150 47480
rect 18350 47410 18360 47480
rect 18140 47360 18360 47410
rect 18640 47480 18860 47500
rect 18640 47410 18650 47480
rect 18850 47410 18860 47480
rect 18640 47360 18860 47410
rect 19140 47480 19360 47500
rect 19140 47410 19150 47480
rect 19350 47410 19360 47480
rect 19140 47360 19360 47410
rect 19640 47480 19860 47500
rect 19640 47410 19650 47480
rect 19850 47410 19860 47480
rect 19640 47360 19860 47410
rect 20140 47480 20360 47500
rect 20140 47410 20150 47480
rect 20350 47410 20360 47480
rect 20140 47360 20360 47410
rect 20640 47480 20860 47500
rect 20640 47410 20650 47480
rect 20850 47410 20860 47480
rect 20640 47360 20860 47410
rect 21140 47480 21360 47500
rect 21140 47410 21150 47480
rect 21350 47410 21360 47480
rect 21140 47360 21360 47410
rect 21640 47480 21860 47500
rect 21640 47410 21650 47480
rect 21850 47410 21860 47480
rect 21640 47360 21860 47410
rect 22140 47480 22360 47500
rect 22140 47410 22150 47480
rect 22350 47410 22360 47480
rect 22140 47360 22360 47410
rect 22640 47480 22860 47500
rect 22640 47410 22650 47480
rect 22850 47410 22860 47480
rect 22640 47360 22860 47410
rect 23140 47480 23360 47500
rect 23140 47410 23150 47480
rect 23350 47410 23360 47480
rect 23140 47360 23360 47410
rect 23640 47480 23860 47500
rect 23640 47410 23650 47480
rect 23850 47410 23860 47480
rect 23640 47360 23860 47410
rect 24140 47480 24360 47500
rect 24140 47410 24150 47480
rect 24350 47410 24360 47480
rect 24140 47360 24360 47410
rect 24640 47480 24860 47500
rect 24640 47410 24650 47480
rect 24850 47410 24860 47480
rect 24640 47360 24860 47410
rect 25140 47480 25360 47500
rect 25140 47410 25150 47480
rect 25350 47410 25360 47480
rect 25140 47360 25360 47410
rect 25640 47480 25860 47500
rect 25640 47410 25650 47480
rect 25850 47410 25860 47480
rect 25640 47360 25860 47410
rect 26140 47480 26360 47500
rect 26140 47410 26150 47480
rect 26350 47410 26360 47480
rect 26140 47360 26360 47410
rect 0 47350 26500 47360
rect 0 47150 20 47350
rect 90 47150 410 47350
rect 480 47150 520 47350
rect 590 47150 910 47350
rect 980 47150 1020 47350
rect 1090 47150 1410 47350
rect 1480 47150 1520 47350
rect 1590 47150 1910 47350
rect 1980 47150 2020 47350
rect 2090 47150 2410 47350
rect 2480 47150 2520 47350
rect 2590 47150 2910 47350
rect 2980 47150 3020 47350
rect 3090 47150 3410 47350
rect 3480 47150 3520 47350
rect 3590 47150 3910 47350
rect 3980 47150 4020 47350
rect 4090 47150 4410 47350
rect 4480 47150 4520 47350
rect 4590 47150 4910 47350
rect 4980 47150 5020 47350
rect 5090 47150 5410 47350
rect 5480 47150 5520 47350
rect 5590 47150 5910 47350
rect 5980 47150 6020 47350
rect 6090 47150 6410 47350
rect 6480 47150 6520 47350
rect 6590 47150 6910 47350
rect 6980 47150 7020 47350
rect 7090 47150 7410 47350
rect 7480 47150 7520 47350
rect 7590 47150 7910 47350
rect 7980 47150 8020 47350
rect 8090 47150 8410 47350
rect 8480 47150 8520 47350
rect 8590 47150 8910 47350
rect 8980 47150 9020 47350
rect 9090 47150 9410 47350
rect 9480 47150 9520 47350
rect 9590 47150 9910 47350
rect 9980 47150 10020 47350
rect 10090 47150 10410 47350
rect 10480 47150 10520 47350
rect 10590 47150 10910 47350
rect 10980 47150 11020 47350
rect 11090 47150 11410 47350
rect 11480 47150 11520 47350
rect 11590 47150 11910 47350
rect 11980 47150 12020 47350
rect 12090 47150 12410 47350
rect 12480 47150 12520 47350
rect 12590 47150 12910 47350
rect 12980 47150 13020 47350
rect 13090 47150 13410 47350
rect 13480 47150 13520 47350
rect 13590 47150 13910 47350
rect 13980 47150 14020 47350
rect 14090 47150 14410 47350
rect 14480 47150 14520 47350
rect 14590 47150 14910 47350
rect 14980 47150 15020 47350
rect 15090 47150 15410 47350
rect 15480 47150 15520 47350
rect 15590 47150 15910 47350
rect 15980 47150 16020 47350
rect 16090 47150 16410 47350
rect 16480 47150 16520 47350
rect 16590 47150 16910 47350
rect 16980 47150 17020 47350
rect 17090 47150 17410 47350
rect 17480 47150 17520 47350
rect 17590 47150 17910 47350
rect 17980 47150 18020 47350
rect 18090 47150 18410 47350
rect 18480 47150 18520 47350
rect 18590 47150 18910 47350
rect 18980 47150 19020 47350
rect 19090 47150 19410 47350
rect 19480 47150 19520 47350
rect 19590 47150 19910 47350
rect 19980 47150 20020 47350
rect 20090 47150 20410 47350
rect 20480 47150 20520 47350
rect 20590 47150 20910 47350
rect 20980 47150 21020 47350
rect 21090 47150 21410 47350
rect 21480 47150 21520 47350
rect 21590 47150 21910 47350
rect 21980 47150 22020 47350
rect 22090 47150 22410 47350
rect 22480 47150 22520 47350
rect 22590 47150 22910 47350
rect 22980 47150 23020 47350
rect 23090 47150 23410 47350
rect 23480 47150 23520 47350
rect 23590 47150 23910 47350
rect 23980 47150 24020 47350
rect 24090 47150 24410 47350
rect 24480 47150 24520 47350
rect 24590 47150 24910 47350
rect 24980 47150 25020 47350
rect 25090 47150 25410 47350
rect 25480 47150 25520 47350
rect 25590 47150 25910 47350
rect 25980 47150 26020 47350
rect 26090 47150 26410 47350
rect 26480 47150 26500 47350
rect 0 47140 26500 47150
rect 140 47090 360 47140
rect 140 47020 150 47090
rect 350 47020 360 47090
rect 140 46980 360 47020
rect 140 46910 150 46980
rect 350 46910 360 46980
rect 140 46860 360 46910
rect 640 47090 860 47140
rect 640 47020 650 47090
rect 850 47020 860 47090
rect 640 46980 860 47020
rect 640 46910 650 46980
rect 850 46910 860 46980
rect 640 46860 860 46910
rect 1140 47090 1360 47140
rect 1140 47020 1150 47090
rect 1350 47020 1360 47090
rect 1140 46980 1360 47020
rect 1140 46910 1150 46980
rect 1350 46910 1360 46980
rect 1140 46860 1360 46910
rect 1640 47090 1860 47140
rect 1640 47020 1650 47090
rect 1850 47020 1860 47090
rect 1640 46980 1860 47020
rect 1640 46910 1650 46980
rect 1850 46910 1860 46980
rect 1640 46860 1860 46910
rect 2140 47090 2360 47140
rect 2140 47020 2150 47090
rect 2350 47020 2360 47090
rect 2140 46980 2360 47020
rect 2140 46910 2150 46980
rect 2350 46910 2360 46980
rect 2140 46860 2360 46910
rect 2640 47090 2860 47140
rect 2640 47020 2650 47090
rect 2850 47020 2860 47090
rect 2640 46980 2860 47020
rect 2640 46910 2650 46980
rect 2850 46910 2860 46980
rect 2640 46860 2860 46910
rect 3140 47090 3360 47140
rect 3140 47020 3150 47090
rect 3350 47020 3360 47090
rect 3140 46980 3360 47020
rect 3140 46910 3150 46980
rect 3350 46910 3360 46980
rect 3140 46860 3360 46910
rect 3640 47090 3860 47140
rect 3640 47020 3650 47090
rect 3850 47020 3860 47090
rect 3640 46980 3860 47020
rect 3640 46910 3650 46980
rect 3850 46910 3860 46980
rect 3640 46860 3860 46910
rect 4140 47090 4360 47140
rect 4140 47020 4150 47090
rect 4350 47020 4360 47090
rect 4140 46980 4360 47020
rect 4140 46910 4150 46980
rect 4350 46910 4360 46980
rect 4140 46860 4360 46910
rect 4640 47090 4860 47140
rect 4640 47020 4650 47090
rect 4850 47020 4860 47090
rect 4640 46980 4860 47020
rect 4640 46910 4650 46980
rect 4850 46910 4860 46980
rect 4640 46860 4860 46910
rect 5140 47090 5360 47140
rect 5140 47020 5150 47090
rect 5350 47020 5360 47090
rect 5140 46980 5360 47020
rect 5140 46910 5150 46980
rect 5350 46910 5360 46980
rect 5140 46860 5360 46910
rect 5640 47090 5860 47140
rect 5640 47020 5650 47090
rect 5850 47020 5860 47090
rect 5640 46980 5860 47020
rect 5640 46910 5650 46980
rect 5850 46910 5860 46980
rect 5640 46860 5860 46910
rect 6140 47090 6360 47140
rect 6140 47020 6150 47090
rect 6350 47020 6360 47090
rect 6140 46980 6360 47020
rect 6140 46910 6150 46980
rect 6350 46910 6360 46980
rect 6140 46860 6360 46910
rect 6640 47090 6860 47140
rect 6640 47020 6650 47090
rect 6850 47020 6860 47090
rect 6640 46980 6860 47020
rect 6640 46910 6650 46980
rect 6850 46910 6860 46980
rect 6640 46860 6860 46910
rect 7140 47090 7360 47140
rect 7140 47020 7150 47090
rect 7350 47020 7360 47090
rect 7140 46980 7360 47020
rect 7140 46910 7150 46980
rect 7350 46910 7360 46980
rect 7140 46860 7360 46910
rect 7640 47090 7860 47140
rect 7640 47020 7650 47090
rect 7850 47020 7860 47090
rect 7640 46980 7860 47020
rect 7640 46910 7650 46980
rect 7850 46910 7860 46980
rect 7640 46860 7860 46910
rect 8140 47090 8360 47140
rect 8140 47020 8150 47090
rect 8350 47020 8360 47090
rect 8140 46980 8360 47020
rect 8140 46910 8150 46980
rect 8350 46910 8360 46980
rect 8140 46860 8360 46910
rect 8640 47090 8860 47140
rect 8640 47020 8650 47090
rect 8850 47020 8860 47090
rect 8640 46980 8860 47020
rect 8640 46910 8650 46980
rect 8850 46910 8860 46980
rect 8640 46860 8860 46910
rect 9140 47090 9360 47140
rect 9140 47020 9150 47090
rect 9350 47020 9360 47090
rect 9140 46980 9360 47020
rect 9140 46910 9150 46980
rect 9350 46910 9360 46980
rect 9140 46860 9360 46910
rect 9640 47090 9860 47140
rect 9640 47020 9650 47090
rect 9850 47020 9860 47090
rect 9640 46980 9860 47020
rect 9640 46910 9650 46980
rect 9850 46910 9860 46980
rect 9640 46860 9860 46910
rect 10140 47090 10360 47140
rect 10140 47020 10150 47090
rect 10350 47020 10360 47090
rect 10140 46980 10360 47020
rect 10140 46910 10150 46980
rect 10350 46910 10360 46980
rect 10140 46860 10360 46910
rect 10640 47090 10860 47140
rect 10640 47020 10650 47090
rect 10850 47020 10860 47090
rect 10640 46980 10860 47020
rect 10640 46910 10650 46980
rect 10850 46910 10860 46980
rect 10640 46860 10860 46910
rect 11140 47090 11360 47140
rect 11140 47020 11150 47090
rect 11350 47020 11360 47090
rect 11140 46980 11360 47020
rect 11140 46910 11150 46980
rect 11350 46910 11360 46980
rect 11140 46860 11360 46910
rect 11640 47090 11860 47140
rect 11640 47020 11650 47090
rect 11850 47020 11860 47090
rect 11640 46980 11860 47020
rect 11640 46910 11650 46980
rect 11850 46910 11860 46980
rect 11640 46860 11860 46910
rect 12140 47090 12360 47140
rect 12140 47020 12150 47090
rect 12350 47020 12360 47090
rect 12140 46980 12360 47020
rect 12140 46910 12150 46980
rect 12350 46910 12360 46980
rect 12140 46860 12360 46910
rect 12640 47090 12860 47140
rect 12640 47020 12650 47090
rect 12850 47020 12860 47090
rect 12640 46980 12860 47020
rect 12640 46910 12650 46980
rect 12850 46910 12860 46980
rect 12640 46860 12860 46910
rect 13140 47090 13360 47140
rect 13140 47020 13150 47090
rect 13350 47020 13360 47090
rect 13140 46980 13360 47020
rect 13140 46910 13150 46980
rect 13350 46910 13360 46980
rect 13140 46860 13360 46910
rect 13640 47090 13860 47140
rect 13640 47020 13650 47090
rect 13850 47020 13860 47090
rect 13640 46980 13860 47020
rect 13640 46910 13650 46980
rect 13850 46910 13860 46980
rect 13640 46860 13860 46910
rect 14140 47090 14360 47140
rect 14140 47020 14150 47090
rect 14350 47020 14360 47090
rect 14140 46980 14360 47020
rect 14140 46910 14150 46980
rect 14350 46910 14360 46980
rect 14140 46860 14360 46910
rect 14640 47090 14860 47140
rect 14640 47020 14650 47090
rect 14850 47020 14860 47090
rect 14640 46980 14860 47020
rect 14640 46910 14650 46980
rect 14850 46910 14860 46980
rect 14640 46860 14860 46910
rect 15140 47090 15360 47140
rect 15140 47020 15150 47090
rect 15350 47020 15360 47090
rect 15140 46980 15360 47020
rect 15140 46910 15150 46980
rect 15350 46910 15360 46980
rect 15140 46860 15360 46910
rect 15640 47090 15860 47140
rect 15640 47020 15650 47090
rect 15850 47020 15860 47090
rect 15640 46980 15860 47020
rect 15640 46910 15650 46980
rect 15850 46910 15860 46980
rect 15640 46860 15860 46910
rect 16140 47090 16360 47140
rect 16140 47020 16150 47090
rect 16350 47020 16360 47090
rect 16140 46980 16360 47020
rect 16140 46910 16150 46980
rect 16350 46910 16360 46980
rect 16140 46860 16360 46910
rect 16640 47090 16860 47140
rect 16640 47020 16650 47090
rect 16850 47020 16860 47090
rect 16640 46980 16860 47020
rect 16640 46910 16650 46980
rect 16850 46910 16860 46980
rect 16640 46860 16860 46910
rect 17140 47090 17360 47140
rect 17140 47020 17150 47090
rect 17350 47020 17360 47090
rect 17140 46980 17360 47020
rect 17140 46910 17150 46980
rect 17350 46910 17360 46980
rect 17140 46860 17360 46910
rect 17640 47090 17860 47140
rect 17640 47020 17650 47090
rect 17850 47020 17860 47090
rect 17640 46980 17860 47020
rect 17640 46910 17650 46980
rect 17850 46910 17860 46980
rect 17640 46860 17860 46910
rect 18140 47090 18360 47140
rect 18140 47020 18150 47090
rect 18350 47020 18360 47090
rect 18140 46980 18360 47020
rect 18140 46910 18150 46980
rect 18350 46910 18360 46980
rect 18140 46860 18360 46910
rect 18640 47090 18860 47140
rect 18640 47020 18650 47090
rect 18850 47020 18860 47090
rect 18640 46980 18860 47020
rect 18640 46910 18650 46980
rect 18850 46910 18860 46980
rect 18640 46860 18860 46910
rect 19140 47090 19360 47140
rect 19140 47020 19150 47090
rect 19350 47020 19360 47090
rect 19140 46980 19360 47020
rect 19140 46910 19150 46980
rect 19350 46910 19360 46980
rect 19140 46860 19360 46910
rect 19640 47090 19860 47140
rect 19640 47020 19650 47090
rect 19850 47020 19860 47090
rect 19640 46980 19860 47020
rect 19640 46910 19650 46980
rect 19850 46910 19860 46980
rect 19640 46860 19860 46910
rect 20140 47090 20360 47140
rect 20140 47020 20150 47090
rect 20350 47020 20360 47090
rect 20140 46980 20360 47020
rect 20140 46910 20150 46980
rect 20350 46910 20360 46980
rect 20140 46860 20360 46910
rect 20640 47090 20860 47140
rect 20640 47020 20650 47090
rect 20850 47020 20860 47090
rect 20640 46980 20860 47020
rect 20640 46910 20650 46980
rect 20850 46910 20860 46980
rect 20640 46860 20860 46910
rect 21140 47090 21360 47140
rect 21140 47020 21150 47090
rect 21350 47020 21360 47090
rect 21140 46980 21360 47020
rect 21140 46910 21150 46980
rect 21350 46910 21360 46980
rect 21140 46860 21360 46910
rect 21640 47090 21860 47140
rect 21640 47020 21650 47090
rect 21850 47020 21860 47090
rect 21640 46980 21860 47020
rect 21640 46910 21650 46980
rect 21850 46910 21860 46980
rect 21640 46860 21860 46910
rect 22140 47090 22360 47140
rect 22140 47020 22150 47090
rect 22350 47020 22360 47090
rect 22140 46980 22360 47020
rect 22140 46910 22150 46980
rect 22350 46910 22360 46980
rect 22140 46860 22360 46910
rect 22640 47090 22860 47140
rect 22640 47020 22650 47090
rect 22850 47020 22860 47090
rect 22640 46980 22860 47020
rect 22640 46910 22650 46980
rect 22850 46910 22860 46980
rect 22640 46860 22860 46910
rect 23140 47090 23360 47140
rect 23140 47020 23150 47090
rect 23350 47020 23360 47090
rect 23140 46980 23360 47020
rect 23140 46910 23150 46980
rect 23350 46910 23360 46980
rect 23140 46860 23360 46910
rect 23640 47090 23860 47140
rect 23640 47020 23650 47090
rect 23850 47020 23860 47090
rect 23640 46980 23860 47020
rect 23640 46910 23650 46980
rect 23850 46910 23860 46980
rect 23640 46860 23860 46910
rect 24140 47090 24360 47140
rect 24140 47020 24150 47090
rect 24350 47020 24360 47090
rect 24140 46980 24360 47020
rect 24140 46910 24150 46980
rect 24350 46910 24360 46980
rect 24140 46860 24360 46910
rect 24640 47090 24860 47140
rect 24640 47020 24650 47090
rect 24850 47020 24860 47090
rect 24640 46980 24860 47020
rect 24640 46910 24650 46980
rect 24850 46910 24860 46980
rect 24640 46860 24860 46910
rect 25140 47090 25360 47140
rect 25140 47020 25150 47090
rect 25350 47020 25360 47090
rect 25140 46980 25360 47020
rect 25140 46910 25150 46980
rect 25350 46910 25360 46980
rect 25140 46860 25360 46910
rect 25640 47090 25860 47140
rect 25640 47020 25650 47090
rect 25850 47020 25860 47090
rect 25640 46980 25860 47020
rect 25640 46910 25650 46980
rect 25850 46910 25860 46980
rect 25640 46860 25860 46910
rect 26140 47090 26360 47140
rect 26140 47020 26150 47090
rect 26350 47020 26360 47090
rect 26140 46980 26360 47020
rect 26140 46910 26150 46980
rect 26350 46910 26360 46980
rect 26140 46860 26360 46910
rect 0 46850 26500 46860
rect 0 46650 20 46850
rect 90 46650 410 46850
rect 480 46650 520 46850
rect 590 46650 910 46850
rect 980 46650 1020 46850
rect 1090 46650 1410 46850
rect 1480 46650 1520 46850
rect 1590 46650 1910 46850
rect 1980 46650 2020 46850
rect 2090 46650 2410 46850
rect 2480 46650 2520 46850
rect 2590 46650 2910 46850
rect 2980 46650 3020 46850
rect 3090 46650 3410 46850
rect 3480 46650 3520 46850
rect 3590 46650 3910 46850
rect 3980 46650 4020 46850
rect 4090 46650 4410 46850
rect 4480 46650 4520 46850
rect 4590 46650 4910 46850
rect 4980 46650 5020 46850
rect 5090 46650 5410 46850
rect 5480 46650 5520 46850
rect 5590 46650 5910 46850
rect 5980 46650 6020 46850
rect 6090 46650 6410 46850
rect 6480 46650 6520 46850
rect 6590 46650 6910 46850
rect 6980 46650 7020 46850
rect 7090 46650 7410 46850
rect 7480 46650 7520 46850
rect 7590 46650 7910 46850
rect 7980 46650 8020 46850
rect 8090 46650 8410 46850
rect 8480 46650 8520 46850
rect 8590 46650 8910 46850
rect 8980 46650 9020 46850
rect 9090 46650 9410 46850
rect 9480 46650 9520 46850
rect 9590 46650 9910 46850
rect 9980 46650 10020 46850
rect 10090 46650 10410 46850
rect 10480 46650 10520 46850
rect 10590 46650 10910 46850
rect 10980 46650 11020 46850
rect 11090 46650 11410 46850
rect 11480 46650 11520 46850
rect 11590 46650 11910 46850
rect 11980 46650 12020 46850
rect 12090 46650 12410 46850
rect 12480 46650 12520 46850
rect 12590 46650 12910 46850
rect 12980 46650 13020 46850
rect 13090 46650 13410 46850
rect 13480 46650 13520 46850
rect 13590 46650 13910 46850
rect 13980 46650 14020 46850
rect 14090 46650 14410 46850
rect 14480 46650 14520 46850
rect 14590 46650 14910 46850
rect 14980 46650 15020 46850
rect 15090 46650 15410 46850
rect 15480 46650 15520 46850
rect 15590 46650 15910 46850
rect 15980 46650 16020 46850
rect 16090 46650 16410 46850
rect 16480 46650 16520 46850
rect 16590 46650 16910 46850
rect 16980 46650 17020 46850
rect 17090 46650 17410 46850
rect 17480 46650 17520 46850
rect 17590 46650 17910 46850
rect 17980 46650 18020 46850
rect 18090 46650 18410 46850
rect 18480 46650 18520 46850
rect 18590 46650 18910 46850
rect 18980 46650 19020 46850
rect 19090 46650 19410 46850
rect 19480 46650 19520 46850
rect 19590 46650 19910 46850
rect 19980 46650 20020 46850
rect 20090 46650 20410 46850
rect 20480 46650 20520 46850
rect 20590 46650 20910 46850
rect 20980 46650 21020 46850
rect 21090 46650 21410 46850
rect 21480 46650 21520 46850
rect 21590 46650 21910 46850
rect 21980 46650 22020 46850
rect 22090 46650 22410 46850
rect 22480 46650 22520 46850
rect 22590 46650 22910 46850
rect 22980 46650 23020 46850
rect 23090 46650 23410 46850
rect 23480 46650 23520 46850
rect 23590 46650 23910 46850
rect 23980 46650 24020 46850
rect 24090 46650 24410 46850
rect 24480 46650 24520 46850
rect 24590 46650 24910 46850
rect 24980 46650 25020 46850
rect 25090 46650 25410 46850
rect 25480 46650 25520 46850
rect 25590 46650 25910 46850
rect 25980 46650 26020 46850
rect 26090 46650 26410 46850
rect 26480 46650 26500 46850
rect 0 46640 26500 46650
rect 140 46590 360 46640
rect 140 46520 150 46590
rect 350 46520 360 46590
rect 140 46480 360 46520
rect 140 46410 150 46480
rect 350 46410 360 46480
rect 140 46360 360 46410
rect 640 46590 860 46640
rect 640 46520 650 46590
rect 850 46520 860 46590
rect 640 46480 860 46520
rect 1140 46590 1360 46640
rect 1140 46520 1150 46590
rect 1350 46520 1360 46590
rect 1140 46500 1360 46520
rect 1640 46590 1860 46640
rect 1640 46520 1650 46590
rect 1850 46520 1860 46590
rect 1640 46500 1860 46520
rect 2140 46590 2360 46640
rect 2140 46520 2150 46590
rect 2350 46520 2360 46590
rect 2140 46500 2360 46520
rect 2640 46590 2860 46640
rect 2640 46520 2650 46590
rect 2850 46520 2860 46590
rect 2640 46500 2860 46520
rect 3140 46590 3360 46640
rect 3140 46520 3150 46590
rect 3350 46520 3360 46590
rect 3140 46500 3360 46520
rect 3640 46590 3860 46640
rect 3640 46520 3650 46590
rect 3850 46520 3860 46590
rect 3640 46500 3860 46520
rect 4140 46590 4360 46640
rect 4140 46520 4150 46590
rect 4350 46520 4360 46590
rect 4140 46500 4360 46520
rect 4640 46590 4860 46640
rect 4640 46520 4650 46590
rect 4850 46520 4860 46590
rect 4640 46500 4860 46520
rect 5140 46590 5360 46640
rect 5140 46520 5150 46590
rect 5350 46520 5360 46590
rect 5140 46500 5360 46520
rect 5640 46590 5860 46640
rect 5640 46520 5650 46590
rect 5850 46520 5860 46590
rect 5640 46500 5860 46520
rect 6140 46590 6360 46640
rect 6140 46520 6150 46590
rect 6350 46520 6360 46590
rect 6140 46500 6360 46520
rect 6640 46590 6860 46640
rect 6640 46520 6650 46590
rect 6850 46520 6860 46590
rect 640 46410 650 46480
rect 850 46410 860 46480
rect 640 46360 860 46410
rect 6640 46480 6860 46520
rect 6640 46410 6650 46480
rect 6850 46410 6860 46480
rect 6640 46360 6860 46410
rect 7140 46590 7360 46640
rect 7140 46520 7150 46590
rect 7350 46520 7360 46590
rect 7140 46480 7360 46520
rect 7640 46590 7860 46640
rect 7640 46520 7650 46590
rect 7850 46520 7860 46590
rect 7640 46500 7860 46520
rect 8140 46590 8360 46640
rect 8140 46520 8150 46590
rect 8350 46520 8360 46590
rect 8140 46500 8360 46520
rect 8640 46590 8860 46640
rect 8640 46520 8650 46590
rect 8850 46520 8860 46590
rect 8640 46500 8860 46520
rect 9140 46590 9360 46640
rect 9140 46520 9150 46590
rect 9350 46520 9360 46590
rect 9140 46500 9360 46520
rect 9640 46590 9860 46640
rect 9640 46520 9650 46590
rect 9850 46520 9860 46590
rect 9640 46500 9860 46520
rect 10140 46590 10360 46640
rect 10140 46520 10150 46590
rect 10350 46520 10360 46590
rect 10140 46500 10360 46520
rect 10640 46590 10860 46640
rect 10640 46520 10650 46590
rect 10850 46520 10860 46590
rect 10640 46500 10860 46520
rect 11140 46590 11360 46640
rect 11140 46520 11150 46590
rect 11350 46520 11360 46590
rect 11140 46500 11360 46520
rect 11640 46590 11860 46640
rect 11640 46520 11650 46590
rect 11850 46520 11860 46590
rect 11640 46500 11860 46520
rect 12140 46590 12360 46640
rect 12140 46520 12150 46590
rect 12350 46520 12360 46590
rect 12140 46500 12360 46520
rect 12640 46590 12860 46640
rect 12640 46520 12650 46590
rect 12850 46520 12860 46590
rect 12640 46500 12860 46520
rect 13140 46590 13360 46640
rect 13140 46520 13150 46590
rect 13350 46520 13360 46590
rect 7140 46410 7150 46480
rect 7350 46410 7360 46480
rect 7140 46360 7360 46410
rect 13140 46480 13360 46520
rect 13140 46410 13150 46480
rect 13350 46410 13360 46480
rect 13140 46360 13360 46410
rect 13640 46590 13860 46640
rect 13640 46520 13650 46590
rect 13850 46520 13860 46590
rect 13640 46480 13860 46520
rect 14140 46590 14360 46640
rect 14140 46520 14150 46590
rect 14350 46520 14360 46590
rect 14140 46500 14360 46520
rect 14640 46590 14860 46640
rect 14640 46520 14650 46590
rect 14850 46520 14860 46590
rect 14640 46500 14860 46520
rect 15140 46590 15360 46640
rect 15140 46520 15150 46590
rect 15350 46520 15360 46590
rect 15140 46500 15360 46520
rect 15640 46590 15860 46640
rect 15640 46520 15650 46590
rect 15850 46520 15860 46590
rect 15640 46500 15860 46520
rect 16140 46590 16360 46640
rect 16140 46520 16150 46590
rect 16350 46520 16360 46590
rect 16140 46500 16360 46520
rect 16640 46590 16860 46640
rect 16640 46520 16650 46590
rect 16850 46520 16860 46590
rect 16640 46500 16860 46520
rect 17140 46590 17360 46640
rect 17140 46520 17150 46590
rect 17350 46520 17360 46590
rect 17140 46500 17360 46520
rect 17640 46590 17860 46640
rect 17640 46520 17650 46590
rect 17850 46520 17860 46590
rect 17640 46500 17860 46520
rect 18140 46590 18360 46640
rect 18140 46520 18150 46590
rect 18350 46520 18360 46590
rect 18140 46500 18360 46520
rect 18640 46590 18860 46640
rect 18640 46520 18650 46590
rect 18850 46520 18860 46590
rect 18640 46500 18860 46520
rect 19140 46590 19360 46640
rect 19140 46520 19150 46590
rect 19350 46520 19360 46590
rect 13640 46410 13650 46480
rect 13850 46410 13860 46480
rect 13640 46360 13860 46410
rect 19140 46480 19360 46520
rect 19140 46410 19150 46480
rect 19350 46410 19360 46480
rect 19140 46360 19360 46410
rect 19640 46590 19860 46640
rect 19640 46520 19650 46590
rect 19850 46520 19860 46590
rect 19640 46480 19860 46520
rect 20140 46590 20360 46640
rect 20140 46520 20150 46590
rect 20350 46520 20360 46590
rect 20140 46500 20360 46520
rect 20640 46590 20860 46640
rect 20640 46520 20650 46590
rect 20850 46520 20860 46590
rect 20640 46500 20860 46520
rect 21140 46590 21360 46640
rect 21140 46520 21150 46590
rect 21350 46520 21360 46590
rect 21140 46500 21360 46520
rect 21640 46590 21860 46640
rect 21640 46520 21650 46590
rect 21850 46520 21860 46590
rect 21640 46500 21860 46520
rect 22140 46590 22360 46640
rect 22140 46520 22150 46590
rect 22350 46520 22360 46590
rect 22140 46500 22360 46520
rect 22640 46590 22860 46640
rect 22640 46520 22650 46590
rect 22850 46520 22860 46590
rect 22640 46500 22860 46520
rect 23140 46590 23360 46640
rect 23140 46520 23150 46590
rect 23350 46520 23360 46590
rect 23140 46500 23360 46520
rect 23640 46590 23860 46640
rect 23640 46520 23650 46590
rect 23850 46520 23860 46590
rect 23640 46500 23860 46520
rect 24140 46590 24360 46640
rect 24140 46520 24150 46590
rect 24350 46520 24360 46590
rect 24140 46500 24360 46520
rect 24640 46590 24860 46640
rect 24640 46520 24650 46590
rect 24850 46520 24860 46590
rect 24640 46500 24860 46520
rect 25140 46590 25360 46640
rect 25140 46520 25150 46590
rect 25350 46520 25360 46590
rect 25140 46500 25360 46520
rect 25640 46590 25860 46640
rect 25640 46520 25650 46590
rect 25850 46520 25860 46590
rect 19640 46410 19650 46480
rect 19850 46410 19860 46480
rect 19640 46360 19860 46410
rect 25640 46480 25860 46520
rect 25640 46410 25650 46480
rect 25850 46410 25860 46480
rect 25640 46360 25860 46410
rect 26140 46590 26360 46640
rect 26140 46520 26150 46590
rect 26350 46520 26360 46590
rect 26140 46480 26360 46520
rect 26140 46410 26150 46480
rect 26350 46410 26360 46480
rect 26140 46360 26360 46410
rect 0 46350 1000 46360
rect 0 46150 20 46350
rect 90 46150 410 46350
rect 480 46150 520 46350
rect 590 46150 910 46350
rect 980 46150 1000 46350
rect 6500 46350 7500 46360
rect 6500 46200 6520 46350
rect 6400 46180 6520 46200
rect 0 46140 1000 46150
rect 140 46090 360 46140
rect 140 46020 150 46090
rect 350 46020 360 46090
rect 140 45980 360 46020
rect 140 45910 150 45980
rect 350 45910 360 45980
rect 140 45860 360 45910
rect 640 46090 860 46140
rect 640 46020 650 46090
rect 850 46020 860 46090
rect 640 45980 860 46020
rect 640 45910 650 45980
rect 850 45910 860 45980
rect 640 45860 860 45910
rect 1330 46120 1400 46180
rect 0 45850 1000 45860
rect 0 45650 20 45850
rect 90 45650 410 45850
rect 480 45650 520 45850
rect 590 45650 910 45850
rect 980 45650 1000 45850
rect 0 45640 1000 45650
rect 140 45590 360 45640
rect 140 45520 150 45590
rect 350 45520 360 45590
rect 140 45480 360 45520
rect 140 45410 150 45480
rect 350 45410 360 45480
rect 140 45360 360 45410
rect 640 45590 860 45640
rect 640 45520 650 45590
rect 850 45520 860 45590
rect 640 45480 860 45520
rect 640 45410 650 45480
rect 850 45410 860 45480
rect 640 45360 860 45410
rect 0 45350 1000 45360
rect 0 45150 20 45350
rect 90 45150 410 45350
rect 480 45150 520 45350
rect 590 45150 910 45350
rect 980 45150 1000 45350
rect 0 45140 1000 45150
rect 140 45090 360 45140
rect 140 45020 150 45090
rect 350 45020 360 45090
rect 140 44980 360 45020
rect 140 44910 150 44980
rect 350 44910 360 44980
rect 140 44860 360 44910
rect 640 45090 860 45140
rect 640 45020 650 45090
rect 850 45020 860 45090
rect 640 44980 860 45020
rect 640 44910 650 44980
rect 850 44910 860 44980
rect 640 44860 860 44910
rect 0 44850 1000 44860
rect 0 44650 20 44850
rect 90 44650 410 44850
rect 480 44650 520 44850
rect 590 44650 910 44850
rect 980 44650 1000 44850
rect 0 44640 1000 44650
rect 140 44590 360 44640
rect 140 44520 150 44590
rect 350 44520 360 44590
rect 140 44480 360 44520
rect 140 44410 150 44480
rect 350 44410 360 44480
rect 140 44360 360 44410
rect 640 44590 860 44640
rect 640 44520 650 44590
rect 850 44520 860 44590
rect 640 44480 860 44520
rect 640 44410 650 44480
rect 850 44410 860 44480
rect 640 44360 860 44410
rect 0 44350 1000 44360
rect 0 44150 20 44350
rect 90 44150 410 44350
rect 480 44150 520 44350
rect 590 44150 910 44350
rect 980 44150 1000 44350
rect 0 44140 1000 44150
rect 140 44090 360 44140
rect 140 44020 150 44090
rect 350 44020 360 44090
rect 140 43980 360 44020
rect 140 43910 150 43980
rect 350 43910 360 43980
rect 140 43860 360 43910
rect 640 44090 860 44140
rect 640 44020 650 44090
rect 850 44020 860 44090
rect 640 43980 860 44020
rect 640 43910 650 43980
rect 850 43910 860 43980
rect 640 43860 860 43910
rect 0 43850 1000 43860
rect 0 43650 20 43850
rect 90 43650 410 43850
rect 480 43650 520 43850
rect 590 43650 910 43850
rect 980 43650 1000 43850
rect 0 43640 1000 43650
rect 140 43590 360 43640
rect 140 43520 150 43590
rect 350 43520 360 43590
rect 140 43480 360 43520
rect 140 43410 150 43480
rect 350 43410 360 43480
rect 140 43360 360 43410
rect 640 43590 860 43640
rect 640 43520 650 43590
rect 850 43520 860 43590
rect 640 43480 860 43520
rect 640 43410 650 43480
rect 850 43410 860 43480
rect 640 43360 860 43410
rect 0 43350 1000 43360
rect 0 43150 20 43350
rect 90 43150 410 43350
rect 480 43150 520 43350
rect 590 43150 910 43350
rect 980 43150 1000 43350
rect 0 43140 1000 43150
rect 140 43090 360 43140
rect 140 43020 150 43090
rect 350 43020 360 43090
rect 140 42980 360 43020
rect 140 42910 150 42980
rect 350 42910 360 42980
rect 140 42860 360 42910
rect 640 43090 860 43140
rect 640 43020 650 43090
rect 850 43020 860 43090
rect 640 42980 860 43020
rect 640 42910 650 42980
rect 850 42910 860 42980
rect 640 42860 860 42910
rect 0 42850 1000 42860
rect 0 42650 20 42850
rect 90 42650 410 42850
rect 480 42650 520 42850
rect 590 42650 910 42850
rect 980 42650 1000 42850
rect 0 42640 1000 42650
rect 140 42590 360 42640
rect 140 42520 150 42590
rect 350 42520 360 42590
rect 140 42480 360 42520
rect 140 42410 150 42480
rect 350 42410 360 42480
rect 140 42360 360 42410
rect 640 42590 860 42640
rect 640 42520 650 42590
rect 850 42520 860 42590
rect 640 42480 860 42520
rect 640 42410 650 42480
rect 850 42410 860 42480
rect 640 42360 860 42410
rect 0 42350 1000 42360
rect 0 42150 20 42350
rect 90 42150 410 42350
rect 480 42150 520 42350
rect 590 42150 910 42350
rect 980 42150 1000 42350
rect 0 42140 1000 42150
rect 140 42090 360 42140
rect 140 42020 150 42090
rect 350 42020 360 42090
rect 140 41980 360 42020
rect 140 41910 150 41980
rect 350 41910 360 41980
rect 140 41860 360 41910
rect 640 42090 860 42140
rect 640 42020 650 42090
rect 850 42020 860 42090
rect 640 41980 860 42020
rect 640 41910 650 41980
rect 850 41910 860 41980
rect 640 41860 860 41910
rect 0 41850 1000 41860
rect 0 41650 20 41850
rect 90 41650 410 41850
rect 480 41650 520 41850
rect 590 41650 910 41850
rect 980 41650 1000 41850
rect 0 41640 1000 41650
rect 140 41590 360 41640
rect 140 41520 150 41590
rect 350 41520 360 41590
rect 140 41480 360 41520
rect 140 41410 150 41480
rect 350 41410 360 41480
rect 140 41360 360 41410
rect 640 41590 860 41640
rect 640 41520 650 41590
rect 850 41520 860 41590
rect 640 41480 860 41520
rect 640 41410 650 41480
rect 850 41410 860 41480
rect 640 41360 860 41410
rect 0 41350 1000 41360
rect 0 41150 20 41350
rect 90 41150 410 41350
rect 480 41150 520 41350
rect 590 41150 910 41350
rect 980 41150 1000 41350
rect 0 41140 1000 41150
rect 140 41090 360 41140
rect 140 41020 150 41090
rect 350 41020 360 41090
rect 140 40980 360 41020
rect 140 40910 150 40980
rect 350 40910 360 40980
rect 140 40860 360 40910
rect 640 41090 860 41140
rect 640 41020 650 41090
rect 850 41020 860 41090
rect 640 40980 860 41020
rect 640 40910 650 40980
rect 850 40910 860 40980
rect 640 40860 860 40910
rect 0 40850 1000 40860
rect 0 40650 20 40850
rect 90 40650 410 40850
rect 480 40650 520 40850
rect 590 40650 910 40850
rect 980 40650 1000 40850
rect 0 40640 1000 40650
rect 140 40590 360 40640
rect 140 40520 150 40590
rect 350 40520 360 40590
rect 140 40480 360 40520
rect -3300 40450 -3100 40460
rect -3300 40190 -3290 40450
rect -3110 40190 -3100 40450
rect 140 40410 150 40480
rect 350 40410 360 40480
rect 140 40360 360 40410
rect 640 40590 860 40640
rect 640 40520 650 40590
rect 850 40520 860 40590
rect 640 40480 860 40520
rect 640 40410 650 40480
rect 850 40410 860 40480
rect 640 40360 860 40410
rect -3300 40180 -3100 40190
rect 0 40350 1000 40360
rect 0 40150 20 40350
rect 90 40150 410 40350
rect 480 40150 520 40350
rect 590 40150 910 40350
rect 980 40150 1000 40350
rect 0 40140 1000 40150
rect 140 40090 360 40140
rect 140 40020 150 40090
rect 350 40020 360 40090
rect -2860 39980 -2640 40000
rect -2860 39910 -2850 39980
rect -2650 39910 -2640 39980
rect -2860 39860 -2640 39910
rect -2360 39980 -2140 40000
rect -2360 39910 -2350 39980
rect -2150 39910 -2140 39980
rect -2360 39860 -2140 39910
rect -1860 39980 -1640 40000
rect -1860 39910 -1850 39980
rect -1650 39910 -1640 39980
rect -1860 39860 -1640 39910
rect -1360 39980 -1140 40000
rect -1360 39910 -1350 39980
rect -1150 39910 -1140 39980
rect -1360 39860 -1140 39910
rect -860 39980 -640 40000
rect -860 39910 -850 39980
rect -650 39910 -640 39980
rect -860 39860 -640 39910
rect -360 39980 -140 40000
rect -360 39910 -350 39980
rect -150 39910 -140 39980
rect -360 39860 -140 39910
rect 140 39980 360 40020
rect 140 39910 150 39980
rect 350 39910 360 39980
rect 140 39860 360 39910
rect 640 40090 860 40140
rect 640 40020 650 40090
rect 850 40020 860 40090
rect 640 39980 860 40020
rect 640 39910 650 39980
rect 850 39910 860 39980
rect 640 39860 860 39910
rect -3000 39850 1000 39860
rect -3000 39650 -2980 39850
rect -2910 39650 -2590 39850
rect -2520 39650 -2480 39850
rect -2410 39650 -2090 39850
rect -2020 39650 -1980 39850
rect -1910 39650 -1590 39850
rect -1520 39650 -1480 39850
rect -1410 39650 -1090 39850
rect -1020 39650 -980 39850
rect -910 39650 -590 39850
rect -520 39650 -480 39850
rect -410 39650 -90 39850
rect -20 39650 20 39850
rect 90 39650 410 39850
rect 480 39650 520 39850
rect 590 39650 910 39850
rect 980 39650 1000 39850
rect 6340 46150 6520 46180
rect 6590 46150 6910 46350
rect 6980 46150 7020 46350
rect 7090 46150 7410 46350
rect 7480 46200 7500 46350
rect 13000 46350 14000 46360
rect 13000 46300 13020 46350
rect 7480 46150 7700 46200
rect 12700 46180 13020 46300
rect 6340 46120 7700 46150
rect 1532 46080 1552 46090
rect 6186 46080 6206 46090
rect 1532 46010 1540 46080
rect 6200 46010 6206 46080
rect 1532 45990 1552 46010
rect 6186 45990 6206 46010
rect 1465 45938 1531 45958
rect 1465 39958 1531 39978
rect 1623 45938 1689 45958
rect 1623 39958 1689 39978
rect 1781 45938 1847 45958
rect 1781 39958 1847 39978
rect 1939 45938 2005 45958
rect 1939 39958 2005 39978
rect 2097 45938 2163 45958
rect 2097 39958 2163 39978
rect 2255 45938 2321 45958
rect 2255 39958 2321 39978
rect 2413 45938 2479 45958
rect 2413 39958 2479 39978
rect 2571 45938 2637 45958
rect 2571 39958 2637 39978
rect 2729 45938 2795 45958
rect 2729 39958 2795 39978
rect 2887 45938 2953 45958
rect 2887 39958 2953 39978
rect 3045 45938 3111 45958
rect 3045 39958 3111 39978
rect 3203 45938 3269 45958
rect 3203 39958 3269 39978
rect 3361 45938 3427 45958
rect 3361 39958 3427 39978
rect 3519 45938 3585 45958
rect 3519 39958 3585 39978
rect 3677 45938 3743 45958
rect 3677 39958 3743 39978
rect 3835 45938 3901 45958
rect 3835 39958 3901 39978
rect 3993 45938 4059 45958
rect 3993 39958 4059 39978
rect 4151 45938 4217 45958
rect 4151 39958 4217 39978
rect 4309 45938 4375 45958
rect 4309 39958 4375 39978
rect 4467 45938 4533 45958
rect 4467 39958 4533 39978
rect 4625 45938 4691 45958
rect 4625 39958 4691 39978
rect 4783 45938 4849 45958
rect 4783 39958 4849 39978
rect 4941 45938 5007 45958
rect 4941 39958 5007 39978
rect 5099 45938 5165 45958
rect 5099 39958 5165 39978
rect 5257 45938 5323 45958
rect 5257 39958 5323 39978
rect 5415 45938 5481 45958
rect 5415 39958 5481 39978
rect 5573 45938 5639 45958
rect 5573 39958 5639 39978
rect 5731 45938 5797 45958
rect 5731 39958 5797 39978
rect 5889 45938 5955 45958
rect 5889 39958 5955 39978
rect 6047 45938 6113 45958
rect 6047 39958 6113 39978
rect 6205 45938 6271 45958
rect 6205 39958 6271 39978
rect 1532 39910 1552 39926
rect 6186 39910 6206 39926
rect 1532 39840 1540 39910
rect 6190 39840 6206 39910
rect 1532 39826 1552 39840
rect 6186 39826 6206 39840
rect 1330 39730 1400 39800
rect 6410 46090 7630 46120
rect 6410 46020 6650 46090
rect 6850 46020 7150 46090
rect 7350 46020 7630 46090
rect 6410 45800 7630 46020
rect 6410 45200 7630 45600
rect 6410 44600 7630 45000
rect 6410 44000 7630 44400
rect 6410 43400 7630 43800
rect 6410 42800 7630 43200
rect 6410 42200 7630 42600
rect 6410 41600 7630 42000
rect 6410 41000 7630 41400
rect 6410 40400 7630 40800
rect 6410 39800 7630 40200
rect 12640 46150 13020 46180
rect 13090 46150 13410 46350
rect 13480 46150 13520 46350
rect 13590 46150 13910 46350
rect 13980 46150 14000 46350
rect 19000 46350 20000 46360
rect 19000 46180 19020 46350
rect 12640 46120 14000 46150
rect 7832 46080 7852 46090
rect 12486 46080 12506 46090
rect 7832 46010 7840 46080
rect 12500 46010 12506 46080
rect 7832 45990 7852 46010
rect 12486 45990 12506 46010
rect 7765 45938 7831 45958
rect 7765 39958 7831 39978
rect 7923 45938 7989 45958
rect 7923 39958 7989 39978
rect 8081 45938 8147 45958
rect 8081 39958 8147 39978
rect 8239 45938 8305 45958
rect 8239 39958 8305 39978
rect 8397 45938 8463 45958
rect 8397 39958 8463 39978
rect 8555 45938 8621 45958
rect 8555 39958 8621 39978
rect 8713 45938 8779 45958
rect 8713 39958 8779 39978
rect 8871 45938 8937 45958
rect 8871 39958 8937 39978
rect 9029 45938 9095 45958
rect 9029 39958 9095 39978
rect 9187 45938 9253 45958
rect 9187 39958 9253 39978
rect 9345 45938 9411 45958
rect 9345 39958 9411 39978
rect 9503 45938 9569 45958
rect 9503 39958 9569 39978
rect 9661 45938 9727 45958
rect 9661 39958 9727 39978
rect 9819 45938 9885 45958
rect 9819 39958 9885 39978
rect 9977 45938 10043 45958
rect 9977 39958 10043 39978
rect 10135 45938 10201 45958
rect 10135 39958 10201 39978
rect 10293 45938 10359 45958
rect 10293 39958 10359 39978
rect 10451 45938 10517 45958
rect 10451 39958 10517 39978
rect 10609 45938 10675 45958
rect 10609 39958 10675 39978
rect 10767 45938 10833 45958
rect 10767 39958 10833 39978
rect 10925 45938 10991 45958
rect 10925 39958 10991 39978
rect 11083 45938 11149 45958
rect 11083 39958 11149 39978
rect 11241 45938 11307 45958
rect 11241 39958 11307 39978
rect 11399 45938 11465 45958
rect 11399 39958 11465 39978
rect 11557 45938 11623 45958
rect 11557 39958 11623 39978
rect 11715 45938 11781 45958
rect 11715 39958 11781 39978
rect 11873 45938 11939 45958
rect 11873 39958 11939 39978
rect 12031 45938 12097 45958
rect 12031 39958 12097 39978
rect 12189 45938 12255 45958
rect 12189 39958 12255 39978
rect 12347 45938 12413 45958
rect 12347 39958 12413 39978
rect 12505 45938 12571 45958
rect 12505 39958 12571 39978
rect 7832 39910 7852 39926
rect 12486 39910 12506 39926
rect 7832 39840 7840 39910
rect 12490 39840 12506 39910
rect 7832 39826 7852 39840
rect 12486 39826 12506 39840
rect 6340 39730 6410 39800
rect -3000 39640 1000 39650
rect -2860 39590 -2640 39640
rect -2860 39520 -2850 39590
rect -2650 39520 -2640 39590
rect -2860 39480 -2640 39520
rect -2860 39410 -2850 39480
rect -2650 39410 -2640 39480
rect -2860 39360 -2640 39410
rect -2360 39590 -2140 39640
rect -2360 39520 -2350 39590
rect -2150 39520 -2140 39590
rect -2360 39480 -2140 39520
rect -2360 39410 -2350 39480
rect -2150 39410 -2140 39480
rect -2360 39360 -2140 39410
rect -1860 39590 -1640 39640
rect -1860 39520 -1850 39590
rect -1650 39520 -1640 39590
rect -1860 39480 -1640 39520
rect -1860 39410 -1850 39480
rect -1650 39410 -1640 39480
rect -1860 39360 -1640 39410
rect -1360 39590 -1140 39640
rect -1360 39520 -1350 39590
rect -1150 39520 -1140 39590
rect -1360 39480 -1140 39520
rect -1360 39410 -1350 39480
rect -1150 39410 -1140 39480
rect -1360 39360 -1140 39410
rect -860 39590 -640 39640
rect -860 39520 -850 39590
rect -650 39520 -640 39590
rect -860 39480 -640 39520
rect -860 39410 -850 39480
rect -650 39410 -640 39480
rect -860 39360 -640 39410
rect -360 39590 -140 39640
rect -360 39520 -350 39590
rect -150 39520 -140 39590
rect -360 39480 -140 39520
rect -360 39410 -350 39480
rect -150 39410 -140 39480
rect -360 39360 -140 39410
rect 140 39590 360 39640
rect 140 39520 150 39590
rect 350 39520 360 39590
rect 140 39480 360 39520
rect 140 39410 150 39480
rect 350 39410 360 39480
rect 140 39360 360 39410
rect 640 39590 860 39640
rect 640 39520 650 39590
rect 850 39520 860 39590
rect 640 39480 860 39520
rect 640 39410 650 39480
rect 850 39410 860 39480
rect 640 39360 860 39410
rect -3000 39350 1000 39360
rect -3000 39150 -2980 39350
rect -2910 39150 -2590 39350
rect -2520 39150 -2480 39350
rect -2410 39150 -2090 39350
rect -2020 39150 -1980 39350
rect -1910 39150 -1590 39350
rect -1520 39150 -1480 39350
rect -1410 39150 -1090 39350
rect -1020 39150 -980 39350
rect -910 39150 -590 39350
rect -520 39150 -480 39350
rect -410 39150 -90 39350
rect -20 39150 20 39350
rect 90 39150 410 39350
rect 480 39150 520 39350
rect 590 39150 910 39350
rect 980 39150 1000 39350
rect 6800 39200 7300 39800
rect 7630 39730 7700 39800
rect 12710 46090 13930 46120
rect 12710 46020 13150 46090
rect 13350 46020 13650 46090
rect 13850 46020 13930 46090
rect 12710 45900 13930 46020
rect 12710 45300 13930 45700
rect 12710 44700 13930 45100
rect 12710 44100 13930 44500
rect 12710 43500 13930 43900
rect 12710 42900 13930 43300
rect 12710 42300 13930 42700
rect 12710 41700 13930 42100
rect 12710 41100 13930 41500
rect 12710 40500 13930 40900
rect 12710 39900 13930 40300
rect 12640 39730 12710 39800
rect 13100 39200 13600 39900
rect 18940 46150 19020 46180
rect 19090 46150 19410 46350
rect 19480 46150 19520 46350
rect 19590 46150 19910 46350
rect 19980 46200 20000 46350
rect 25500 46350 26500 46360
rect 19980 46150 20300 46200
rect 18940 46120 20300 46150
rect 14132 46080 14152 46090
rect 18786 46080 18806 46090
rect 14132 46010 14140 46080
rect 18800 46010 18806 46080
rect 14132 45990 14152 46010
rect 18786 45990 18806 46010
rect 14065 45938 14131 45958
rect 14065 39958 14131 39978
rect 14223 45938 14289 45958
rect 14223 39958 14289 39978
rect 14381 45938 14447 45958
rect 14381 39958 14447 39978
rect 14539 45938 14605 45958
rect 14539 39958 14605 39978
rect 14697 45938 14763 45958
rect 14697 39958 14763 39978
rect 14855 45938 14921 45958
rect 14855 39958 14921 39978
rect 15013 45938 15079 45958
rect 15013 39958 15079 39978
rect 15171 45938 15237 45958
rect 15171 39958 15237 39978
rect 15329 45938 15395 45958
rect 15329 39958 15395 39978
rect 15487 45938 15553 45958
rect 15487 39958 15553 39978
rect 15645 45938 15711 45958
rect 15645 39958 15711 39978
rect 15803 45938 15869 45958
rect 15803 39958 15869 39978
rect 15961 45938 16027 45958
rect 15961 39958 16027 39978
rect 16119 45938 16185 45958
rect 16119 39958 16185 39978
rect 16277 45938 16343 45958
rect 16277 39958 16343 39978
rect 16435 45938 16501 45958
rect 16435 39958 16501 39978
rect 16593 45938 16659 45958
rect 16593 39958 16659 39978
rect 16751 45938 16817 45958
rect 16751 39958 16817 39978
rect 16909 45938 16975 45958
rect 16909 39958 16975 39978
rect 17067 45938 17133 45958
rect 17067 39958 17133 39978
rect 17225 45938 17291 45958
rect 17225 39958 17291 39978
rect 17383 45938 17449 45958
rect 17383 39958 17449 39978
rect 17541 45938 17607 45958
rect 17541 39958 17607 39978
rect 17699 45938 17765 45958
rect 17699 39958 17765 39978
rect 17857 45938 17923 45958
rect 17857 39958 17923 39978
rect 18015 45938 18081 45958
rect 18015 39958 18081 39978
rect 18173 45938 18239 45958
rect 18173 39958 18239 39978
rect 18331 45938 18397 45958
rect 18331 39958 18397 39978
rect 18489 45938 18555 45958
rect 18489 39958 18555 39978
rect 18647 45938 18713 45958
rect 18647 39958 18713 39978
rect 18805 45938 18871 45958
rect 18805 39958 18871 39978
rect 14132 39910 14152 39926
rect 18786 39910 18806 39926
rect 14132 39840 14140 39910
rect 18790 39840 18806 39910
rect 14132 39826 14152 39840
rect 18786 39826 18806 39840
rect 13930 39730 14000 39800
rect 19010 46090 20230 46120
rect 19010 46020 19150 46090
rect 19350 46020 19650 46090
rect 19850 46020 20230 46090
rect 19010 45800 20230 46020
rect 19010 45200 20230 45600
rect 19010 44600 20230 45000
rect 19010 44000 20230 44400
rect 19010 43400 20230 43800
rect 19010 42800 20230 43200
rect 19010 42200 20230 42600
rect 19010 41600 20230 42000
rect 19010 41000 20230 41400
rect 19010 40400 20230 40800
rect 19010 39800 20230 40200
rect 25240 46120 25310 46180
rect 25500 46150 25520 46350
rect 25590 46150 25910 46350
rect 25980 46150 26020 46350
rect 26090 46150 26410 46350
rect 26480 46150 26500 46350
rect 25500 46140 26500 46150
rect 20432 46080 20452 46090
rect 25086 46080 25106 46090
rect 20432 46010 20440 46080
rect 25100 46010 25106 46080
rect 20432 45990 20452 46010
rect 25086 45990 25106 46010
rect 20365 45938 20431 45958
rect 20365 39958 20431 39978
rect 20523 45938 20589 45958
rect 20523 39958 20589 39978
rect 20681 45938 20747 45958
rect 20681 39958 20747 39978
rect 20839 45938 20905 45958
rect 20839 39958 20905 39978
rect 20997 45938 21063 45958
rect 20997 39958 21063 39978
rect 21155 45938 21221 45958
rect 21155 39958 21221 39978
rect 21313 45938 21379 45958
rect 21313 39958 21379 39978
rect 21471 45938 21537 45958
rect 21471 39958 21537 39978
rect 21629 45938 21695 45958
rect 21629 39958 21695 39978
rect 21787 45938 21853 45958
rect 21787 39958 21853 39978
rect 21945 45938 22011 45958
rect 21945 39958 22011 39978
rect 22103 45938 22169 45958
rect 22103 39958 22169 39978
rect 22261 45938 22327 45958
rect 22261 39958 22327 39978
rect 22419 45938 22485 45958
rect 22419 39958 22485 39978
rect 22577 45938 22643 45958
rect 22577 39958 22643 39978
rect 22735 45938 22801 45958
rect 22735 39958 22801 39978
rect 22893 45938 22959 45958
rect 22893 39958 22959 39978
rect 23051 45938 23117 45958
rect 23051 39958 23117 39978
rect 23209 45938 23275 45958
rect 23209 39958 23275 39978
rect 23367 45938 23433 45958
rect 23367 39958 23433 39978
rect 23525 45938 23591 45958
rect 23525 39958 23591 39978
rect 23683 45938 23749 45958
rect 23683 39958 23749 39978
rect 23841 45938 23907 45958
rect 23841 39958 23907 39978
rect 23999 45938 24065 45958
rect 23999 39958 24065 39978
rect 24157 45938 24223 45958
rect 24157 39958 24223 39978
rect 24315 45938 24381 45958
rect 24315 39958 24381 39978
rect 24473 45938 24539 45958
rect 24473 39958 24539 39978
rect 24631 45938 24697 45958
rect 24631 39958 24697 39978
rect 24789 45938 24855 45958
rect 24789 39958 24855 39978
rect 24947 45938 25013 45958
rect 24947 39958 25013 39978
rect 25105 45938 25171 45958
rect 25105 39958 25171 39978
rect 20432 39910 20452 39926
rect 25086 39910 25106 39926
rect 20432 39840 20440 39910
rect 25090 39840 25106 39910
rect 20432 39826 20452 39840
rect 25086 39826 25106 39840
rect 18940 39730 19010 39800
rect 19400 39200 19900 39800
rect 20230 39730 20300 39800
rect 25640 46090 25860 46140
rect 25640 46020 25650 46090
rect 25850 46020 25860 46090
rect 25640 45980 25860 46020
rect 25640 45910 25650 45980
rect 25850 45910 25860 45980
rect 25640 45860 25860 45910
rect 26140 46090 26360 46140
rect 26140 46020 26150 46090
rect 26350 46020 26360 46090
rect 26140 45980 26360 46020
rect 26140 45910 26150 45980
rect 26350 45910 26360 45980
rect 26140 45860 26360 45910
rect 25500 45850 26500 45860
rect 25500 45650 25520 45850
rect 25590 45650 25910 45850
rect 25980 45650 26020 45850
rect 26090 45650 26410 45850
rect 26480 45650 26500 45850
rect 25500 45640 26500 45650
rect 25640 45590 25860 45640
rect 25640 45520 25650 45590
rect 25850 45520 25860 45590
rect 25640 45480 25860 45520
rect 25640 45410 25650 45480
rect 25850 45410 25860 45480
rect 25640 45360 25860 45410
rect 26140 45590 26360 45640
rect 26140 45520 26150 45590
rect 26350 45520 26360 45590
rect 26140 45480 26360 45520
rect 26140 45410 26150 45480
rect 26350 45410 26360 45480
rect 26140 45360 26360 45410
rect 25500 45350 26500 45360
rect 25500 45150 25520 45350
rect 25590 45150 25910 45350
rect 25980 45150 26020 45350
rect 26090 45150 26410 45350
rect 26480 45150 26500 45350
rect 25500 45140 26500 45150
rect 25640 45090 25860 45140
rect 25640 45020 25650 45090
rect 25850 45020 25860 45090
rect 25640 44980 25860 45020
rect 25640 44910 25650 44980
rect 25850 44910 25860 44980
rect 25640 44860 25860 44910
rect 26140 45090 26360 45140
rect 26140 45020 26150 45090
rect 26350 45020 26360 45090
rect 26140 44980 26360 45020
rect 26140 44910 26150 44980
rect 26350 44910 26360 44980
rect 26140 44860 26360 44910
rect 25500 44850 26500 44860
rect 25500 44650 25520 44850
rect 25590 44650 25910 44850
rect 25980 44650 26020 44850
rect 26090 44650 26410 44850
rect 26480 44650 26500 44850
rect 25500 44640 26500 44650
rect 25640 44590 25860 44640
rect 25640 44520 25650 44590
rect 25850 44520 25860 44590
rect 25640 44480 25860 44520
rect 25640 44410 25650 44480
rect 25850 44410 25860 44480
rect 25640 44360 25860 44410
rect 26140 44590 26360 44640
rect 26140 44520 26150 44590
rect 26350 44520 26360 44590
rect 26140 44480 26360 44520
rect 26140 44410 26150 44480
rect 26350 44410 26360 44480
rect 26140 44360 26360 44410
rect 25500 44350 26500 44360
rect 25500 44150 25520 44350
rect 25590 44150 25910 44350
rect 25980 44150 26020 44350
rect 26090 44150 26410 44350
rect 26480 44150 26500 44350
rect 25500 44140 26500 44150
rect 25640 44090 25860 44140
rect 25640 44020 25650 44090
rect 25850 44020 25860 44090
rect 25640 43980 25860 44020
rect 25640 43910 25650 43980
rect 25850 43910 25860 43980
rect 25640 43860 25860 43910
rect 26140 44090 26360 44140
rect 26140 44020 26150 44090
rect 26350 44020 26360 44090
rect 26140 43980 26360 44020
rect 26140 43910 26150 43980
rect 26350 43910 26360 43980
rect 26140 43860 26360 43910
rect 25500 43850 26500 43860
rect 25500 43650 25520 43850
rect 25590 43650 25910 43850
rect 25980 43650 26020 43850
rect 26090 43650 26410 43850
rect 26480 43650 26500 43850
rect 25500 43640 26500 43650
rect 25640 43590 25860 43640
rect 25640 43520 25650 43590
rect 25850 43520 25860 43590
rect 25640 43480 25860 43520
rect 25640 43410 25650 43480
rect 25850 43410 25860 43480
rect 25640 43360 25860 43410
rect 26140 43590 26360 43640
rect 26140 43520 26150 43590
rect 26350 43520 26360 43590
rect 26140 43480 26360 43520
rect 26140 43410 26150 43480
rect 26350 43410 26360 43480
rect 26140 43360 26360 43410
rect 25500 43350 26500 43360
rect 25500 43150 25520 43350
rect 25590 43150 25910 43350
rect 25980 43150 26020 43350
rect 26090 43150 26410 43350
rect 26480 43150 26500 43350
rect 25500 43140 26500 43150
rect 25640 43090 25860 43140
rect 25640 43020 25650 43090
rect 25850 43020 25860 43090
rect 25640 42980 25860 43020
rect 25640 42910 25650 42980
rect 25850 42910 25860 42980
rect 25640 42860 25860 42910
rect 26140 43090 26360 43140
rect 26140 43020 26150 43090
rect 26350 43020 26360 43090
rect 26140 42980 26360 43020
rect 26140 42910 26150 42980
rect 26350 42910 26360 42980
rect 26140 42860 26360 42910
rect 25500 42850 26500 42860
rect 25500 42650 25520 42850
rect 25590 42650 25910 42850
rect 25980 42650 26020 42850
rect 26090 42650 26410 42850
rect 26480 42650 26500 42850
rect 25500 42640 26500 42650
rect 25640 42590 25860 42640
rect 25640 42520 25650 42590
rect 25850 42520 25860 42590
rect 25640 42480 25860 42520
rect 25640 42410 25650 42480
rect 25850 42410 25860 42480
rect 25640 42360 25860 42410
rect 26140 42590 26360 42640
rect 26140 42520 26150 42590
rect 26350 42520 26360 42590
rect 26140 42480 26360 42520
rect 26140 42410 26150 42480
rect 26350 42410 26360 42480
rect 26140 42360 26360 42410
rect 25500 42350 26500 42360
rect 25500 42150 25520 42350
rect 25590 42150 25910 42350
rect 25980 42150 26020 42350
rect 26090 42150 26410 42350
rect 26480 42150 26500 42350
rect 25500 42140 26500 42150
rect 25640 42090 25860 42140
rect 25640 42020 25650 42090
rect 25850 42020 25860 42090
rect 25640 41980 25860 42020
rect 25640 41910 25650 41980
rect 25850 41910 25860 41980
rect 25640 41860 25860 41910
rect 26140 42090 26360 42140
rect 26140 42020 26150 42090
rect 26350 42020 26360 42090
rect 26140 41980 26360 42020
rect 26140 41910 26150 41980
rect 26350 41910 26360 41980
rect 26140 41860 26360 41910
rect 25500 41850 26500 41860
rect 25500 41650 25520 41850
rect 25590 41650 25910 41850
rect 25980 41650 26020 41850
rect 26090 41650 26410 41850
rect 26480 41650 26500 41850
rect 25500 41640 26500 41650
rect 25640 41590 25860 41640
rect 25640 41520 25650 41590
rect 25850 41520 25860 41590
rect 25640 41480 25860 41520
rect 25640 41410 25650 41480
rect 25850 41410 25860 41480
rect 25640 41360 25860 41410
rect 26140 41590 26360 41640
rect 26140 41520 26150 41590
rect 26350 41520 26360 41590
rect 26140 41480 26360 41520
rect 26140 41410 26150 41480
rect 26350 41410 26360 41480
rect 26140 41360 26360 41410
rect 25500 41350 26500 41360
rect 25500 41150 25520 41350
rect 25590 41150 25910 41350
rect 25980 41150 26020 41350
rect 26090 41150 26410 41350
rect 26480 41150 26500 41350
rect 25500 41140 26500 41150
rect 25640 41090 25860 41140
rect 25640 41020 25650 41090
rect 25850 41020 25860 41090
rect 25640 40980 25860 41020
rect 25640 40910 25650 40980
rect 25850 40910 25860 40980
rect 25640 40860 25860 40910
rect 26140 41090 26360 41140
rect 26140 41020 26150 41090
rect 26350 41020 26360 41090
rect 26140 40980 26360 41020
rect 26140 40910 26150 40980
rect 26350 40910 26360 40980
rect 26140 40860 26360 40910
rect 25500 40850 26500 40860
rect 25500 40650 25520 40850
rect 25590 40650 25910 40850
rect 25980 40650 26020 40850
rect 26090 40650 26410 40850
rect 26480 40650 26500 40850
rect 25500 40640 26500 40650
rect 25640 40590 25860 40640
rect 25640 40520 25650 40590
rect 25850 40520 25860 40590
rect 25640 40480 25860 40520
rect 25640 40410 25650 40480
rect 25850 40410 25860 40480
rect 25640 40360 25860 40410
rect 26140 40590 26360 40640
rect 26140 40520 26150 40590
rect 26350 40520 26360 40590
rect 26140 40480 26360 40520
rect 26140 40410 26150 40480
rect 26350 40410 26360 40480
rect 26140 40360 26360 40410
rect 29900 40450 30100 40460
rect 25500 40350 26500 40360
rect 25500 40150 25520 40350
rect 25590 40150 25910 40350
rect 25980 40150 26020 40350
rect 26090 40150 26410 40350
rect 26480 40150 26500 40350
rect 29900 40190 29910 40450
rect 30090 40190 30100 40450
rect 29900 40180 30100 40190
rect 25500 40140 26500 40150
rect 25640 40090 25860 40140
rect 25640 40020 25650 40090
rect 25850 40020 25860 40090
rect 25640 39980 25860 40020
rect 25640 39910 25650 39980
rect 25850 39910 25860 39980
rect 25640 39860 25860 39910
rect 26140 40090 26360 40140
rect 26140 40020 26150 40090
rect 26350 40020 26360 40090
rect 26140 39980 26360 40020
rect 26140 39910 26150 39980
rect 26350 39910 26360 39980
rect 26140 39860 26360 39910
rect 26640 39980 26860 40000
rect 26640 39910 26650 39980
rect 26850 39910 26860 39980
rect 26640 39860 26860 39910
rect 27140 39980 27360 40000
rect 27140 39910 27150 39980
rect 27350 39910 27360 39980
rect 27140 39860 27360 39910
rect 27640 39980 27860 40000
rect 27640 39910 27650 39980
rect 27850 39910 27860 39980
rect 27640 39860 27860 39910
rect 28140 39980 28360 40000
rect 28140 39910 28150 39980
rect 28350 39910 28360 39980
rect 28140 39860 28360 39910
rect 28640 39980 28860 40000
rect 28640 39910 28650 39980
rect 28850 39910 28860 39980
rect 28640 39860 28860 39910
rect 29140 39980 29360 40000
rect 29140 39910 29150 39980
rect 29350 39910 29360 39980
rect 29140 39860 29360 39910
rect 25240 39730 25310 39800
rect 25500 39850 29500 39860
rect 25500 39650 25520 39850
rect 25590 39650 25910 39850
rect 25980 39650 26020 39850
rect 26090 39650 26410 39850
rect 26480 39650 26520 39850
rect 26590 39650 26910 39850
rect 26980 39650 27020 39850
rect 27090 39650 27410 39850
rect 27480 39650 27520 39850
rect 27590 39650 27910 39850
rect 27980 39650 28020 39850
rect 28090 39650 28410 39850
rect 28480 39650 28520 39850
rect 28590 39650 28910 39850
rect 28980 39650 29020 39850
rect 29090 39650 29410 39850
rect 29480 39650 29500 39850
rect 25500 39640 29500 39650
rect 25640 39590 25860 39640
rect 25640 39520 25650 39590
rect 25850 39520 25860 39590
rect 25640 39480 25860 39520
rect 25640 39410 25650 39480
rect 25850 39410 25860 39480
rect 25640 39360 25860 39410
rect 26140 39590 26360 39640
rect 26140 39520 26150 39590
rect 26350 39520 26360 39590
rect 26140 39480 26360 39520
rect 26140 39410 26150 39480
rect 26350 39410 26360 39480
rect 26140 39360 26360 39410
rect 26640 39590 26860 39640
rect 26640 39520 26650 39590
rect 26850 39520 26860 39590
rect 26640 39480 26860 39520
rect 26640 39410 26650 39480
rect 26850 39410 26860 39480
rect 26640 39360 26860 39410
rect 27140 39590 27360 39640
rect 27140 39520 27150 39590
rect 27350 39520 27360 39590
rect 27140 39480 27360 39520
rect 27140 39410 27150 39480
rect 27350 39410 27360 39480
rect 27140 39360 27360 39410
rect 27640 39590 27860 39640
rect 27640 39520 27650 39590
rect 27850 39520 27860 39590
rect 27640 39480 27860 39520
rect 27640 39410 27650 39480
rect 27850 39410 27860 39480
rect 27640 39360 27860 39410
rect 28140 39590 28360 39640
rect 28140 39520 28150 39590
rect 28350 39520 28360 39590
rect 28140 39480 28360 39520
rect 28140 39410 28150 39480
rect 28350 39410 28360 39480
rect 28140 39360 28360 39410
rect 28640 39590 28860 39640
rect 28640 39520 28650 39590
rect 28850 39520 28860 39590
rect 28640 39480 28860 39520
rect 28640 39410 28650 39480
rect 28850 39410 28860 39480
rect 28640 39360 28860 39410
rect 29140 39590 29360 39640
rect 29140 39520 29150 39590
rect 29350 39520 29360 39590
rect 29140 39480 29360 39520
rect 29140 39410 29150 39480
rect 29350 39410 29360 39480
rect 29140 39360 29360 39410
rect 25500 39350 29500 39360
rect 6400 39180 7700 39200
rect 12700 39180 14000 39200
rect 19000 39180 20300 39200
rect -3000 39140 1000 39150
rect -2860 39090 -2640 39140
rect -2860 39020 -2850 39090
rect -2650 39020 -2640 39090
rect -2860 39000 -2640 39020
rect -2360 39090 -2140 39140
rect -2360 39020 -2350 39090
rect -2150 39020 -2140 39090
rect -2360 39000 -2140 39020
rect -1860 39090 -1640 39140
rect -1860 39020 -1850 39090
rect -1650 39020 -1640 39090
rect -1860 39000 -1640 39020
rect -1360 39090 -1140 39140
rect -1360 39020 -1350 39090
rect -1150 39020 -1140 39090
rect -1360 39000 -1140 39020
rect -860 39090 -640 39140
rect -860 39020 -850 39090
rect -650 39020 -640 39090
rect -860 39000 -640 39020
rect -360 39090 -140 39140
rect -360 39020 -350 39090
rect -150 39020 -140 39090
rect -360 39000 -140 39020
rect 140 39090 360 39140
rect 140 39020 150 39090
rect 350 39020 360 39090
rect 140 38980 360 39020
rect -3300 38910 -3100 38920
rect -3300 38690 -3290 38910
rect -3110 38690 -3100 38910
rect 140 38910 150 38980
rect 350 38910 360 38980
rect 140 38860 360 38910
rect 640 39090 860 39140
rect 640 39020 650 39090
rect 850 39020 860 39090
rect 640 38980 860 39020
rect 640 38910 650 38980
rect 850 38910 860 38980
rect 640 38860 860 38910
rect 1330 39120 1400 39180
rect -3300 38680 -3100 38690
rect 0 38850 1000 38860
rect 0 38650 20 38850
rect 90 38650 410 38850
rect 480 38650 520 38850
rect 590 38650 910 38850
rect 980 38650 1000 38850
rect 0 38640 1000 38650
rect 140 38590 360 38640
rect 140 38520 150 38590
rect 350 38520 360 38590
rect 140 38480 360 38520
rect 140 38410 150 38480
rect 350 38410 360 38480
rect 140 38360 360 38410
rect 640 38590 860 38640
rect 640 38520 650 38590
rect 850 38520 860 38590
rect 640 38480 860 38520
rect 640 38410 650 38480
rect 850 38410 860 38480
rect 640 38360 860 38410
rect 0 38350 1000 38360
rect 0 38150 20 38350
rect 90 38150 410 38350
rect 480 38150 520 38350
rect 590 38150 910 38350
rect 980 38150 1000 38350
rect 0 38140 1000 38150
rect 140 38090 360 38140
rect 140 38020 150 38090
rect 350 38020 360 38090
rect 140 37980 360 38020
rect 140 37910 150 37980
rect 350 37910 360 37980
rect 140 37860 360 37910
rect 640 38090 860 38140
rect 640 38020 650 38090
rect 850 38020 860 38090
rect 640 37980 860 38020
rect 640 37910 650 37980
rect 850 37910 860 37980
rect 640 37860 860 37910
rect 0 37850 1000 37860
rect 0 37650 20 37850
rect 90 37650 410 37850
rect 480 37650 520 37850
rect 590 37650 910 37850
rect 980 37650 1000 37850
rect 0 37640 1000 37650
rect 140 37590 360 37640
rect 140 37520 150 37590
rect 350 37520 360 37590
rect 140 37480 360 37520
rect 140 37410 150 37480
rect 350 37410 360 37480
rect 140 37360 360 37410
rect 640 37590 860 37640
rect 640 37520 650 37590
rect 850 37520 860 37590
rect 640 37480 860 37520
rect 640 37410 650 37480
rect 850 37410 860 37480
rect 640 37360 860 37410
rect 0 37350 1000 37360
rect 0 37150 20 37350
rect 90 37150 410 37350
rect 480 37150 520 37350
rect 590 37150 910 37350
rect 980 37150 1000 37350
rect 0 37140 1000 37150
rect 140 37090 360 37140
rect 140 37020 150 37090
rect 350 37020 360 37090
rect 140 36980 360 37020
rect 140 36910 150 36980
rect 350 36910 360 36980
rect 140 36860 360 36910
rect 640 37090 860 37140
rect 640 37020 650 37090
rect 850 37020 860 37090
rect 640 36980 860 37020
rect 640 36910 650 36980
rect 850 36910 860 36980
rect 640 36860 860 36910
rect 0 36850 1000 36860
rect 0 36650 20 36850
rect 90 36650 410 36850
rect 480 36650 520 36850
rect 590 36650 910 36850
rect 980 36650 1000 36850
rect 0 36640 1000 36650
rect 140 36590 360 36640
rect 140 36520 150 36590
rect 350 36520 360 36590
rect 140 36480 360 36520
rect 140 36410 150 36480
rect 350 36410 360 36480
rect 140 36360 360 36410
rect 640 36590 860 36640
rect 640 36520 650 36590
rect 850 36520 860 36590
rect 640 36480 860 36520
rect 640 36410 650 36480
rect 850 36410 860 36480
rect 640 36360 860 36410
rect 0 36350 1000 36360
rect 0 36150 20 36350
rect 90 36150 410 36350
rect 480 36150 520 36350
rect 590 36150 910 36350
rect 980 36150 1000 36350
rect 0 36140 1000 36150
rect 140 36090 360 36140
rect 140 36020 150 36090
rect 350 36020 360 36090
rect 140 35980 360 36020
rect 140 35910 150 35980
rect 350 35910 360 35980
rect 140 35860 360 35910
rect 640 36090 860 36140
rect 640 36020 650 36090
rect 850 36020 860 36090
rect 640 35980 860 36020
rect 640 35910 650 35980
rect 850 35910 860 35980
rect 640 35860 860 35910
rect 0 35850 1000 35860
rect 0 35650 20 35850
rect 90 35650 410 35850
rect 480 35650 520 35850
rect 590 35650 910 35850
rect 980 35650 1000 35850
rect 0 35640 1000 35650
rect 140 35590 360 35640
rect 140 35520 150 35590
rect 350 35520 360 35590
rect 140 35480 360 35520
rect 140 35410 150 35480
rect 350 35410 360 35480
rect 140 35360 360 35410
rect 640 35590 860 35640
rect 640 35520 650 35590
rect 850 35520 860 35590
rect 640 35480 860 35520
rect 640 35410 650 35480
rect 850 35410 860 35480
rect 640 35360 860 35410
rect 0 35350 1000 35360
rect 0 35150 20 35350
rect 90 35150 410 35350
rect 480 35150 520 35350
rect 590 35150 910 35350
rect 980 35150 1000 35350
rect 0 35140 1000 35150
rect 140 35090 360 35140
rect 140 35020 150 35090
rect 350 35020 360 35090
rect 140 34980 360 35020
rect 140 34910 150 34980
rect 350 34910 360 34980
rect 140 34860 360 34910
rect 640 35090 860 35140
rect 640 35020 650 35090
rect 850 35020 860 35090
rect 640 34980 860 35020
rect 640 34910 650 34980
rect 850 34910 860 34980
rect 640 34860 860 34910
rect 0 34850 1000 34860
rect 0 34650 20 34850
rect 90 34650 410 34850
rect 480 34650 520 34850
rect 590 34650 910 34850
rect 980 34650 1000 34850
rect 0 34640 1000 34650
rect 140 34590 360 34640
rect 140 34520 150 34590
rect 350 34520 360 34590
rect 140 34480 360 34520
rect 140 34410 150 34480
rect 350 34410 360 34480
rect 140 34360 360 34410
rect 640 34590 860 34640
rect 640 34520 650 34590
rect 850 34520 860 34590
rect 640 34480 860 34520
rect 640 34410 650 34480
rect 850 34410 860 34480
rect 640 34360 860 34410
rect 0 34350 1000 34360
rect 0 34150 20 34350
rect 90 34150 410 34350
rect 480 34150 520 34350
rect 590 34150 910 34350
rect 980 34150 1000 34350
rect 0 34140 1000 34150
rect 140 34090 360 34140
rect 140 34020 150 34090
rect 350 34020 360 34090
rect 140 33980 360 34020
rect 140 33910 150 33980
rect 350 33910 360 33980
rect 140 33860 360 33910
rect 640 34090 860 34140
rect 640 34020 650 34090
rect 850 34020 860 34090
rect 640 33980 860 34020
rect 640 33910 650 33980
rect 850 33910 860 33980
rect 640 33860 860 33910
rect 0 33850 1000 33860
rect 0 33650 20 33850
rect 90 33650 410 33850
rect 480 33650 520 33850
rect 590 33650 910 33850
rect 980 33650 1000 33850
rect 0 33640 1000 33650
rect 140 33590 360 33640
rect 140 33520 150 33590
rect 350 33520 360 33590
rect 140 33480 360 33520
rect 140 33410 150 33480
rect 350 33410 360 33480
rect 140 33360 360 33410
rect 640 33590 860 33640
rect 640 33520 650 33590
rect 850 33520 860 33590
rect 640 33480 860 33520
rect 640 33410 650 33480
rect 850 33410 860 33480
rect 640 33360 860 33410
rect 0 33350 1000 33360
rect 0 33150 20 33350
rect 90 33150 410 33350
rect 480 33150 520 33350
rect 590 33150 910 33350
rect 980 33150 1000 33350
rect 0 33140 1000 33150
rect 140 33090 360 33140
rect 140 33020 150 33090
rect 350 33020 360 33090
rect 140 32980 360 33020
rect 140 32910 150 32980
rect 350 32910 360 32980
rect 140 32860 360 32910
rect 640 33090 860 33140
rect 640 33020 650 33090
rect 850 33020 860 33090
rect 640 32980 860 33020
rect 640 32910 650 32980
rect 850 32910 860 32980
rect 640 32860 860 32910
rect 0 32850 1000 32860
rect 0 32650 20 32850
rect 90 32650 410 32850
rect 480 32650 520 32850
rect 590 32650 910 32850
rect 980 32650 1000 32850
rect 6340 39120 7700 39180
rect 1532 39080 1552 39090
rect 6186 39080 6206 39090
rect 1532 39010 1540 39080
rect 6200 39010 6206 39080
rect 1532 38990 1552 39010
rect 6186 38990 6206 39010
rect 1465 38938 1531 38958
rect 1465 32958 1531 32978
rect 1623 38938 1689 38958
rect 1623 32958 1689 32978
rect 1781 38938 1847 38958
rect 1781 32958 1847 32978
rect 1939 38938 2005 38958
rect 1939 32958 2005 32978
rect 2097 38938 2163 38958
rect 2097 32958 2163 32978
rect 2255 38938 2321 38958
rect 2255 32958 2321 32978
rect 2413 38938 2479 38958
rect 2413 32958 2479 32978
rect 2571 38938 2637 38958
rect 2571 32958 2637 32978
rect 2729 38938 2795 38958
rect 2729 32958 2795 32978
rect 2887 38938 2953 38958
rect 2887 32958 2953 32978
rect 3045 38938 3111 38958
rect 3045 32958 3111 32978
rect 3203 38938 3269 38958
rect 3203 32958 3269 32978
rect 3361 38938 3427 38958
rect 3361 32958 3427 32978
rect 3519 38938 3585 38958
rect 3519 32958 3585 32978
rect 3677 38938 3743 38958
rect 3677 32958 3743 32978
rect 3835 38938 3901 38958
rect 3835 32958 3901 32978
rect 3993 38938 4059 38958
rect 3993 32958 4059 32978
rect 4151 38938 4217 38958
rect 4151 32958 4217 32978
rect 4309 38938 4375 38958
rect 4309 32958 4375 32978
rect 4467 38938 4533 38958
rect 4467 32958 4533 32978
rect 4625 38938 4691 38958
rect 4625 32958 4691 32978
rect 4783 38938 4849 38958
rect 4783 32958 4849 32978
rect 4941 38938 5007 38958
rect 4941 32958 5007 32978
rect 5099 38938 5165 38958
rect 5099 32958 5165 32978
rect 5257 38938 5323 38958
rect 5257 32958 5323 32978
rect 5415 38938 5481 38958
rect 5415 32958 5481 32978
rect 5573 38938 5639 38958
rect 5573 32958 5639 32978
rect 5731 38938 5797 38958
rect 5731 32958 5797 32978
rect 5889 38938 5955 38958
rect 5889 32958 5955 32978
rect 6047 38938 6113 38958
rect 6047 32958 6113 32978
rect 6205 38938 6271 38958
rect 6205 32958 6271 32978
rect 1532 32910 1552 32926
rect 6186 32910 6206 32926
rect 1532 32840 1540 32910
rect 6190 32840 6206 32910
rect 1532 32826 1552 32840
rect 6186 32826 6206 32840
rect 1330 32730 1400 32800
rect 6410 38800 7630 39120
rect 6410 38200 7630 38600
rect 6410 37600 7630 38000
rect 6410 37000 7630 37400
rect 6410 36400 7630 36800
rect 6410 35800 7630 36200
rect 6410 35200 7630 35600
rect 6410 34600 7630 35000
rect 6410 34000 7630 34400
rect 6410 33400 7630 33800
rect 6410 32980 7630 33200
rect 6410 32910 6650 32980
rect 6850 32910 7150 32980
rect 7350 32910 7630 32980
rect 6410 32850 7630 32910
rect 6410 32800 6520 32850
rect 6340 32730 6410 32800
rect 0 32640 1000 32650
rect 6500 32650 6520 32800
rect 6590 32650 6910 32850
rect 6980 32650 7020 32850
rect 7090 32650 7410 32850
rect 7480 32800 7630 32850
rect 12640 39120 14000 39180
rect 7832 39080 7852 39090
rect 12486 39080 12506 39090
rect 7832 39010 7840 39080
rect 12500 39010 12506 39080
rect 7832 38990 7852 39010
rect 12486 38990 12506 39010
rect 7765 38938 7831 38958
rect 7765 32958 7831 32978
rect 7923 38938 7989 38958
rect 7923 32958 7989 32978
rect 8081 38938 8147 38958
rect 8081 32958 8147 32978
rect 8239 38938 8305 38958
rect 8239 32958 8305 32978
rect 8397 38938 8463 38958
rect 8397 32958 8463 32978
rect 8555 38938 8621 38958
rect 8555 32958 8621 32978
rect 8713 38938 8779 38958
rect 8713 32958 8779 32978
rect 8871 38938 8937 38958
rect 8871 32958 8937 32978
rect 9029 38938 9095 38958
rect 9029 32958 9095 32978
rect 9187 38938 9253 38958
rect 9187 32958 9253 32978
rect 9345 38938 9411 38958
rect 9345 32958 9411 32978
rect 9503 38938 9569 38958
rect 9503 32958 9569 32978
rect 9661 38938 9727 38958
rect 9661 32958 9727 32978
rect 9819 38938 9885 38958
rect 9819 32958 9885 32978
rect 9977 38938 10043 38958
rect 9977 32958 10043 32978
rect 10135 38938 10201 38958
rect 10135 32958 10201 32978
rect 10293 38938 10359 38958
rect 10293 32958 10359 32978
rect 10451 38938 10517 38958
rect 10451 32958 10517 32978
rect 10609 38938 10675 38958
rect 10609 32958 10675 32978
rect 10767 38938 10833 38958
rect 10767 32958 10833 32978
rect 10925 38938 10991 38958
rect 10925 32958 10991 32978
rect 11083 38938 11149 38958
rect 11083 32958 11149 32978
rect 11241 38938 11307 38958
rect 11241 32958 11307 32978
rect 11399 38938 11465 38958
rect 11399 32958 11465 32978
rect 11557 38938 11623 38958
rect 11557 32958 11623 32978
rect 11715 38938 11781 38958
rect 11715 32958 11781 32978
rect 11873 38938 11939 38958
rect 11873 32958 11939 32978
rect 12031 38938 12097 38958
rect 12031 32958 12097 32978
rect 12189 38938 12255 38958
rect 12189 32958 12255 32978
rect 12347 38938 12413 38958
rect 12347 32958 12413 32978
rect 12505 38938 12571 38958
rect 12505 32958 12571 32978
rect 7832 32910 7852 32926
rect 12486 32910 12506 32926
rect 7832 32840 7840 32910
rect 12490 32840 12506 32910
rect 7832 32826 7852 32840
rect 12486 32826 12506 32840
rect 7480 32650 7500 32800
rect 7630 32730 7700 32800
rect 12710 38800 13930 39120
rect 12710 38200 13930 38600
rect 12710 37600 13930 38000
rect 12710 37000 13930 37400
rect 12710 36400 13930 36800
rect 12710 35800 13930 36200
rect 12710 35200 13930 35600
rect 12710 34600 13930 35000
rect 12710 34000 13930 34400
rect 12710 33400 13930 33800
rect 12710 32980 13930 33200
rect 12710 32910 13150 32980
rect 13350 32910 13930 32980
rect 12710 32850 13930 32910
rect 12710 32800 13020 32850
rect 12640 32730 12710 32800
rect 6500 32640 7500 32650
rect 13000 32650 13020 32800
rect 13090 32650 13410 32850
rect 13480 32800 13930 32850
rect 18940 39120 20300 39180
rect 14132 39080 14152 39090
rect 18786 39080 18806 39090
rect 14132 39010 14140 39080
rect 18800 39010 18806 39080
rect 14132 38990 14152 39010
rect 18786 38990 18806 39010
rect 14065 38938 14131 38958
rect 14065 32958 14131 32978
rect 14223 38938 14289 38958
rect 14223 32958 14289 32978
rect 14381 38938 14447 38958
rect 14381 32958 14447 32978
rect 14539 38938 14605 38958
rect 14539 32958 14605 32978
rect 14697 38938 14763 38958
rect 14697 32958 14763 32978
rect 14855 38938 14921 38958
rect 14855 32958 14921 32978
rect 15013 38938 15079 38958
rect 15013 32958 15079 32978
rect 15171 38938 15237 38958
rect 15171 32958 15237 32978
rect 15329 38938 15395 38958
rect 15329 32958 15395 32978
rect 15487 38938 15553 38958
rect 15487 32958 15553 32978
rect 15645 38938 15711 38958
rect 15645 32958 15711 32978
rect 15803 38938 15869 38958
rect 15803 32958 15869 32978
rect 15961 38938 16027 38958
rect 15961 32958 16027 32978
rect 16119 38938 16185 38958
rect 16119 32958 16185 32978
rect 16277 38938 16343 38958
rect 16277 32958 16343 32978
rect 16435 38938 16501 38958
rect 16435 32958 16501 32978
rect 16593 38938 16659 38958
rect 16593 32958 16659 32978
rect 16751 38938 16817 38958
rect 16751 32958 16817 32978
rect 16909 38938 16975 38958
rect 16909 32958 16975 32978
rect 17067 38938 17133 38958
rect 17067 32958 17133 32978
rect 17225 38938 17291 38958
rect 17225 32958 17291 32978
rect 17383 38938 17449 38958
rect 17383 32958 17449 32978
rect 17541 38938 17607 38958
rect 17541 32958 17607 32978
rect 17699 38938 17765 38958
rect 17699 32958 17765 32978
rect 17857 38938 17923 38958
rect 17857 32958 17923 32978
rect 18015 38938 18081 38958
rect 18015 32958 18081 32978
rect 18173 38938 18239 38958
rect 18173 32958 18239 32978
rect 18331 38938 18397 38958
rect 18331 32958 18397 32978
rect 18489 38938 18555 38958
rect 18489 32958 18555 32978
rect 18647 38938 18713 38958
rect 18647 32958 18713 32978
rect 18805 38938 18871 38958
rect 18805 32958 18871 32978
rect 14132 32910 14152 32926
rect 18786 32910 18806 32926
rect 14132 32840 14140 32910
rect 18790 32840 18806 32910
rect 14132 32826 14152 32840
rect 18786 32826 18806 32840
rect 13480 32650 13500 32800
rect 13930 32730 14000 32800
rect 19010 38800 20230 39120
rect 19010 38200 20230 38600
rect 19010 37600 20230 38000
rect 19010 37000 20230 37400
rect 19010 36400 20230 36800
rect 19010 35800 20230 36200
rect 19010 35200 20230 35600
rect 19010 34600 20230 35000
rect 19010 34000 20230 34400
rect 19010 33400 20230 33800
rect 19010 32980 20230 33200
rect 19010 32910 19650 32980
rect 19850 32910 20230 32980
rect 19010 32850 20230 32910
rect 19010 32800 19520 32850
rect 18940 32730 19010 32800
rect 13000 32640 13500 32650
rect 19500 32650 19520 32800
rect 19590 32650 19910 32850
rect 19980 32800 20230 32850
rect 25240 39120 25310 39180
rect 25500 39150 25520 39350
rect 25590 39150 25910 39350
rect 25980 39150 26020 39350
rect 26090 39150 26410 39350
rect 26480 39150 26520 39350
rect 26590 39150 26910 39350
rect 26980 39150 27020 39350
rect 27090 39150 27410 39350
rect 27480 39150 27520 39350
rect 27590 39150 27910 39350
rect 27980 39150 28020 39350
rect 28090 39150 28410 39350
rect 28480 39150 28520 39350
rect 28590 39150 28910 39350
rect 28980 39150 29020 39350
rect 29090 39150 29410 39350
rect 29480 39150 29500 39350
rect 25500 39140 29500 39150
rect 20432 39080 20452 39090
rect 25086 39080 25106 39090
rect 20432 39010 20440 39080
rect 25100 39010 25106 39080
rect 20432 38990 20452 39010
rect 25086 38990 25106 39010
rect 20365 38938 20431 38958
rect 20365 32958 20431 32978
rect 20523 38938 20589 38958
rect 20523 32958 20589 32978
rect 20681 38938 20747 38958
rect 20681 32958 20747 32978
rect 20839 38938 20905 38958
rect 20839 32958 20905 32978
rect 20997 38938 21063 38958
rect 20997 32958 21063 32978
rect 21155 38938 21221 38958
rect 21155 32958 21221 32978
rect 21313 38938 21379 38958
rect 21313 32958 21379 32978
rect 21471 38938 21537 38958
rect 21471 32958 21537 32978
rect 21629 38938 21695 38958
rect 21629 32958 21695 32978
rect 21787 38938 21853 38958
rect 21787 32958 21853 32978
rect 21945 38938 22011 38958
rect 21945 32958 22011 32978
rect 22103 38938 22169 38958
rect 22103 32958 22169 32978
rect 22261 38938 22327 38958
rect 22261 32958 22327 32978
rect 22419 38938 22485 38958
rect 22419 32958 22485 32978
rect 22577 38938 22643 38958
rect 22577 32958 22643 32978
rect 22735 38938 22801 38958
rect 22735 32958 22801 32978
rect 22893 38938 22959 38958
rect 22893 32958 22959 32978
rect 23051 38938 23117 38958
rect 23051 32958 23117 32978
rect 23209 38938 23275 38958
rect 23209 32958 23275 32978
rect 23367 38938 23433 38958
rect 23367 32958 23433 32978
rect 23525 38938 23591 38958
rect 23525 32958 23591 32978
rect 23683 38938 23749 38958
rect 23683 32958 23749 32978
rect 23841 38938 23907 38958
rect 23841 32958 23907 32978
rect 23999 38938 24065 38958
rect 23999 32958 24065 32978
rect 24157 38938 24223 38958
rect 24157 32958 24223 32978
rect 24315 38938 24381 38958
rect 24315 32958 24381 32978
rect 24473 38938 24539 38958
rect 24473 32958 24539 32978
rect 24631 38938 24697 38958
rect 24631 32958 24697 32978
rect 24789 38938 24855 38958
rect 24789 32958 24855 32978
rect 24947 38938 25013 38958
rect 24947 32958 25013 32978
rect 25105 38938 25171 38958
rect 25105 32958 25171 32978
rect 20432 32910 20452 32926
rect 25086 32910 25106 32926
rect 20432 32840 20440 32910
rect 25090 32840 25106 32910
rect 20432 32826 20452 32840
rect 25086 32826 25106 32840
rect 19980 32650 20000 32800
rect 20230 32730 20300 32800
rect 25640 39090 25860 39140
rect 25640 39020 25650 39090
rect 25850 39020 25860 39090
rect 25640 38980 25860 39020
rect 25640 38910 25650 38980
rect 25850 38910 25860 38980
rect 25640 38860 25860 38910
rect 26140 39090 26360 39140
rect 26140 39020 26150 39090
rect 26350 39020 26360 39090
rect 26140 38980 26360 39020
rect 26640 39090 26860 39140
rect 26640 39020 26650 39090
rect 26850 39020 26860 39090
rect 26640 39000 26860 39020
rect 27140 39090 27360 39140
rect 27140 39020 27150 39090
rect 27350 39020 27360 39090
rect 27140 39000 27360 39020
rect 27640 39090 27860 39140
rect 27640 39020 27650 39090
rect 27850 39020 27860 39090
rect 27640 39000 27860 39020
rect 28140 39090 28360 39140
rect 28140 39020 28150 39090
rect 28350 39020 28360 39090
rect 28140 39000 28360 39020
rect 28640 39090 28860 39140
rect 28640 39020 28650 39090
rect 28850 39020 28860 39090
rect 28640 39000 28860 39020
rect 29140 39090 29360 39140
rect 29140 39020 29150 39090
rect 29350 39020 29360 39090
rect 29140 39000 29360 39020
rect 26140 38910 26150 38980
rect 26350 38910 26360 38980
rect 26140 38860 26360 38910
rect 29900 38910 30100 38920
rect 25500 38850 26500 38860
rect 25500 38650 25520 38850
rect 25590 38650 25910 38850
rect 25980 38650 26020 38850
rect 26090 38650 26410 38850
rect 26480 38650 26500 38850
rect 29900 38690 29910 38910
rect 30090 38690 30100 38910
rect 29900 38680 30100 38690
rect 25500 38640 26500 38650
rect 25640 38590 25860 38640
rect 25640 38520 25650 38590
rect 25850 38520 25860 38590
rect 25640 38480 25860 38520
rect 25640 38410 25650 38480
rect 25850 38410 25860 38480
rect 25640 38360 25860 38410
rect 26140 38590 26360 38640
rect 26140 38520 26150 38590
rect 26350 38520 26360 38590
rect 26140 38480 26360 38520
rect 26140 38410 26150 38480
rect 26350 38410 26360 38480
rect 26140 38360 26360 38410
rect 25500 38350 26500 38360
rect 25500 38150 25520 38350
rect 25590 38150 25910 38350
rect 25980 38150 26020 38350
rect 26090 38150 26410 38350
rect 26480 38150 26500 38350
rect 25500 38140 26500 38150
rect 25640 38090 25860 38140
rect 25640 38020 25650 38090
rect 25850 38020 25860 38090
rect 25640 37980 25860 38020
rect 25640 37910 25650 37980
rect 25850 37910 25860 37980
rect 25640 37860 25860 37910
rect 26140 38090 26360 38140
rect 26140 38020 26150 38090
rect 26350 38020 26360 38090
rect 26140 37980 26360 38020
rect 26140 37910 26150 37980
rect 26350 37910 26360 37980
rect 26140 37860 26360 37910
rect 25500 37850 26500 37860
rect 25500 37650 25520 37850
rect 25590 37650 25910 37850
rect 25980 37650 26020 37850
rect 26090 37650 26410 37850
rect 26480 37650 26500 37850
rect 25500 37640 26500 37650
rect 25640 37590 25860 37640
rect 25640 37520 25650 37590
rect 25850 37520 25860 37590
rect 25640 37480 25860 37520
rect 25640 37410 25650 37480
rect 25850 37410 25860 37480
rect 25640 37360 25860 37410
rect 26140 37590 26360 37640
rect 26140 37520 26150 37590
rect 26350 37520 26360 37590
rect 26140 37480 26360 37520
rect 26140 37410 26150 37480
rect 26350 37410 26360 37480
rect 26140 37360 26360 37410
rect 25500 37350 26500 37360
rect 25500 37150 25520 37350
rect 25590 37150 25910 37350
rect 25980 37150 26020 37350
rect 26090 37150 26410 37350
rect 26480 37150 26500 37350
rect 25500 37140 26500 37150
rect 25640 37090 25860 37140
rect 25640 37020 25650 37090
rect 25850 37020 25860 37090
rect 25640 36980 25860 37020
rect 25640 36910 25650 36980
rect 25850 36910 25860 36980
rect 25640 36860 25860 36910
rect 26140 37090 26360 37140
rect 26140 37020 26150 37090
rect 26350 37020 26360 37090
rect 26140 36980 26360 37020
rect 26140 36910 26150 36980
rect 26350 36910 26360 36980
rect 26140 36860 26360 36910
rect 25500 36850 26500 36860
rect 25500 36650 25520 36850
rect 25590 36650 25910 36850
rect 25980 36650 26020 36850
rect 26090 36650 26410 36850
rect 26480 36650 26500 36850
rect 25500 36640 26500 36650
rect 25640 36590 25860 36640
rect 25640 36520 25650 36590
rect 25850 36520 25860 36590
rect 25640 36480 25860 36520
rect 25640 36410 25650 36480
rect 25850 36410 25860 36480
rect 25640 36360 25860 36410
rect 26140 36590 26360 36640
rect 26140 36520 26150 36590
rect 26350 36520 26360 36590
rect 26140 36480 26360 36520
rect 26140 36410 26150 36480
rect 26350 36410 26360 36480
rect 26140 36360 26360 36410
rect 25500 36350 26500 36360
rect 25500 36150 25520 36350
rect 25590 36150 25910 36350
rect 25980 36150 26020 36350
rect 26090 36150 26410 36350
rect 26480 36150 26500 36350
rect 25500 36140 26500 36150
rect 25640 36090 25860 36140
rect 25640 36020 25650 36090
rect 25850 36020 25860 36090
rect 25640 35980 25860 36020
rect 25640 35910 25650 35980
rect 25850 35910 25860 35980
rect 25640 35860 25860 35910
rect 26140 36090 26360 36140
rect 26140 36020 26150 36090
rect 26350 36020 26360 36090
rect 26140 35980 26360 36020
rect 26140 35910 26150 35980
rect 26350 35910 26360 35980
rect 26140 35860 26360 35910
rect 25500 35850 26500 35860
rect 25500 35650 25520 35850
rect 25590 35650 25910 35850
rect 25980 35650 26020 35850
rect 26090 35650 26410 35850
rect 26480 35650 26500 35850
rect 25500 35640 26500 35650
rect 25640 35590 25860 35640
rect 25640 35520 25650 35590
rect 25850 35520 25860 35590
rect 25640 35480 25860 35520
rect 25640 35410 25650 35480
rect 25850 35410 25860 35480
rect 25640 35360 25860 35410
rect 26140 35590 26360 35640
rect 26140 35520 26150 35590
rect 26350 35520 26360 35590
rect 26140 35480 26360 35520
rect 26140 35410 26150 35480
rect 26350 35410 26360 35480
rect 26140 35360 26360 35410
rect 25500 35350 26500 35360
rect 25500 35150 25520 35350
rect 25590 35150 25910 35350
rect 25980 35150 26020 35350
rect 26090 35150 26410 35350
rect 26480 35150 26500 35350
rect 25500 35140 26500 35150
rect 25640 35090 25860 35140
rect 25640 35020 25650 35090
rect 25850 35020 25860 35090
rect 25640 34980 25860 35020
rect 25640 34910 25650 34980
rect 25850 34910 25860 34980
rect 25640 34860 25860 34910
rect 26140 35090 26360 35140
rect 26140 35020 26150 35090
rect 26350 35020 26360 35090
rect 26140 34980 26360 35020
rect 26140 34910 26150 34980
rect 26350 34910 26360 34980
rect 26140 34860 26360 34910
rect 25500 34850 26500 34860
rect 25500 34650 25520 34850
rect 25590 34650 25910 34850
rect 25980 34650 26020 34850
rect 26090 34650 26410 34850
rect 26480 34650 26500 34850
rect 25500 34640 26500 34650
rect 25640 34590 25860 34640
rect 25640 34520 25650 34590
rect 25850 34520 25860 34590
rect 25640 34480 25860 34520
rect 25640 34410 25650 34480
rect 25850 34410 25860 34480
rect 25640 34360 25860 34410
rect 26140 34590 26360 34640
rect 26140 34520 26150 34590
rect 26350 34520 26360 34590
rect 26140 34480 26360 34520
rect 26140 34410 26150 34480
rect 26350 34410 26360 34480
rect 26140 34360 26360 34410
rect 25500 34350 26500 34360
rect 25500 34150 25520 34350
rect 25590 34150 25910 34350
rect 25980 34150 26020 34350
rect 26090 34150 26410 34350
rect 26480 34150 26500 34350
rect 25500 34140 26500 34150
rect 25640 34090 25860 34140
rect 25640 34020 25650 34090
rect 25850 34020 25860 34090
rect 25640 33980 25860 34020
rect 25640 33910 25650 33980
rect 25850 33910 25860 33980
rect 25640 33860 25860 33910
rect 26140 34090 26360 34140
rect 26140 34020 26150 34090
rect 26350 34020 26360 34090
rect 26140 33980 26360 34020
rect 26140 33910 26150 33980
rect 26350 33910 26360 33980
rect 26140 33860 26360 33910
rect 25500 33850 26500 33860
rect 25500 33650 25520 33850
rect 25590 33650 25910 33850
rect 25980 33650 26020 33850
rect 26090 33650 26410 33850
rect 26480 33650 26500 33850
rect 25500 33640 26500 33650
rect 25640 33590 25860 33640
rect 25640 33520 25650 33590
rect 25850 33520 25860 33590
rect 25640 33480 25860 33520
rect 25640 33410 25650 33480
rect 25850 33410 25860 33480
rect 25640 33360 25860 33410
rect 26140 33590 26360 33640
rect 26140 33520 26150 33590
rect 26350 33520 26360 33590
rect 26140 33480 26360 33520
rect 26140 33410 26150 33480
rect 26350 33410 26360 33480
rect 26140 33360 26360 33410
rect 25500 33350 26500 33360
rect 25500 33150 25520 33350
rect 25590 33150 25910 33350
rect 25980 33150 26020 33350
rect 26090 33150 26410 33350
rect 26480 33150 26500 33350
rect 25500 33140 26500 33150
rect 25640 33090 25860 33140
rect 25640 33020 25650 33090
rect 25850 33020 25860 33090
rect 25640 32980 25860 33020
rect 25640 32910 25650 32980
rect 25850 32910 25860 32980
rect 25640 32860 25860 32910
rect 26140 33090 26360 33140
rect 26140 33020 26150 33090
rect 26350 33020 26360 33090
rect 26140 32980 26360 33020
rect 26140 32910 26150 32980
rect 26350 32910 26360 32980
rect 26140 32860 26360 32910
rect 25240 32730 25310 32800
rect 25500 32850 26500 32860
rect 19500 32640 20000 32650
rect 25500 32650 25520 32850
rect 25590 32650 25910 32850
rect 25980 32650 26020 32850
rect 26090 32650 26410 32850
rect 26480 32650 26500 32850
rect 25500 32640 26500 32650
rect 140 32590 360 32640
rect 140 32520 150 32590
rect 350 32520 360 32590
rect 140 32480 360 32520
rect 140 32410 150 32480
rect 350 32410 360 32480
rect 140 32360 360 32410
rect 640 32590 860 32640
rect 640 32520 650 32590
rect 850 32520 860 32590
rect 640 32480 860 32520
rect 6640 32590 6860 32640
rect 6640 32520 6650 32590
rect 6850 32520 6860 32590
rect 640 32410 650 32480
rect 850 32410 860 32480
rect 640 32360 860 32410
rect 1140 32480 1360 32500
rect 1140 32410 1150 32480
rect 1350 32410 1360 32480
rect 1140 32360 1360 32410
rect 1640 32480 1860 32500
rect 1640 32410 1650 32480
rect 1850 32410 1860 32480
rect 1640 32360 1860 32410
rect 2140 32480 2360 32500
rect 2140 32410 2150 32480
rect 2350 32410 2360 32480
rect 2140 32360 2360 32410
rect 2640 32480 2860 32500
rect 2640 32410 2650 32480
rect 2850 32410 2860 32480
rect 2640 32360 2860 32410
rect 3140 32480 3360 32500
rect 3140 32410 3150 32480
rect 3350 32410 3360 32480
rect 3140 32360 3360 32410
rect 3640 32480 3860 32500
rect 3640 32410 3650 32480
rect 3850 32410 3860 32480
rect 3640 32360 3860 32410
rect 4140 32480 4360 32500
rect 4140 32410 4150 32480
rect 4350 32410 4360 32480
rect 4140 32360 4360 32410
rect 4640 32480 4860 32500
rect 4640 32410 4650 32480
rect 4850 32410 4860 32480
rect 4640 32360 4860 32410
rect 5140 32480 5360 32500
rect 5140 32410 5150 32480
rect 5350 32410 5360 32480
rect 5140 32360 5360 32410
rect 5640 32480 5860 32500
rect 5640 32410 5650 32480
rect 5850 32410 5860 32480
rect 5640 32360 5860 32410
rect 6140 32480 6360 32500
rect 6140 32410 6150 32480
rect 6350 32410 6360 32480
rect 6140 32360 6360 32410
rect 6640 32480 6860 32520
rect 6640 32410 6650 32480
rect 6850 32410 6860 32480
rect 6640 32360 6860 32410
rect 7140 32590 7360 32640
rect 7140 32520 7150 32590
rect 7350 32520 7360 32590
rect 7140 32480 7360 32520
rect 13140 32590 13360 32640
rect 13140 32520 13150 32590
rect 13350 32520 13360 32590
rect 7140 32410 7150 32480
rect 7350 32410 7360 32480
rect 7140 32360 7360 32410
rect 7640 32480 7860 32500
rect 7640 32410 7650 32480
rect 7850 32410 7860 32480
rect 7640 32360 7860 32410
rect 8140 32480 8360 32500
rect 8140 32410 8150 32480
rect 8350 32410 8360 32480
rect 8140 32360 8360 32410
rect 8640 32480 8860 32500
rect 8640 32410 8650 32480
rect 8850 32410 8860 32480
rect 8640 32360 8860 32410
rect 9140 32480 9360 32500
rect 9140 32410 9150 32480
rect 9350 32410 9360 32480
rect 9140 32360 9360 32410
rect 9640 32480 9860 32500
rect 9640 32410 9650 32480
rect 9850 32410 9860 32480
rect 9640 32360 9860 32410
rect 10140 32480 10360 32500
rect 10140 32410 10150 32480
rect 10350 32410 10360 32480
rect 10140 32360 10360 32410
rect 10640 32480 10860 32500
rect 10640 32410 10650 32480
rect 10850 32410 10860 32480
rect 10640 32360 10860 32410
rect 11140 32480 11360 32500
rect 11140 32410 11150 32480
rect 11350 32410 11360 32480
rect 11140 32360 11360 32410
rect 11640 32480 11860 32500
rect 11640 32410 11650 32480
rect 11850 32410 11860 32480
rect 11640 32360 11860 32410
rect 12140 32480 12360 32500
rect 12140 32410 12150 32480
rect 12350 32410 12360 32480
rect 12140 32360 12360 32410
rect 12640 32480 12860 32500
rect 12640 32410 12650 32480
rect 12850 32410 12860 32480
rect 12640 32360 12860 32410
rect 13140 32480 13360 32520
rect 19640 32590 19860 32640
rect 19640 32520 19650 32590
rect 19850 32520 19860 32590
rect 13140 32410 13150 32480
rect 13350 32410 13360 32480
rect 13140 32360 13360 32410
rect 13640 32480 13860 32500
rect 13640 32410 13650 32480
rect 13850 32410 13860 32480
rect 13640 32360 13860 32410
rect 14140 32480 14360 32500
rect 14140 32410 14150 32480
rect 14350 32410 14360 32480
rect 14140 32360 14360 32410
rect 14640 32480 14860 32500
rect 14640 32410 14650 32480
rect 14850 32410 14860 32480
rect 14640 32360 14860 32410
rect 15140 32480 15360 32500
rect 15140 32410 15150 32480
rect 15350 32410 15360 32480
rect 15140 32360 15360 32410
rect 15640 32480 15860 32500
rect 15640 32410 15650 32480
rect 15850 32410 15860 32480
rect 15640 32360 15860 32410
rect 16140 32480 16360 32500
rect 16140 32410 16150 32480
rect 16350 32410 16360 32480
rect 16140 32360 16360 32410
rect 16640 32480 16860 32500
rect 16640 32410 16650 32480
rect 16850 32410 16860 32480
rect 16640 32360 16860 32410
rect 17140 32480 17360 32500
rect 17140 32410 17150 32480
rect 17350 32410 17360 32480
rect 17140 32360 17360 32410
rect 17640 32480 17860 32500
rect 17640 32410 17650 32480
rect 17850 32410 17860 32480
rect 17640 32360 17860 32410
rect 18140 32480 18360 32500
rect 18140 32410 18150 32480
rect 18350 32410 18360 32480
rect 18140 32360 18360 32410
rect 18640 32480 18860 32500
rect 18640 32410 18650 32480
rect 18850 32410 18860 32480
rect 18640 32360 18860 32410
rect 19140 32480 19360 32500
rect 19140 32410 19150 32480
rect 19350 32410 19360 32480
rect 19140 32360 19360 32410
rect 19640 32480 19860 32520
rect 25640 32590 25860 32640
rect 25640 32520 25650 32590
rect 25850 32520 25860 32590
rect 19640 32410 19650 32480
rect 19850 32410 19860 32480
rect 19640 32360 19860 32410
rect 20140 32480 20360 32500
rect 20140 32410 20150 32480
rect 20350 32410 20360 32480
rect 20140 32360 20360 32410
rect 20640 32480 20860 32500
rect 20640 32410 20650 32480
rect 20850 32410 20860 32480
rect 20640 32360 20860 32410
rect 21140 32480 21360 32500
rect 21140 32410 21150 32480
rect 21350 32410 21360 32480
rect 21140 32360 21360 32410
rect 21640 32480 21860 32500
rect 21640 32410 21650 32480
rect 21850 32410 21860 32480
rect 21640 32360 21860 32410
rect 22140 32480 22360 32500
rect 22140 32410 22150 32480
rect 22350 32410 22360 32480
rect 22140 32360 22360 32410
rect 22640 32480 22860 32500
rect 22640 32410 22650 32480
rect 22850 32410 22860 32480
rect 22640 32360 22860 32410
rect 23140 32480 23360 32500
rect 23140 32410 23150 32480
rect 23350 32410 23360 32480
rect 23140 32360 23360 32410
rect 23640 32480 23860 32500
rect 23640 32410 23650 32480
rect 23850 32410 23860 32480
rect 23640 32360 23860 32410
rect 24140 32480 24360 32500
rect 24140 32410 24150 32480
rect 24350 32410 24360 32480
rect 24140 32360 24360 32410
rect 24640 32480 24860 32500
rect 24640 32410 24650 32480
rect 24850 32410 24860 32480
rect 24640 32360 24860 32410
rect 25140 32480 25360 32500
rect 25140 32410 25150 32480
rect 25350 32410 25360 32480
rect 25140 32360 25360 32410
rect 25640 32480 25860 32520
rect 25640 32410 25650 32480
rect 25850 32410 25860 32480
rect 25640 32360 25860 32410
rect 26140 32590 26360 32640
rect 26140 32520 26150 32590
rect 26350 32520 26360 32590
rect 26140 32480 26360 32520
rect 26140 32410 26150 32480
rect 26350 32410 26360 32480
rect 26140 32360 26360 32410
rect 0 32350 26500 32360
rect 0 32150 20 32350
rect 90 32150 410 32350
rect 480 32150 520 32350
rect 590 32150 910 32350
rect 980 32150 1020 32350
rect 1090 32150 1410 32350
rect 1480 32150 1520 32350
rect 1590 32150 1910 32350
rect 1980 32150 2020 32350
rect 2090 32150 2410 32350
rect 2480 32150 2520 32350
rect 2590 32150 2910 32350
rect 2980 32150 3020 32350
rect 3090 32150 3410 32350
rect 3480 32150 3520 32350
rect 3590 32150 3910 32350
rect 3980 32150 4020 32350
rect 4090 32150 4410 32350
rect 4480 32150 4520 32350
rect 4590 32150 4910 32350
rect 4980 32150 5020 32350
rect 5090 32150 5410 32350
rect 5480 32150 5520 32350
rect 5590 32150 5910 32350
rect 5980 32150 6020 32350
rect 6090 32150 6410 32350
rect 6480 32150 6520 32350
rect 6590 32150 6910 32350
rect 6980 32150 7020 32350
rect 7090 32150 7410 32350
rect 7480 32150 7520 32350
rect 7590 32150 7910 32350
rect 7980 32150 8020 32350
rect 8090 32150 8410 32350
rect 8480 32150 8520 32350
rect 8590 32150 8910 32350
rect 8980 32150 9020 32350
rect 9090 32150 9410 32350
rect 9480 32150 9520 32350
rect 9590 32150 9910 32350
rect 9980 32150 10020 32350
rect 10090 32150 10410 32350
rect 10480 32150 10520 32350
rect 10590 32150 10910 32350
rect 10980 32150 11020 32350
rect 11090 32150 11410 32350
rect 11480 32150 11520 32350
rect 11590 32150 11910 32350
rect 11980 32150 12020 32350
rect 12090 32150 12410 32350
rect 12480 32150 12520 32350
rect 12590 32150 12910 32350
rect 12980 32150 13020 32350
rect 13090 32150 13410 32350
rect 13480 32150 13520 32350
rect 13590 32150 13910 32350
rect 13980 32150 14020 32350
rect 14090 32150 14410 32350
rect 14480 32150 14520 32350
rect 14590 32150 14910 32350
rect 14980 32150 15020 32350
rect 15090 32150 15410 32350
rect 15480 32150 15520 32350
rect 15590 32150 15910 32350
rect 15980 32150 16020 32350
rect 16090 32150 16410 32350
rect 16480 32150 16520 32350
rect 16590 32150 16910 32350
rect 16980 32150 17020 32350
rect 17090 32150 17410 32350
rect 17480 32150 17520 32350
rect 17590 32150 17910 32350
rect 17980 32150 18020 32350
rect 18090 32150 18410 32350
rect 18480 32150 18520 32350
rect 18590 32150 18910 32350
rect 18980 32150 19020 32350
rect 19090 32150 19410 32350
rect 19480 32150 19520 32350
rect 19590 32150 19910 32350
rect 19980 32150 20020 32350
rect 20090 32150 20410 32350
rect 20480 32150 20520 32350
rect 20590 32150 20910 32350
rect 20980 32150 21020 32350
rect 21090 32150 21410 32350
rect 21480 32150 21520 32350
rect 21590 32150 21910 32350
rect 21980 32150 22020 32350
rect 22090 32150 22410 32350
rect 22480 32150 22520 32350
rect 22590 32150 22910 32350
rect 22980 32150 23020 32350
rect 23090 32150 23410 32350
rect 23480 32150 23520 32350
rect 23590 32150 23910 32350
rect 23980 32150 24020 32350
rect 24090 32150 24410 32350
rect 24480 32150 24520 32350
rect 24590 32150 24910 32350
rect 24980 32150 25020 32350
rect 25090 32150 25410 32350
rect 25480 32150 25520 32350
rect 25590 32150 25910 32350
rect 25980 32150 26020 32350
rect 26090 32150 26410 32350
rect 26480 32150 26500 32350
rect 0 32140 26500 32150
rect 140 32090 360 32140
rect 140 32020 150 32090
rect 350 32020 360 32090
rect 140 31980 360 32020
rect 140 31910 150 31980
rect 350 31910 360 31980
rect 140 31860 360 31910
rect 640 32090 860 32140
rect 640 32020 650 32090
rect 850 32020 860 32090
rect 640 31980 860 32020
rect 640 31910 650 31980
rect 850 31910 860 31980
rect 640 31860 860 31910
rect 1140 32090 1360 32140
rect 1140 32020 1150 32090
rect 1350 32020 1360 32090
rect 1140 31980 1360 32020
rect 1140 31910 1150 31980
rect 1350 31910 1360 31980
rect 1140 31860 1360 31910
rect 1640 32090 1860 32140
rect 1640 32020 1650 32090
rect 1850 32020 1860 32090
rect 1640 31980 1860 32020
rect 1640 31910 1650 31980
rect 1850 31910 1860 31980
rect 1640 31860 1860 31910
rect 2140 32090 2360 32140
rect 2140 32020 2150 32090
rect 2350 32020 2360 32090
rect 2140 31980 2360 32020
rect 2140 31910 2150 31980
rect 2350 31910 2360 31980
rect 2140 31860 2360 31910
rect 2640 32090 2860 32140
rect 2640 32020 2650 32090
rect 2850 32020 2860 32090
rect 2640 31980 2860 32020
rect 2640 31910 2650 31980
rect 2850 31910 2860 31980
rect 2640 31860 2860 31910
rect 3140 32090 3360 32140
rect 3140 32020 3150 32090
rect 3350 32020 3360 32090
rect 3140 31980 3360 32020
rect 3140 31910 3150 31980
rect 3350 31910 3360 31980
rect 3140 31860 3360 31910
rect 3640 32090 3860 32140
rect 3640 32020 3650 32090
rect 3850 32020 3860 32090
rect 3640 31980 3860 32020
rect 3640 31910 3650 31980
rect 3850 31910 3860 31980
rect 3640 31860 3860 31910
rect 4140 32090 4360 32140
rect 4140 32020 4150 32090
rect 4350 32020 4360 32090
rect 4140 31980 4360 32020
rect 4140 31910 4150 31980
rect 4350 31910 4360 31980
rect 4140 31860 4360 31910
rect 4640 32090 4860 32140
rect 4640 32020 4650 32090
rect 4850 32020 4860 32090
rect 4640 31980 4860 32020
rect 4640 31910 4650 31980
rect 4850 31910 4860 31980
rect 4640 31860 4860 31910
rect 5140 32090 5360 32140
rect 5140 32020 5150 32090
rect 5350 32020 5360 32090
rect 5140 31980 5360 32020
rect 5140 31910 5150 31980
rect 5350 31910 5360 31980
rect 5140 31860 5360 31910
rect 5640 32090 5860 32140
rect 5640 32020 5650 32090
rect 5850 32020 5860 32090
rect 5640 31980 5860 32020
rect 5640 31910 5650 31980
rect 5850 31910 5860 31980
rect 5640 31860 5860 31910
rect 6140 32090 6360 32140
rect 6140 32020 6150 32090
rect 6350 32020 6360 32090
rect 6140 31980 6360 32020
rect 6140 31910 6150 31980
rect 6350 31910 6360 31980
rect 6140 31860 6360 31910
rect 6640 32090 6860 32140
rect 6640 32020 6650 32090
rect 6850 32020 6860 32090
rect 6640 31980 6860 32020
rect 6640 31910 6650 31980
rect 6850 31910 6860 31980
rect 6640 31860 6860 31910
rect 7140 32090 7360 32140
rect 7140 32020 7150 32090
rect 7350 32020 7360 32090
rect 7140 31980 7360 32020
rect 7140 31910 7150 31980
rect 7350 31910 7360 31980
rect 7140 31860 7360 31910
rect 7640 32090 7860 32140
rect 7640 32020 7650 32090
rect 7850 32020 7860 32090
rect 7640 31980 7860 32020
rect 7640 31910 7650 31980
rect 7850 31910 7860 31980
rect 7640 31860 7860 31910
rect 8140 32090 8360 32140
rect 8140 32020 8150 32090
rect 8350 32020 8360 32090
rect 8140 31980 8360 32020
rect 8140 31910 8150 31980
rect 8350 31910 8360 31980
rect 8140 31860 8360 31910
rect 8640 32090 8860 32140
rect 8640 32020 8650 32090
rect 8850 32020 8860 32090
rect 8640 31980 8860 32020
rect 8640 31910 8650 31980
rect 8850 31910 8860 31980
rect 8640 31860 8860 31910
rect 9140 32090 9360 32140
rect 9140 32020 9150 32090
rect 9350 32020 9360 32090
rect 9140 31980 9360 32020
rect 9140 31910 9150 31980
rect 9350 31910 9360 31980
rect 9140 31860 9360 31910
rect 9640 32090 9860 32140
rect 9640 32020 9650 32090
rect 9850 32020 9860 32090
rect 9640 31980 9860 32020
rect 9640 31910 9650 31980
rect 9850 31910 9860 31980
rect 9640 31860 9860 31910
rect 10140 32090 10360 32140
rect 10140 32020 10150 32090
rect 10350 32020 10360 32090
rect 10140 31980 10360 32020
rect 10140 31910 10150 31980
rect 10350 31910 10360 31980
rect 10140 31860 10360 31910
rect 10640 32090 10860 32140
rect 10640 32020 10650 32090
rect 10850 32020 10860 32090
rect 10640 31980 10860 32020
rect 10640 31910 10650 31980
rect 10850 31910 10860 31980
rect 10640 31860 10860 31910
rect 11140 32090 11360 32140
rect 11140 32020 11150 32090
rect 11350 32020 11360 32090
rect 11140 31980 11360 32020
rect 11140 31910 11150 31980
rect 11350 31910 11360 31980
rect 11140 31860 11360 31910
rect 11640 32090 11860 32140
rect 11640 32020 11650 32090
rect 11850 32020 11860 32090
rect 11640 31980 11860 32020
rect 11640 31910 11650 31980
rect 11850 31910 11860 31980
rect 11640 31860 11860 31910
rect 12140 32090 12360 32140
rect 12140 32020 12150 32090
rect 12350 32020 12360 32090
rect 12140 31980 12360 32020
rect 12140 31910 12150 31980
rect 12350 31910 12360 31980
rect 12140 31860 12360 31910
rect 12640 32090 12860 32140
rect 12640 32020 12650 32090
rect 12850 32020 12860 32090
rect 12640 31980 12860 32020
rect 12640 31910 12650 31980
rect 12850 31910 12860 31980
rect 12640 31860 12860 31910
rect 13140 32090 13360 32140
rect 13140 32020 13150 32090
rect 13350 32020 13360 32090
rect 13140 31980 13360 32020
rect 13140 31910 13150 31980
rect 13350 31910 13360 31980
rect 13140 31860 13360 31910
rect 13640 32090 13860 32140
rect 13640 32020 13650 32090
rect 13850 32020 13860 32090
rect 13640 31980 13860 32020
rect 13640 31910 13650 31980
rect 13850 31910 13860 31980
rect 13640 31860 13860 31910
rect 14140 32090 14360 32140
rect 14140 32020 14150 32090
rect 14350 32020 14360 32090
rect 14140 31980 14360 32020
rect 14140 31910 14150 31980
rect 14350 31910 14360 31980
rect 14140 31860 14360 31910
rect 14640 32090 14860 32140
rect 14640 32020 14650 32090
rect 14850 32020 14860 32090
rect 14640 31980 14860 32020
rect 14640 31910 14650 31980
rect 14850 31910 14860 31980
rect 14640 31860 14860 31910
rect 15140 32090 15360 32140
rect 15140 32020 15150 32090
rect 15350 32020 15360 32090
rect 15140 31980 15360 32020
rect 15140 31910 15150 31980
rect 15350 31910 15360 31980
rect 15140 31860 15360 31910
rect 15640 32090 15860 32140
rect 15640 32020 15650 32090
rect 15850 32020 15860 32090
rect 15640 31980 15860 32020
rect 15640 31910 15650 31980
rect 15850 31910 15860 31980
rect 15640 31860 15860 31910
rect 16140 32090 16360 32140
rect 16140 32020 16150 32090
rect 16350 32020 16360 32090
rect 16140 31980 16360 32020
rect 16140 31910 16150 31980
rect 16350 31910 16360 31980
rect 16140 31860 16360 31910
rect 16640 32090 16860 32140
rect 16640 32020 16650 32090
rect 16850 32020 16860 32090
rect 16640 31980 16860 32020
rect 16640 31910 16650 31980
rect 16850 31910 16860 31980
rect 16640 31860 16860 31910
rect 17140 32090 17360 32140
rect 17140 32020 17150 32090
rect 17350 32020 17360 32090
rect 17140 31980 17360 32020
rect 17140 31910 17150 31980
rect 17350 31910 17360 31980
rect 17140 31860 17360 31910
rect 17640 32090 17860 32140
rect 17640 32020 17650 32090
rect 17850 32020 17860 32090
rect 17640 31980 17860 32020
rect 17640 31910 17650 31980
rect 17850 31910 17860 31980
rect 17640 31860 17860 31910
rect 18140 32090 18360 32140
rect 18140 32020 18150 32090
rect 18350 32020 18360 32090
rect 18140 31980 18360 32020
rect 18140 31910 18150 31980
rect 18350 31910 18360 31980
rect 18140 31860 18360 31910
rect 18640 32090 18860 32140
rect 18640 32020 18650 32090
rect 18850 32020 18860 32090
rect 18640 31980 18860 32020
rect 18640 31910 18650 31980
rect 18850 31910 18860 31980
rect 18640 31860 18860 31910
rect 19140 32090 19360 32140
rect 19140 32020 19150 32090
rect 19350 32020 19360 32090
rect 19140 31980 19360 32020
rect 19140 31910 19150 31980
rect 19350 31910 19360 31980
rect 19140 31860 19360 31910
rect 19640 32090 19860 32140
rect 19640 32020 19650 32090
rect 19850 32020 19860 32090
rect 19640 31980 19860 32020
rect 19640 31910 19650 31980
rect 19850 31910 19860 31980
rect 19640 31860 19860 31910
rect 20140 32090 20360 32140
rect 20140 32020 20150 32090
rect 20350 32020 20360 32090
rect 20140 31980 20360 32020
rect 20140 31910 20150 31980
rect 20350 31910 20360 31980
rect 20140 31860 20360 31910
rect 20640 32090 20860 32140
rect 20640 32020 20650 32090
rect 20850 32020 20860 32090
rect 20640 31980 20860 32020
rect 20640 31910 20650 31980
rect 20850 31910 20860 31980
rect 20640 31860 20860 31910
rect 21140 32090 21360 32140
rect 21140 32020 21150 32090
rect 21350 32020 21360 32090
rect 21140 31980 21360 32020
rect 21140 31910 21150 31980
rect 21350 31910 21360 31980
rect 21140 31860 21360 31910
rect 21640 32090 21860 32140
rect 21640 32020 21650 32090
rect 21850 32020 21860 32090
rect 21640 31980 21860 32020
rect 21640 31910 21650 31980
rect 21850 31910 21860 31980
rect 21640 31860 21860 31910
rect 22140 32090 22360 32140
rect 22140 32020 22150 32090
rect 22350 32020 22360 32090
rect 22140 31980 22360 32020
rect 22140 31910 22150 31980
rect 22350 31910 22360 31980
rect 22140 31860 22360 31910
rect 22640 32090 22860 32140
rect 22640 32020 22650 32090
rect 22850 32020 22860 32090
rect 22640 31980 22860 32020
rect 22640 31910 22650 31980
rect 22850 31910 22860 31980
rect 22640 31860 22860 31910
rect 23140 32090 23360 32140
rect 23140 32020 23150 32090
rect 23350 32020 23360 32090
rect 23140 31980 23360 32020
rect 23140 31910 23150 31980
rect 23350 31910 23360 31980
rect 23140 31860 23360 31910
rect 23640 32090 23860 32140
rect 23640 32020 23650 32090
rect 23850 32020 23860 32090
rect 23640 31980 23860 32020
rect 23640 31910 23650 31980
rect 23850 31910 23860 31980
rect 23640 31860 23860 31910
rect 24140 32090 24360 32140
rect 24140 32020 24150 32090
rect 24350 32020 24360 32090
rect 24140 31980 24360 32020
rect 24140 31910 24150 31980
rect 24350 31910 24360 31980
rect 24140 31860 24360 31910
rect 24640 32090 24860 32140
rect 24640 32020 24650 32090
rect 24850 32020 24860 32090
rect 24640 31980 24860 32020
rect 24640 31910 24650 31980
rect 24850 31910 24860 31980
rect 24640 31860 24860 31910
rect 25140 32090 25360 32140
rect 25140 32020 25150 32090
rect 25350 32020 25360 32090
rect 25140 31980 25360 32020
rect 25140 31910 25150 31980
rect 25350 31910 25360 31980
rect 25140 31860 25360 31910
rect 25640 32090 25860 32140
rect 25640 32020 25650 32090
rect 25850 32020 25860 32090
rect 25640 31980 25860 32020
rect 25640 31910 25650 31980
rect 25850 31910 25860 31980
rect 25640 31860 25860 31910
rect 26140 32090 26360 32140
rect 26140 32020 26150 32090
rect 26350 32020 26360 32090
rect 26140 31980 26360 32020
rect 26140 31910 26150 31980
rect 26350 31910 26360 31980
rect 26140 31860 26360 31910
rect 0 31850 26500 31860
rect 0 31650 20 31850
rect 90 31650 410 31850
rect 480 31650 520 31850
rect 590 31650 910 31850
rect 980 31650 1020 31850
rect 1090 31650 1410 31850
rect 1480 31650 1520 31850
rect 1590 31650 1910 31850
rect 1980 31650 2020 31850
rect 2090 31650 2410 31850
rect 2480 31650 2520 31850
rect 2590 31650 2910 31850
rect 2980 31650 3020 31850
rect 3090 31650 3410 31850
rect 3480 31650 3520 31850
rect 3590 31650 3910 31850
rect 3980 31650 4020 31850
rect 4090 31650 4410 31850
rect 4480 31650 4520 31850
rect 4590 31650 4910 31850
rect 4980 31650 5020 31850
rect 5090 31650 5410 31850
rect 5480 31650 5520 31850
rect 5590 31650 5910 31850
rect 5980 31650 6020 31850
rect 6090 31650 6410 31850
rect 6480 31650 6520 31850
rect 6590 31650 6910 31850
rect 6980 31650 7020 31850
rect 7090 31650 7410 31850
rect 7480 31650 7520 31850
rect 7590 31650 7910 31850
rect 7980 31650 8020 31850
rect 8090 31650 8410 31850
rect 8480 31650 8520 31850
rect 8590 31650 8910 31850
rect 8980 31650 9020 31850
rect 9090 31650 9410 31850
rect 9480 31650 9520 31850
rect 9590 31650 9910 31850
rect 9980 31650 10020 31850
rect 10090 31650 10410 31850
rect 10480 31650 10520 31850
rect 10590 31650 10910 31850
rect 10980 31650 11020 31850
rect 11090 31650 11410 31850
rect 11480 31650 11520 31850
rect 11590 31650 11910 31850
rect 11980 31650 12020 31850
rect 12090 31650 12410 31850
rect 12480 31650 12520 31850
rect 12590 31650 12910 31850
rect 12980 31650 13020 31850
rect 13090 31650 13410 31850
rect 13480 31650 13520 31850
rect 13590 31650 13910 31850
rect 13980 31650 14020 31850
rect 14090 31650 14410 31850
rect 14480 31650 14520 31850
rect 14590 31650 14910 31850
rect 14980 31650 15020 31850
rect 15090 31650 15410 31850
rect 15480 31650 15520 31850
rect 15590 31650 15910 31850
rect 15980 31650 16020 31850
rect 16090 31650 16410 31850
rect 16480 31650 16520 31850
rect 16590 31650 16910 31850
rect 16980 31650 17020 31850
rect 17090 31650 17410 31850
rect 17480 31650 17520 31850
rect 17590 31650 17910 31850
rect 17980 31650 18020 31850
rect 18090 31650 18410 31850
rect 18480 31650 18520 31850
rect 18590 31650 18910 31850
rect 18980 31650 19020 31850
rect 19090 31650 19410 31850
rect 19480 31650 19520 31850
rect 19590 31650 19910 31850
rect 19980 31650 20020 31850
rect 20090 31650 20410 31850
rect 20480 31650 20520 31850
rect 20590 31650 20910 31850
rect 20980 31650 21020 31850
rect 21090 31650 21410 31850
rect 21480 31650 21520 31850
rect 21590 31650 21910 31850
rect 21980 31650 22020 31850
rect 22090 31650 22410 31850
rect 22480 31650 22520 31850
rect 22590 31650 22910 31850
rect 22980 31650 23020 31850
rect 23090 31650 23410 31850
rect 23480 31650 23520 31850
rect 23590 31650 23910 31850
rect 23980 31650 24020 31850
rect 24090 31650 24410 31850
rect 24480 31650 24520 31850
rect 24590 31650 24910 31850
rect 24980 31650 25020 31850
rect 25090 31650 25410 31850
rect 25480 31650 25520 31850
rect 25590 31650 25910 31850
rect 25980 31650 26020 31850
rect 26090 31650 26410 31850
rect 26480 31650 26500 31850
rect 0 31640 26500 31650
rect 140 31590 360 31640
rect 140 31520 150 31590
rect 350 31520 360 31590
rect 140 31480 360 31520
rect 140 31410 150 31480
rect 350 31410 360 31480
rect 140 31360 360 31410
rect 640 31590 860 31640
rect 640 31520 650 31590
rect 850 31520 860 31590
rect 640 31480 860 31520
rect 1140 31590 1360 31640
rect 1140 31520 1150 31590
rect 1350 31520 1360 31590
rect 1140 31500 1360 31520
rect 1640 31590 1860 31640
rect 1640 31520 1650 31590
rect 1850 31520 1860 31590
rect 1640 31500 1860 31520
rect 2140 31590 2360 31640
rect 2140 31520 2150 31590
rect 2350 31520 2360 31590
rect 2140 31500 2360 31520
rect 2640 31590 2860 31640
rect 2640 31520 2650 31590
rect 2850 31520 2860 31590
rect 2640 31500 2860 31520
rect 3140 31590 3360 31640
rect 3140 31520 3150 31590
rect 3350 31520 3360 31590
rect 3140 31500 3360 31520
rect 3640 31590 3860 31640
rect 3640 31520 3650 31590
rect 3850 31520 3860 31590
rect 3640 31500 3860 31520
rect 4140 31590 4360 31640
rect 4140 31520 4150 31590
rect 4350 31520 4360 31590
rect 4140 31500 4360 31520
rect 4640 31590 4860 31640
rect 4640 31520 4650 31590
rect 4850 31520 4860 31590
rect 4640 31500 4860 31520
rect 5140 31590 5360 31640
rect 5140 31520 5150 31590
rect 5350 31520 5360 31590
rect 5140 31500 5360 31520
rect 5640 31590 5860 31640
rect 5640 31520 5650 31590
rect 5850 31520 5860 31590
rect 5640 31500 5860 31520
rect 6140 31590 6360 31640
rect 6140 31520 6150 31590
rect 6350 31520 6360 31590
rect 6140 31500 6360 31520
rect 6640 31590 6860 31640
rect 6640 31520 6650 31590
rect 6850 31520 6860 31590
rect 640 31410 650 31480
rect 850 31410 860 31480
rect 640 31360 860 31410
rect 6640 31480 6860 31520
rect 6640 31410 6650 31480
rect 6850 31410 6860 31480
rect 6640 31360 6860 31410
rect 7140 31590 7360 31640
rect 7140 31520 7150 31590
rect 7350 31520 7360 31590
rect 7140 31480 7360 31520
rect 7640 31590 7860 31640
rect 7640 31520 7650 31590
rect 7850 31520 7860 31590
rect 7640 31500 7860 31520
rect 8140 31590 8360 31640
rect 8140 31520 8150 31590
rect 8350 31520 8360 31590
rect 8140 31500 8360 31520
rect 8640 31590 8860 31640
rect 8640 31520 8650 31590
rect 8850 31520 8860 31590
rect 8640 31500 8860 31520
rect 9140 31590 9360 31640
rect 9140 31520 9150 31590
rect 9350 31520 9360 31590
rect 9140 31500 9360 31520
rect 9640 31590 9860 31640
rect 9640 31520 9650 31590
rect 9850 31520 9860 31590
rect 9640 31500 9860 31520
rect 10140 31590 10360 31640
rect 10140 31520 10150 31590
rect 10350 31520 10360 31590
rect 10140 31500 10360 31520
rect 10640 31590 10860 31640
rect 10640 31520 10650 31590
rect 10850 31520 10860 31590
rect 10640 31500 10860 31520
rect 11140 31590 11360 31640
rect 11140 31520 11150 31590
rect 11350 31520 11360 31590
rect 11140 31500 11360 31520
rect 11640 31590 11860 31640
rect 11640 31520 11650 31590
rect 11850 31520 11860 31590
rect 11640 31500 11860 31520
rect 12140 31590 12360 31640
rect 12140 31520 12150 31590
rect 12350 31520 12360 31590
rect 12140 31500 12360 31520
rect 12640 31590 12860 31640
rect 12640 31520 12650 31590
rect 12850 31520 12860 31590
rect 12640 31500 12860 31520
rect 13140 31590 13360 31640
rect 13140 31520 13150 31590
rect 13350 31520 13360 31590
rect 7140 31410 7150 31480
rect 7350 31410 7360 31480
rect 7140 31360 7360 31410
rect 13140 31480 13360 31520
rect 13640 31590 13860 31640
rect 13640 31520 13650 31590
rect 13850 31520 13860 31590
rect 13640 31500 13860 31520
rect 14140 31590 14360 31640
rect 14140 31520 14150 31590
rect 14350 31520 14360 31590
rect 14140 31500 14360 31520
rect 14640 31590 14860 31640
rect 14640 31520 14650 31590
rect 14850 31520 14860 31590
rect 14640 31500 14860 31520
rect 15140 31590 15360 31640
rect 15140 31520 15150 31590
rect 15350 31520 15360 31590
rect 15140 31500 15360 31520
rect 15640 31590 15860 31640
rect 15640 31520 15650 31590
rect 15850 31520 15860 31590
rect 15640 31500 15860 31520
rect 16140 31590 16360 31640
rect 16140 31520 16150 31590
rect 16350 31520 16360 31590
rect 16140 31500 16360 31520
rect 16640 31590 16860 31640
rect 16640 31520 16650 31590
rect 16850 31520 16860 31590
rect 16640 31500 16860 31520
rect 17140 31590 17360 31640
rect 17140 31520 17150 31590
rect 17350 31520 17360 31590
rect 17140 31500 17360 31520
rect 17640 31590 17860 31640
rect 17640 31520 17650 31590
rect 17850 31520 17860 31590
rect 17640 31500 17860 31520
rect 18140 31590 18360 31640
rect 18140 31520 18150 31590
rect 18350 31520 18360 31590
rect 18140 31500 18360 31520
rect 18640 31590 18860 31640
rect 18640 31520 18650 31590
rect 18850 31520 18860 31590
rect 18640 31500 18860 31520
rect 19140 31590 19360 31640
rect 19140 31520 19150 31590
rect 19350 31520 19360 31590
rect 19140 31500 19360 31520
rect 19640 31590 19860 31640
rect 19640 31520 19650 31590
rect 19850 31520 19860 31590
rect 13140 31410 13150 31480
rect 13350 31410 13360 31480
rect 13140 31360 13360 31410
rect 19640 31480 19860 31520
rect 20140 31590 20360 31640
rect 20140 31520 20150 31590
rect 20350 31520 20360 31590
rect 20140 31500 20360 31520
rect 20640 31590 20860 31640
rect 20640 31520 20650 31590
rect 20850 31520 20860 31590
rect 20640 31500 20860 31520
rect 21140 31590 21360 31640
rect 21140 31520 21150 31590
rect 21350 31520 21360 31590
rect 21140 31500 21360 31520
rect 21640 31590 21860 31640
rect 21640 31520 21650 31590
rect 21850 31520 21860 31590
rect 21640 31500 21860 31520
rect 22140 31590 22360 31640
rect 22140 31520 22150 31590
rect 22350 31520 22360 31590
rect 22140 31500 22360 31520
rect 22640 31590 22860 31640
rect 22640 31520 22650 31590
rect 22850 31520 22860 31590
rect 22640 31500 22860 31520
rect 23140 31590 23360 31640
rect 23140 31520 23150 31590
rect 23350 31520 23360 31590
rect 23140 31500 23360 31520
rect 23640 31590 23860 31640
rect 23640 31520 23650 31590
rect 23850 31520 23860 31590
rect 23640 31500 23860 31520
rect 24140 31590 24360 31640
rect 24140 31520 24150 31590
rect 24350 31520 24360 31590
rect 24140 31500 24360 31520
rect 24640 31590 24860 31640
rect 24640 31520 24650 31590
rect 24850 31520 24860 31590
rect 24640 31500 24860 31520
rect 25140 31590 25360 31640
rect 25140 31520 25150 31590
rect 25350 31520 25360 31590
rect 25140 31500 25360 31520
rect 25640 31590 25860 31640
rect 25640 31520 25650 31590
rect 25850 31520 25860 31590
rect 19640 31410 19650 31480
rect 19850 31410 19860 31480
rect 19640 31360 19860 31410
rect 25640 31480 25860 31520
rect 25640 31410 25650 31480
rect 25850 31410 25860 31480
rect 25640 31360 25860 31410
rect 26140 31590 26360 31640
rect 26140 31520 26150 31590
rect 26350 31520 26360 31590
rect 26140 31480 26360 31520
rect 26140 31410 26150 31480
rect 26350 31410 26360 31480
rect 26140 31360 26360 31410
rect 0 31350 1000 31360
rect 0 31150 20 31350
rect 90 31150 410 31350
rect 480 31150 520 31350
rect 590 31150 910 31350
rect 980 31150 1000 31350
rect 0 31140 1000 31150
rect 6500 31350 7500 31360
rect 6500 31150 6520 31350
rect 6590 31150 6910 31350
rect 6980 31150 7020 31350
rect 7090 31150 7410 31350
rect 7480 31150 7500 31350
rect 6500 31140 7500 31150
rect 13000 31350 13500 31360
rect 13000 31150 13020 31350
rect 13090 31150 13410 31350
rect 13480 31150 13500 31350
rect 13000 31140 13500 31150
rect 19500 31350 20000 31360
rect 19500 31150 19520 31350
rect 19590 31150 19910 31350
rect 19980 31150 20000 31350
rect 19500 31140 20000 31150
rect 25500 31350 26500 31360
rect 25500 31150 25520 31350
rect 25590 31150 25910 31350
rect 25980 31150 26020 31350
rect 26090 31150 26410 31350
rect 26480 31150 26500 31350
rect 25500 31140 26500 31150
rect 140 31090 360 31140
rect 140 31020 150 31090
rect 350 31020 360 31090
rect 140 30980 360 31020
rect 140 30910 150 30980
rect 350 30910 360 30980
rect 140 30860 360 30910
rect 640 31090 860 31140
rect 640 31020 650 31090
rect 850 31020 860 31090
rect 640 30980 860 31020
rect 640 30910 650 30980
rect 850 30910 860 30980
rect 640 30860 860 30910
rect 6640 31090 6860 31140
rect 6640 31020 6650 31090
rect 6850 31020 6860 31090
rect 6640 30980 6860 31020
rect 6640 30910 6650 30980
rect 6850 30910 6860 30980
rect 6640 30900 6860 30910
rect 7140 31090 7360 31140
rect 7140 31020 7150 31090
rect 7350 31020 7360 31090
rect 7140 30980 7360 31020
rect 13140 31090 13360 31140
rect 13140 31020 13150 31090
rect 13350 31020 13360 31090
rect 13140 31000 13360 31020
rect 19640 31090 19860 31140
rect 19640 31020 19650 31090
rect 19850 31020 19860 31090
rect 7140 30910 7150 30980
rect 7350 30910 7360 30980
rect 7140 30900 7360 30910
rect 6400 30880 7700 30900
rect 12700 30880 14000 31000
rect 19640 30980 19860 31020
rect 19640 30910 19650 30980
rect 19850 30910 19860 30980
rect 19640 30900 19860 30910
rect 25640 31090 25860 31140
rect 25640 31020 25650 31090
rect 25850 31020 25860 31090
rect 25640 30980 25860 31020
rect 25640 30910 25650 30980
rect 25850 30910 25860 30980
rect 19000 30880 20300 30900
rect 0 30850 1000 30860
rect 0 30650 20 30850
rect 90 30650 410 30850
rect 480 30650 520 30850
rect 590 30650 910 30850
rect 980 30650 1000 30850
rect 0 30640 1000 30650
rect 1330 30820 1400 30880
rect 140 30590 360 30640
rect 140 30520 150 30590
rect 350 30520 360 30590
rect 140 30480 360 30520
rect 140 30410 150 30480
rect 350 30410 360 30480
rect 140 30360 360 30410
rect 640 30590 860 30640
rect 640 30520 650 30590
rect 850 30520 860 30590
rect 640 30480 860 30520
rect 640 30410 650 30480
rect 850 30410 860 30480
rect 640 30360 860 30410
rect 0 30350 1000 30360
rect 0 30150 20 30350
rect 90 30150 410 30350
rect 480 30150 520 30350
rect 590 30150 910 30350
rect 980 30150 1000 30350
rect 0 30140 1000 30150
rect 140 30090 360 30140
rect 140 30020 150 30090
rect 350 30020 360 30090
rect 140 29980 360 30020
rect 140 29910 150 29980
rect 350 29910 360 29980
rect 140 29860 360 29910
rect 640 30090 860 30140
rect 640 30020 650 30090
rect 850 30020 860 30090
rect 640 29980 860 30020
rect 640 29910 650 29980
rect 850 29910 860 29980
rect 640 29860 860 29910
rect 0 29850 1000 29860
rect 0 29650 20 29850
rect 90 29650 410 29850
rect 480 29650 520 29850
rect 590 29650 910 29850
rect 980 29650 1000 29850
rect 0 29640 1000 29650
rect 140 29590 360 29640
rect 140 29520 150 29590
rect 350 29520 360 29590
rect 140 29480 360 29520
rect 140 29410 150 29480
rect 350 29410 360 29480
rect 140 29360 360 29410
rect 640 29590 860 29640
rect 640 29520 650 29590
rect 850 29520 860 29590
rect 640 29480 860 29520
rect 640 29410 650 29480
rect 850 29410 860 29480
rect 640 29360 860 29410
rect 0 29350 1000 29360
rect 0 29150 20 29350
rect 90 29150 410 29350
rect 480 29150 520 29350
rect 590 29150 910 29350
rect 980 29150 1000 29350
rect 0 29140 1000 29150
rect 140 29090 360 29140
rect 140 29020 150 29090
rect 350 29020 360 29090
rect 140 28980 360 29020
rect 140 28910 150 28980
rect 350 28910 360 28980
rect 140 28860 360 28910
rect 640 29090 860 29140
rect 640 29020 650 29090
rect 850 29020 860 29090
rect 640 28980 860 29020
rect 640 28910 650 28980
rect 850 28910 860 28980
rect 640 28860 860 28910
rect 0 28850 1000 28860
rect 0 28650 20 28850
rect 90 28650 410 28850
rect 480 28650 520 28850
rect 590 28650 910 28850
rect 980 28650 1000 28850
rect 0 28640 1000 28650
rect 140 28590 360 28640
rect 140 28520 150 28590
rect 350 28520 360 28590
rect 140 28480 360 28520
rect 140 28410 150 28480
rect 350 28410 360 28480
rect 140 28360 360 28410
rect 640 28590 860 28640
rect 640 28520 650 28590
rect 850 28520 860 28590
rect 640 28480 860 28520
rect 640 28410 650 28480
rect 850 28410 860 28480
rect 640 28360 860 28410
rect 0 28350 1000 28360
rect 0 28150 20 28350
rect 90 28150 410 28350
rect 480 28150 520 28350
rect 590 28150 910 28350
rect 980 28150 1000 28350
rect 0 28140 1000 28150
rect 140 28090 360 28140
rect 140 28020 150 28090
rect 350 28020 360 28090
rect 140 27980 360 28020
rect 140 27910 150 27980
rect 350 27910 360 27980
rect 140 27860 360 27910
rect 640 28090 860 28140
rect 640 28020 650 28090
rect 850 28020 860 28090
rect 640 27980 860 28020
rect 640 27910 650 27980
rect 850 27910 860 27980
rect 640 27860 860 27910
rect 0 27850 1000 27860
rect 0 27650 20 27850
rect 90 27650 410 27850
rect 480 27650 520 27850
rect 590 27650 910 27850
rect 980 27650 1000 27850
rect 0 27640 1000 27650
rect 140 27590 360 27640
rect 140 27520 150 27590
rect 350 27520 360 27590
rect 140 27480 360 27520
rect 140 27410 150 27480
rect 350 27410 360 27480
rect 140 27360 360 27410
rect 640 27590 860 27640
rect 640 27520 650 27590
rect 850 27520 860 27590
rect 640 27480 860 27520
rect 640 27410 650 27480
rect 850 27410 860 27480
rect 640 27360 860 27410
rect 0 27350 1000 27360
rect -4300 27250 -4100 27260
rect -4300 27030 -4290 27250
rect -4110 27030 -4100 27250
rect 0 27150 20 27350
rect 90 27150 410 27350
rect 480 27150 520 27350
rect 590 27150 910 27350
rect 980 27150 1000 27350
rect 0 27140 1000 27150
rect -4300 27020 -4100 27030
rect 140 27090 360 27140
rect 140 27020 150 27090
rect 350 27020 360 27090
rect -3860 26980 -3640 27000
rect -3860 26910 -3850 26980
rect -3650 26910 -3640 26980
rect -3860 26860 -3640 26910
rect -3360 26980 -3140 27000
rect -3360 26910 -3350 26980
rect -3150 26910 -3140 26980
rect -3360 26860 -3140 26910
rect -2860 26980 -2640 27000
rect -2860 26910 -2850 26980
rect -2650 26910 -2640 26980
rect -2860 26860 -2640 26910
rect -2360 26980 -2140 27000
rect -2360 26910 -2350 26980
rect -2150 26910 -2140 26980
rect -2360 26860 -2140 26910
rect -1860 26980 -1640 27000
rect -1860 26910 -1850 26980
rect -1650 26910 -1640 26980
rect -1860 26860 -1640 26910
rect -1360 26980 -1140 27000
rect -1360 26910 -1350 26980
rect -1150 26910 -1140 26980
rect -1360 26860 -1140 26910
rect -860 26980 -640 27000
rect -860 26910 -850 26980
rect -650 26910 -640 26980
rect -860 26860 -640 26910
rect -360 26980 -140 27000
rect -360 26910 -350 26980
rect -150 26910 -140 26980
rect -360 26860 -140 26910
rect 140 26980 360 27020
rect 140 26910 150 26980
rect 350 26910 360 26980
rect 140 26860 360 26910
rect 640 27090 860 27140
rect 640 27020 650 27090
rect 850 27020 860 27090
rect 640 26980 860 27020
rect 640 26910 650 26980
rect 850 26910 860 26980
rect 640 26860 860 26910
rect -4000 26850 1000 26860
rect -4000 26650 -3980 26850
rect -3910 26650 -3590 26850
rect -3520 26650 -3480 26850
rect -3410 26650 -3090 26850
rect -3020 26650 -2980 26850
rect -2910 26650 -2590 26850
rect -2520 26650 -2480 26850
rect -2410 26650 -2090 26850
rect -2020 26650 -1980 26850
rect -1910 26650 -1590 26850
rect -1520 26650 -1480 26850
rect -1410 26650 -1090 26850
rect -1020 26650 -980 26850
rect -910 26650 -590 26850
rect -520 26650 -480 26850
rect -410 26650 -90 26850
rect -20 26650 20 26850
rect 90 26650 410 26850
rect 480 26650 520 26850
rect 590 26650 910 26850
rect 980 26650 1000 26850
rect -4000 26640 1000 26650
rect -3860 26590 -3640 26640
rect -3860 26520 -3850 26590
rect -3650 26520 -3640 26590
rect -3860 26480 -3640 26520
rect -3860 26410 -3850 26480
rect -3650 26410 -3640 26480
rect -3860 26360 -3640 26410
rect -3360 26590 -3140 26640
rect -3360 26520 -3350 26590
rect -3150 26520 -3140 26590
rect -3360 26480 -3140 26520
rect -3360 26410 -3350 26480
rect -3150 26410 -3140 26480
rect -3360 26360 -3140 26410
rect -2860 26590 -2640 26640
rect -2860 26520 -2850 26590
rect -2650 26520 -2640 26590
rect -2860 26480 -2640 26520
rect -2860 26410 -2850 26480
rect -2650 26410 -2640 26480
rect -2860 26360 -2640 26410
rect -2360 26590 -2140 26640
rect -2360 26520 -2350 26590
rect -2150 26520 -2140 26590
rect -2360 26480 -2140 26520
rect -2360 26410 -2350 26480
rect -2150 26410 -2140 26480
rect -2360 26360 -2140 26410
rect -1860 26590 -1640 26640
rect -1860 26520 -1850 26590
rect -1650 26520 -1640 26590
rect -1860 26480 -1640 26520
rect -1860 26410 -1850 26480
rect -1650 26410 -1640 26480
rect -1860 26360 -1640 26410
rect -1360 26590 -1140 26640
rect -1360 26520 -1350 26590
rect -1150 26520 -1140 26590
rect -1360 26480 -1140 26520
rect -1360 26410 -1350 26480
rect -1150 26410 -1140 26480
rect -1360 26360 -1140 26410
rect -860 26590 -640 26640
rect -860 26520 -850 26590
rect -650 26520 -640 26590
rect -860 26480 -640 26520
rect -860 26410 -850 26480
rect -650 26410 -640 26480
rect -860 26360 -640 26410
rect -360 26590 -140 26640
rect -360 26520 -350 26590
rect -150 26520 -140 26590
rect -360 26480 -140 26520
rect -360 26410 -350 26480
rect -150 26410 -140 26480
rect -360 26360 -140 26410
rect 140 26590 360 26640
rect 140 26520 150 26590
rect 350 26520 360 26590
rect 140 26480 360 26520
rect 140 26410 150 26480
rect 350 26410 360 26480
rect 140 26360 360 26410
rect 640 26590 860 26640
rect 640 26520 650 26590
rect 850 26520 860 26590
rect 640 26480 860 26520
rect 640 26410 650 26480
rect 850 26410 860 26480
rect 640 26360 860 26410
rect -4000 26350 1000 26360
rect -4000 26150 -3980 26350
rect -3910 26150 -3590 26350
rect -3520 26150 -3480 26350
rect -3410 26150 -3090 26350
rect -3020 26150 -2980 26350
rect -2910 26150 -2590 26350
rect -2520 26150 -2480 26350
rect -2410 26150 -2090 26350
rect -2020 26150 -1980 26350
rect -1910 26150 -1590 26350
rect -1520 26150 -1480 26350
rect -1410 26150 -1090 26350
rect -1020 26150 -980 26350
rect -910 26150 -590 26350
rect -520 26150 -480 26350
rect -410 26150 -90 26350
rect -20 26150 20 26350
rect 90 26150 410 26350
rect 480 26150 520 26350
rect 590 26150 910 26350
rect 980 26150 1000 26350
rect -4000 26140 1000 26150
rect -3860 26090 -3640 26140
rect -3860 26020 -3850 26090
rect -3650 26020 -3640 26090
rect -3860 26000 -3640 26020
rect -3360 26090 -3140 26140
rect -3360 26020 -3350 26090
rect -3150 26020 -3140 26090
rect -3360 26000 -3140 26020
rect -2860 26090 -2640 26140
rect -2860 26020 -2850 26090
rect -2650 26020 -2640 26090
rect -2860 26000 -2640 26020
rect -2360 26090 -2140 26140
rect -2360 26020 -2350 26090
rect -2150 26020 -2140 26090
rect -2360 26000 -2140 26020
rect -1860 26090 -1640 26140
rect -1860 26020 -1850 26090
rect -1650 26020 -1640 26090
rect -1860 26000 -1640 26020
rect -1360 26090 -1140 26140
rect -1360 26020 -1350 26090
rect -1150 26020 -1140 26090
rect -1360 26000 -1140 26020
rect -860 26090 -640 26140
rect -860 26020 -850 26090
rect -650 26020 -640 26090
rect -860 26000 -640 26020
rect -360 26090 -140 26140
rect -360 26020 -350 26090
rect -150 26020 -140 26090
rect -360 26000 -140 26020
rect 140 26090 360 26140
rect 140 26020 150 26090
rect 350 26020 360 26090
rect 140 25980 360 26020
rect 140 25910 150 25980
rect 350 25910 360 25980
rect 140 25860 360 25910
rect 640 26090 860 26140
rect 640 26020 650 26090
rect 850 26020 860 26090
rect 640 25980 860 26020
rect 640 25910 650 25980
rect 850 25910 860 25980
rect 640 25860 860 25910
rect 0 25850 1000 25860
rect -4300 25710 -4100 25720
rect -4300 25490 -4290 25710
rect -4110 25490 -4100 25710
rect 0 25650 20 25850
rect 90 25650 410 25850
rect 480 25650 520 25850
rect 590 25650 910 25850
rect 980 25650 1000 25850
rect 0 25640 1000 25650
rect -4300 25480 -4100 25490
rect 140 25590 360 25640
rect 140 25520 150 25590
rect 350 25520 360 25590
rect 140 25480 360 25520
rect 140 25410 150 25480
rect 350 25410 360 25480
rect 140 25360 360 25410
rect 640 25590 860 25640
rect 640 25520 650 25590
rect 850 25520 860 25590
rect 640 25480 860 25520
rect 640 25410 650 25480
rect 850 25410 860 25480
rect 640 25360 860 25410
rect 0 25350 1000 25360
rect 0 25150 20 25350
rect 90 25150 410 25350
rect 480 25150 520 25350
rect 590 25150 910 25350
rect 980 25150 1000 25350
rect 0 25140 1000 25150
rect 140 25090 360 25140
rect 140 25020 150 25090
rect 350 25020 360 25090
rect 140 24980 360 25020
rect 140 24910 150 24980
rect 350 24910 360 24980
rect 140 24860 360 24910
rect 640 25090 860 25140
rect 640 25020 650 25090
rect 850 25020 860 25090
rect 640 24980 860 25020
rect 640 24910 650 24980
rect 850 24910 860 24980
rect 640 24860 860 24910
rect 0 24850 1000 24860
rect 0 24650 20 24850
rect 90 24650 410 24850
rect 480 24650 520 24850
rect 590 24650 910 24850
rect 980 24650 1000 24850
rect 0 24640 1000 24650
rect 140 24590 360 24640
rect 140 24520 150 24590
rect 350 24520 360 24590
rect 140 24480 360 24520
rect 140 24410 150 24480
rect 350 24410 360 24480
rect 140 24360 360 24410
rect 640 24590 860 24640
rect 640 24520 650 24590
rect 850 24520 860 24590
rect 640 24480 860 24520
rect 640 24410 650 24480
rect 850 24410 860 24480
rect 6340 30850 7700 30880
rect 6340 30820 6520 30850
rect 1532 30780 1552 30790
rect 6186 30780 6206 30790
rect 1532 30710 1540 30780
rect 6200 30710 6206 30780
rect 1532 30690 1552 30710
rect 6186 30690 6206 30710
rect 1465 30638 1531 30658
rect 1465 24658 1531 24678
rect 1623 30638 1689 30658
rect 1623 24658 1689 24678
rect 1781 30638 1847 30658
rect 1781 24658 1847 24678
rect 1939 30638 2005 30658
rect 1939 24658 2005 24678
rect 2097 30638 2163 30658
rect 2097 24658 2163 24678
rect 2255 30638 2321 30658
rect 2255 24658 2321 24678
rect 2413 30638 2479 30658
rect 2413 24658 2479 24678
rect 2571 30638 2637 30658
rect 2571 24658 2637 24678
rect 2729 30638 2795 30658
rect 2729 24658 2795 24678
rect 2887 30638 2953 30658
rect 2887 24658 2953 24678
rect 3045 30638 3111 30658
rect 3045 24658 3111 24678
rect 3203 30638 3269 30658
rect 3203 24658 3269 24678
rect 3361 30638 3427 30658
rect 3361 24658 3427 24678
rect 3519 30638 3585 30658
rect 3519 24658 3585 24678
rect 3677 30638 3743 30658
rect 3677 24658 3743 24678
rect 3835 30638 3901 30658
rect 3835 24658 3901 24678
rect 3993 30638 4059 30658
rect 3993 24658 4059 24678
rect 4151 30638 4217 30658
rect 4151 24658 4217 24678
rect 4309 30638 4375 30658
rect 4309 24658 4375 24678
rect 4467 30638 4533 30658
rect 4467 24658 4533 24678
rect 4625 30638 4691 30658
rect 4625 24658 4691 24678
rect 4783 30638 4849 30658
rect 4783 24658 4849 24678
rect 4941 30638 5007 30658
rect 4941 24658 5007 24678
rect 5099 30638 5165 30658
rect 5099 24658 5165 24678
rect 5257 30638 5323 30658
rect 5257 24658 5323 24678
rect 5415 30638 5481 30658
rect 5415 24658 5481 24678
rect 5573 30638 5639 30658
rect 5573 24658 5639 24678
rect 5731 30638 5797 30658
rect 5731 24658 5797 24678
rect 5889 30638 5955 30658
rect 5889 24658 5955 24678
rect 6047 30638 6113 30658
rect 6047 24658 6113 24678
rect 6205 30638 6271 30658
rect 6205 24658 6271 24678
rect 1532 24610 1552 24626
rect 6186 24610 6206 24626
rect 1532 24540 1540 24610
rect 6190 24540 6206 24610
rect 1532 24526 1552 24540
rect 6186 24526 6206 24540
rect 1330 24430 1400 24500
rect 6410 30650 6520 30820
rect 6590 30650 6910 30850
rect 6980 30650 7020 30850
rect 7090 30650 7410 30850
rect 7480 30820 7700 30850
rect 7480 30650 7630 30820
rect 6410 30590 7630 30650
rect 6410 30520 6650 30590
rect 6850 30520 7150 30590
rect 7350 30520 7630 30590
rect 6410 30500 7630 30520
rect 6410 29900 7630 30300
rect 6410 29300 7630 29700
rect 6410 28700 7630 29100
rect 6410 28100 7630 28500
rect 6410 27500 7630 27900
rect 6410 26900 7630 27300
rect 6410 26300 7630 26700
rect 6410 25700 7630 26100
rect 6410 25100 7630 25500
rect 6410 24500 7630 24900
rect 12640 30820 14000 30880
rect 7832 30780 7852 30790
rect 12486 30780 12506 30790
rect 7832 30710 7840 30780
rect 12500 30710 12506 30780
rect 7832 30690 7852 30710
rect 12486 30690 12506 30710
rect 7765 30638 7831 30658
rect 7765 24658 7831 24678
rect 7923 30638 7989 30658
rect 7923 24658 7989 24678
rect 8081 30638 8147 30658
rect 8081 24658 8147 24678
rect 8239 30638 8305 30658
rect 8239 24658 8305 24678
rect 8397 30638 8463 30658
rect 8397 24658 8463 24678
rect 8555 30638 8621 30658
rect 8555 24658 8621 24678
rect 8713 30638 8779 30658
rect 8713 24658 8779 24678
rect 8871 30638 8937 30658
rect 8871 24658 8937 24678
rect 9029 30638 9095 30658
rect 9029 24658 9095 24678
rect 9187 30638 9253 30658
rect 9187 24658 9253 24678
rect 9345 30638 9411 30658
rect 9345 24658 9411 24678
rect 9503 30638 9569 30658
rect 9503 24658 9569 24678
rect 9661 30638 9727 30658
rect 9661 24658 9727 24678
rect 9819 30638 9885 30658
rect 9819 24658 9885 24678
rect 9977 30638 10043 30658
rect 9977 24658 10043 24678
rect 10135 30638 10201 30658
rect 10135 24658 10201 24678
rect 10293 30638 10359 30658
rect 10293 24658 10359 24678
rect 10451 30638 10517 30658
rect 10451 24658 10517 24678
rect 10609 30638 10675 30658
rect 10609 24658 10675 24678
rect 10767 30638 10833 30658
rect 10767 24658 10833 24678
rect 10925 30638 10991 30658
rect 10925 24658 10991 24678
rect 11083 30638 11149 30658
rect 11083 24658 11149 24678
rect 11241 30638 11307 30658
rect 11241 24658 11307 24678
rect 11399 30638 11465 30658
rect 11399 24658 11465 24678
rect 11557 30638 11623 30658
rect 11557 24658 11623 24678
rect 11715 30638 11781 30658
rect 11715 24658 11781 24678
rect 11873 30638 11939 30658
rect 11873 24658 11939 24678
rect 12031 30638 12097 30658
rect 12031 24658 12097 24678
rect 12189 30638 12255 30658
rect 12189 24658 12255 24678
rect 12347 30638 12413 30658
rect 12347 24658 12413 24678
rect 12505 30638 12571 30658
rect 12505 24658 12571 24678
rect 7832 24610 7852 24626
rect 12486 24610 12506 24626
rect 7832 24540 7840 24610
rect 12490 24540 12506 24610
rect 7832 24526 7852 24540
rect 12486 24526 12506 24540
rect 6340 24430 6410 24500
rect 640 24360 860 24410
rect 0 24350 1000 24360
rect 0 24150 20 24350
rect 90 24150 410 24350
rect 480 24150 520 24350
rect 590 24150 910 24350
rect 980 24150 1000 24350
rect 0 24140 1000 24150
rect 140 24090 360 24140
rect 140 24020 150 24090
rect 350 24020 360 24090
rect 140 23980 360 24020
rect 140 23910 150 23980
rect 350 23910 360 23980
rect 140 23860 360 23910
rect 640 24090 860 24140
rect 640 24020 650 24090
rect 850 24020 860 24090
rect 640 23980 860 24020
rect 640 23910 650 23980
rect 850 23910 860 23980
rect 640 23860 860 23910
rect 6800 23900 7300 24500
rect 7630 24430 7700 24500
rect 12710 30600 13930 30820
rect 12710 30000 13930 30400
rect 12710 29400 13930 29800
rect 12710 28800 13930 29200
rect 12710 28200 13930 28600
rect 12710 27600 13930 28000
rect 12710 27000 13930 27400
rect 12710 26400 13930 26800
rect 12710 25800 13930 26200
rect 12710 25200 13930 25600
rect 12710 24600 13930 25000
rect 12640 24430 12710 24500
rect 13100 23900 13600 24600
rect 18940 30850 20300 30880
rect 18940 30820 19520 30850
rect 14132 30780 14152 30790
rect 18786 30780 18806 30790
rect 14132 30710 14140 30780
rect 18800 30710 18806 30780
rect 14132 30690 14152 30710
rect 18786 30690 18806 30710
rect 14065 30638 14131 30658
rect 14065 24658 14131 24678
rect 14223 30638 14289 30658
rect 14223 24658 14289 24678
rect 14381 30638 14447 30658
rect 14381 24658 14447 24678
rect 14539 30638 14605 30658
rect 14539 24658 14605 24678
rect 14697 30638 14763 30658
rect 14697 24658 14763 24678
rect 14855 30638 14921 30658
rect 14855 24658 14921 24678
rect 15013 30638 15079 30658
rect 15013 24658 15079 24678
rect 15171 30638 15237 30658
rect 15171 24658 15237 24678
rect 15329 30638 15395 30658
rect 15329 24658 15395 24678
rect 15487 30638 15553 30658
rect 15487 24658 15553 24678
rect 15645 30638 15711 30658
rect 15645 24658 15711 24678
rect 15803 30638 15869 30658
rect 15803 24658 15869 24678
rect 15961 30638 16027 30658
rect 15961 24658 16027 24678
rect 16119 30638 16185 30658
rect 16119 24658 16185 24678
rect 16277 30638 16343 30658
rect 16277 24658 16343 24678
rect 16435 30638 16501 30658
rect 16435 24658 16501 24678
rect 16593 30638 16659 30658
rect 16593 24658 16659 24678
rect 16751 30638 16817 30658
rect 16751 24658 16817 24678
rect 16909 30638 16975 30658
rect 16909 24658 16975 24678
rect 17067 30638 17133 30658
rect 17067 24658 17133 24678
rect 17225 30638 17291 30658
rect 17225 24658 17291 24678
rect 17383 30638 17449 30658
rect 17383 24658 17449 24678
rect 17541 30638 17607 30658
rect 17541 24658 17607 24678
rect 17699 30638 17765 30658
rect 17699 24658 17765 24678
rect 17857 30638 17923 30658
rect 17857 24658 17923 24678
rect 18015 30638 18081 30658
rect 18015 24658 18081 24678
rect 18173 30638 18239 30658
rect 18173 24658 18239 24678
rect 18331 30638 18397 30658
rect 18331 24658 18397 24678
rect 18489 30638 18555 30658
rect 18489 24658 18555 24678
rect 18647 30638 18713 30658
rect 18647 24658 18713 24678
rect 18805 30638 18871 30658
rect 18805 24658 18871 24678
rect 14132 24610 14152 24626
rect 18786 24610 18806 24626
rect 14132 24540 14140 24610
rect 18790 24540 18806 24610
rect 14132 24526 14152 24540
rect 18786 24526 18806 24540
rect 13930 24430 14000 24500
rect 19010 30650 19520 30820
rect 19590 30650 19910 30850
rect 19980 30820 20300 30850
rect 19980 30650 20230 30820
rect 19010 30590 20230 30650
rect 19010 30520 19650 30590
rect 19850 30520 20230 30590
rect 19010 30500 20230 30520
rect 19010 29900 20230 30300
rect 19010 29300 20230 29700
rect 19010 28700 20230 29100
rect 19010 28100 20230 28500
rect 19010 27500 20230 27900
rect 19010 26900 20230 27300
rect 19010 26300 20230 26700
rect 19010 25700 20230 26100
rect 19010 25100 20230 25500
rect 19010 24500 20230 24900
rect 25240 30820 25310 30880
rect 25640 30860 25860 30910
rect 26140 31090 26360 31140
rect 26140 31020 26150 31090
rect 26350 31020 26360 31090
rect 26140 30980 26360 31020
rect 26140 30910 26150 30980
rect 26350 30910 26360 30980
rect 26140 30860 26360 30910
rect 20432 30780 20452 30790
rect 25086 30780 25106 30790
rect 20432 30710 20440 30780
rect 25100 30710 25106 30780
rect 20432 30690 20452 30710
rect 25086 30690 25106 30710
rect 20365 30638 20431 30658
rect 20365 24658 20431 24678
rect 20523 30638 20589 30658
rect 20523 24658 20589 24678
rect 20681 30638 20747 30658
rect 20681 24658 20747 24678
rect 20839 30638 20905 30658
rect 20839 24658 20905 24678
rect 20997 30638 21063 30658
rect 20997 24658 21063 24678
rect 21155 30638 21221 30658
rect 21155 24658 21221 24678
rect 21313 30638 21379 30658
rect 21313 24658 21379 24678
rect 21471 30638 21537 30658
rect 21471 24658 21537 24678
rect 21629 30638 21695 30658
rect 21629 24658 21695 24678
rect 21787 30638 21853 30658
rect 21787 24658 21853 24678
rect 21945 30638 22011 30658
rect 21945 24658 22011 24678
rect 22103 30638 22169 30658
rect 22103 24658 22169 24678
rect 22261 30638 22327 30658
rect 22261 24658 22327 24678
rect 22419 30638 22485 30658
rect 22419 24658 22485 24678
rect 22577 30638 22643 30658
rect 22577 24658 22643 24678
rect 22735 30638 22801 30658
rect 22735 24658 22801 24678
rect 22893 30638 22959 30658
rect 22893 24658 22959 24678
rect 23051 30638 23117 30658
rect 23051 24658 23117 24678
rect 23209 30638 23275 30658
rect 23209 24658 23275 24678
rect 23367 30638 23433 30658
rect 23367 24658 23433 24678
rect 23525 30638 23591 30658
rect 23525 24658 23591 24678
rect 23683 30638 23749 30658
rect 23683 24658 23749 24678
rect 23841 30638 23907 30658
rect 23841 24658 23907 24678
rect 23999 30638 24065 30658
rect 23999 24658 24065 24678
rect 24157 30638 24223 30658
rect 24157 24658 24223 24678
rect 24315 30638 24381 30658
rect 24315 24658 24381 24678
rect 24473 30638 24539 30658
rect 24473 24658 24539 24678
rect 24631 30638 24697 30658
rect 24631 24658 24697 24678
rect 24789 30638 24855 30658
rect 24789 24658 24855 24678
rect 24947 30638 25013 30658
rect 24947 24658 25013 24678
rect 25105 30638 25171 30658
rect 25105 24658 25171 24678
rect 20432 24610 20452 24626
rect 25086 24610 25106 24626
rect 20432 24540 20440 24610
rect 25090 24540 25106 24610
rect 20432 24526 20452 24540
rect 25086 24526 25106 24540
rect 18940 24430 19010 24500
rect 19400 23900 19900 24500
rect 20230 24430 20300 24500
rect 25500 30850 26500 30860
rect 25500 30650 25520 30850
rect 25590 30650 25910 30850
rect 25980 30650 26020 30850
rect 26090 30650 26410 30850
rect 26480 30650 26500 30850
rect 25500 30640 26500 30650
rect 25640 30590 25860 30640
rect 25640 30520 25650 30590
rect 25850 30520 25860 30590
rect 25640 30480 25860 30520
rect 25640 30410 25650 30480
rect 25850 30410 25860 30480
rect 25640 30360 25860 30410
rect 26140 30590 26360 30640
rect 26140 30520 26150 30590
rect 26350 30520 26360 30590
rect 26140 30480 26360 30520
rect 26140 30410 26150 30480
rect 26350 30410 26360 30480
rect 26140 30360 26360 30410
rect 25500 30350 26500 30360
rect 25500 30150 25520 30350
rect 25590 30150 25910 30350
rect 25980 30150 26020 30350
rect 26090 30150 26410 30350
rect 26480 30150 26500 30350
rect 25500 30140 26500 30150
rect 25640 30090 25860 30140
rect 25640 30020 25650 30090
rect 25850 30020 25860 30090
rect 25640 29980 25860 30020
rect 25640 29910 25650 29980
rect 25850 29910 25860 29980
rect 25640 29860 25860 29910
rect 26140 30090 26360 30140
rect 26140 30020 26150 30090
rect 26350 30020 26360 30090
rect 26140 29980 26360 30020
rect 26140 29910 26150 29980
rect 26350 29910 26360 29980
rect 26140 29860 26360 29910
rect 25500 29850 26500 29860
rect 25500 29650 25520 29850
rect 25590 29650 25910 29850
rect 25980 29650 26020 29850
rect 26090 29650 26410 29850
rect 26480 29650 26500 29850
rect 25500 29640 26500 29650
rect 25640 29590 25860 29640
rect 25640 29520 25650 29590
rect 25850 29520 25860 29590
rect 25640 29480 25860 29520
rect 25640 29410 25650 29480
rect 25850 29410 25860 29480
rect 25640 29360 25860 29410
rect 26140 29590 26360 29640
rect 26140 29520 26150 29590
rect 26350 29520 26360 29590
rect 26140 29480 26360 29520
rect 26140 29410 26150 29480
rect 26350 29410 26360 29480
rect 26140 29360 26360 29410
rect 25500 29350 26500 29360
rect 25500 29150 25520 29350
rect 25590 29150 25910 29350
rect 25980 29150 26020 29350
rect 26090 29150 26410 29350
rect 26480 29150 26500 29350
rect 25500 29140 26500 29150
rect 25640 29090 25860 29140
rect 25640 29020 25650 29090
rect 25850 29020 25860 29090
rect 25640 28980 25860 29020
rect 25640 28910 25650 28980
rect 25850 28910 25860 28980
rect 25640 28860 25860 28910
rect 26140 29090 26360 29140
rect 26140 29020 26150 29090
rect 26350 29020 26360 29090
rect 26140 28980 26360 29020
rect 26140 28910 26150 28980
rect 26350 28910 26360 28980
rect 26140 28860 26360 28910
rect 25500 28850 26500 28860
rect 25500 28650 25520 28850
rect 25590 28650 25910 28850
rect 25980 28650 26020 28850
rect 26090 28650 26410 28850
rect 26480 28650 26500 28850
rect 25500 28640 26500 28650
rect 25640 28590 25860 28640
rect 25640 28520 25650 28590
rect 25850 28520 25860 28590
rect 25640 28480 25860 28520
rect 25640 28410 25650 28480
rect 25850 28410 25860 28480
rect 25640 28360 25860 28410
rect 26140 28590 26360 28640
rect 26140 28520 26150 28590
rect 26350 28520 26360 28590
rect 26140 28480 26360 28520
rect 26140 28410 26150 28480
rect 26350 28410 26360 28480
rect 26140 28360 26360 28410
rect 25500 28350 26500 28360
rect 25500 28150 25520 28350
rect 25590 28150 25910 28350
rect 25980 28150 26020 28350
rect 26090 28150 26410 28350
rect 26480 28150 26500 28350
rect 25500 28140 26500 28150
rect 25640 28090 25860 28140
rect 25640 28020 25650 28090
rect 25850 28020 25860 28090
rect 25640 27980 25860 28020
rect 25640 27910 25650 27980
rect 25850 27910 25860 27980
rect 25640 27860 25860 27910
rect 26140 28090 26360 28140
rect 26140 28020 26150 28090
rect 26350 28020 26360 28090
rect 26140 27980 26360 28020
rect 26140 27910 26150 27980
rect 26350 27910 26360 27980
rect 26140 27860 26360 27910
rect 25500 27850 26500 27860
rect 25500 27650 25520 27850
rect 25590 27650 25910 27850
rect 25980 27650 26020 27850
rect 26090 27650 26410 27850
rect 26480 27650 26500 27850
rect 25500 27640 26500 27650
rect 25640 27590 25860 27640
rect 25640 27520 25650 27590
rect 25850 27520 25860 27590
rect 25640 27480 25860 27520
rect 25640 27410 25650 27480
rect 25850 27410 25860 27480
rect 25640 27360 25860 27410
rect 26140 27590 26360 27640
rect 26140 27520 26150 27590
rect 26350 27520 26360 27590
rect 26140 27480 26360 27520
rect 26140 27410 26150 27480
rect 26350 27410 26360 27480
rect 26140 27360 26360 27410
rect 25500 27350 26500 27360
rect 25500 27150 25520 27350
rect 25590 27150 25910 27350
rect 25980 27150 26020 27350
rect 26090 27150 26410 27350
rect 26480 27150 26500 27350
rect 25500 27140 26500 27150
rect 30900 27250 31100 27260
rect 25640 27090 25860 27140
rect 25640 27020 25650 27090
rect 25850 27020 25860 27090
rect 25640 26980 25860 27020
rect 25640 26910 25650 26980
rect 25850 26910 25860 26980
rect 25640 26860 25860 26910
rect 26140 27090 26360 27140
rect 26140 27020 26150 27090
rect 26350 27020 26360 27090
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect 26140 26980 26360 27020
rect 26140 26910 26150 26980
rect 26350 26910 26360 26980
rect 26140 26860 26360 26910
rect 26640 26980 26860 27000
rect 26640 26910 26650 26980
rect 26850 26910 26860 26980
rect 26640 26860 26860 26910
rect 27140 26980 27360 27000
rect 27140 26910 27150 26980
rect 27350 26910 27360 26980
rect 27140 26860 27360 26910
rect 27640 26980 27860 27000
rect 27640 26910 27650 26980
rect 27850 26910 27860 26980
rect 27640 26860 27860 26910
rect 28140 26980 28360 27000
rect 28140 26910 28150 26980
rect 28350 26910 28360 26980
rect 28140 26860 28360 26910
rect 28640 26980 28860 27000
rect 28640 26910 28650 26980
rect 28850 26910 28860 26980
rect 28640 26860 28860 26910
rect 29140 26980 29360 27000
rect 29140 26910 29150 26980
rect 29350 26910 29360 26980
rect 29140 26860 29360 26910
rect 29640 26980 29860 27000
rect 29640 26910 29650 26980
rect 29850 26910 29860 26980
rect 29640 26860 29860 26910
rect 30140 26980 30360 27000
rect 30140 26910 30150 26980
rect 30350 26910 30360 26980
rect 30140 26860 30360 26910
rect 25500 26850 30500 26860
rect 25500 26650 25520 26850
rect 25590 26650 25910 26850
rect 25980 26650 26020 26850
rect 26090 26650 26410 26850
rect 26480 26650 26520 26850
rect 26590 26650 26910 26850
rect 26980 26650 27020 26850
rect 27090 26650 27410 26850
rect 27480 26650 27520 26850
rect 27590 26650 27910 26850
rect 27980 26650 28020 26850
rect 28090 26650 28410 26850
rect 28480 26650 28520 26850
rect 28590 26650 28910 26850
rect 28980 26650 29020 26850
rect 29090 26650 29410 26850
rect 29480 26650 29520 26850
rect 29590 26650 29910 26850
rect 29980 26650 30020 26850
rect 30090 26650 30410 26850
rect 30480 26650 30500 26850
rect 25500 26640 30500 26650
rect 25640 26590 25860 26640
rect 25640 26520 25650 26590
rect 25850 26520 25860 26590
rect 25640 26480 25860 26520
rect 25640 26410 25650 26480
rect 25850 26410 25860 26480
rect 25640 26360 25860 26410
rect 26140 26590 26360 26640
rect 26140 26520 26150 26590
rect 26350 26520 26360 26590
rect 26140 26480 26360 26520
rect 26140 26410 26150 26480
rect 26350 26410 26360 26480
rect 26140 26360 26360 26410
rect 26640 26590 26860 26640
rect 26640 26520 26650 26590
rect 26850 26520 26860 26590
rect 26640 26480 26860 26520
rect 26640 26410 26650 26480
rect 26850 26410 26860 26480
rect 26640 26360 26860 26410
rect 27140 26590 27360 26640
rect 27140 26520 27150 26590
rect 27350 26520 27360 26590
rect 27140 26480 27360 26520
rect 27140 26410 27150 26480
rect 27350 26410 27360 26480
rect 27140 26360 27360 26410
rect 27640 26590 27860 26640
rect 27640 26520 27650 26590
rect 27850 26520 27860 26590
rect 27640 26480 27860 26520
rect 27640 26410 27650 26480
rect 27850 26410 27860 26480
rect 27640 26360 27860 26410
rect 28140 26590 28360 26640
rect 28140 26520 28150 26590
rect 28350 26520 28360 26590
rect 28140 26480 28360 26520
rect 28140 26410 28150 26480
rect 28350 26410 28360 26480
rect 28140 26360 28360 26410
rect 28640 26590 28860 26640
rect 28640 26520 28650 26590
rect 28850 26520 28860 26590
rect 28640 26480 28860 26520
rect 28640 26410 28650 26480
rect 28850 26410 28860 26480
rect 28640 26360 28860 26410
rect 29140 26590 29360 26640
rect 29140 26520 29150 26590
rect 29350 26520 29360 26590
rect 29140 26480 29360 26520
rect 29140 26410 29150 26480
rect 29350 26410 29360 26480
rect 29140 26360 29360 26410
rect 29640 26590 29860 26640
rect 29640 26520 29650 26590
rect 29850 26520 29860 26590
rect 29640 26480 29860 26520
rect 29640 26410 29650 26480
rect 29850 26410 29860 26480
rect 29640 26360 29860 26410
rect 30140 26590 30360 26640
rect 30140 26520 30150 26590
rect 30350 26520 30360 26590
rect 30140 26480 30360 26520
rect 30140 26410 30150 26480
rect 30350 26410 30360 26480
rect 30140 26360 30360 26410
rect 25500 26350 30500 26360
rect 25500 26150 25520 26350
rect 25590 26150 25910 26350
rect 25980 26150 26020 26350
rect 26090 26150 26410 26350
rect 26480 26150 26520 26350
rect 26590 26150 26910 26350
rect 26980 26150 27020 26350
rect 27090 26150 27410 26350
rect 27480 26150 27520 26350
rect 27590 26150 27910 26350
rect 27980 26150 28020 26350
rect 28090 26150 28410 26350
rect 28480 26150 28520 26350
rect 28590 26150 28910 26350
rect 28980 26150 29020 26350
rect 29090 26150 29410 26350
rect 29480 26150 29520 26350
rect 29590 26150 29910 26350
rect 29980 26150 30020 26350
rect 30090 26150 30410 26350
rect 30480 26150 30500 26350
rect 25500 26140 30500 26150
rect 25640 26090 25860 26140
rect 25640 26020 25650 26090
rect 25850 26020 25860 26090
rect 25640 25980 25860 26020
rect 25640 25910 25650 25980
rect 25850 25910 25860 25980
rect 25640 25860 25860 25910
rect 26140 26090 26360 26140
rect 26140 26020 26150 26090
rect 26350 26020 26360 26090
rect 26140 25980 26360 26020
rect 26640 26090 26860 26140
rect 26640 26020 26650 26090
rect 26850 26020 26860 26090
rect 26640 26000 26860 26020
rect 27140 26090 27360 26140
rect 27140 26020 27150 26090
rect 27350 26020 27360 26090
rect 27140 26000 27360 26020
rect 27640 26090 27860 26140
rect 27640 26020 27650 26090
rect 27850 26020 27860 26090
rect 27640 26000 27860 26020
rect 28140 26090 28360 26140
rect 28140 26020 28150 26090
rect 28350 26020 28360 26090
rect 28140 26000 28360 26020
rect 28640 26090 28860 26140
rect 28640 26020 28650 26090
rect 28850 26020 28860 26090
rect 28640 26000 28860 26020
rect 29140 26090 29360 26140
rect 29140 26020 29150 26090
rect 29350 26020 29360 26090
rect 29140 26000 29360 26020
rect 29640 26090 29860 26140
rect 29640 26020 29650 26090
rect 29850 26020 29860 26090
rect 29640 26000 29860 26020
rect 30140 26090 30360 26140
rect 30140 26020 30150 26090
rect 30350 26020 30360 26090
rect 30140 26000 30360 26020
rect 26140 25910 26150 25980
rect 26350 25910 26360 25980
rect 26140 25860 26360 25910
rect 25500 25850 26500 25860
rect 25500 25650 25520 25850
rect 25590 25650 25910 25850
rect 25980 25650 26020 25850
rect 26090 25650 26410 25850
rect 26480 25650 26500 25850
rect 25500 25640 26500 25650
rect 30900 25710 31100 25720
rect 25640 25590 25860 25640
rect 25640 25520 25650 25590
rect 25850 25520 25860 25590
rect 25640 25480 25860 25520
rect 25640 25410 25650 25480
rect 25850 25410 25860 25480
rect 25640 25360 25860 25410
rect 26140 25590 26360 25640
rect 26140 25520 26150 25590
rect 26350 25520 26360 25590
rect 26140 25480 26360 25520
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect 26140 25410 26150 25480
rect 26350 25410 26360 25480
rect 26140 25360 26360 25410
rect 25500 25350 26500 25360
rect 25500 25150 25520 25350
rect 25590 25150 25910 25350
rect 25980 25150 26020 25350
rect 26090 25150 26410 25350
rect 26480 25150 26500 25350
rect 25500 25140 26500 25150
rect 25640 25090 25860 25140
rect 25640 25020 25650 25090
rect 25850 25020 25860 25090
rect 25640 24980 25860 25020
rect 25640 24910 25650 24980
rect 25850 24910 25860 24980
rect 25640 24860 25860 24910
rect 26140 25090 26360 25140
rect 26140 25020 26150 25090
rect 26350 25020 26360 25090
rect 26140 24980 26360 25020
rect 26140 24910 26150 24980
rect 26350 24910 26360 24980
rect 26140 24860 26360 24910
rect 25500 24850 26500 24860
rect 25500 24650 25520 24850
rect 25590 24650 25910 24850
rect 25980 24650 26020 24850
rect 26090 24650 26410 24850
rect 26480 24650 26500 24850
rect 25500 24640 26500 24650
rect 25240 24430 25310 24500
rect 25640 24590 25860 24640
rect 25640 24520 25650 24590
rect 25850 24520 25860 24590
rect 25640 24480 25860 24520
rect 25640 24410 25650 24480
rect 25850 24410 25860 24480
rect 25640 24360 25860 24410
rect 26140 24590 26360 24640
rect 26140 24520 26150 24590
rect 26350 24520 26360 24590
rect 26140 24480 26360 24520
rect 26140 24410 26150 24480
rect 26350 24410 26360 24480
rect 26140 24360 26360 24410
rect 25500 24350 26500 24360
rect 25500 24150 25520 24350
rect 25590 24150 25910 24350
rect 25980 24150 26020 24350
rect 26090 24150 26410 24350
rect 26480 24150 26500 24350
rect 25500 24140 26500 24150
rect 25640 24090 25860 24140
rect 25640 24020 25650 24090
rect 25850 24020 25860 24090
rect 25640 23980 25860 24020
rect 25640 23910 25650 23980
rect 25850 23910 25860 23980
rect 6400 23880 7700 23900
rect 12700 23880 14000 23900
rect 19000 23880 20300 23900
rect 0 23850 1000 23860
rect 0 23650 20 23850
rect 90 23650 410 23850
rect 480 23650 520 23850
rect 590 23650 910 23850
rect 980 23650 1000 23850
rect 0 23640 1000 23650
rect 1330 23820 1400 23880
rect 140 23590 360 23640
rect 140 23520 150 23590
rect 350 23520 360 23590
rect 140 23480 360 23520
rect 140 23410 150 23480
rect 350 23410 360 23480
rect 140 23360 360 23410
rect 640 23590 860 23640
rect 640 23520 650 23590
rect 850 23520 860 23590
rect 640 23480 860 23520
rect 640 23410 650 23480
rect 850 23410 860 23480
rect 640 23360 860 23410
rect 0 23350 1000 23360
rect 0 23150 20 23350
rect 90 23150 410 23350
rect 480 23150 520 23350
rect 590 23150 910 23350
rect 980 23150 1000 23350
rect 0 23140 1000 23150
rect 140 23090 360 23140
rect 140 23020 150 23090
rect 350 23020 360 23090
rect 140 22980 360 23020
rect 140 22910 150 22980
rect 350 22910 360 22980
rect 140 22860 360 22910
rect 640 23090 860 23140
rect 640 23020 650 23090
rect 850 23020 860 23090
rect 640 22980 860 23020
rect 640 22910 650 22980
rect 850 22910 860 22980
rect 640 22860 860 22910
rect 0 22850 1000 22860
rect 0 22650 20 22850
rect 90 22650 410 22850
rect 480 22650 520 22850
rect 590 22650 910 22850
rect 980 22650 1000 22850
rect 0 22640 1000 22650
rect 140 22590 360 22640
rect 140 22520 150 22590
rect 350 22520 360 22590
rect 140 22480 360 22520
rect 140 22410 150 22480
rect 350 22410 360 22480
rect 140 22360 360 22410
rect 640 22590 860 22640
rect 640 22520 650 22590
rect 850 22520 860 22590
rect 640 22480 860 22520
rect 640 22410 650 22480
rect 850 22410 860 22480
rect 640 22360 860 22410
rect 0 22350 1000 22360
rect 0 22150 20 22350
rect 90 22150 410 22350
rect 480 22150 520 22350
rect 590 22150 910 22350
rect 980 22150 1000 22350
rect 0 22140 1000 22150
rect 140 22090 360 22140
rect 140 22020 150 22090
rect 350 22020 360 22090
rect 140 21980 360 22020
rect 140 21910 150 21980
rect 350 21910 360 21980
rect 140 21860 360 21910
rect 640 22090 860 22140
rect 640 22020 650 22090
rect 850 22020 860 22090
rect 640 21980 860 22020
rect 640 21910 650 21980
rect 850 21910 860 21980
rect 640 21860 860 21910
rect 0 21850 1000 21860
rect 0 21650 20 21850
rect 90 21650 410 21850
rect 480 21650 520 21850
rect 590 21650 910 21850
rect 980 21650 1000 21850
rect 0 21640 1000 21650
rect 140 21590 360 21640
rect 140 21520 150 21590
rect 350 21520 360 21590
rect 140 21480 360 21520
rect 140 21410 150 21480
rect 350 21410 360 21480
rect 140 21360 360 21410
rect 640 21590 860 21640
rect 640 21520 650 21590
rect 850 21520 860 21590
rect 640 21480 860 21520
rect 640 21410 650 21480
rect 850 21410 860 21480
rect 640 21360 860 21410
rect 0 21350 1000 21360
rect 0 21150 20 21350
rect 90 21150 410 21350
rect 480 21150 520 21350
rect 590 21150 910 21350
rect 980 21150 1000 21350
rect 0 21140 1000 21150
rect 140 21090 360 21140
rect 140 21020 150 21090
rect 350 21020 360 21090
rect 140 20980 360 21020
rect 140 20910 150 20980
rect 350 20910 360 20980
rect 140 20860 360 20910
rect 640 21090 860 21140
rect 640 21020 650 21090
rect 850 21020 860 21090
rect 640 20980 860 21020
rect 640 20910 650 20980
rect 850 20910 860 20980
rect 640 20860 860 20910
rect 0 20850 1000 20860
rect 0 20650 20 20850
rect 90 20650 410 20850
rect 480 20650 520 20850
rect 590 20650 910 20850
rect 980 20650 1000 20850
rect 0 20640 1000 20650
rect 140 20590 360 20640
rect 140 20520 150 20590
rect 350 20520 360 20590
rect 140 20480 360 20520
rect 140 20410 150 20480
rect 350 20410 360 20480
rect 140 20360 360 20410
rect 640 20590 860 20640
rect 640 20520 650 20590
rect 850 20520 860 20590
rect 640 20480 860 20520
rect 640 20410 650 20480
rect 850 20410 860 20480
rect 640 20360 860 20410
rect 0 20350 1000 20360
rect 0 20150 20 20350
rect 90 20150 410 20350
rect 480 20150 520 20350
rect 590 20150 910 20350
rect 980 20150 1000 20350
rect 0 20140 1000 20150
rect 140 20090 360 20140
rect 140 20020 150 20090
rect 350 20020 360 20090
rect 140 19980 360 20020
rect 140 19910 150 19980
rect 350 19910 360 19980
rect 140 19860 360 19910
rect 640 20090 860 20140
rect 640 20020 650 20090
rect 850 20020 860 20090
rect 640 19980 860 20020
rect 640 19910 650 19980
rect 850 19910 860 19980
rect 640 19860 860 19910
rect 0 19850 1000 19860
rect 0 19650 20 19850
rect 90 19650 410 19850
rect 480 19650 520 19850
rect 590 19650 910 19850
rect 980 19650 1000 19850
rect 0 19640 1000 19650
rect 140 19590 360 19640
rect 140 19520 150 19590
rect 350 19520 360 19590
rect 140 19480 360 19520
rect 140 19410 150 19480
rect 350 19410 360 19480
rect 140 19360 360 19410
rect 640 19590 860 19640
rect 640 19520 650 19590
rect 850 19520 860 19590
rect 640 19480 860 19520
rect 640 19410 650 19480
rect 850 19410 860 19480
rect 640 19360 860 19410
rect 0 19350 1000 19360
rect 0 19150 20 19350
rect 90 19150 410 19350
rect 480 19150 520 19350
rect 590 19150 910 19350
rect 980 19150 1000 19350
rect 0 19140 1000 19150
rect 140 19090 360 19140
rect 140 19020 150 19090
rect 350 19020 360 19090
rect 140 18980 360 19020
rect 140 18910 150 18980
rect 350 18910 360 18980
rect 140 18860 360 18910
rect 640 19090 860 19140
rect 640 19020 650 19090
rect 850 19020 860 19090
rect 640 18980 860 19020
rect 640 18910 650 18980
rect 850 18910 860 18980
rect 640 18860 860 18910
rect 0 18850 1000 18860
rect 0 18650 20 18850
rect 90 18650 410 18850
rect 480 18650 520 18850
rect 590 18650 910 18850
rect 980 18650 1000 18850
rect 0 18640 1000 18650
rect 140 18590 360 18640
rect 140 18520 150 18590
rect 350 18520 360 18590
rect 140 18480 360 18520
rect 140 18410 150 18480
rect 350 18410 360 18480
rect 140 18360 360 18410
rect 640 18590 860 18640
rect 640 18520 650 18590
rect 850 18520 860 18590
rect 640 18480 860 18520
rect 640 18410 650 18480
rect 850 18410 860 18480
rect 640 18360 860 18410
rect 0 18350 1000 18360
rect 0 18150 20 18350
rect 90 18150 410 18350
rect 480 18150 520 18350
rect 590 18150 910 18350
rect 980 18150 1000 18350
rect 0 18140 1000 18150
rect 140 18090 360 18140
rect 140 18020 150 18090
rect 350 18020 360 18090
rect 140 17980 360 18020
rect 140 17910 150 17980
rect 350 17910 360 17980
rect 140 17860 360 17910
rect 640 18090 860 18140
rect 640 18020 650 18090
rect 850 18020 860 18090
rect 640 17980 860 18020
rect 640 17910 650 17980
rect 850 17910 860 17980
rect 640 17860 860 17910
rect 0 17850 1000 17860
rect 0 17650 20 17850
rect 90 17650 410 17850
rect 480 17650 520 17850
rect 590 17650 910 17850
rect 980 17650 1000 17850
rect 0 17640 1000 17650
rect 140 17590 360 17640
rect 140 17520 150 17590
rect 350 17520 360 17590
rect 140 17480 360 17520
rect 140 17410 150 17480
rect 350 17410 360 17480
rect 140 17360 360 17410
rect 640 17590 860 17640
rect 640 17520 650 17590
rect 850 17520 860 17590
rect 640 17480 860 17520
rect 640 17410 650 17480
rect 850 17410 860 17480
rect 6340 23820 7700 23880
rect 1532 23780 1552 23790
rect 6186 23780 6206 23790
rect 1532 23710 1540 23780
rect 6200 23710 6206 23780
rect 1532 23690 1552 23710
rect 6186 23690 6206 23710
rect 1465 23638 1531 23658
rect 1465 17658 1531 17678
rect 1623 23638 1689 23658
rect 1623 17658 1689 17678
rect 1781 23638 1847 23658
rect 1781 17658 1847 17678
rect 1939 23638 2005 23658
rect 1939 17658 2005 17678
rect 2097 23638 2163 23658
rect 2097 17658 2163 17678
rect 2255 23638 2321 23658
rect 2255 17658 2321 17678
rect 2413 23638 2479 23658
rect 2413 17658 2479 17678
rect 2571 23638 2637 23658
rect 2571 17658 2637 17678
rect 2729 23638 2795 23658
rect 2729 17658 2795 17678
rect 2887 23638 2953 23658
rect 2887 17658 2953 17678
rect 3045 23638 3111 23658
rect 3045 17658 3111 17678
rect 3203 23638 3269 23658
rect 3203 17658 3269 17678
rect 3361 23638 3427 23658
rect 3361 17658 3427 17678
rect 3519 23638 3585 23658
rect 3519 17658 3585 17678
rect 3677 23638 3743 23658
rect 3677 17658 3743 17678
rect 3835 23638 3901 23658
rect 3835 17658 3901 17678
rect 3993 23638 4059 23658
rect 3993 17658 4059 17678
rect 4151 23638 4217 23658
rect 4151 17658 4217 17678
rect 4309 23638 4375 23658
rect 4309 17658 4375 17678
rect 4467 23638 4533 23658
rect 4467 17658 4533 17678
rect 4625 23638 4691 23658
rect 4625 17658 4691 17678
rect 4783 23638 4849 23658
rect 4783 17658 4849 17678
rect 4941 23638 5007 23658
rect 4941 17658 5007 17678
rect 5099 23638 5165 23658
rect 5099 17658 5165 17678
rect 5257 23638 5323 23658
rect 5257 17658 5323 17678
rect 5415 23638 5481 23658
rect 5415 17658 5481 17678
rect 5573 23638 5639 23658
rect 5573 17658 5639 17678
rect 5731 23638 5797 23658
rect 5731 17658 5797 17678
rect 5889 23638 5955 23658
rect 5889 17658 5955 17678
rect 6047 23638 6113 23658
rect 6047 17658 6113 17678
rect 6205 23638 6271 23658
rect 6205 17658 6271 17678
rect 1532 17610 1552 17626
rect 6186 17610 6206 17626
rect 1532 17540 1540 17610
rect 6190 17540 6206 17610
rect 1532 17526 1552 17540
rect 6186 17526 6206 17540
rect 1330 17430 1400 17500
rect 6410 23500 7630 23820
rect 6410 22900 7630 23300
rect 6410 22300 7630 22700
rect 6410 21700 7630 22100
rect 6410 21100 7630 21500
rect 6410 20500 7630 20900
rect 6410 19900 7630 20300
rect 6410 19300 7630 19700
rect 6410 18700 7630 19100
rect 6410 18100 7630 18500
rect 6410 17500 7630 17900
rect 12640 23820 14000 23880
rect 7832 23780 7852 23790
rect 12486 23780 12506 23790
rect 7832 23710 7840 23780
rect 12500 23710 12506 23780
rect 7832 23690 7852 23710
rect 12486 23690 12506 23710
rect 7765 23638 7831 23658
rect 7765 17658 7831 17678
rect 7923 23638 7989 23658
rect 7923 17658 7989 17678
rect 8081 23638 8147 23658
rect 8081 17658 8147 17678
rect 8239 23638 8305 23658
rect 8239 17658 8305 17678
rect 8397 23638 8463 23658
rect 8397 17658 8463 17678
rect 8555 23638 8621 23658
rect 8555 17658 8621 17678
rect 8713 23638 8779 23658
rect 8713 17658 8779 17678
rect 8871 23638 8937 23658
rect 8871 17658 8937 17678
rect 9029 23638 9095 23658
rect 9029 17658 9095 17678
rect 9187 23638 9253 23658
rect 9187 17658 9253 17678
rect 9345 23638 9411 23658
rect 9345 17658 9411 17678
rect 9503 23638 9569 23658
rect 9503 17658 9569 17678
rect 9661 23638 9727 23658
rect 9661 17658 9727 17678
rect 9819 23638 9885 23658
rect 9819 17658 9885 17678
rect 9977 23638 10043 23658
rect 9977 17658 10043 17678
rect 10135 23638 10201 23658
rect 10135 17658 10201 17678
rect 10293 23638 10359 23658
rect 10293 17658 10359 17678
rect 10451 23638 10517 23658
rect 10451 17658 10517 17678
rect 10609 23638 10675 23658
rect 10609 17658 10675 17678
rect 10767 23638 10833 23658
rect 10767 17658 10833 17678
rect 10925 23638 10991 23658
rect 10925 17658 10991 17678
rect 11083 23638 11149 23658
rect 11083 17658 11149 17678
rect 11241 23638 11307 23658
rect 11241 17658 11307 17678
rect 11399 23638 11465 23658
rect 11399 17658 11465 17678
rect 11557 23638 11623 23658
rect 11557 17658 11623 17678
rect 11715 23638 11781 23658
rect 11715 17658 11781 17678
rect 11873 23638 11939 23658
rect 11873 17658 11939 17678
rect 12031 23638 12097 23658
rect 12031 17658 12097 17678
rect 12189 23638 12255 23658
rect 12189 17658 12255 17678
rect 12347 23638 12413 23658
rect 12347 17658 12413 17678
rect 12505 23638 12571 23658
rect 12505 17658 12571 17678
rect 7832 17610 7852 17626
rect 12486 17610 12506 17626
rect 7832 17540 7840 17610
rect 12490 17540 12506 17610
rect 7832 17526 7852 17540
rect 12486 17526 12506 17540
rect 6340 17430 6410 17500
rect 6640 17480 6860 17500
rect 640 17360 860 17410
rect 6640 17410 6650 17480
rect 6850 17410 6860 17480
rect 6640 17360 6860 17410
rect 7140 17480 7360 17500
rect 7140 17410 7150 17480
rect 7350 17410 7360 17480
rect 7630 17430 7700 17500
rect 12710 23500 13930 23820
rect 12710 22900 13930 23300
rect 12710 22300 13930 22700
rect 12710 21700 13930 22100
rect 12710 21100 13930 21500
rect 12710 20500 13930 20900
rect 12710 19900 13930 20300
rect 12710 19300 13930 19700
rect 12710 18700 13930 19100
rect 12710 18100 13930 18500
rect 12710 17500 13930 17900
rect 18940 23820 20300 23880
rect 14132 23780 14152 23790
rect 18786 23780 18806 23790
rect 14132 23710 14140 23780
rect 18800 23710 18806 23780
rect 14132 23690 14152 23710
rect 18786 23690 18806 23710
rect 14065 23638 14131 23658
rect 14065 17658 14131 17678
rect 14223 23638 14289 23658
rect 14223 17658 14289 17678
rect 14381 23638 14447 23658
rect 14381 17658 14447 17678
rect 14539 23638 14605 23658
rect 14539 17658 14605 17678
rect 14697 23638 14763 23658
rect 14697 17658 14763 17678
rect 14855 23638 14921 23658
rect 14855 17658 14921 17678
rect 15013 23638 15079 23658
rect 15013 17658 15079 17678
rect 15171 23638 15237 23658
rect 15171 17658 15237 17678
rect 15329 23638 15395 23658
rect 15329 17658 15395 17678
rect 15487 23638 15553 23658
rect 15487 17658 15553 17678
rect 15645 23638 15711 23658
rect 15645 17658 15711 17678
rect 15803 23638 15869 23658
rect 15803 17658 15869 17678
rect 15961 23638 16027 23658
rect 15961 17658 16027 17678
rect 16119 23638 16185 23658
rect 16119 17658 16185 17678
rect 16277 23638 16343 23658
rect 16277 17658 16343 17678
rect 16435 23638 16501 23658
rect 16435 17658 16501 17678
rect 16593 23638 16659 23658
rect 16593 17658 16659 17678
rect 16751 23638 16817 23658
rect 16751 17658 16817 17678
rect 16909 23638 16975 23658
rect 16909 17658 16975 17678
rect 17067 23638 17133 23658
rect 17067 17658 17133 17678
rect 17225 23638 17291 23658
rect 17225 17658 17291 17678
rect 17383 23638 17449 23658
rect 17383 17658 17449 17678
rect 17541 23638 17607 23658
rect 17541 17658 17607 17678
rect 17699 23638 17765 23658
rect 17699 17658 17765 17678
rect 17857 23638 17923 23658
rect 17857 17658 17923 17678
rect 18015 23638 18081 23658
rect 18015 17658 18081 17678
rect 18173 23638 18239 23658
rect 18173 17658 18239 17678
rect 18331 23638 18397 23658
rect 18331 17658 18397 17678
rect 18489 23638 18555 23658
rect 18489 17658 18555 17678
rect 18647 23638 18713 23658
rect 18647 17658 18713 17678
rect 18805 23638 18871 23658
rect 18805 17658 18871 17678
rect 14132 17610 14152 17626
rect 18786 17610 18806 17626
rect 14132 17540 14140 17610
rect 18790 17540 18806 17610
rect 14132 17526 14152 17540
rect 18786 17526 18806 17540
rect 12640 17430 12710 17500
rect 13140 17480 13360 17500
rect 7140 17360 7360 17410
rect 13140 17410 13150 17480
rect 13350 17410 13360 17480
rect 13140 17360 13360 17410
rect 13640 17480 13860 17500
rect 13640 17410 13650 17480
rect 13850 17410 13860 17480
rect 13930 17430 14000 17500
rect 19010 23500 20230 23820
rect 19010 22900 20230 23300
rect 19010 22300 20230 22700
rect 19010 21700 20230 22100
rect 19010 21100 20230 21500
rect 19010 20500 20230 20900
rect 19010 19900 20230 20300
rect 19010 19300 20230 19700
rect 19010 18700 20230 19100
rect 19010 18100 20230 18500
rect 19010 17500 20230 17900
rect 25240 23820 25310 23880
rect 25640 23860 25860 23910
rect 26140 24090 26360 24140
rect 26140 24020 26150 24090
rect 26350 24020 26360 24090
rect 26140 23980 26360 24020
rect 26140 23910 26150 23980
rect 26350 23910 26360 23980
rect 26140 23860 26360 23910
rect 20432 23780 20452 23790
rect 25086 23780 25106 23790
rect 20432 23710 20440 23780
rect 25100 23710 25106 23780
rect 20432 23690 20452 23710
rect 25086 23690 25106 23710
rect 20365 23638 20431 23658
rect 20365 17658 20431 17678
rect 20523 23638 20589 23658
rect 20523 17658 20589 17678
rect 20681 23638 20747 23658
rect 20681 17658 20747 17678
rect 20839 23638 20905 23658
rect 20839 17658 20905 17678
rect 20997 23638 21063 23658
rect 20997 17658 21063 17678
rect 21155 23638 21221 23658
rect 21155 17658 21221 17678
rect 21313 23638 21379 23658
rect 21313 17658 21379 17678
rect 21471 23638 21537 23658
rect 21471 17658 21537 17678
rect 21629 23638 21695 23658
rect 21629 17658 21695 17678
rect 21787 23638 21853 23658
rect 21787 17658 21853 17678
rect 21945 23638 22011 23658
rect 21945 17658 22011 17678
rect 22103 23638 22169 23658
rect 22103 17658 22169 17678
rect 22261 23638 22327 23658
rect 22261 17658 22327 17678
rect 22419 23638 22485 23658
rect 22419 17658 22485 17678
rect 22577 23638 22643 23658
rect 22577 17658 22643 17678
rect 22735 23638 22801 23658
rect 22735 17658 22801 17678
rect 22893 23638 22959 23658
rect 22893 17658 22959 17678
rect 23051 23638 23117 23658
rect 23051 17658 23117 17678
rect 23209 23638 23275 23658
rect 23209 17658 23275 17678
rect 23367 23638 23433 23658
rect 23367 17658 23433 17678
rect 23525 23638 23591 23658
rect 23525 17658 23591 17678
rect 23683 23638 23749 23658
rect 23683 17658 23749 17678
rect 23841 23638 23907 23658
rect 23841 17658 23907 17678
rect 23999 23638 24065 23658
rect 23999 17658 24065 17678
rect 24157 23638 24223 23658
rect 24157 17658 24223 17678
rect 24315 23638 24381 23658
rect 24315 17658 24381 17678
rect 24473 23638 24539 23658
rect 24473 17658 24539 17678
rect 24631 23638 24697 23658
rect 24631 17658 24697 17678
rect 24789 23638 24855 23658
rect 24789 17658 24855 17678
rect 24947 23638 25013 23658
rect 24947 17658 25013 17678
rect 25105 23638 25171 23658
rect 25105 17658 25171 17678
rect 20432 17610 20452 17626
rect 25086 17610 25106 17626
rect 20432 17540 20440 17610
rect 25090 17540 25106 17610
rect 20432 17526 20452 17540
rect 25086 17526 25106 17540
rect 18940 17430 19010 17500
rect 19140 17480 19360 17500
rect 13640 17360 13860 17410
rect 19140 17410 19150 17480
rect 19350 17410 19360 17480
rect 19140 17360 19360 17410
rect 19640 17480 19860 17500
rect 19640 17410 19650 17480
rect 19850 17410 19860 17480
rect 20230 17430 20300 17500
rect 25500 23850 26500 23860
rect 25500 23650 25520 23850
rect 25590 23650 25910 23850
rect 25980 23650 26020 23850
rect 26090 23650 26410 23850
rect 26480 23650 26500 23850
rect 25500 23640 26500 23650
rect 25640 23590 25860 23640
rect 25640 23520 25650 23590
rect 25850 23520 25860 23590
rect 25640 23480 25860 23520
rect 25640 23410 25650 23480
rect 25850 23410 25860 23480
rect 25640 23360 25860 23410
rect 26140 23590 26360 23640
rect 26140 23520 26150 23590
rect 26350 23520 26360 23590
rect 26140 23480 26360 23520
rect 26140 23410 26150 23480
rect 26350 23410 26360 23480
rect 26140 23360 26360 23410
rect 25500 23350 26500 23360
rect 25500 23150 25520 23350
rect 25590 23150 25910 23350
rect 25980 23150 26020 23350
rect 26090 23150 26410 23350
rect 26480 23150 26500 23350
rect 25500 23140 26500 23150
rect 25640 23090 25860 23140
rect 25640 23020 25650 23090
rect 25850 23020 25860 23090
rect 25640 22980 25860 23020
rect 25640 22910 25650 22980
rect 25850 22910 25860 22980
rect 25640 22860 25860 22910
rect 26140 23090 26360 23140
rect 26140 23020 26150 23090
rect 26350 23020 26360 23090
rect 26140 22980 26360 23020
rect 26140 22910 26150 22980
rect 26350 22910 26360 22980
rect 26140 22860 26360 22910
rect 25500 22850 26500 22860
rect 25500 22650 25520 22850
rect 25590 22650 25910 22850
rect 25980 22650 26020 22850
rect 26090 22650 26410 22850
rect 26480 22650 26500 22850
rect 25500 22640 26500 22650
rect 25640 22590 25860 22640
rect 25640 22520 25650 22590
rect 25850 22520 25860 22590
rect 25640 22480 25860 22520
rect 25640 22410 25650 22480
rect 25850 22410 25860 22480
rect 25640 22360 25860 22410
rect 26140 22590 26360 22640
rect 26140 22520 26150 22590
rect 26350 22520 26360 22590
rect 26140 22480 26360 22520
rect 26140 22410 26150 22480
rect 26350 22410 26360 22480
rect 26140 22360 26360 22410
rect 25500 22350 26500 22360
rect 25500 22150 25520 22350
rect 25590 22150 25910 22350
rect 25980 22150 26020 22350
rect 26090 22150 26410 22350
rect 26480 22150 26500 22350
rect 25500 22140 26500 22150
rect 25640 22090 25860 22140
rect 25640 22020 25650 22090
rect 25850 22020 25860 22090
rect 25640 21980 25860 22020
rect 25640 21910 25650 21980
rect 25850 21910 25860 21980
rect 25640 21860 25860 21910
rect 26140 22090 26360 22140
rect 26140 22020 26150 22090
rect 26350 22020 26360 22090
rect 26140 21980 26360 22020
rect 26140 21910 26150 21980
rect 26350 21910 26360 21980
rect 26140 21860 26360 21910
rect 25500 21850 26500 21860
rect 25500 21650 25520 21850
rect 25590 21650 25910 21850
rect 25980 21650 26020 21850
rect 26090 21650 26410 21850
rect 26480 21650 26500 21850
rect 25500 21640 26500 21650
rect 25640 21590 25860 21640
rect 25640 21520 25650 21590
rect 25850 21520 25860 21590
rect 25640 21480 25860 21520
rect 25640 21410 25650 21480
rect 25850 21410 25860 21480
rect 25640 21360 25860 21410
rect 26140 21590 26360 21640
rect 26140 21520 26150 21590
rect 26350 21520 26360 21590
rect 26140 21480 26360 21520
rect 26140 21410 26150 21480
rect 26350 21410 26360 21480
rect 26140 21360 26360 21410
rect 25500 21350 26500 21360
rect 25500 21150 25520 21350
rect 25590 21150 25910 21350
rect 25980 21150 26020 21350
rect 26090 21150 26410 21350
rect 26480 21150 26500 21350
rect 25500 21140 26500 21150
rect 25640 21090 25860 21140
rect 25640 21020 25650 21090
rect 25850 21020 25860 21090
rect 25640 20980 25860 21020
rect 25640 20910 25650 20980
rect 25850 20910 25860 20980
rect 25640 20860 25860 20910
rect 26140 21090 26360 21140
rect 26140 21020 26150 21090
rect 26350 21020 26360 21090
rect 26140 20980 26360 21020
rect 26140 20910 26150 20980
rect 26350 20910 26360 20980
rect 26140 20860 26360 20910
rect 25500 20850 26500 20860
rect 25500 20650 25520 20850
rect 25590 20650 25910 20850
rect 25980 20650 26020 20850
rect 26090 20650 26410 20850
rect 26480 20650 26500 20850
rect 25500 20640 26500 20650
rect 25640 20590 25860 20640
rect 25640 20520 25650 20590
rect 25850 20520 25860 20590
rect 25640 20480 25860 20520
rect 25640 20410 25650 20480
rect 25850 20410 25860 20480
rect 25640 20360 25860 20410
rect 26140 20590 26360 20640
rect 26140 20520 26150 20590
rect 26350 20520 26360 20590
rect 26140 20480 26360 20520
rect 26140 20410 26150 20480
rect 26350 20410 26360 20480
rect 26140 20360 26360 20410
rect 25500 20350 26500 20360
rect 25500 20150 25520 20350
rect 25590 20150 25910 20350
rect 25980 20150 26020 20350
rect 26090 20150 26410 20350
rect 26480 20150 26500 20350
rect 25500 20140 26500 20150
rect 25640 20090 25860 20140
rect 25640 20020 25650 20090
rect 25850 20020 25860 20090
rect 25640 19980 25860 20020
rect 25640 19910 25650 19980
rect 25850 19910 25860 19980
rect 25640 19860 25860 19910
rect 26140 20090 26360 20140
rect 26140 20020 26150 20090
rect 26350 20020 26360 20090
rect 26140 19980 26360 20020
rect 26140 19910 26150 19980
rect 26350 19910 26360 19980
rect 26140 19860 26360 19910
rect 25500 19850 26500 19860
rect 25500 19650 25520 19850
rect 25590 19650 25910 19850
rect 25980 19650 26020 19850
rect 26090 19650 26410 19850
rect 26480 19650 26500 19850
rect 25500 19640 26500 19650
rect 25640 19590 25860 19640
rect 25640 19520 25650 19590
rect 25850 19520 25860 19590
rect 25640 19480 25860 19520
rect 25640 19410 25650 19480
rect 25850 19410 25860 19480
rect 25640 19360 25860 19410
rect 26140 19590 26360 19640
rect 26140 19520 26150 19590
rect 26350 19520 26360 19590
rect 26140 19480 26360 19520
rect 26140 19410 26150 19480
rect 26350 19410 26360 19480
rect 26140 19360 26360 19410
rect 25500 19350 26500 19360
rect 25500 19150 25520 19350
rect 25590 19150 25910 19350
rect 25980 19150 26020 19350
rect 26090 19150 26410 19350
rect 26480 19150 26500 19350
rect 25500 19140 26500 19150
rect 25640 19090 25860 19140
rect 25640 19020 25650 19090
rect 25850 19020 25860 19090
rect 25640 18980 25860 19020
rect 25640 18910 25650 18980
rect 25850 18910 25860 18980
rect 25640 18860 25860 18910
rect 26140 19090 26360 19140
rect 26140 19020 26150 19090
rect 26350 19020 26360 19090
rect 26140 18980 26360 19020
rect 26140 18910 26150 18980
rect 26350 18910 26360 18980
rect 26140 18860 26360 18910
rect 25500 18850 26500 18860
rect 25500 18650 25520 18850
rect 25590 18650 25910 18850
rect 25980 18650 26020 18850
rect 26090 18650 26410 18850
rect 26480 18650 26500 18850
rect 25500 18640 26500 18650
rect 25640 18590 25860 18640
rect 25640 18520 25650 18590
rect 25850 18520 25860 18590
rect 25640 18480 25860 18520
rect 25640 18410 25650 18480
rect 25850 18410 25860 18480
rect 25640 18360 25860 18410
rect 26140 18590 26360 18640
rect 26140 18520 26150 18590
rect 26350 18520 26360 18590
rect 26140 18480 26360 18520
rect 26140 18410 26150 18480
rect 26350 18410 26360 18480
rect 26140 18360 26360 18410
rect 25500 18350 26500 18360
rect 25500 18150 25520 18350
rect 25590 18150 25910 18350
rect 25980 18150 26020 18350
rect 26090 18150 26410 18350
rect 26480 18150 26500 18350
rect 25500 18140 26500 18150
rect 25640 18090 25860 18140
rect 25640 18020 25650 18090
rect 25850 18020 25860 18090
rect 25640 17980 25860 18020
rect 25640 17910 25650 17980
rect 25850 17910 25860 17980
rect 25640 17860 25860 17910
rect 26140 18090 26360 18140
rect 26140 18020 26150 18090
rect 26350 18020 26360 18090
rect 26140 17980 26360 18020
rect 26140 17910 26150 17980
rect 26350 17910 26360 17980
rect 26140 17860 26360 17910
rect 25500 17850 26500 17860
rect 25500 17650 25520 17850
rect 25590 17650 25910 17850
rect 25980 17650 26020 17850
rect 26090 17650 26410 17850
rect 26480 17650 26500 17850
rect 25500 17640 26500 17650
rect 25240 17430 25310 17500
rect 25640 17590 25860 17640
rect 25640 17520 25650 17590
rect 25850 17520 25860 17590
rect 25640 17480 25860 17520
rect 19640 17360 19860 17410
rect 25640 17410 25650 17480
rect 25850 17410 25860 17480
rect 25640 17360 25860 17410
rect 26140 17590 26360 17640
rect 26140 17520 26150 17590
rect 26350 17520 26360 17590
rect 26140 17480 26360 17520
rect 26140 17410 26150 17480
rect 26350 17410 26360 17480
rect 26140 17360 26360 17410
rect 0 17350 1000 17360
rect 0 17150 20 17350
rect 90 17150 410 17350
rect 480 17150 520 17350
rect 590 17150 910 17350
rect 980 17150 1000 17350
rect 0 17140 1000 17150
rect 6500 17350 7500 17360
rect 6500 17150 6520 17350
rect 6590 17150 6910 17350
rect 6980 17150 7020 17350
rect 7090 17150 7410 17350
rect 7480 17150 7500 17350
rect 6500 17140 7500 17150
rect 13000 17350 14000 17360
rect 13000 17150 13020 17350
rect 13090 17150 13410 17350
rect 13480 17150 13520 17350
rect 13590 17150 13910 17350
rect 13980 17150 14000 17350
rect 13000 17140 14000 17150
rect 19000 17350 20000 17360
rect 19000 17150 19020 17350
rect 19090 17150 19410 17350
rect 19480 17150 19520 17350
rect 19590 17150 19910 17350
rect 19980 17150 20000 17350
rect 19000 17140 20000 17150
rect 25500 17350 26500 17360
rect 25500 17150 25520 17350
rect 25590 17150 25910 17350
rect 25980 17150 26020 17350
rect 26090 17150 26410 17350
rect 26480 17150 26500 17350
rect 25500 17140 26500 17150
rect 140 17090 360 17140
rect 140 17020 150 17090
rect 350 17020 360 17090
rect 140 16980 360 17020
rect 140 16910 150 16980
rect 350 16910 360 16980
rect 140 16860 360 16910
rect 640 17090 860 17140
rect 640 17020 650 17090
rect 850 17020 860 17090
rect 640 16980 860 17020
rect 6640 17090 6860 17140
rect 6640 17020 6650 17090
rect 6850 17020 6860 17090
rect 640 16910 650 16980
rect 850 16910 860 16980
rect 640 16860 860 16910
rect 1140 16980 1360 17000
rect 1140 16910 1150 16980
rect 1350 16910 1360 16980
rect 1140 16860 1360 16910
rect 1640 16980 1860 17000
rect 1640 16910 1650 16980
rect 1850 16910 1860 16980
rect 1640 16860 1860 16910
rect 2140 16980 2360 17000
rect 2140 16910 2150 16980
rect 2350 16910 2360 16980
rect 2140 16860 2360 16910
rect 2640 16980 2860 17000
rect 2640 16910 2650 16980
rect 2850 16910 2860 16980
rect 2640 16860 2860 16910
rect 3140 16980 3360 17000
rect 3140 16910 3150 16980
rect 3350 16910 3360 16980
rect 3140 16860 3360 16910
rect 3640 16980 3860 17000
rect 3640 16910 3650 16980
rect 3850 16910 3860 16980
rect 3640 16860 3860 16910
rect 4140 16980 4360 17000
rect 4140 16910 4150 16980
rect 4350 16910 4360 16980
rect 4140 16860 4360 16910
rect 4640 16980 4860 17000
rect 4640 16910 4650 16980
rect 4850 16910 4860 16980
rect 4640 16860 4860 16910
rect 5140 16980 5360 17000
rect 5140 16910 5150 16980
rect 5350 16910 5360 16980
rect 5140 16860 5360 16910
rect 5640 16980 5860 17000
rect 5640 16910 5650 16980
rect 5850 16910 5860 16980
rect 5640 16860 5860 16910
rect 6140 16980 6360 17000
rect 6140 16910 6150 16980
rect 6350 16910 6360 16980
rect 6140 16860 6360 16910
rect 6640 16980 6860 17020
rect 6640 16910 6650 16980
rect 6850 16910 6860 16980
rect 6640 16860 6860 16910
rect 7140 17090 7360 17140
rect 7140 17020 7150 17090
rect 7350 17020 7360 17090
rect 7140 16980 7360 17020
rect 13140 17090 13360 17140
rect 13140 17020 13150 17090
rect 13350 17020 13360 17090
rect 7140 16910 7150 16980
rect 7350 16910 7360 16980
rect 7140 16860 7360 16910
rect 7640 16980 7860 17000
rect 7640 16910 7650 16980
rect 7850 16910 7860 16980
rect 7640 16860 7860 16910
rect 8140 16980 8360 17000
rect 8140 16910 8150 16980
rect 8350 16910 8360 16980
rect 8140 16860 8360 16910
rect 8640 16980 8860 17000
rect 8640 16910 8650 16980
rect 8850 16910 8860 16980
rect 8640 16860 8860 16910
rect 9140 16980 9360 17000
rect 9140 16910 9150 16980
rect 9350 16910 9360 16980
rect 9140 16860 9360 16910
rect 9640 16980 9860 17000
rect 9640 16910 9650 16980
rect 9850 16910 9860 16980
rect 9640 16860 9860 16910
rect 10140 16980 10360 17000
rect 10140 16910 10150 16980
rect 10350 16910 10360 16980
rect 10140 16860 10360 16910
rect 10640 16980 10860 17000
rect 10640 16910 10650 16980
rect 10850 16910 10860 16980
rect 10640 16860 10860 16910
rect 11140 16980 11360 17000
rect 11140 16910 11150 16980
rect 11350 16910 11360 16980
rect 11140 16860 11360 16910
rect 11640 16980 11860 17000
rect 11640 16910 11650 16980
rect 11850 16910 11860 16980
rect 11640 16860 11860 16910
rect 12140 16980 12360 17000
rect 12140 16910 12150 16980
rect 12350 16910 12360 16980
rect 12140 16860 12360 16910
rect 12640 16980 12860 17000
rect 12640 16910 12650 16980
rect 12850 16910 12860 16980
rect 12640 16860 12860 16910
rect 13140 16980 13360 17020
rect 13140 16910 13150 16980
rect 13350 16910 13360 16980
rect 13140 16860 13360 16910
rect 13640 17090 13860 17140
rect 13640 17020 13650 17090
rect 13850 17020 13860 17090
rect 13640 16980 13860 17020
rect 19140 17090 19360 17140
rect 19140 17020 19150 17090
rect 19350 17020 19360 17090
rect 13640 16910 13650 16980
rect 13850 16910 13860 16980
rect 13640 16860 13860 16910
rect 14140 16980 14360 17000
rect 14140 16910 14150 16980
rect 14350 16910 14360 16980
rect 14140 16860 14360 16910
rect 14640 16980 14860 17000
rect 14640 16910 14650 16980
rect 14850 16910 14860 16980
rect 14640 16860 14860 16910
rect 15140 16980 15360 17000
rect 15140 16910 15150 16980
rect 15350 16910 15360 16980
rect 15140 16860 15360 16910
rect 15640 16980 15860 17000
rect 15640 16910 15650 16980
rect 15850 16910 15860 16980
rect 15640 16860 15860 16910
rect 16140 16980 16360 17000
rect 16140 16910 16150 16980
rect 16350 16910 16360 16980
rect 16140 16860 16360 16910
rect 16640 16980 16860 17000
rect 16640 16910 16650 16980
rect 16850 16910 16860 16980
rect 16640 16860 16860 16910
rect 17140 16980 17360 17000
rect 17140 16910 17150 16980
rect 17350 16910 17360 16980
rect 17140 16860 17360 16910
rect 17640 16980 17860 17000
rect 17640 16910 17650 16980
rect 17850 16910 17860 16980
rect 17640 16860 17860 16910
rect 18140 16980 18360 17000
rect 18140 16910 18150 16980
rect 18350 16910 18360 16980
rect 18140 16860 18360 16910
rect 18640 16980 18860 17000
rect 18640 16910 18650 16980
rect 18850 16910 18860 16980
rect 18640 16860 18860 16910
rect 19140 16980 19360 17020
rect 19140 16910 19150 16980
rect 19350 16910 19360 16980
rect 19140 16860 19360 16910
rect 19640 17090 19860 17140
rect 19640 17020 19650 17090
rect 19850 17020 19860 17090
rect 19640 16980 19860 17020
rect 25640 17090 25860 17140
rect 25640 17020 25650 17090
rect 25850 17020 25860 17090
rect 19640 16910 19650 16980
rect 19850 16910 19860 16980
rect 19640 16860 19860 16910
rect 20140 16980 20360 17000
rect 20140 16910 20150 16980
rect 20350 16910 20360 16980
rect 20140 16860 20360 16910
rect 20640 16980 20860 17000
rect 20640 16910 20650 16980
rect 20850 16910 20860 16980
rect 20640 16860 20860 16910
rect 21140 16980 21360 17000
rect 21140 16910 21150 16980
rect 21350 16910 21360 16980
rect 21140 16860 21360 16910
rect 21640 16980 21860 17000
rect 21640 16910 21650 16980
rect 21850 16910 21860 16980
rect 21640 16860 21860 16910
rect 22140 16980 22360 17000
rect 22140 16910 22150 16980
rect 22350 16910 22360 16980
rect 22140 16860 22360 16910
rect 22640 16980 22860 17000
rect 22640 16910 22650 16980
rect 22850 16910 22860 16980
rect 22640 16860 22860 16910
rect 23140 16980 23360 17000
rect 23140 16910 23150 16980
rect 23350 16910 23360 16980
rect 23140 16860 23360 16910
rect 23640 16980 23860 17000
rect 23640 16910 23650 16980
rect 23850 16910 23860 16980
rect 23640 16860 23860 16910
rect 24140 16980 24360 17000
rect 24140 16910 24150 16980
rect 24350 16910 24360 16980
rect 24140 16860 24360 16910
rect 24640 16980 24860 17000
rect 24640 16910 24650 16980
rect 24850 16910 24860 16980
rect 24640 16860 24860 16910
rect 25140 16980 25360 17000
rect 25140 16910 25150 16980
rect 25350 16910 25360 16980
rect 25140 16860 25360 16910
rect 25640 16980 25860 17020
rect 25640 16910 25650 16980
rect 25850 16910 25860 16980
rect 25640 16860 25860 16910
rect 26140 17090 26360 17140
rect 26140 17020 26150 17090
rect 26350 17020 26360 17090
rect 26140 16980 26360 17020
rect 26140 16910 26150 16980
rect 26350 16910 26360 16980
rect 26140 16860 26360 16910
rect 0 16850 26500 16860
rect 0 16650 20 16850
rect 90 16650 410 16850
rect 480 16650 520 16850
rect 590 16650 910 16850
rect 980 16650 1020 16850
rect 1090 16650 1410 16850
rect 1480 16650 1520 16850
rect 1590 16650 1910 16850
rect 1980 16650 2020 16850
rect 2090 16650 2410 16850
rect 2480 16650 2520 16850
rect 2590 16650 2910 16850
rect 2980 16650 3020 16850
rect 3090 16650 3410 16850
rect 3480 16650 3520 16850
rect 3590 16650 3910 16850
rect 3980 16650 4020 16850
rect 4090 16650 4410 16850
rect 4480 16650 4520 16850
rect 4590 16650 4910 16850
rect 4980 16650 5020 16850
rect 5090 16650 5410 16850
rect 5480 16650 5520 16850
rect 5590 16650 5910 16850
rect 5980 16650 6020 16850
rect 6090 16650 6410 16850
rect 6480 16650 6520 16850
rect 6590 16650 6910 16850
rect 6980 16650 7020 16850
rect 7090 16650 7410 16850
rect 7480 16650 7520 16850
rect 7590 16650 7910 16850
rect 7980 16650 8020 16850
rect 8090 16650 8410 16850
rect 8480 16650 8520 16850
rect 8590 16650 8910 16850
rect 8980 16650 9020 16850
rect 9090 16650 9410 16850
rect 9480 16650 9520 16850
rect 9590 16650 9910 16850
rect 9980 16650 10020 16850
rect 10090 16650 10410 16850
rect 10480 16650 10520 16850
rect 10590 16650 10910 16850
rect 10980 16650 11020 16850
rect 11090 16650 11410 16850
rect 11480 16650 11520 16850
rect 11590 16650 11910 16850
rect 11980 16650 12020 16850
rect 12090 16650 12410 16850
rect 12480 16650 12520 16850
rect 12590 16650 12910 16850
rect 12980 16650 13020 16850
rect 13090 16650 13410 16850
rect 13480 16650 13520 16850
rect 13590 16650 13910 16850
rect 13980 16650 14020 16850
rect 14090 16650 14410 16850
rect 14480 16650 14520 16850
rect 14590 16650 14910 16850
rect 14980 16650 15020 16850
rect 15090 16650 15410 16850
rect 15480 16650 15520 16850
rect 15590 16650 15910 16850
rect 15980 16650 16020 16850
rect 16090 16650 16410 16850
rect 16480 16650 16520 16850
rect 16590 16650 16910 16850
rect 16980 16650 17020 16850
rect 17090 16650 17410 16850
rect 17480 16650 17520 16850
rect 17590 16650 17910 16850
rect 17980 16650 18020 16850
rect 18090 16650 18410 16850
rect 18480 16650 18520 16850
rect 18590 16650 18910 16850
rect 18980 16650 19020 16850
rect 19090 16650 19410 16850
rect 19480 16650 19520 16850
rect 19590 16650 19910 16850
rect 19980 16650 20020 16850
rect 20090 16650 20410 16850
rect 20480 16650 20520 16850
rect 20590 16650 20910 16850
rect 20980 16650 21020 16850
rect 21090 16650 21410 16850
rect 21480 16650 21520 16850
rect 21590 16650 21910 16850
rect 21980 16650 22020 16850
rect 22090 16650 22410 16850
rect 22480 16650 22520 16850
rect 22590 16650 22910 16850
rect 22980 16650 23020 16850
rect 23090 16650 23410 16850
rect 23480 16650 23520 16850
rect 23590 16650 23910 16850
rect 23980 16650 24020 16850
rect 24090 16650 24410 16850
rect 24480 16650 24520 16850
rect 24590 16650 24910 16850
rect 24980 16650 25020 16850
rect 25090 16650 25410 16850
rect 25480 16650 25520 16850
rect 25590 16650 25910 16850
rect 25980 16650 26020 16850
rect 26090 16650 26410 16850
rect 26480 16650 26500 16850
rect 0 16640 26500 16650
rect 140 16590 360 16640
rect 140 16520 150 16590
rect 350 16520 360 16590
rect 140 16480 360 16520
rect 140 16410 150 16480
rect 350 16410 360 16480
rect 140 16360 360 16410
rect 640 16590 860 16640
rect 640 16520 650 16590
rect 850 16520 860 16590
rect 640 16480 860 16520
rect 640 16410 650 16480
rect 850 16410 860 16480
rect 640 16360 860 16410
rect 1140 16590 1360 16640
rect 1140 16520 1150 16590
rect 1350 16520 1360 16590
rect 1140 16480 1360 16520
rect 1140 16410 1150 16480
rect 1350 16410 1360 16480
rect 1140 16360 1360 16410
rect 1640 16590 1860 16640
rect 1640 16520 1650 16590
rect 1850 16520 1860 16590
rect 1640 16480 1860 16520
rect 1640 16410 1650 16480
rect 1850 16410 1860 16480
rect 1640 16360 1860 16410
rect 2140 16590 2360 16640
rect 2140 16520 2150 16590
rect 2350 16520 2360 16590
rect 2140 16480 2360 16520
rect 2140 16410 2150 16480
rect 2350 16410 2360 16480
rect 2140 16360 2360 16410
rect 2640 16590 2860 16640
rect 2640 16520 2650 16590
rect 2850 16520 2860 16590
rect 2640 16480 2860 16520
rect 2640 16410 2650 16480
rect 2850 16410 2860 16480
rect 2640 16360 2860 16410
rect 3140 16590 3360 16640
rect 3140 16520 3150 16590
rect 3350 16520 3360 16590
rect 3140 16480 3360 16520
rect 3140 16410 3150 16480
rect 3350 16410 3360 16480
rect 3140 16360 3360 16410
rect 3640 16590 3860 16640
rect 3640 16520 3650 16590
rect 3850 16520 3860 16590
rect 3640 16480 3860 16520
rect 3640 16410 3650 16480
rect 3850 16410 3860 16480
rect 3640 16360 3860 16410
rect 4140 16590 4360 16640
rect 4140 16520 4150 16590
rect 4350 16520 4360 16590
rect 4140 16480 4360 16520
rect 4140 16410 4150 16480
rect 4350 16410 4360 16480
rect 4140 16360 4360 16410
rect 4640 16590 4860 16640
rect 4640 16520 4650 16590
rect 4850 16520 4860 16590
rect 4640 16480 4860 16520
rect 4640 16410 4650 16480
rect 4850 16410 4860 16480
rect 4640 16360 4860 16410
rect 5140 16590 5360 16640
rect 5140 16520 5150 16590
rect 5350 16520 5360 16590
rect 5140 16480 5360 16520
rect 5140 16410 5150 16480
rect 5350 16410 5360 16480
rect 5140 16360 5360 16410
rect 5640 16590 5860 16640
rect 5640 16520 5650 16590
rect 5850 16520 5860 16590
rect 5640 16480 5860 16520
rect 5640 16410 5650 16480
rect 5850 16410 5860 16480
rect 5640 16360 5860 16410
rect 6140 16590 6360 16640
rect 6140 16520 6150 16590
rect 6350 16520 6360 16590
rect 6140 16480 6360 16520
rect 6140 16410 6150 16480
rect 6350 16410 6360 16480
rect 6140 16360 6360 16410
rect 6640 16590 6860 16640
rect 6640 16520 6650 16590
rect 6850 16520 6860 16590
rect 6640 16480 6860 16520
rect 6640 16410 6650 16480
rect 6850 16410 6860 16480
rect 6640 16360 6860 16410
rect 7140 16590 7360 16640
rect 7140 16520 7150 16590
rect 7350 16520 7360 16590
rect 7140 16480 7360 16520
rect 7140 16410 7150 16480
rect 7350 16410 7360 16480
rect 7140 16360 7360 16410
rect 7640 16590 7860 16640
rect 7640 16520 7650 16590
rect 7850 16520 7860 16590
rect 7640 16480 7860 16520
rect 7640 16410 7650 16480
rect 7850 16410 7860 16480
rect 7640 16360 7860 16410
rect 8140 16590 8360 16640
rect 8140 16520 8150 16590
rect 8350 16520 8360 16590
rect 8140 16480 8360 16520
rect 8140 16410 8150 16480
rect 8350 16410 8360 16480
rect 8140 16360 8360 16410
rect 8640 16590 8860 16640
rect 8640 16520 8650 16590
rect 8850 16520 8860 16590
rect 8640 16480 8860 16520
rect 8640 16410 8650 16480
rect 8850 16410 8860 16480
rect 8640 16360 8860 16410
rect 9140 16590 9360 16640
rect 9140 16520 9150 16590
rect 9350 16520 9360 16590
rect 9140 16480 9360 16520
rect 9140 16410 9150 16480
rect 9350 16410 9360 16480
rect 9140 16360 9360 16410
rect 9640 16590 9860 16640
rect 9640 16520 9650 16590
rect 9850 16520 9860 16590
rect 9640 16480 9860 16520
rect 9640 16410 9650 16480
rect 9850 16410 9860 16480
rect 9640 16360 9860 16410
rect 10140 16590 10360 16640
rect 10140 16520 10150 16590
rect 10350 16520 10360 16590
rect 10140 16480 10360 16520
rect 10140 16410 10150 16480
rect 10350 16410 10360 16480
rect 10140 16360 10360 16410
rect 10640 16590 10860 16640
rect 10640 16520 10650 16590
rect 10850 16520 10860 16590
rect 10640 16480 10860 16520
rect 10640 16410 10650 16480
rect 10850 16410 10860 16480
rect 10640 16360 10860 16410
rect 11140 16590 11360 16640
rect 11140 16520 11150 16590
rect 11350 16520 11360 16590
rect 11140 16480 11360 16520
rect 11140 16410 11150 16480
rect 11350 16410 11360 16480
rect 11140 16360 11360 16410
rect 11640 16590 11860 16640
rect 11640 16520 11650 16590
rect 11850 16520 11860 16590
rect 11640 16480 11860 16520
rect 11640 16410 11650 16480
rect 11850 16410 11860 16480
rect 11640 16360 11860 16410
rect 12140 16590 12360 16640
rect 12140 16520 12150 16590
rect 12350 16520 12360 16590
rect 12140 16480 12360 16520
rect 12140 16410 12150 16480
rect 12350 16410 12360 16480
rect 12140 16360 12360 16410
rect 12640 16590 12860 16640
rect 12640 16520 12650 16590
rect 12850 16520 12860 16590
rect 12640 16480 12860 16520
rect 12640 16410 12650 16480
rect 12850 16410 12860 16480
rect 12640 16360 12860 16410
rect 13140 16590 13360 16640
rect 13140 16520 13150 16590
rect 13350 16520 13360 16590
rect 13140 16480 13360 16520
rect 13140 16410 13150 16480
rect 13350 16410 13360 16480
rect 13140 16360 13360 16410
rect 13640 16590 13860 16640
rect 13640 16520 13650 16590
rect 13850 16520 13860 16590
rect 13640 16480 13860 16520
rect 13640 16410 13650 16480
rect 13850 16410 13860 16480
rect 13640 16360 13860 16410
rect 14140 16590 14360 16640
rect 14140 16520 14150 16590
rect 14350 16520 14360 16590
rect 14140 16480 14360 16520
rect 14140 16410 14150 16480
rect 14350 16410 14360 16480
rect 14140 16360 14360 16410
rect 14640 16590 14860 16640
rect 14640 16520 14650 16590
rect 14850 16520 14860 16590
rect 14640 16480 14860 16520
rect 14640 16410 14650 16480
rect 14850 16410 14860 16480
rect 14640 16360 14860 16410
rect 15140 16590 15360 16640
rect 15140 16520 15150 16590
rect 15350 16520 15360 16590
rect 15140 16480 15360 16520
rect 15140 16410 15150 16480
rect 15350 16410 15360 16480
rect 15140 16360 15360 16410
rect 15640 16590 15860 16640
rect 15640 16520 15650 16590
rect 15850 16520 15860 16590
rect 15640 16480 15860 16520
rect 15640 16410 15650 16480
rect 15850 16410 15860 16480
rect 15640 16360 15860 16410
rect 16140 16590 16360 16640
rect 16140 16520 16150 16590
rect 16350 16520 16360 16590
rect 16140 16480 16360 16520
rect 16140 16410 16150 16480
rect 16350 16410 16360 16480
rect 16140 16360 16360 16410
rect 16640 16590 16860 16640
rect 16640 16520 16650 16590
rect 16850 16520 16860 16590
rect 16640 16480 16860 16520
rect 16640 16410 16650 16480
rect 16850 16410 16860 16480
rect 16640 16360 16860 16410
rect 17140 16590 17360 16640
rect 17140 16520 17150 16590
rect 17350 16520 17360 16590
rect 17140 16480 17360 16520
rect 17140 16410 17150 16480
rect 17350 16410 17360 16480
rect 17140 16360 17360 16410
rect 17640 16590 17860 16640
rect 17640 16520 17650 16590
rect 17850 16520 17860 16590
rect 17640 16480 17860 16520
rect 17640 16410 17650 16480
rect 17850 16410 17860 16480
rect 17640 16360 17860 16410
rect 18140 16590 18360 16640
rect 18140 16520 18150 16590
rect 18350 16520 18360 16590
rect 18140 16480 18360 16520
rect 18140 16410 18150 16480
rect 18350 16410 18360 16480
rect 18140 16360 18360 16410
rect 18640 16590 18860 16640
rect 18640 16520 18650 16590
rect 18850 16520 18860 16590
rect 18640 16480 18860 16520
rect 18640 16410 18650 16480
rect 18850 16410 18860 16480
rect 18640 16360 18860 16410
rect 19140 16590 19360 16640
rect 19140 16520 19150 16590
rect 19350 16520 19360 16590
rect 19140 16480 19360 16520
rect 19140 16410 19150 16480
rect 19350 16410 19360 16480
rect 19140 16360 19360 16410
rect 19640 16590 19860 16640
rect 19640 16520 19650 16590
rect 19850 16520 19860 16590
rect 19640 16480 19860 16520
rect 19640 16410 19650 16480
rect 19850 16410 19860 16480
rect 19640 16360 19860 16410
rect 20140 16590 20360 16640
rect 20140 16520 20150 16590
rect 20350 16520 20360 16590
rect 20140 16480 20360 16520
rect 20140 16410 20150 16480
rect 20350 16410 20360 16480
rect 20140 16360 20360 16410
rect 20640 16590 20860 16640
rect 20640 16520 20650 16590
rect 20850 16520 20860 16590
rect 20640 16480 20860 16520
rect 20640 16410 20650 16480
rect 20850 16410 20860 16480
rect 20640 16360 20860 16410
rect 21140 16590 21360 16640
rect 21140 16520 21150 16590
rect 21350 16520 21360 16590
rect 21140 16480 21360 16520
rect 21140 16410 21150 16480
rect 21350 16410 21360 16480
rect 21140 16360 21360 16410
rect 21640 16590 21860 16640
rect 21640 16520 21650 16590
rect 21850 16520 21860 16590
rect 21640 16480 21860 16520
rect 21640 16410 21650 16480
rect 21850 16410 21860 16480
rect 21640 16360 21860 16410
rect 22140 16590 22360 16640
rect 22140 16520 22150 16590
rect 22350 16520 22360 16590
rect 22140 16480 22360 16520
rect 22140 16410 22150 16480
rect 22350 16410 22360 16480
rect 22140 16360 22360 16410
rect 22640 16590 22860 16640
rect 22640 16520 22650 16590
rect 22850 16520 22860 16590
rect 22640 16480 22860 16520
rect 22640 16410 22650 16480
rect 22850 16410 22860 16480
rect 22640 16360 22860 16410
rect 23140 16590 23360 16640
rect 23140 16520 23150 16590
rect 23350 16520 23360 16590
rect 23140 16480 23360 16520
rect 23140 16410 23150 16480
rect 23350 16410 23360 16480
rect 23140 16360 23360 16410
rect 23640 16590 23860 16640
rect 23640 16520 23650 16590
rect 23850 16520 23860 16590
rect 23640 16480 23860 16520
rect 23640 16410 23650 16480
rect 23850 16410 23860 16480
rect 23640 16360 23860 16410
rect 24140 16590 24360 16640
rect 24140 16520 24150 16590
rect 24350 16520 24360 16590
rect 24140 16480 24360 16520
rect 24140 16410 24150 16480
rect 24350 16410 24360 16480
rect 24140 16360 24360 16410
rect 24640 16590 24860 16640
rect 24640 16520 24650 16590
rect 24850 16520 24860 16590
rect 24640 16480 24860 16520
rect 24640 16410 24650 16480
rect 24850 16410 24860 16480
rect 24640 16360 24860 16410
rect 25140 16590 25360 16640
rect 25140 16520 25150 16590
rect 25350 16520 25360 16590
rect 25140 16480 25360 16520
rect 25140 16410 25150 16480
rect 25350 16410 25360 16480
rect 25140 16360 25360 16410
rect 25640 16590 25860 16640
rect 25640 16520 25650 16590
rect 25850 16520 25860 16590
rect 25640 16480 25860 16520
rect 25640 16410 25650 16480
rect 25850 16410 25860 16480
rect 25640 16360 25860 16410
rect 26140 16590 26360 16640
rect 26140 16520 26150 16590
rect 26350 16520 26360 16590
rect 26140 16480 26360 16520
rect 26140 16410 26150 16480
rect 26350 16410 26360 16480
rect 26140 16360 26360 16410
rect 0 16350 26500 16360
rect 0 16150 20 16350
rect 90 16150 410 16350
rect 480 16150 520 16350
rect 590 16150 910 16350
rect 980 16150 1020 16350
rect 1090 16150 1410 16350
rect 1480 16150 1520 16350
rect 1590 16150 1910 16350
rect 1980 16150 2020 16350
rect 2090 16150 2410 16350
rect 2480 16150 2520 16350
rect 2590 16150 2910 16350
rect 2980 16150 3020 16350
rect 3090 16150 3410 16350
rect 3480 16150 3520 16350
rect 3590 16150 3910 16350
rect 3980 16150 4020 16350
rect 4090 16150 4410 16350
rect 4480 16150 4520 16350
rect 4590 16150 4910 16350
rect 4980 16150 5020 16350
rect 5090 16150 5410 16350
rect 5480 16150 5520 16350
rect 5590 16150 5910 16350
rect 5980 16150 6020 16350
rect 6090 16150 6410 16350
rect 6480 16150 6520 16350
rect 6590 16150 6910 16350
rect 6980 16150 7020 16350
rect 7090 16150 7410 16350
rect 7480 16150 7520 16350
rect 7590 16150 7910 16350
rect 7980 16150 8020 16350
rect 8090 16150 8410 16350
rect 8480 16150 8520 16350
rect 8590 16150 8910 16350
rect 8980 16150 9020 16350
rect 9090 16150 9410 16350
rect 9480 16150 9520 16350
rect 9590 16150 9910 16350
rect 9980 16150 10020 16350
rect 10090 16150 10410 16350
rect 10480 16150 10520 16350
rect 10590 16150 10910 16350
rect 10980 16150 11020 16350
rect 11090 16150 11410 16350
rect 11480 16150 11520 16350
rect 11590 16150 11910 16350
rect 11980 16150 12020 16350
rect 12090 16150 12410 16350
rect 12480 16150 12520 16350
rect 12590 16150 12910 16350
rect 12980 16150 13020 16350
rect 13090 16150 13410 16350
rect 13480 16150 13520 16350
rect 13590 16150 13910 16350
rect 13980 16150 14020 16350
rect 14090 16150 14410 16350
rect 14480 16150 14520 16350
rect 14590 16150 14910 16350
rect 14980 16150 15020 16350
rect 15090 16150 15410 16350
rect 15480 16150 15520 16350
rect 15590 16150 15910 16350
rect 15980 16150 16020 16350
rect 16090 16150 16410 16350
rect 16480 16150 16520 16350
rect 16590 16150 16910 16350
rect 16980 16150 17020 16350
rect 17090 16150 17410 16350
rect 17480 16150 17520 16350
rect 17590 16150 17910 16350
rect 17980 16150 18020 16350
rect 18090 16150 18410 16350
rect 18480 16150 18520 16350
rect 18590 16150 18910 16350
rect 18980 16150 19020 16350
rect 19090 16150 19410 16350
rect 19480 16150 19520 16350
rect 19590 16150 19910 16350
rect 19980 16150 20020 16350
rect 20090 16150 20410 16350
rect 20480 16150 20520 16350
rect 20590 16150 20910 16350
rect 20980 16150 21020 16350
rect 21090 16150 21410 16350
rect 21480 16150 21520 16350
rect 21590 16150 21910 16350
rect 21980 16150 22020 16350
rect 22090 16150 22410 16350
rect 22480 16150 22520 16350
rect 22590 16150 22910 16350
rect 22980 16150 23020 16350
rect 23090 16150 23410 16350
rect 23480 16150 23520 16350
rect 23590 16150 23910 16350
rect 23980 16150 24020 16350
rect 24090 16150 24410 16350
rect 24480 16150 24520 16350
rect 24590 16150 24910 16350
rect 24980 16150 25020 16350
rect 25090 16150 25410 16350
rect 25480 16150 25520 16350
rect 25590 16150 25910 16350
rect 25980 16150 26020 16350
rect 26090 16150 26410 16350
rect 26480 16150 26500 16350
rect 0 16140 26500 16150
rect 140 16090 360 16140
rect 140 16020 150 16090
rect 350 16020 360 16090
rect 140 15980 360 16020
rect 140 15910 150 15980
rect 350 15910 360 15980
rect 140 15860 360 15910
rect 640 16090 860 16140
rect 640 16020 650 16090
rect 850 16020 860 16090
rect 640 15980 860 16020
rect 1140 16090 1360 16140
rect 1140 16020 1150 16090
rect 1350 16020 1360 16090
rect 1140 16000 1360 16020
rect 1640 16090 1860 16140
rect 1640 16020 1650 16090
rect 1850 16020 1860 16090
rect 1640 16000 1860 16020
rect 2140 16090 2360 16140
rect 2140 16020 2150 16090
rect 2350 16020 2360 16090
rect 2140 16000 2360 16020
rect 2640 16090 2860 16140
rect 2640 16020 2650 16090
rect 2850 16020 2860 16090
rect 2640 16000 2860 16020
rect 3140 16090 3360 16140
rect 3140 16020 3150 16090
rect 3350 16020 3360 16090
rect 3140 16000 3360 16020
rect 3640 16090 3860 16140
rect 3640 16020 3650 16090
rect 3850 16020 3860 16090
rect 3640 16000 3860 16020
rect 4140 16090 4360 16140
rect 4140 16020 4150 16090
rect 4350 16020 4360 16090
rect 4140 16000 4360 16020
rect 4640 16090 4860 16140
rect 4640 16020 4650 16090
rect 4850 16020 4860 16090
rect 4640 16000 4860 16020
rect 5140 16090 5360 16140
rect 5140 16020 5150 16090
rect 5350 16020 5360 16090
rect 5140 16000 5360 16020
rect 5640 16090 5860 16140
rect 5640 16020 5650 16090
rect 5850 16020 5860 16090
rect 5640 16000 5860 16020
rect 6140 16090 6360 16140
rect 6140 16020 6150 16090
rect 6350 16020 6360 16090
rect 6140 16000 6360 16020
rect 6640 16090 6860 16140
rect 6640 16020 6650 16090
rect 6850 16020 6860 16090
rect 640 15910 650 15980
rect 850 15910 860 15980
rect 640 15860 860 15910
rect 6640 15980 6860 16020
rect 6640 15910 6650 15980
rect 6850 15910 6860 15980
rect 6640 15860 6860 15910
rect 7140 16090 7360 16140
rect 7140 16020 7150 16090
rect 7350 16020 7360 16090
rect 7140 15980 7360 16020
rect 7640 16090 7860 16140
rect 7640 16020 7650 16090
rect 7850 16020 7860 16090
rect 7640 16000 7860 16020
rect 8140 16090 8360 16140
rect 8140 16020 8150 16090
rect 8350 16020 8360 16090
rect 8140 16000 8360 16020
rect 8640 16090 8860 16140
rect 8640 16020 8650 16090
rect 8850 16020 8860 16090
rect 8640 16000 8860 16020
rect 9140 16090 9360 16140
rect 9140 16020 9150 16090
rect 9350 16020 9360 16090
rect 9140 16000 9360 16020
rect 9640 16090 9860 16140
rect 9640 16020 9650 16090
rect 9850 16020 9860 16090
rect 9640 16000 9860 16020
rect 10140 16090 10360 16140
rect 10140 16020 10150 16090
rect 10350 16020 10360 16090
rect 10140 16000 10360 16020
rect 10640 16090 10860 16140
rect 10640 16020 10650 16090
rect 10850 16020 10860 16090
rect 10640 16000 10860 16020
rect 11140 16090 11360 16140
rect 11140 16020 11150 16090
rect 11350 16020 11360 16090
rect 11140 16000 11360 16020
rect 11640 16090 11860 16140
rect 11640 16020 11650 16090
rect 11850 16020 11860 16090
rect 11640 16000 11860 16020
rect 12140 16090 12360 16140
rect 12140 16020 12150 16090
rect 12350 16020 12360 16090
rect 12140 16000 12360 16020
rect 12640 16090 12860 16140
rect 12640 16020 12650 16090
rect 12850 16020 12860 16090
rect 12640 16000 12860 16020
rect 13140 16090 13360 16140
rect 13140 16020 13150 16090
rect 13350 16020 13360 16090
rect 7140 15910 7150 15980
rect 7350 15910 7360 15980
rect 7140 15860 7360 15910
rect 13140 15980 13360 16020
rect 13140 15910 13150 15980
rect 13350 15910 13360 15980
rect 13140 15860 13360 15910
rect 13640 16090 13860 16140
rect 13640 16020 13650 16090
rect 13850 16020 13860 16090
rect 13640 15980 13860 16020
rect 14140 16090 14360 16140
rect 14140 16020 14150 16090
rect 14350 16020 14360 16090
rect 14140 16000 14360 16020
rect 14640 16090 14860 16140
rect 14640 16020 14650 16090
rect 14850 16020 14860 16090
rect 14640 16000 14860 16020
rect 15140 16090 15360 16140
rect 15140 16020 15150 16090
rect 15350 16020 15360 16090
rect 15140 16000 15360 16020
rect 15640 16090 15860 16140
rect 15640 16020 15650 16090
rect 15850 16020 15860 16090
rect 15640 16000 15860 16020
rect 16140 16090 16360 16140
rect 16140 16020 16150 16090
rect 16350 16020 16360 16090
rect 16140 16000 16360 16020
rect 16640 16090 16860 16140
rect 16640 16020 16650 16090
rect 16850 16020 16860 16090
rect 16640 16000 16860 16020
rect 17140 16090 17360 16140
rect 17140 16020 17150 16090
rect 17350 16020 17360 16090
rect 17140 16000 17360 16020
rect 17640 16090 17860 16140
rect 17640 16020 17650 16090
rect 17850 16020 17860 16090
rect 17640 16000 17860 16020
rect 18140 16090 18360 16140
rect 18140 16020 18150 16090
rect 18350 16020 18360 16090
rect 18140 16000 18360 16020
rect 18640 16090 18860 16140
rect 18640 16020 18650 16090
rect 18850 16020 18860 16090
rect 18640 16000 18860 16020
rect 19140 16090 19360 16140
rect 19140 16020 19150 16090
rect 19350 16020 19360 16090
rect 13640 15910 13650 15980
rect 13850 15910 13860 15980
rect 13640 15860 13860 15910
rect 19140 15980 19360 16020
rect 19140 15910 19150 15980
rect 19350 15910 19360 15980
rect 19140 15860 19360 15910
rect 19640 16090 19860 16140
rect 19640 16020 19650 16090
rect 19850 16020 19860 16090
rect 19640 15980 19860 16020
rect 20140 16090 20360 16140
rect 20140 16020 20150 16090
rect 20350 16020 20360 16090
rect 20140 16000 20360 16020
rect 20640 16090 20860 16140
rect 20640 16020 20650 16090
rect 20850 16020 20860 16090
rect 20640 16000 20860 16020
rect 21140 16090 21360 16140
rect 21140 16020 21150 16090
rect 21350 16020 21360 16090
rect 21140 16000 21360 16020
rect 21640 16090 21860 16140
rect 21640 16020 21650 16090
rect 21850 16020 21860 16090
rect 21640 16000 21860 16020
rect 22140 16090 22360 16140
rect 22140 16020 22150 16090
rect 22350 16020 22360 16090
rect 22140 16000 22360 16020
rect 22640 16090 22860 16140
rect 22640 16020 22650 16090
rect 22850 16020 22860 16090
rect 22640 16000 22860 16020
rect 23140 16090 23360 16140
rect 23140 16020 23150 16090
rect 23350 16020 23360 16090
rect 23140 16000 23360 16020
rect 23640 16090 23860 16140
rect 23640 16020 23650 16090
rect 23850 16020 23860 16090
rect 23640 16000 23860 16020
rect 24140 16090 24360 16140
rect 24140 16020 24150 16090
rect 24350 16020 24360 16090
rect 24140 16000 24360 16020
rect 24640 16090 24860 16140
rect 24640 16020 24650 16090
rect 24850 16020 24860 16090
rect 24640 16000 24860 16020
rect 25140 16090 25360 16140
rect 25140 16020 25150 16090
rect 25350 16020 25360 16090
rect 25140 16000 25360 16020
rect 25640 16090 25860 16140
rect 25640 16020 25650 16090
rect 25850 16020 25860 16090
rect 19640 15910 19650 15980
rect 19850 15910 19860 15980
rect 19640 15860 19860 15910
rect 25640 15980 25860 16020
rect 25640 15910 25650 15980
rect 25850 15910 25860 15980
rect 25640 15860 25860 15910
rect 26140 16090 26360 16140
rect 26140 16020 26150 16090
rect 26350 16020 26360 16090
rect 26140 15980 26360 16020
rect 26140 15910 26150 15980
rect 26350 15910 26360 15980
rect 26140 15860 26360 15910
rect 0 15850 1000 15860
rect 0 15650 20 15850
rect 90 15650 410 15850
rect 480 15650 520 15850
rect 590 15650 910 15850
rect 980 15650 1000 15850
rect 0 15640 1000 15650
rect 6500 15850 7500 15860
rect 6500 15650 6520 15850
rect 6590 15650 6910 15850
rect 6980 15650 7020 15850
rect 7090 15650 7410 15850
rect 7480 15650 7500 15850
rect 13000 15850 14000 15860
rect 13000 15700 13020 15850
rect 6500 15640 7500 15650
rect 12700 15650 13020 15700
rect 13090 15650 13410 15850
rect 13480 15650 13520 15850
rect 13590 15650 13910 15850
rect 13980 15650 14000 15850
rect 140 15590 360 15640
rect 140 15520 150 15590
rect 350 15520 360 15590
rect 140 15480 360 15520
rect 140 15410 150 15480
rect 350 15410 360 15480
rect 140 15360 360 15410
rect 640 15590 860 15640
rect 6640 15600 6860 15640
rect 7140 15600 7360 15640
rect 640 15520 650 15590
rect 850 15520 860 15590
rect 6400 15590 7700 15600
rect 6400 15580 6650 15590
rect 640 15480 860 15520
rect 640 15410 650 15480
rect 850 15410 860 15480
rect 640 15360 860 15410
rect 1330 15520 1400 15580
rect 0 15350 1000 15360
rect 0 15150 20 15350
rect 90 15150 410 15350
rect 480 15150 520 15350
rect 590 15150 910 15350
rect 980 15150 1000 15350
rect 0 15140 1000 15150
rect 140 15090 360 15140
rect 140 15020 150 15090
rect 350 15020 360 15090
rect 140 14980 360 15020
rect 140 14910 150 14980
rect 350 14910 360 14980
rect 140 14860 360 14910
rect 640 15090 860 15140
rect 640 15020 650 15090
rect 850 15020 860 15090
rect 640 14980 860 15020
rect 640 14910 650 14980
rect 850 14910 860 14980
rect 640 14860 860 14910
rect 0 14850 1000 14860
rect 0 14650 20 14850
rect 90 14650 410 14850
rect 480 14650 520 14850
rect 590 14650 910 14850
rect 980 14650 1000 14850
rect 0 14640 1000 14650
rect 140 14590 360 14640
rect 140 14520 150 14590
rect 350 14520 360 14590
rect 140 14480 360 14520
rect 140 14410 150 14480
rect 350 14410 360 14480
rect 140 14360 360 14410
rect 640 14590 860 14640
rect 640 14520 650 14590
rect 850 14520 860 14590
rect 640 14480 860 14520
rect 640 14410 650 14480
rect 850 14410 860 14480
rect 640 14360 860 14410
rect 0 14350 1000 14360
rect 0 14150 20 14350
rect 90 14150 410 14350
rect 480 14150 520 14350
rect 590 14150 910 14350
rect 980 14150 1000 14350
rect 0 14140 1000 14150
rect 140 14090 360 14140
rect 140 14020 150 14090
rect 350 14020 360 14090
rect -3860 13980 -3640 14000
rect -3860 13910 -3850 13980
rect -3650 13910 -3640 13980
rect -4300 13900 -4100 13910
rect -4300 13420 -4290 13900
rect -4110 13420 -4100 13900
rect -3860 13860 -3640 13910
rect -3360 13980 -3140 14000
rect -3360 13910 -3350 13980
rect -3150 13910 -3140 13980
rect -3360 13860 -3140 13910
rect -2860 13980 -2640 14000
rect -2860 13910 -2850 13980
rect -2650 13910 -2640 13980
rect -2860 13860 -2640 13910
rect -2360 13980 -2140 14000
rect -2360 13910 -2350 13980
rect -2150 13910 -2140 13980
rect -2360 13860 -2140 13910
rect -1860 13980 -1640 14000
rect -1860 13910 -1850 13980
rect -1650 13910 -1640 13980
rect -1860 13860 -1640 13910
rect -1360 13980 -1140 14000
rect -1360 13910 -1350 13980
rect -1150 13910 -1140 13980
rect -1360 13860 -1140 13910
rect -860 13980 -640 14000
rect -860 13910 -850 13980
rect -650 13910 -640 13980
rect -860 13860 -640 13910
rect -360 13980 -140 14000
rect -360 13910 -350 13980
rect -150 13910 -140 13980
rect -360 13860 -140 13910
rect 140 13980 360 14020
rect 140 13910 150 13980
rect 350 13910 360 13980
rect 140 13860 360 13910
rect 640 14090 860 14140
rect 640 14020 650 14090
rect 850 14020 860 14090
rect 640 13980 860 14020
rect 640 13910 650 13980
rect 850 13910 860 13980
rect 640 13860 860 13910
rect -4000 13850 1000 13860
rect -4000 13650 -3980 13850
rect -3910 13650 -3590 13850
rect -3520 13650 -3480 13850
rect -3410 13650 -3090 13850
rect -3020 13650 -2980 13850
rect -2910 13650 -2590 13850
rect -2520 13650 -2480 13850
rect -2410 13650 -2090 13850
rect -2020 13650 -1980 13850
rect -1910 13650 -1590 13850
rect -1520 13650 -1480 13850
rect -1410 13650 -1090 13850
rect -1020 13650 -980 13850
rect -910 13650 -590 13850
rect -520 13650 -480 13850
rect -410 13650 -90 13850
rect -20 13650 20 13850
rect 90 13650 410 13850
rect 480 13650 520 13850
rect 590 13650 910 13850
rect 980 13650 1000 13850
rect -4000 13640 1000 13650
rect -4300 13410 -4100 13420
rect -3860 13590 -3640 13640
rect -3860 13520 -3850 13590
rect -3650 13520 -3640 13590
rect -3860 13480 -3640 13520
rect -3860 13410 -3850 13480
rect -3650 13410 -3640 13480
rect -3860 13360 -3640 13410
rect -3360 13590 -3140 13640
rect -3360 13520 -3350 13590
rect -3150 13520 -3140 13590
rect -3360 13480 -3140 13520
rect -3360 13410 -3350 13480
rect -3150 13410 -3140 13480
rect -3360 13360 -3140 13410
rect -2860 13590 -2640 13640
rect -2860 13520 -2850 13590
rect -2650 13520 -2640 13590
rect -2860 13480 -2640 13520
rect -2860 13410 -2850 13480
rect -2650 13410 -2640 13480
rect -2860 13360 -2640 13410
rect -2360 13590 -2140 13640
rect -2360 13520 -2350 13590
rect -2150 13520 -2140 13590
rect -2360 13480 -2140 13520
rect -2360 13410 -2350 13480
rect -2150 13410 -2140 13480
rect -2360 13360 -2140 13410
rect -1860 13590 -1640 13640
rect -1860 13520 -1850 13590
rect -1650 13520 -1640 13590
rect -1860 13480 -1640 13520
rect -1860 13410 -1850 13480
rect -1650 13410 -1640 13480
rect -1860 13360 -1640 13410
rect -1360 13590 -1140 13640
rect -1360 13520 -1350 13590
rect -1150 13520 -1140 13590
rect -1360 13480 -1140 13520
rect -1360 13410 -1350 13480
rect -1150 13410 -1140 13480
rect -1360 13360 -1140 13410
rect -860 13590 -640 13640
rect -860 13520 -850 13590
rect -650 13520 -640 13590
rect -860 13480 -640 13520
rect -860 13410 -850 13480
rect -650 13410 -640 13480
rect -860 13360 -640 13410
rect -360 13590 -140 13640
rect -360 13520 -350 13590
rect -150 13520 -140 13590
rect -360 13480 -140 13520
rect -360 13410 -350 13480
rect -150 13410 -140 13480
rect -360 13360 -140 13410
rect 140 13590 360 13640
rect 140 13520 150 13590
rect 350 13520 360 13590
rect 140 13480 360 13520
rect 140 13410 150 13480
rect 350 13410 360 13480
rect 140 13360 360 13410
rect 640 13590 860 13640
rect 640 13520 650 13590
rect 850 13520 860 13590
rect 640 13480 860 13520
rect 640 13410 650 13480
rect 850 13410 860 13480
rect 640 13360 860 13410
rect -4000 13350 1000 13360
rect -4000 13150 -3980 13350
rect -3910 13150 -3590 13350
rect -3520 13150 -3480 13350
rect -3410 13150 -3090 13350
rect -3020 13150 -2980 13350
rect -2910 13150 -2590 13350
rect -2520 13150 -2480 13350
rect -2410 13150 -2090 13350
rect -2020 13150 -1980 13350
rect -1910 13150 -1590 13350
rect -1520 13150 -1480 13350
rect -1410 13150 -1090 13350
rect -1020 13150 -980 13350
rect -910 13150 -590 13350
rect -520 13150 -480 13350
rect -410 13150 -90 13350
rect -20 13150 20 13350
rect 90 13150 410 13350
rect 480 13150 520 13350
rect 590 13150 910 13350
rect 980 13150 1000 13350
rect -4000 13140 1000 13150
rect -4300 13090 -4100 13100
rect -4300 12610 -4290 13090
rect -4110 12610 -4100 13090
rect -3860 13090 -3640 13140
rect -3860 13020 -3850 13090
rect -3650 13020 -3640 13090
rect -3860 13000 -3640 13020
rect -3360 13090 -3140 13140
rect -3360 13020 -3350 13090
rect -3150 13020 -3140 13090
rect -3360 13000 -3140 13020
rect -2860 13090 -2640 13140
rect -2860 13020 -2850 13090
rect -2650 13020 -2640 13090
rect -2860 13000 -2640 13020
rect -2360 13090 -2140 13140
rect -2360 13020 -2350 13090
rect -2150 13020 -2140 13090
rect -2360 13000 -2140 13020
rect -1860 13090 -1640 13140
rect -1860 13020 -1850 13090
rect -1650 13020 -1640 13090
rect -1860 13000 -1640 13020
rect -1360 13090 -1140 13140
rect -1360 13020 -1350 13090
rect -1150 13020 -1140 13090
rect -1360 13000 -1140 13020
rect -860 13090 -640 13140
rect -860 13020 -850 13090
rect -650 13020 -640 13090
rect -860 13000 -640 13020
rect -360 13090 -140 13140
rect -360 13020 -350 13090
rect -150 13020 -140 13090
rect -360 13000 -140 13020
rect 140 13090 360 13140
rect 140 13020 150 13090
rect 350 13020 360 13090
rect 140 12980 360 13020
rect 140 12910 150 12980
rect 350 12910 360 12980
rect 140 12860 360 12910
rect 640 13090 860 13140
rect 640 13020 650 13090
rect 850 13020 860 13090
rect 640 12980 860 13020
rect 640 12910 650 12980
rect 850 12910 860 12980
rect 640 12860 860 12910
rect 0 12850 1000 12860
rect 0 12650 20 12850
rect 90 12650 410 12850
rect 480 12650 520 12850
rect 590 12650 910 12850
rect 980 12650 1000 12850
rect 0 12640 1000 12650
rect -4300 12600 -4100 12610
rect 140 12590 360 12640
rect 140 12520 150 12590
rect 350 12520 360 12590
rect 140 12480 360 12520
rect 140 12410 150 12480
rect 350 12410 360 12480
rect 140 12360 360 12410
rect 640 12590 860 12640
rect 640 12520 650 12590
rect 850 12520 860 12590
rect 640 12480 860 12520
rect 640 12410 650 12480
rect 850 12410 860 12480
rect 640 12360 860 12410
rect 0 12350 1000 12360
rect 0 12150 20 12350
rect 90 12150 410 12350
rect 480 12150 520 12350
rect 590 12150 910 12350
rect 980 12150 1000 12350
rect 0 12140 1000 12150
rect 140 12090 360 12140
rect 140 12020 150 12090
rect 350 12020 360 12090
rect 140 11980 360 12020
rect 140 11910 150 11980
rect 350 11910 360 11980
rect 140 11860 360 11910
rect 640 12090 860 12140
rect 640 12020 650 12090
rect 850 12020 860 12090
rect 640 11980 860 12020
rect 640 11910 650 11980
rect 850 11910 860 11980
rect 640 11860 860 11910
rect 0 11850 1000 11860
rect 0 11650 20 11850
rect 90 11650 410 11850
rect 480 11650 520 11850
rect 590 11650 910 11850
rect 980 11650 1000 11850
rect 0 11640 1000 11650
rect 140 11590 360 11640
rect 140 11520 150 11590
rect 350 11520 360 11590
rect 140 11480 360 11520
rect 140 11410 150 11480
rect 350 11410 360 11480
rect 140 11360 360 11410
rect 640 11590 860 11640
rect 640 11520 650 11590
rect 850 11520 860 11590
rect 640 11480 860 11520
rect 640 11410 650 11480
rect 850 11410 860 11480
rect 640 11360 860 11410
rect 0 11350 1000 11360
rect 0 11150 20 11350
rect 90 11150 410 11350
rect 480 11150 520 11350
rect 590 11150 910 11350
rect 980 11150 1000 11350
rect 0 11140 1000 11150
rect 140 11090 360 11140
rect 140 11020 150 11090
rect 350 11020 360 11090
rect 140 10980 360 11020
rect 140 10910 150 10980
rect 350 10910 360 10980
rect 140 10860 360 10910
rect 640 11090 860 11140
rect 640 11020 650 11090
rect 850 11020 860 11090
rect 640 10980 860 11020
rect 640 10910 650 10980
rect 850 10910 860 10980
rect 640 10860 860 10910
rect 0 10850 1000 10860
rect 0 10650 20 10850
rect 90 10650 410 10850
rect 480 10650 520 10850
rect 590 10650 910 10850
rect 980 10650 1000 10850
rect 0 10640 1000 10650
rect 140 10590 360 10640
rect 140 10520 150 10590
rect 350 10520 360 10590
rect 140 10480 360 10520
rect 140 10410 150 10480
rect 350 10410 360 10480
rect 140 10360 360 10410
rect 640 10590 860 10640
rect 640 10520 650 10590
rect 850 10520 860 10590
rect 640 10480 860 10520
rect 640 10410 650 10480
rect 850 10410 860 10480
rect 640 10360 860 10410
rect 0 10350 1000 10360
rect 0 10150 20 10350
rect 90 10150 410 10350
rect 480 10150 520 10350
rect 590 10150 910 10350
rect 980 10150 1000 10350
rect 0 10140 1000 10150
rect 140 10090 360 10140
rect 140 10020 150 10090
rect 350 10020 360 10090
rect 140 9980 360 10020
rect 140 9910 150 9980
rect 350 9910 360 9980
rect 140 9860 360 9910
rect 640 10090 860 10140
rect 640 10020 650 10090
rect 850 10020 860 10090
rect 640 9980 860 10020
rect 640 9910 650 9980
rect 850 9910 860 9980
rect 640 9860 860 9910
rect 0 9850 1000 9860
rect 0 9650 20 9850
rect 90 9650 410 9850
rect 480 9650 520 9850
rect 590 9650 910 9850
rect 980 9650 1000 9850
rect 0 9640 1000 9650
rect 140 9590 360 9640
rect 140 9520 150 9590
rect 350 9520 360 9590
rect 140 9480 360 9520
rect 140 9410 150 9480
rect 350 9410 360 9480
rect 140 9360 360 9410
rect 640 9590 860 9640
rect 640 9520 650 9590
rect 850 9520 860 9590
rect 640 9480 860 9520
rect 640 9410 650 9480
rect 850 9410 860 9480
rect 640 9360 860 9410
rect 0 9350 1000 9360
rect 0 9150 20 9350
rect 90 9150 410 9350
rect 480 9150 520 9350
rect 590 9150 910 9350
rect 980 9150 1000 9350
rect 0 9140 1000 9150
rect 6340 15520 6650 15580
rect 6850 15520 7150 15590
rect 7350 15520 7700 15590
rect 12700 15590 14000 15650
rect 19000 15850 20000 15860
rect 19000 15650 19020 15850
rect 19090 15650 19410 15850
rect 19480 15650 19520 15850
rect 19590 15650 19910 15850
rect 19980 15650 20000 15850
rect 19000 15640 20000 15650
rect 25500 15850 26500 15860
rect 25500 15650 25520 15850
rect 25590 15650 25910 15850
rect 25980 15650 26020 15850
rect 26090 15650 26410 15850
rect 26480 15650 26500 15850
rect 25500 15640 26500 15650
rect 19140 15600 19360 15640
rect 19640 15600 19860 15640
rect 12700 15580 13150 15590
rect 1532 15480 1552 15490
rect 6186 15480 6206 15490
rect 1532 15410 1540 15480
rect 6200 15410 6206 15480
rect 1532 15390 1552 15410
rect 6186 15390 6206 15410
rect 1465 15338 1531 15358
rect 1465 9358 1531 9378
rect 1623 15338 1689 15358
rect 1623 9358 1689 9378
rect 1781 15338 1847 15358
rect 1781 9358 1847 9378
rect 1939 15338 2005 15358
rect 1939 9358 2005 9378
rect 2097 15338 2163 15358
rect 2097 9358 2163 9378
rect 2255 15338 2321 15358
rect 2255 9358 2321 9378
rect 2413 15338 2479 15358
rect 2413 9358 2479 9378
rect 2571 15338 2637 15358
rect 2571 9358 2637 9378
rect 2729 15338 2795 15358
rect 2729 9358 2795 9378
rect 2887 15338 2953 15358
rect 2887 9358 2953 9378
rect 3045 15338 3111 15358
rect 3045 9358 3111 9378
rect 3203 15338 3269 15358
rect 3203 9358 3269 9378
rect 3361 15338 3427 15358
rect 3361 9358 3427 9378
rect 3519 15338 3585 15358
rect 3519 9358 3585 9378
rect 3677 15338 3743 15358
rect 3677 9358 3743 9378
rect 3835 15338 3901 15358
rect 3835 9358 3901 9378
rect 3993 15338 4059 15358
rect 3993 9358 4059 9378
rect 4151 15338 4217 15358
rect 4151 9358 4217 9378
rect 4309 15338 4375 15358
rect 4309 9358 4375 9378
rect 4467 15338 4533 15358
rect 4467 9358 4533 9378
rect 4625 15338 4691 15358
rect 4625 9358 4691 9378
rect 4783 15338 4849 15358
rect 4783 9358 4849 9378
rect 4941 15338 5007 15358
rect 4941 9358 5007 9378
rect 5099 15338 5165 15358
rect 5099 9358 5165 9378
rect 5257 15338 5323 15358
rect 5257 9358 5323 9378
rect 5415 15338 5481 15358
rect 5415 9358 5481 9378
rect 5573 15338 5639 15358
rect 5573 9358 5639 9378
rect 5731 15338 5797 15358
rect 5731 9358 5797 9378
rect 5889 15338 5955 15358
rect 5889 9358 5955 9378
rect 6047 15338 6113 15358
rect 6047 9358 6113 9378
rect 6205 15338 6271 15358
rect 6205 9358 6271 9378
rect 1532 9310 1552 9326
rect 6186 9310 6206 9326
rect 1532 9240 1540 9310
rect 6190 9240 6206 9310
rect 1532 9226 1552 9240
rect 6186 9226 6206 9240
rect 140 9090 360 9140
rect 140 9020 150 9090
rect 350 9020 360 9090
rect 140 8980 360 9020
rect 140 8910 150 8980
rect 350 8910 360 8980
rect 140 8860 360 8910
rect 640 9090 860 9140
rect 1330 9130 1400 9200
rect 6410 15200 7630 15520
rect 6410 14600 7630 15000
rect 6410 14000 7630 14400
rect 6410 13400 7630 13800
rect 6410 12800 7630 13200
rect 6410 12200 7630 12600
rect 6410 11600 7630 12000
rect 6410 11000 7630 11400
rect 6410 10400 7630 10800
rect 6410 9800 7630 10200
rect 6410 9200 7630 9600
rect 12640 15520 13150 15580
rect 13350 15520 13650 15590
rect 13850 15520 14000 15590
rect 19000 15590 20300 15600
rect 19000 15580 19150 15590
rect 7832 15480 7852 15490
rect 12486 15480 12506 15490
rect 7832 15410 7840 15480
rect 12500 15410 12506 15480
rect 7832 15390 7852 15410
rect 12486 15390 12506 15410
rect 7765 15338 7831 15358
rect 7765 9358 7831 9378
rect 7923 15338 7989 15358
rect 7923 9358 7989 9378
rect 8081 15338 8147 15358
rect 8081 9358 8147 9378
rect 8239 15338 8305 15358
rect 8239 9358 8305 9378
rect 8397 15338 8463 15358
rect 8397 9358 8463 9378
rect 8555 15338 8621 15358
rect 8555 9358 8621 9378
rect 8713 15338 8779 15358
rect 8713 9358 8779 9378
rect 8871 15338 8937 15358
rect 8871 9358 8937 9378
rect 9029 15338 9095 15358
rect 9029 9358 9095 9378
rect 9187 15338 9253 15358
rect 9187 9358 9253 9378
rect 9345 15338 9411 15358
rect 9345 9358 9411 9378
rect 9503 15338 9569 15358
rect 9503 9358 9569 9378
rect 9661 15338 9727 15358
rect 9661 9358 9727 9378
rect 9819 15338 9885 15358
rect 9819 9358 9885 9378
rect 9977 15338 10043 15358
rect 9977 9358 10043 9378
rect 10135 15338 10201 15358
rect 10135 9358 10201 9378
rect 10293 15338 10359 15358
rect 10293 9358 10359 9378
rect 10451 15338 10517 15358
rect 10451 9358 10517 9378
rect 10609 15338 10675 15358
rect 10609 9358 10675 9378
rect 10767 15338 10833 15358
rect 10767 9358 10833 9378
rect 10925 15338 10991 15358
rect 10925 9358 10991 9378
rect 11083 15338 11149 15358
rect 11083 9358 11149 9378
rect 11241 15338 11307 15358
rect 11241 9358 11307 9378
rect 11399 15338 11465 15358
rect 11399 9358 11465 9378
rect 11557 15338 11623 15358
rect 11557 9358 11623 9378
rect 11715 15338 11781 15358
rect 11715 9358 11781 9378
rect 11873 15338 11939 15358
rect 11873 9358 11939 9378
rect 12031 15338 12097 15358
rect 12031 9358 12097 9378
rect 12189 15338 12255 15358
rect 12189 9358 12255 9378
rect 12347 15338 12413 15358
rect 12347 9358 12413 9378
rect 12505 15338 12571 15358
rect 12505 9358 12571 9378
rect 7832 9310 7852 9326
rect 12486 9310 12506 9326
rect 7832 9240 7840 9310
rect 12490 9240 12506 9310
rect 7832 9226 7852 9240
rect 12486 9226 12506 9240
rect 6340 9130 6410 9200
rect 640 9020 650 9090
rect 850 9020 860 9090
rect 640 8980 860 9020
rect 640 8910 650 8980
rect 850 8910 860 8980
rect 640 8860 860 8910
rect 0 8850 1000 8860
rect 0 8650 20 8850
rect 90 8650 410 8850
rect 480 8650 520 8850
rect 590 8650 910 8850
rect 980 8650 1000 8850
rect 0 8640 1000 8650
rect 140 8590 360 8640
rect 140 8520 150 8590
rect 350 8520 360 8590
rect 140 8480 360 8520
rect 140 8410 150 8480
rect 350 8410 360 8480
rect 140 8360 360 8410
rect 640 8590 860 8640
rect 6800 8600 7300 9200
rect 7630 9130 7700 9200
rect 12710 15300 13930 15520
rect 12710 14700 13930 15100
rect 12710 14100 13930 14500
rect 12710 13500 13930 13900
rect 12710 12900 13930 13300
rect 12710 12300 13930 12700
rect 12710 11700 13930 12100
rect 12710 11100 13930 11500
rect 12710 10500 13930 10900
rect 12710 9900 13930 10300
rect 12710 9300 13930 9700
rect 12640 9130 12710 9200
rect 13100 8600 13600 9300
rect 18940 15520 19150 15580
rect 19350 15520 19650 15590
rect 19850 15520 20300 15590
rect 25640 15590 25860 15640
rect 14132 15480 14152 15490
rect 18786 15480 18806 15490
rect 14132 15410 14140 15480
rect 18800 15410 18806 15480
rect 14132 15390 14152 15410
rect 18786 15390 18806 15410
rect 14065 15338 14131 15358
rect 14065 9358 14131 9378
rect 14223 15338 14289 15358
rect 14223 9358 14289 9378
rect 14381 15338 14447 15358
rect 14381 9358 14447 9378
rect 14539 15338 14605 15358
rect 14539 9358 14605 9378
rect 14697 15338 14763 15358
rect 14697 9358 14763 9378
rect 14855 15338 14921 15358
rect 14855 9358 14921 9378
rect 15013 15338 15079 15358
rect 15013 9358 15079 9378
rect 15171 15338 15237 15358
rect 15171 9358 15237 9378
rect 15329 15338 15395 15358
rect 15329 9358 15395 9378
rect 15487 15338 15553 15358
rect 15487 9358 15553 9378
rect 15645 15338 15711 15358
rect 15645 9358 15711 9378
rect 15803 15338 15869 15358
rect 15803 9358 15869 9378
rect 15961 15338 16027 15358
rect 15961 9358 16027 9378
rect 16119 15338 16185 15358
rect 16119 9358 16185 9378
rect 16277 15338 16343 15358
rect 16277 9358 16343 9378
rect 16435 15338 16501 15358
rect 16435 9358 16501 9378
rect 16593 15338 16659 15358
rect 16593 9358 16659 9378
rect 16751 15338 16817 15358
rect 16751 9358 16817 9378
rect 16909 15338 16975 15358
rect 16909 9358 16975 9378
rect 17067 15338 17133 15358
rect 17067 9358 17133 9378
rect 17225 15338 17291 15358
rect 17225 9358 17291 9378
rect 17383 15338 17449 15358
rect 17383 9358 17449 9378
rect 17541 15338 17607 15358
rect 17541 9358 17607 9378
rect 17699 15338 17765 15358
rect 17699 9358 17765 9378
rect 17857 15338 17923 15358
rect 17857 9358 17923 9378
rect 18015 15338 18081 15358
rect 18015 9358 18081 9378
rect 18173 15338 18239 15358
rect 18173 9358 18239 9378
rect 18331 15338 18397 15358
rect 18331 9358 18397 9378
rect 18489 15338 18555 15358
rect 18489 9358 18555 9378
rect 18647 15338 18713 15358
rect 18647 9358 18713 9378
rect 18805 15338 18871 15358
rect 18805 9358 18871 9378
rect 14132 9310 14152 9326
rect 18786 9310 18806 9326
rect 14132 9240 14140 9310
rect 18790 9240 18806 9310
rect 14132 9226 14152 9240
rect 18786 9226 18806 9240
rect 13930 9130 14000 9200
rect 19010 15200 20230 15520
rect 19010 14600 20230 15000
rect 19010 14000 20230 14400
rect 19010 13400 20230 13800
rect 19010 12800 20230 13200
rect 19010 12200 20230 12600
rect 19010 11600 20230 12000
rect 19010 11000 20230 11400
rect 19010 10400 20230 10800
rect 19010 9800 20230 10200
rect 19010 9200 20230 9600
rect 25240 15520 25310 15580
rect 20432 15480 20452 15490
rect 25086 15480 25106 15490
rect 20432 15410 20440 15480
rect 25100 15410 25106 15480
rect 20432 15390 20452 15410
rect 25086 15390 25106 15410
rect 20365 15338 20431 15358
rect 20365 9358 20431 9378
rect 20523 15338 20589 15358
rect 20523 9358 20589 9378
rect 20681 15338 20747 15358
rect 20681 9358 20747 9378
rect 20839 15338 20905 15358
rect 20839 9358 20905 9378
rect 20997 15338 21063 15358
rect 20997 9358 21063 9378
rect 21155 15338 21221 15358
rect 21155 9358 21221 9378
rect 21313 15338 21379 15358
rect 21313 9358 21379 9378
rect 21471 15338 21537 15358
rect 21471 9358 21537 9378
rect 21629 15338 21695 15358
rect 21629 9358 21695 9378
rect 21787 15338 21853 15358
rect 21787 9358 21853 9378
rect 21945 15338 22011 15358
rect 21945 9358 22011 9378
rect 22103 15338 22169 15358
rect 22103 9358 22169 9378
rect 22261 15338 22327 15358
rect 22261 9358 22327 9378
rect 22419 15338 22485 15358
rect 22419 9358 22485 9378
rect 22577 15338 22643 15358
rect 22577 9358 22643 9378
rect 22735 15338 22801 15358
rect 22735 9358 22801 9378
rect 22893 15338 22959 15358
rect 22893 9358 22959 9378
rect 23051 15338 23117 15358
rect 23051 9358 23117 9378
rect 23209 15338 23275 15358
rect 23209 9358 23275 9378
rect 23367 15338 23433 15358
rect 23367 9358 23433 9378
rect 23525 15338 23591 15358
rect 23525 9358 23591 9378
rect 23683 15338 23749 15358
rect 23683 9358 23749 9378
rect 23841 15338 23907 15358
rect 23841 9358 23907 9378
rect 23999 15338 24065 15358
rect 23999 9358 24065 9378
rect 24157 15338 24223 15358
rect 24157 9358 24223 9378
rect 24315 15338 24381 15358
rect 24315 9358 24381 9378
rect 24473 15338 24539 15358
rect 24473 9358 24539 9378
rect 24631 15338 24697 15358
rect 24631 9358 24697 9378
rect 24789 15338 24855 15358
rect 24789 9358 24855 9378
rect 24947 15338 25013 15358
rect 24947 9358 25013 9378
rect 25105 15338 25171 15358
rect 25105 9358 25171 9378
rect 20432 9310 20452 9326
rect 25086 9310 25106 9326
rect 20432 9240 20440 9310
rect 25090 9240 25106 9310
rect 20432 9226 20452 9240
rect 25086 9226 25106 9240
rect 18940 9130 19010 9200
rect 19400 8600 19900 9200
rect 20230 9130 20300 9200
rect 25640 15520 25650 15590
rect 25850 15520 25860 15590
rect 25640 15480 25860 15520
rect 25640 15410 25650 15480
rect 25850 15410 25860 15480
rect 25640 15360 25860 15410
rect 26140 15590 26360 15640
rect 26140 15520 26150 15590
rect 26350 15520 26360 15590
rect 26140 15480 26360 15520
rect 26140 15410 26150 15480
rect 26350 15410 26360 15480
rect 26140 15360 26360 15410
rect 25500 15350 26500 15360
rect 25500 15150 25520 15350
rect 25590 15150 25910 15350
rect 25980 15150 26020 15350
rect 26090 15150 26410 15350
rect 26480 15150 26500 15350
rect 25500 15140 26500 15150
rect 25640 15090 25860 15140
rect 25640 15020 25650 15090
rect 25850 15020 25860 15090
rect 25640 14980 25860 15020
rect 25640 14910 25650 14980
rect 25850 14910 25860 14980
rect 25640 14860 25860 14910
rect 26140 15090 26360 15140
rect 26140 15020 26150 15090
rect 26350 15020 26360 15090
rect 26140 14980 26360 15020
rect 26140 14910 26150 14980
rect 26350 14910 26360 14980
rect 26140 14860 26360 14910
rect 25500 14850 26500 14860
rect 25500 14650 25520 14850
rect 25590 14650 25910 14850
rect 25980 14650 26020 14850
rect 26090 14650 26410 14850
rect 26480 14650 26500 14850
rect 25500 14640 26500 14650
rect 25640 14590 25860 14640
rect 25640 14520 25650 14590
rect 25850 14520 25860 14590
rect 25640 14480 25860 14520
rect 25640 14410 25650 14480
rect 25850 14410 25860 14480
rect 25640 14360 25860 14410
rect 26140 14590 26360 14640
rect 26140 14520 26150 14590
rect 26350 14520 26360 14590
rect 26140 14480 26360 14520
rect 26140 14410 26150 14480
rect 26350 14410 26360 14480
rect 26140 14360 26360 14410
rect 25500 14350 26500 14360
rect 25500 14150 25520 14350
rect 25590 14150 25910 14350
rect 25980 14150 26020 14350
rect 26090 14150 26410 14350
rect 26480 14150 26500 14350
rect 25500 14140 26500 14150
rect 25640 14090 25860 14140
rect 25640 14020 25650 14090
rect 25850 14020 25860 14090
rect 25640 13980 25860 14020
rect 25640 13910 25650 13980
rect 25850 13910 25860 13980
rect 25640 13860 25860 13910
rect 26140 14090 26360 14140
rect 26140 14020 26150 14090
rect 26350 14020 26360 14090
rect 26140 13980 26360 14020
rect 26140 13910 26150 13980
rect 26350 13910 26360 13980
rect 26140 13860 26360 13910
rect 26640 13980 26860 14000
rect 26640 13910 26650 13980
rect 26850 13910 26860 13980
rect 26640 13860 26860 13910
rect 27140 13980 27360 14000
rect 27140 13910 27150 13980
rect 27350 13910 27360 13980
rect 27140 13860 27360 13910
rect 27640 13980 27860 14000
rect 27640 13910 27650 13980
rect 27850 13910 27860 13980
rect 27640 13860 27860 13910
rect 28140 13980 28360 14000
rect 28140 13910 28150 13980
rect 28350 13910 28360 13980
rect 28140 13860 28360 13910
rect 28640 13980 28860 14000
rect 28640 13910 28650 13980
rect 28850 13910 28860 13980
rect 28640 13860 28860 13910
rect 29140 13980 29360 14000
rect 29140 13910 29150 13980
rect 29350 13910 29360 13980
rect 29140 13860 29360 13910
rect 29640 13980 29860 14000
rect 29640 13910 29650 13980
rect 29850 13910 29860 13980
rect 29640 13860 29860 13910
rect 30140 13980 30360 14000
rect 30140 13910 30150 13980
rect 30350 13910 30360 13980
rect 30140 13860 30360 13910
rect 30900 13900 31100 13910
rect 25500 13850 30500 13860
rect 25500 13650 25520 13850
rect 25590 13650 25910 13850
rect 25980 13650 26020 13850
rect 26090 13650 26410 13850
rect 26480 13650 26520 13850
rect 26590 13650 26910 13850
rect 26980 13650 27020 13850
rect 27090 13650 27410 13850
rect 27480 13650 27520 13850
rect 27590 13650 27910 13850
rect 27980 13650 28020 13850
rect 28090 13650 28410 13850
rect 28480 13650 28520 13850
rect 28590 13650 28910 13850
rect 28980 13650 29020 13850
rect 29090 13650 29410 13850
rect 29480 13650 29520 13850
rect 29590 13650 29910 13850
rect 29980 13650 30020 13850
rect 30090 13650 30410 13850
rect 30480 13650 30500 13850
rect 25500 13640 30500 13650
rect 25640 13590 25860 13640
rect 25640 13520 25650 13590
rect 25850 13520 25860 13590
rect 25640 13480 25860 13520
rect 25640 13410 25650 13480
rect 25850 13410 25860 13480
rect 25640 13360 25860 13410
rect 26140 13590 26360 13640
rect 26140 13520 26150 13590
rect 26350 13520 26360 13590
rect 26140 13480 26360 13520
rect 26140 13410 26150 13480
rect 26350 13410 26360 13480
rect 26140 13360 26360 13410
rect 26640 13590 26860 13640
rect 26640 13520 26650 13590
rect 26850 13520 26860 13590
rect 26640 13480 26860 13520
rect 26640 13410 26650 13480
rect 26850 13410 26860 13480
rect 26640 13360 26860 13410
rect 27140 13590 27360 13640
rect 27140 13520 27150 13590
rect 27350 13520 27360 13590
rect 27140 13480 27360 13520
rect 27140 13410 27150 13480
rect 27350 13410 27360 13480
rect 27140 13360 27360 13410
rect 27640 13590 27860 13640
rect 27640 13520 27650 13590
rect 27850 13520 27860 13590
rect 27640 13480 27860 13520
rect 27640 13410 27650 13480
rect 27850 13410 27860 13480
rect 27640 13360 27860 13410
rect 28140 13590 28360 13640
rect 28140 13520 28150 13590
rect 28350 13520 28360 13590
rect 28140 13480 28360 13520
rect 28140 13410 28150 13480
rect 28350 13410 28360 13480
rect 28140 13360 28360 13410
rect 28640 13590 28860 13640
rect 28640 13520 28650 13590
rect 28850 13520 28860 13590
rect 28640 13480 28860 13520
rect 28640 13410 28650 13480
rect 28850 13410 28860 13480
rect 28640 13360 28860 13410
rect 29140 13590 29360 13640
rect 29140 13520 29150 13590
rect 29350 13520 29360 13590
rect 29140 13480 29360 13520
rect 29140 13410 29150 13480
rect 29350 13410 29360 13480
rect 29140 13360 29360 13410
rect 29640 13590 29860 13640
rect 29640 13520 29650 13590
rect 29850 13520 29860 13590
rect 29640 13480 29860 13520
rect 29640 13410 29650 13480
rect 29850 13410 29860 13480
rect 29640 13360 29860 13410
rect 30140 13590 30360 13640
rect 30140 13520 30150 13590
rect 30350 13520 30360 13590
rect 30140 13480 30360 13520
rect 30140 13410 30150 13480
rect 30350 13410 30360 13480
rect 30900 13420 30910 13900
rect 31090 13420 31100 13900
rect 30900 13410 31100 13420
rect 30140 13360 30360 13410
rect 25500 13350 30500 13360
rect 25500 13150 25520 13350
rect 25590 13150 25910 13350
rect 25980 13150 26020 13350
rect 26090 13150 26410 13350
rect 26480 13150 26520 13350
rect 26590 13150 26910 13350
rect 26980 13150 27020 13350
rect 27090 13150 27410 13350
rect 27480 13150 27520 13350
rect 27590 13150 27910 13350
rect 27980 13150 28020 13350
rect 28090 13150 28410 13350
rect 28480 13150 28520 13350
rect 28590 13150 28910 13350
rect 28980 13150 29020 13350
rect 29090 13150 29410 13350
rect 29480 13150 29520 13350
rect 29590 13150 29910 13350
rect 29980 13150 30020 13350
rect 30090 13150 30410 13350
rect 30480 13150 30500 13350
rect 25500 13140 30500 13150
rect 25640 13090 25860 13140
rect 25640 13020 25650 13090
rect 25850 13020 25860 13090
rect 25640 12980 25860 13020
rect 25640 12910 25650 12980
rect 25850 12910 25860 12980
rect 25640 12860 25860 12910
rect 26140 13090 26360 13140
rect 26140 13020 26150 13090
rect 26350 13020 26360 13090
rect 26140 12980 26360 13020
rect 26640 13090 26860 13140
rect 26640 13020 26650 13090
rect 26850 13020 26860 13090
rect 26640 13000 26860 13020
rect 27140 13090 27360 13140
rect 27140 13020 27150 13090
rect 27350 13020 27360 13090
rect 27140 13000 27360 13020
rect 27640 13090 27860 13140
rect 27640 13020 27650 13090
rect 27850 13020 27860 13090
rect 27640 13000 27860 13020
rect 28140 13090 28360 13140
rect 28140 13020 28150 13090
rect 28350 13020 28360 13090
rect 28140 13000 28360 13020
rect 28640 13090 28860 13140
rect 28640 13020 28650 13090
rect 28850 13020 28860 13090
rect 28640 13000 28860 13020
rect 29140 13090 29360 13140
rect 29140 13020 29150 13090
rect 29350 13020 29360 13090
rect 29140 13000 29360 13020
rect 29640 13090 29860 13140
rect 29640 13020 29650 13090
rect 29850 13020 29860 13090
rect 29640 13000 29860 13020
rect 30140 13090 30360 13140
rect 30140 13020 30150 13090
rect 30350 13020 30360 13090
rect 30140 13000 30360 13020
rect 30900 13090 31100 13100
rect 26140 12910 26150 12980
rect 26350 12910 26360 12980
rect 26140 12860 26360 12910
rect 25500 12850 26500 12860
rect 25500 12650 25520 12850
rect 25590 12650 25910 12850
rect 25980 12650 26020 12850
rect 26090 12650 26410 12850
rect 26480 12650 26500 12850
rect 25500 12640 26500 12650
rect 25640 12590 25860 12640
rect 25640 12520 25650 12590
rect 25850 12520 25860 12590
rect 25640 12480 25860 12520
rect 25640 12410 25650 12480
rect 25850 12410 25860 12480
rect 25640 12360 25860 12410
rect 26140 12590 26360 12640
rect 30900 12610 30910 13090
rect 31090 12610 31100 13090
rect 30900 12600 31100 12610
rect 26140 12520 26150 12590
rect 26350 12520 26360 12590
rect 26140 12480 26360 12520
rect 26140 12410 26150 12480
rect 26350 12410 26360 12480
rect 26140 12360 26360 12410
rect 25500 12350 26500 12360
rect 25500 12150 25520 12350
rect 25590 12150 25910 12350
rect 25980 12150 26020 12350
rect 26090 12150 26410 12350
rect 26480 12150 26500 12350
rect 25500 12140 26500 12150
rect 25640 12090 25860 12140
rect 25640 12020 25650 12090
rect 25850 12020 25860 12090
rect 25640 11980 25860 12020
rect 25640 11910 25650 11980
rect 25850 11910 25860 11980
rect 25640 11860 25860 11910
rect 26140 12090 26360 12140
rect 26140 12020 26150 12090
rect 26350 12020 26360 12090
rect 26140 11980 26360 12020
rect 26140 11910 26150 11980
rect 26350 11910 26360 11980
rect 26140 11860 26360 11910
rect 25500 11850 26500 11860
rect 25500 11650 25520 11850
rect 25590 11650 25910 11850
rect 25980 11650 26020 11850
rect 26090 11650 26410 11850
rect 26480 11650 26500 11850
rect 25500 11640 26500 11650
rect 25640 11590 25860 11640
rect 25640 11520 25650 11590
rect 25850 11520 25860 11590
rect 25640 11480 25860 11520
rect 25640 11410 25650 11480
rect 25850 11410 25860 11480
rect 25640 11360 25860 11410
rect 26140 11590 26360 11640
rect 26140 11520 26150 11590
rect 26350 11520 26360 11590
rect 26140 11480 26360 11520
rect 26140 11410 26150 11480
rect 26350 11410 26360 11480
rect 26140 11360 26360 11410
rect 25500 11350 26500 11360
rect 25500 11150 25520 11350
rect 25590 11150 25910 11350
rect 25980 11150 26020 11350
rect 26090 11150 26410 11350
rect 26480 11150 26500 11350
rect 25500 11140 26500 11150
rect 25640 11090 25860 11140
rect 25640 11020 25650 11090
rect 25850 11020 25860 11090
rect 25640 10980 25860 11020
rect 25640 10910 25650 10980
rect 25850 10910 25860 10980
rect 25640 10860 25860 10910
rect 26140 11090 26360 11140
rect 26140 11020 26150 11090
rect 26350 11020 26360 11090
rect 26140 10980 26360 11020
rect 26140 10910 26150 10980
rect 26350 10910 26360 10980
rect 26140 10860 26360 10910
rect 25500 10850 26500 10860
rect 25500 10650 25520 10850
rect 25590 10650 25910 10850
rect 25980 10650 26020 10850
rect 26090 10650 26410 10850
rect 26480 10650 26500 10850
rect 25500 10640 26500 10650
rect 25640 10590 25860 10640
rect 25640 10520 25650 10590
rect 25850 10520 25860 10590
rect 25640 10480 25860 10520
rect 25640 10410 25650 10480
rect 25850 10410 25860 10480
rect 25640 10360 25860 10410
rect 26140 10590 26360 10640
rect 26140 10520 26150 10590
rect 26350 10520 26360 10590
rect 26140 10480 26360 10520
rect 26140 10410 26150 10480
rect 26350 10410 26360 10480
rect 26140 10360 26360 10410
rect 25500 10350 26500 10360
rect 25500 10150 25520 10350
rect 25590 10150 25910 10350
rect 25980 10150 26020 10350
rect 26090 10150 26410 10350
rect 26480 10150 26500 10350
rect 25500 10140 26500 10150
rect 25640 10090 25860 10140
rect 25640 10020 25650 10090
rect 25850 10020 25860 10090
rect 25640 9980 25860 10020
rect 25640 9910 25650 9980
rect 25850 9910 25860 9980
rect 25640 9860 25860 9910
rect 26140 10090 26360 10140
rect 26140 10020 26150 10090
rect 26350 10020 26360 10090
rect 26140 9980 26360 10020
rect 26140 9910 26150 9980
rect 26350 9910 26360 9980
rect 26140 9860 26360 9910
rect 25500 9850 26500 9860
rect 25500 9650 25520 9850
rect 25590 9650 25910 9850
rect 25980 9650 26020 9850
rect 26090 9650 26410 9850
rect 26480 9650 26500 9850
rect 25500 9640 26500 9650
rect 25640 9590 25860 9640
rect 25640 9520 25650 9590
rect 25850 9520 25860 9590
rect 25640 9480 25860 9520
rect 25640 9410 25650 9480
rect 25850 9410 25860 9480
rect 25640 9360 25860 9410
rect 26140 9590 26360 9640
rect 26140 9520 26150 9590
rect 26350 9520 26360 9590
rect 26140 9480 26360 9520
rect 26140 9410 26150 9480
rect 26350 9410 26360 9480
rect 26140 9360 26360 9410
rect 25240 9130 25310 9200
rect 25500 9350 26500 9360
rect 25500 9150 25520 9350
rect 25590 9150 25910 9350
rect 25980 9150 26020 9350
rect 26090 9150 26410 9350
rect 26480 9150 26500 9350
rect 25500 9140 26500 9150
rect 25640 9090 25860 9140
rect 25640 9020 25650 9090
rect 25850 9020 25860 9090
rect 25640 8980 25860 9020
rect 25640 8910 25650 8980
rect 25850 8910 25860 8980
rect 25640 8860 25860 8910
rect 26140 9090 26360 9140
rect 26140 9020 26150 9090
rect 26350 9020 26360 9090
rect 26140 8980 26360 9020
rect 26140 8910 26150 8980
rect 26350 8910 26360 8980
rect 26140 8860 26360 8910
rect 25500 8850 26500 8860
rect 25500 8650 25520 8850
rect 25590 8650 25910 8850
rect 25980 8650 26020 8850
rect 26090 8650 26410 8850
rect 26480 8650 26500 8850
rect 25500 8640 26500 8650
rect 640 8520 650 8590
rect 850 8520 860 8590
rect 6400 8580 7700 8600
rect 12700 8580 14000 8600
rect 19000 8580 20300 8600
rect 25640 8590 25860 8640
rect 640 8480 860 8520
rect 640 8410 650 8480
rect 850 8410 860 8480
rect 640 8360 860 8410
rect 1330 8520 1400 8580
rect 0 8350 1000 8360
rect 0 8150 20 8350
rect 90 8150 410 8350
rect 480 8150 520 8350
rect 590 8150 910 8350
rect 980 8150 1000 8350
rect 0 8140 1000 8150
rect 140 8090 360 8140
rect 140 8020 150 8090
rect 350 8020 360 8090
rect 140 7980 360 8020
rect 140 7910 150 7980
rect 350 7910 360 7980
rect 140 7860 360 7910
rect 640 8090 860 8140
rect 640 8020 650 8090
rect 850 8020 860 8090
rect 640 7980 860 8020
rect 640 7910 650 7980
rect 850 7910 860 7980
rect 640 7860 860 7910
rect 0 7850 1000 7860
rect 0 7650 20 7850
rect 90 7650 410 7850
rect 480 7650 520 7850
rect 590 7650 910 7850
rect 980 7650 1000 7850
rect 0 7640 1000 7650
rect 140 7590 360 7640
rect 140 7520 150 7590
rect 350 7520 360 7590
rect 140 7480 360 7520
rect 140 7410 150 7480
rect 350 7410 360 7480
rect 140 7360 360 7410
rect 640 7590 860 7640
rect 640 7520 650 7590
rect 850 7520 860 7590
rect 640 7480 860 7520
rect 640 7410 650 7480
rect 850 7410 860 7480
rect 640 7360 860 7410
rect 0 7350 1000 7360
rect 0 7150 20 7350
rect 90 7150 410 7350
rect 480 7150 520 7350
rect 590 7150 910 7350
rect 980 7150 1000 7350
rect 0 7140 1000 7150
rect 140 7090 360 7140
rect 140 7020 150 7090
rect 350 7020 360 7090
rect 140 6980 360 7020
rect 140 6910 150 6980
rect 350 6910 360 6980
rect 140 6860 360 6910
rect 640 7090 860 7140
rect 640 7020 650 7090
rect 850 7020 860 7090
rect 640 6980 860 7020
rect 640 6910 650 6980
rect 850 6910 860 6980
rect 640 6860 860 6910
rect 0 6850 1000 6860
rect 0 6650 20 6850
rect 90 6650 410 6850
rect 480 6650 520 6850
rect 590 6650 910 6850
rect 980 6650 1000 6850
rect 0 6640 1000 6650
rect 140 6590 360 6640
rect 140 6520 150 6590
rect 350 6520 360 6590
rect 140 6480 360 6520
rect 140 6410 150 6480
rect 350 6410 360 6480
rect 140 6360 360 6410
rect 640 6590 860 6640
rect 640 6520 650 6590
rect 850 6520 860 6590
rect 640 6480 860 6520
rect 640 6410 650 6480
rect 850 6410 860 6480
rect 640 6360 860 6410
rect 0 6350 1000 6360
rect 0 6150 20 6350
rect 90 6150 410 6350
rect 480 6150 520 6350
rect 590 6150 910 6350
rect 980 6150 1000 6350
rect 0 6140 1000 6150
rect 140 6090 360 6140
rect 140 6020 150 6090
rect 350 6020 360 6090
rect 140 5980 360 6020
rect 140 5910 150 5980
rect 350 5910 360 5980
rect 140 5860 360 5910
rect 640 6090 860 6140
rect 640 6020 650 6090
rect 850 6020 860 6090
rect 640 5980 860 6020
rect 640 5910 650 5980
rect 850 5910 860 5980
rect 640 5860 860 5910
rect 0 5850 1000 5860
rect 0 5650 20 5850
rect 90 5650 410 5850
rect 480 5650 520 5850
rect 590 5650 910 5850
rect 980 5650 1000 5850
rect 0 5640 1000 5650
rect 140 5590 360 5640
rect 140 5520 150 5590
rect 350 5520 360 5590
rect 140 5480 360 5520
rect 140 5410 150 5480
rect 350 5410 360 5480
rect 140 5360 360 5410
rect 640 5590 860 5640
rect 640 5520 650 5590
rect 850 5520 860 5590
rect 640 5480 860 5520
rect 640 5410 650 5480
rect 850 5410 860 5480
rect 640 5360 860 5410
rect 0 5350 1000 5360
rect 0 5150 20 5350
rect 90 5150 410 5350
rect 480 5150 520 5350
rect 590 5150 910 5350
rect 980 5150 1000 5350
rect 0 5140 1000 5150
rect 140 5090 360 5140
rect 140 5020 150 5090
rect 350 5020 360 5090
rect 140 4980 360 5020
rect 140 4910 150 4980
rect 350 4910 360 4980
rect 140 4860 360 4910
rect 640 5090 860 5140
rect 640 5020 650 5090
rect 850 5020 860 5090
rect 640 4980 860 5020
rect 640 4910 650 4980
rect 850 4910 860 4980
rect 640 4860 860 4910
rect 0 4850 1000 4860
rect 0 4650 20 4850
rect 90 4650 410 4850
rect 480 4650 520 4850
rect 590 4650 910 4850
rect 980 4650 1000 4850
rect 0 4640 1000 4650
rect 140 4590 360 4640
rect 140 4520 150 4590
rect 350 4520 360 4590
rect 140 4480 360 4520
rect 140 4410 150 4480
rect 350 4410 360 4480
rect 140 4360 360 4410
rect 640 4590 860 4640
rect 640 4520 650 4590
rect 850 4520 860 4590
rect 640 4480 860 4520
rect 640 4410 650 4480
rect 850 4410 860 4480
rect 640 4360 860 4410
rect 0 4350 1000 4360
rect 0 4150 20 4350
rect 90 4150 410 4350
rect 480 4150 520 4350
rect 590 4150 910 4350
rect 980 4150 1000 4350
rect 0 4140 1000 4150
rect 140 4090 360 4140
rect 140 4020 150 4090
rect 350 4020 360 4090
rect 140 3980 360 4020
rect 140 3910 150 3980
rect 350 3910 360 3980
rect 140 3860 360 3910
rect 640 4090 860 4140
rect 640 4020 650 4090
rect 850 4020 860 4090
rect 640 3980 860 4020
rect 640 3910 650 3980
rect 850 3910 860 3980
rect 640 3860 860 3910
rect 0 3850 1000 3860
rect 0 3650 20 3850
rect 90 3650 410 3850
rect 480 3650 520 3850
rect 590 3650 910 3850
rect 980 3650 1000 3850
rect 0 3640 1000 3650
rect 140 3590 360 3640
rect 140 3520 150 3590
rect 350 3520 360 3590
rect 140 3480 360 3520
rect 140 3410 150 3480
rect 350 3410 360 3480
rect 140 3360 360 3410
rect 640 3590 860 3640
rect 640 3520 650 3590
rect 850 3520 860 3590
rect 640 3480 860 3520
rect 640 3410 650 3480
rect 850 3410 860 3480
rect 640 3360 860 3410
rect 0 3350 1000 3360
rect 0 3150 20 3350
rect 90 3150 410 3350
rect 480 3150 520 3350
rect 590 3150 910 3350
rect 980 3150 1000 3350
rect 0 3140 1000 3150
rect 140 3090 360 3140
rect 140 3020 150 3090
rect 350 3020 360 3090
rect 140 2980 360 3020
rect 140 2910 150 2980
rect 350 2910 360 2980
rect 140 2860 360 2910
rect 640 3090 860 3140
rect 640 3020 650 3090
rect 850 3020 860 3090
rect 640 2980 860 3020
rect 640 2910 650 2980
rect 850 2910 860 2980
rect 640 2860 860 2910
rect 0 2850 1000 2860
rect 0 2650 20 2850
rect 90 2650 410 2850
rect 480 2650 520 2850
rect 590 2650 910 2850
rect 980 2650 1000 2850
rect 0 2640 1000 2650
rect 140 2590 360 2640
rect 140 2520 150 2590
rect 350 2520 360 2590
rect 140 2480 360 2520
rect 140 2410 150 2480
rect 350 2410 360 2480
rect 140 2360 360 2410
rect 640 2590 860 2640
rect 640 2520 650 2590
rect 850 2520 860 2590
rect 640 2480 860 2520
rect 640 2410 650 2480
rect 850 2410 860 2480
rect 640 2360 860 2410
rect 0 2350 1000 2360
rect 0 2150 20 2350
rect 90 2150 410 2350
rect 480 2150 520 2350
rect 590 2150 910 2350
rect 980 2150 1000 2350
rect 0 2140 1000 2150
rect 6340 8520 7700 8580
rect 1532 8480 1552 8490
rect 6186 8480 6206 8490
rect 1532 8410 1540 8480
rect 6200 8410 6206 8480
rect 1532 8390 1552 8410
rect 6186 8390 6206 8410
rect 1465 8338 1531 8358
rect 1465 2358 1531 2378
rect 1623 8338 1689 8358
rect 1623 2358 1689 2378
rect 1781 8338 1847 8358
rect 1781 2358 1847 2378
rect 1939 8338 2005 8358
rect 1939 2358 2005 2378
rect 2097 8338 2163 8358
rect 2097 2358 2163 2378
rect 2255 8338 2321 8358
rect 2255 2358 2321 2378
rect 2413 8338 2479 8358
rect 2413 2358 2479 2378
rect 2571 8338 2637 8358
rect 2571 2358 2637 2378
rect 2729 8338 2795 8358
rect 2729 2358 2795 2378
rect 2887 8338 2953 8358
rect 2887 2358 2953 2378
rect 3045 8338 3111 8358
rect 3045 2358 3111 2378
rect 3203 8338 3269 8358
rect 3203 2358 3269 2378
rect 3361 8338 3427 8358
rect 3361 2358 3427 2378
rect 3519 8338 3585 8358
rect 3519 2358 3585 2378
rect 3677 8338 3743 8358
rect 3677 2358 3743 2378
rect 3835 8338 3901 8358
rect 3835 2358 3901 2378
rect 3993 8338 4059 8358
rect 3993 2358 4059 2378
rect 4151 8338 4217 8358
rect 4151 2358 4217 2378
rect 4309 8338 4375 8358
rect 4309 2358 4375 2378
rect 4467 8338 4533 8358
rect 4467 2358 4533 2378
rect 4625 8338 4691 8358
rect 4625 2358 4691 2378
rect 4783 8338 4849 8358
rect 4783 2358 4849 2378
rect 4941 8338 5007 8358
rect 4941 2358 5007 2378
rect 5099 8338 5165 8358
rect 5099 2358 5165 2378
rect 5257 8338 5323 8358
rect 5257 2358 5323 2378
rect 5415 8338 5481 8358
rect 5415 2358 5481 2378
rect 5573 8338 5639 8358
rect 5573 2358 5639 2378
rect 5731 8338 5797 8358
rect 5731 2358 5797 2378
rect 5889 8338 5955 8358
rect 5889 2358 5955 2378
rect 6047 8338 6113 8358
rect 6047 2358 6113 2378
rect 6205 8338 6271 8358
rect 6205 2358 6271 2378
rect 1532 2310 1552 2326
rect 6186 2310 6206 2326
rect 1532 2240 1540 2310
rect 6190 2240 6206 2310
rect 1532 2226 1552 2240
rect 6186 2226 6206 2240
rect 140 2090 360 2140
rect 140 2020 150 2090
rect 350 2020 360 2090
rect 140 1980 360 2020
rect 140 1910 150 1980
rect 350 1910 360 1980
rect 140 1860 360 1910
rect 640 2090 860 2140
rect 1330 2130 1400 2200
rect 6410 8200 7630 8520
rect 6410 7600 7630 8000
rect 6410 7000 7630 7400
rect 6410 6400 7630 6800
rect 6410 5800 7630 6200
rect 6410 5200 7630 5600
rect 6410 4600 7630 5000
rect 6410 4000 7630 4400
rect 6410 3400 7630 3800
rect 6410 2800 7630 3200
rect 6410 2480 7630 2600
rect 6410 2410 6650 2480
rect 6850 2410 7150 2480
rect 7350 2410 7630 2480
rect 6410 2350 7630 2410
rect 6410 2200 6520 2350
rect 6340 2130 6410 2200
rect 6500 2150 6520 2200
rect 6590 2150 6910 2350
rect 6980 2150 7020 2350
rect 7090 2150 7410 2350
rect 7480 2200 7630 2350
rect 12640 8520 14000 8580
rect 7832 8480 7852 8490
rect 12486 8480 12506 8490
rect 7832 8410 7840 8480
rect 12500 8410 12506 8480
rect 7832 8390 7852 8410
rect 12486 8390 12506 8410
rect 7765 8338 7831 8358
rect 7765 2358 7831 2378
rect 7923 8338 7989 8358
rect 7923 2358 7989 2378
rect 8081 8338 8147 8358
rect 8081 2358 8147 2378
rect 8239 8338 8305 8358
rect 8239 2358 8305 2378
rect 8397 8338 8463 8358
rect 8397 2358 8463 2378
rect 8555 8338 8621 8358
rect 8555 2358 8621 2378
rect 8713 8338 8779 8358
rect 8713 2358 8779 2378
rect 8871 8338 8937 8358
rect 8871 2358 8937 2378
rect 9029 8338 9095 8358
rect 9029 2358 9095 2378
rect 9187 8338 9253 8358
rect 9187 2358 9253 2378
rect 9345 8338 9411 8358
rect 9345 2358 9411 2378
rect 9503 8338 9569 8358
rect 9503 2358 9569 2378
rect 9661 8338 9727 8358
rect 9661 2358 9727 2378
rect 9819 8338 9885 8358
rect 9819 2358 9885 2378
rect 9977 8338 10043 8358
rect 9977 2358 10043 2378
rect 10135 8338 10201 8358
rect 10135 2358 10201 2378
rect 10293 8338 10359 8358
rect 10293 2358 10359 2378
rect 10451 8338 10517 8358
rect 10451 2358 10517 2378
rect 10609 8338 10675 8358
rect 10609 2358 10675 2378
rect 10767 8338 10833 8358
rect 10767 2358 10833 2378
rect 10925 8338 10991 8358
rect 10925 2358 10991 2378
rect 11083 8338 11149 8358
rect 11083 2358 11149 2378
rect 11241 8338 11307 8358
rect 11241 2358 11307 2378
rect 11399 8338 11465 8358
rect 11399 2358 11465 2378
rect 11557 8338 11623 8358
rect 11557 2358 11623 2378
rect 11715 8338 11781 8358
rect 11715 2358 11781 2378
rect 11873 8338 11939 8358
rect 11873 2358 11939 2378
rect 12031 8338 12097 8358
rect 12031 2358 12097 2378
rect 12189 8338 12255 8358
rect 12189 2358 12255 2378
rect 12347 8338 12413 8358
rect 12347 2358 12413 2378
rect 12505 8338 12571 8358
rect 12505 2358 12571 2378
rect 7832 2310 7852 2326
rect 12486 2310 12506 2326
rect 7832 2240 7840 2310
rect 12490 2240 12506 2310
rect 7832 2226 7852 2240
rect 12486 2226 12506 2240
rect 7480 2150 7500 2200
rect 6500 2140 7500 2150
rect 640 2020 650 2090
rect 850 2020 860 2090
rect 640 1980 860 2020
rect 6640 2090 6860 2140
rect 6640 2020 6650 2090
rect 6850 2020 6860 2090
rect 640 1910 650 1980
rect 850 1910 860 1980
rect 640 1860 860 1910
rect 1140 1980 1360 2000
rect 1140 1910 1150 1980
rect 1350 1910 1360 1980
rect 1140 1860 1360 1910
rect 1640 1980 1860 2000
rect 1640 1910 1650 1980
rect 1850 1910 1860 1980
rect 1640 1860 1860 1910
rect 2140 1980 2360 2000
rect 2140 1910 2150 1980
rect 2350 1910 2360 1980
rect 2140 1860 2360 1910
rect 2640 1980 2860 2000
rect 2640 1910 2650 1980
rect 2850 1910 2860 1980
rect 2640 1860 2860 1910
rect 3140 1980 3360 2000
rect 3140 1910 3150 1980
rect 3350 1910 3360 1980
rect 3140 1860 3360 1910
rect 3640 1980 3860 2000
rect 3640 1910 3650 1980
rect 3850 1910 3860 1980
rect 3640 1860 3860 1910
rect 4140 1980 4360 2000
rect 4140 1910 4150 1980
rect 4350 1910 4360 1980
rect 4140 1860 4360 1910
rect 4640 1980 4860 2000
rect 4640 1910 4650 1980
rect 4850 1910 4860 1980
rect 4640 1860 4860 1910
rect 5140 1980 5360 2000
rect 5140 1910 5150 1980
rect 5350 1910 5360 1980
rect 5140 1860 5360 1910
rect 5640 1980 5860 2000
rect 5640 1910 5650 1980
rect 5850 1910 5860 1980
rect 5640 1860 5860 1910
rect 6140 1980 6360 2000
rect 6140 1910 6150 1980
rect 6350 1910 6360 1980
rect 6140 1860 6360 1910
rect 6640 1980 6860 2020
rect 6640 1910 6650 1980
rect 6850 1910 6860 1980
rect 6640 1860 6860 1910
rect 7140 2090 7360 2140
rect 7630 2130 7700 2200
rect 12710 8200 13930 8520
rect 12710 7600 13930 8000
rect 12710 7000 13930 7400
rect 12710 6400 13930 6800
rect 12710 5800 13930 6200
rect 12710 5200 13930 5600
rect 12710 4600 13930 5000
rect 12710 4000 13930 4400
rect 12710 3400 13930 3800
rect 12710 2800 13930 3200
rect 12710 2480 13930 2600
rect 12710 2410 13150 2480
rect 13350 2410 13930 2480
rect 12710 2350 13930 2410
rect 12710 2200 13020 2350
rect 12640 2130 12710 2200
rect 13000 2150 13020 2200
rect 13090 2150 13410 2350
rect 13480 2200 13930 2350
rect 18940 8520 20300 8580
rect 14132 8480 14152 8490
rect 18786 8480 18806 8490
rect 14132 8410 14140 8480
rect 18800 8410 18806 8480
rect 14132 8390 14152 8410
rect 18786 8390 18806 8410
rect 14065 8338 14131 8358
rect 14065 2358 14131 2378
rect 14223 8338 14289 8358
rect 14223 2358 14289 2378
rect 14381 8338 14447 8358
rect 14381 2358 14447 2378
rect 14539 8338 14605 8358
rect 14539 2358 14605 2378
rect 14697 8338 14763 8358
rect 14697 2358 14763 2378
rect 14855 8338 14921 8358
rect 14855 2358 14921 2378
rect 15013 8338 15079 8358
rect 15013 2358 15079 2378
rect 15171 8338 15237 8358
rect 15171 2358 15237 2378
rect 15329 8338 15395 8358
rect 15329 2358 15395 2378
rect 15487 8338 15553 8358
rect 15487 2358 15553 2378
rect 15645 8338 15711 8358
rect 15645 2358 15711 2378
rect 15803 8338 15869 8358
rect 15803 2358 15869 2378
rect 15961 8338 16027 8358
rect 15961 2358 16027 2378
rect 16119 8338 16185 8358
rect 16119 2358 16185 2378
rect 16277 8338 16343 8358
rect 16277 2358 16343 2378
rect 16435 8338 16501 8358
rect 16435 2358 16501 2378
rect 16593 8338 16659 8358
rect 16593 2358 16659 2378
rect 16751 8338 16817 8358
rect 16751 2358 16817 2378
rect 16909 8338 16975 8358
rect 16909 2358 16975 2378
rect 17067 8338 17133 8358
rect 17067 2358 17133 2378
rect 17225 8338 17291 8358
rect 17225 2358 17291 2378
rect 17383 8338 17449 8358
rect 17383 2358 17449 2378
rect 17541 8338 17607 8358
rect 17541 2358 17607 2378
rect 17699 8338 17765 8358
rect 17699 2358 17765 2378
rect 17857 8338 17923 8358
rect 17857 2358 17923 2378
rect 18015 8338 18081 8358
rect 18015 2358 18081 2378
rect 18173 8338 18239 8358
rect 18173 2358 18239 2378
rect 18331 8338 18397 8358
rect 18331 2358 18397 2378
rect 18489 8338 18555 8358
rect 18489 2358 18555 2378
rect 18647 8338 18713 8358
rect 18647 2358 18713 2378
rect 18805 8338 18871 8358
rect 18805 2358 18871 2378
rect 14132 2310 14152 2326
rect 18786 2310 18806 2326
rect 14132 2240 14140 2310
rect 18790 2240 18806 2310
rect 14132 2226 14152 2240
rect 18786 2226 18806 2240
rect 13480 2150 13500 2200
rect 13000 2140 13500 2150
rect 7140 2020 7150 2090
rect 7350 2020 7360 2090
rect 7140 1980 7360 2020
rect 13140 2090 13360 2140
rect 13930 2130 14000 2200
rect 19010 8200 20230 8520
rect 19010 7600 20230 8000
rect 19010 7000 20230 7400
rect 19010 6400 20230 6800
rect 19010 5800 20230 6200
rect 19010 5200 20230 5600
rect 19010 4600 20230 5000
rect 19010 4000 20230 4400
rect 19010 3400 20230 3800
rect 19010 2800 20230 3200
rect 19010 2480 20230 2600
rect 19010 2410 19650 2480
rect 19850 2410 20230 2480
rect 19010 2350 20230 2410
rect 19010 2200 19520 2350
rect 18940 2130 19010 2200
rect 19500 2150 19520 2200
rect 19590 2150 19910 2350
rect 19980 2200 20230 2350
rect 25240 8520 25310 8580
rect 20432 8480 20452 8490
rect 25086 8480 25106 8490
rect 20432 8410 20440 8480
rect 25100 8410 25106 8480
rect 20432 8390 20452 8410
rect 25086 8390 25106 8410
rect 20365 8338 20431 8358
rect 20365 2358 20431 2378
rect 20523 8338 20589 8358
rect 20523 2358 20589 2378
rect 20681 8338 20747 8358
rect 20681 2358 20747 2378
rect 20839 8338 20905 8358
rect 20839 2358 20905 2378
rect 20997 8338 21063 8358
rect 20997 2358 21063 2378
rect 21155 8338 21221 8358
rect 21155 2358 21221 2378
rect 21313 8338 21379 8358
rect 21313 2358 21379 2378
rect 21471 8338 21537 8358
rect 21471 2358 21537 2378
rect 21629 8338 21695 8358
rect 21629 2358 21695 2378
rect 21787 8338 21853 8358
rect 21787 2358 21853 2378
rect 21945 8338 22011 8358
rect 21945 2358 22011 2378
rect 22103 8338 22169 8358
rect 22103 2358 22169 2378
rect 22261 8338 22327 8358
rect 22261 2358 22327 2378
rect 22419 8338 22485 8358
rect 22419 2358 22485 2378
rect 22577 8338 22643 8358
rect 22577 2358 22643 2378
rect 22735 8338 22801 8358
rect 22735 2358 22801 2378
rect 22893 8338 22959 8358
rect 22893 2358 22959 2378
rect 23051 8338 23117 8358
rect 23051 2358 23117 2378
rect 23209 8338 23275 8358
rect 23209 2358 23275 2378
rect 23367 8338 23433 8358
rect 23367 2358 23433 2378
rect 23525 8338 23591 8358
rect 23525 2358 23591 2378
rect 23683 8338 23749 8358
rect 23683 2358 23749 2378
rect 23841 8338 23907 8358
rect 23841 2358 23907 2378
rect 23999 8338 24065 8358
rect 23999 2358 24065 2378
rect 24157 8338 24223 8358
rect 24157 2358 24223 2378
rect 24315 8338 24381 8358
rect 24315 2358 24381 2378
rect 24473 8338 24539 8358
rect 24473 2358 24539 2378
rect 24631 8338 24697 8358
rect 24631 2358 24697 2378
rect 24789 8338 24855 8358
rect 24789 2358 24855 2378
rect 24947 8338 25013 8358
rect 24947 2358 25013 2378
rect 25105 8338 25171 8358
rect 25105 2358 25171 2378
rect 20432 2310 20452 2326
rect 25086 2310 25106 2326
rect 20432 2240 20440 2310
rect 25090 2240 25106 2310
rect 20432 2226 20452 2240
rect 25086 2226 25106 2240
rect 19980 2150 20000 2200
rect 19500 2140 20000 2150
rect 13140 2020 13150 2090
rect 13350 2020 13360 2090
rect 7140 1910 7150 1980
rect 7350 1910 7360 1980
rect 7140 1860 7360 1910
rect 7640 1980 7860 2000
rect 7640 1910 7650 1980
rect 7850 1910 7860 1980
rect 7640 1860 7860 1910
rect 8140 1980 8360 2000
rect 8140 1910 8150 1980
rect 8350 1910 8360 1980
rect 8140 1860 8360 1910
rect 8640 1980 8860 2000
rect 8640 1910 8650 1980
rect 8850 1910 8860 1980
rect 8640 1860 8860 1910
rect 9140 1980 9360 2000
rect 9140 1910 9150 1980
rect 9350 1910 9360 1980
rect 9140 1860 9360 1910
rect 9640 1980 9860 2000
rect 9640 1910 9650 1980
rect 9850 1910 9860 1980
rect 9640 1860 9860 1910
rect 10140 1980 10360 2000
rect 10140 1910 10150 1980
rect 10350 1910 10360 1980
rect 10140 1860 10360 1910
rect 10640 1980 10860 2000
rect 10640 1910 10650 1980
rect 10850 1910 10860 1980
rect 10640 1860 10860 1910
rect 11140 1980 11360 2000
rect 11140 1910 11150 1980
rect 11350 1910 11360 1980
rect 11140 1860 11360 1910
rect 11640 1980 11860 2000
rect 11640 1910 11650 1980
rect 11850 1910 11860 1980
rect 11640 1860 11860 1910
rect 12140 1980 12360 2000
rect 12140 1910 12150 1980
rect 12350 1910 12360 1980
rect 12140 1860 12360 1910
rect 12640 1980 12860 2000
rect 12640 1910 12650 1980
rect 12850 1910 12860 1980
rect 12640 1860 12860 1910
rect 13140 1980 13360 2020
rect 19640 2090 19860 2140
rect 20230 2130 20300 2200
rect 25640 8520 25650 8590
rect 25850 8520 25860 8590
rect 25640 8480 25860 8520
rect 25640 8410 25650 8480
rect 25850 8410 25860 8480
rect 25640 8360 25860 8410
rect 26140 8590 26360 8640
rect 26140 8520 26150 8590
rect 26350 8520 26360 8590
rect 26140 8480 26360 8520
rect 26140 8410 26150 8480
rect 26350 8410 26360 8480
rect 26140 8360 26360 8410
rect 25500 8350 26500 8360
rect 25500 8150 25520 8350
rect 25590 8150 25910 8350
rect 25980 8150 26020 8350
rect 26090 8150 26410 8350
rect 26480 8150 26500 8350
rect 25500 8140 26500 8150
rect 25640 8090 25860 8140
rect 25640 8020 25650 8090
rect 25850 8020 25860 8090
rect 25640 7980 25860 8020
rect 25640 7910 25650 7980
rect 25850 7910 25860 7980
rect 25640 7860 25860 7910
rect 26140 8090 26360 8140
rect 26140 8020 26150 8090
rect 26350 8020 26360 8090
rect 26140 7980 26360 8020
rect 26140 7910 26150 7980
rect 26350 7910 26360 7980
rect 26140 7860 26360 7910
rect 25500 7850 26500 7860
rect 25500 7650 25520 7850
rect 25590 7650 25910 7850
rect 25980 7650 26020 7850
rect 26090 7650 26410 7850
rect 26480 7650 26500 7850
rect 25500 7640 26500 7650
rect 25640 7590 25860 7640
rect 25640 7520 25650 7590
rect 25850 7520 25860 7590
rect 25640 7480 25860 7520
rect 25640 7410 25650 7480
rect 25850 7410 25860 7480
rect 25640 7360 25860 7410
rect 26140 7590 26360 7640
rect 26140 7520 26150 7590
rect 26350 7520 26360 7590
rect 26140 7480 26360 7520
rect 26140 7410 26150 7480
rect 26350 7410 26360 7480
rect 26140 7360 26360 7410
rect 25500 7350 26500 7360
rect 25500 7150 25520 7350
rect 25590 7150 25910 7350
rect 25980 7150 26020 7350
rect 26090 7150 26410 7350
rect 26480 7150 26500 7350
rect 25500 7140 26500 7150
rect 25640 7090 25860 7140
rect 25640 7020 25650 7090
rect 25850 7020 25860 7090
rect 25640 6980 25860 7020
rect 25640 6910 25650 6980
rect 25850 6910 25860 6980
rect 25640 6860 25860 6910
rect 26140 7090 26360 7140
rect 26140 7020 26150 7090
rect 26350 7020 26360 7090
rect 26140 6980 26360 7020
rect 26140 6910 26150 6980
rect 26350 6910 26360 6980
rect 26140 6860 26360 6910
rect 25500 6850 26500 6860
rect 25500 6650 25520 6850
rect 25590 6650 25910 6850
rect 25980 6650 26020 6850
rect 26090 6650 26410 6850
rect 26480 6650 26500 6850
rect 25500 6640 26500 6650
rect 25640 6590 25860 6640
rect 25640 6520 25650 6590
rect 25850 6520 25860 6590
rect 25640 6480 25860 6520
rect 25640 6410 25650 6480
rect 25850 6410 25860 6480
rect 25640 6360 25860 6410
rect 26140 6590 26360 6640
rect 26140 6520 26150 6590
rect 26350 6520 26360 6590
rect 26140 6480 26360 6520
rect 26140 6410 26150 6480
rect 26350 6410 26360 6480
rect 26140 6360 26360 6410
rect 25500 6350 26500 6360
rect 25500 6150 25520 6350
rect 25590 6150 25910 6350
rect 25980 6150 26020 6350
rect 26090 6150 26410 6350
rect 26480 6150 26500 6350
rect 25500 6140 26500 6150
rect 25640 6090 25860 6140
rect 25640 6020 25650 6090
rect 25850 6020 25860 6090
rect 25640 5980 25860 6020
rect 25640 5910 25650 5980
rect 25850 5910 25860 5980
rect 25640 5860 25860 5910
rect 26140 6090 26360 6140
rect 26140 6020 26150 6090
rect 26350 6020 26360 6090
rect 26140 5980 26360 6020
rect 26140 5910 26150 5980
rect 26350 5910 26360 5980
rect 26140 5860 26360 5910
rect 25500 5850 26500 5860
rect 25500 5650 25520 5850
rect 25590 5650 25910 5850
rect 25980 5650 26020 5850
rect 26090 5650 26410 5850
rect 26480 5650 26500 5850
rect 25500 5640 26500 5650
rect 25640 5590 25860 5640
rect 25640 5520 25650 5590
rect 25850 5520 25860 5590
rect 25640 5480 25860 5520
rect 25640 5410 25650 5480
rect 25850 5410 25860 5480
rect 25640 5360 25860 5410
rect 26140 5590 26360 5640
rect 26140 5520 26150 5590
rect 26350 5520 26360 5590
rect 26140 5480 26360 5520
rect 26140 5410 26150 5480
rect 26350 5410 26360 5480
rect 26140 5360 26360 5410
rect 25500 5350 26500 5360
rect 25500 5150 25520 5350
rect 25590 5150 25910 5350
rect 25980 5150 26020 5350
rect 26090 5150 26410 5350
rect 26480 5150 26500 5350
rect 25500 5140 26500 5150
rect 25640 5090 25860 5140
rect 25640 5020 25650 5090
rect 25850 5020 25860 5090
rect 25640 4980 25860 5020
rect 25640 4910 25650 4980
rect 25850 4910 25860 4980
rect 25640 4860 25860 4910
rect 26140 5090 26360 5140
rect 26140 5020 26150 5090
rect 26350 5020 26360 5090
rect 26140 4980 26360 5020
rect 26140 4910 26150 4980
rect 26350 4910 26360 4980
rect 26140 4860 26360 4910
rect 25500 4850 26500 4860
rect 25500 4650 25520 4850
rect 25590 4650 25910 4850
rect 25980 4650 26020 4850
rect 26090 4650 26410 4850
rect 26480 4650 26500 4850
rect 25500 4640 26500 4650
rect 25640 4590 25860 4640
rect 25640 4520 25650 4590
rect 25850 4520 25860 4590
rect 25640 4480 25860 4520
rect 25640 4410 25650 4480
rect 25850 4410 25860 4480
rect 25640 4360 25860 4410
rect 26140 4590 26360 4640
rect 26140 4520 26150 4590
rect 26350 4520 26360 4590
rect 26140 4480 26360 4520
rect 26140 4410 26150 4480
rect 26350 4410 26360 4480
rect 26140 4360 26360 4410
rect 25500 4350 26500 4360
rect 25500 4150 25520 4350
rect 25590 4150 25910 4350
rect 25980 4150 26020 4350
rect 26090 4150 26410 4350
rect 26480 4150 26500 4350
rect 25500 4140 26500 4150
rect 25640 4090 25860 4140
rect 25640 4020 25650 4090
rect 25850 4020 25860 4090
rect 25640 3980 25860 4020
rect 25640 3910 25650 3980
rect 25850 3910 25860 3980
rect 25640 3860 25860 3910
rect 26140 4090 26360 4140
rect 26140 4020 26150 4090
rect 26350 4020 26360 4090
rect 26140 3980 26360 4020
rect 26140 3910 26150 3980
rect 26350 3910 26360 3980
rect 26140 3860 26360 3910
rect 25500 3850 26500 3860
rect 25500 3650 25520 3850
rect 25590 3650 25910 3850
rect 25980 3650 26020 3850
rect 26090 3650 26410 3850
rect 26480 3650 26500 3850
rect 25500 3640 26500 3650
rect 25640 3590 25860 3640
rect 25640 3520 25650 3590
rect 25850 3520 25860 3590
rect 25640 3480 25860 3520
rect 25640 3410 25650 3480
rect 25850 3410 25860 3480
rect 25640 3360 25860 3410
rect 26140 3590 26360 3640
rect 26140 3520 26150 3590
rect 26350 3520 26360 3590
rect 26140 3480 26360 3520
rect 26140 3410 26150 3480
rect 26350 3410 26360 3480
rect 26140 3360 26360 3410
rect 25500 3350 26500 3360
rect 25500 3150 25520 3350
rect 25590 3150 25910 3350
rect 25980 3150 26020 3350
rect 26090 3150 26410 3350
rect 26480 3150 26500 3350
rect 25500 3140 26500 3150
rect 25640 3090 25860 3140
rect 25640 3020 25650 3090
rect 25850 3020 25860 3090
rect 25640 2980 25860 3020
rect 25640 2910 25650 2980
rect 25850 2910 25860 2980
rect 25640 2860 25860 2910
rect 26140 3090 26360 3140
rect 26140 3020 26150 3090
rect 26350 3020 26360 3090
rect 26140 2980 26360 3020
rect 26140 2910 26150 2980
rect 26350 2910 26360 2980
rect 26140 2860 26360 2910
rect 25500 2850 26500 2860
rect 25500 2650 25520 2850
rect 25590 2650 25910 2850
rect 25980 2650 26020 2850
rect 26090 2650 26410 2850
rect 26480 2650 26500 2850
rect 25500 2640 26500 2650
rect 25640 2590 25860 2640
rect 25640 2520 25650 2590
rect 25850 2520 25860 2590
rect 25640 2480 25860 2520
rect 25640 2410 25650 2480
rect 25850 2410 25860 2480
rect 25640 2360 25860 2410
rect 26140 2590 26360 2640
rect 26140 2520 26150 2590
rect 26350 2520 26360 2590
rect 26140 2480 26360 2520
rect 26140 2410 26150 2480
rect 26350 2410 26360 2480
rect 26140 2360 26360 2410
rect 25240 2130 25310 2200
rect 25500 2350 26500 2360
rect 25500 2150 25520 2350
rect 25590 2150 25910 2350
rect 25980 2150 26020 2350
rect 26090 2150 26410 2350
rect 26480 2150 26500 2350
rect 25500 2140 26500 2150
rect 19640 2020 19650 2090
rect 19850 2020 19860 2090
rect 13140 1910 13150 1980
rect 13350 1910 13360 1980
rect 13140 1860 13360 1910
rect 13640 1980 13860 2000
rect 13640 1910 13650 1980
rect 13850 1910 13860 1980
rect 13640 1860 13860 1910
rect 14140 1980 14360 2000
rect 14140 1910 14150 1980
rect 14350 1910 14360 1980
rect 14140 1860 14360 1910
rect 14640 1980 14860 2000
rect 14640 1910 14650 1980
rect 14850 1910 14860 1980
rect 14640 1860 14860 1910
rect 15140 1980 15360 2000
rect 15140 1910 15150 1980
rect 15350 1910 15360 1980
rect 15140 1860 15360 1910
rect 15640 1980 15860 2000
rect 15640 1910 15650 1980
rect 15850 1910 15860 1980
rect 15640 1860 15860 1910
rect 16140 1980 16360 2000
rect 16140 1910 16150 1980
rect 16350 1910 16360 1980
rect 16140 1860 16360 1910
rect 16640 1980 16860 2000
rect 16640 1910 16650 1980
rect 16850 1910 16860 1980
rect 16640 1860 16860 1910
rect 17140 1980 17360 2000
rect 17140 1910 17150 1980
rect 17350 1910 17360 1980
rect 17140 1860 17360 1910
rect 17640 1980 17860 2000
rect 17640 1910 17650 1980
rect 17850 1910 17860 1980
rect 17640 1860 17860 1910
rect 18140 1980 18360 2000
rect 18140 1910 18150 1980
rect 18350 1910 18360 1980
rect 18140 1860 18360 1910
rect 18640 1980 18860 2000
rect 18640 1910 18650 1980
rect 18850 1910 18860 1980
rect 18640 1860 18860 1910
rect 19140 1980 19360 2000
rect 19140 1910 19150 1980
rect 19350 1910 19360 1980
rect 19140 1860 19360 1910
rect 19640 1980 19860 2020
rect 25640 2090 25860 2140
rect 25640 2020 25650 2090
rect 25850 2020 25860 2090
rect 19640 1910 19650 1980
rect 19850 1910 19860 1980
rect 19640 1860 19860 1910
rect 20140 1980 20360 2000
rect 20140 1910 20150 1980
rect 20350 1910 20360 1980
rect 20140 1860 20360 1910
rect 20640 1980 20860 2000
rect 20640 1910 20650 1980
rect 20850 1910 20860 1980
rect 20640 1860 20860 1910
rect 21140 1980 21360 2000
rect 21140 1910 21150 1980
rect 21350 1910 21360 1980
rect 21140 1860 21360 1910
rect 21640 1980 21860 2000
rect 21640 1910 21650 1980
rect 21850 1910 21860 1980
rect 21640 1860 21860 1910
rect 22140 1980 22360 2000
rect 22140 1910 22150 1980
rect 22350 1910 22360 1980
rect 22140 1860 22360 1910
rect 22640 1980 22860 2000
rect 22640 1910 22650 1980
rect 22850 1910 22860 1980
rect 22640 1860 22860 1910
rect 23140 1980 23360 2000
rect 23140 1910 23150 1980
rect 23350 1910 23360 1980
rect 23140 1860 23360 1910
rect 23640 1980 23860 2000
rect 23640 1910 23650 1980
rect 23850 1910 23860 1980
rect 23640 1860 23860 1910
rect 24140 1980 24360 2000
rect 24140 1910 24150 1980
rect 24350 1910 24360 1980
rect 24140 1860 24360 1910
rect 24640 1980 24860 2000
rect 24640 1910 24650 1980
rect 24850 1910 24860 1980
rect 24640 1860 24860 1910
rect 25140 1980 25360 2000
rect 25140 1910 25150 1980
rect 25350 1910 25360 1980
rect 25140 1860 25360 1910
rect 25640 1980 25860 2020
rect 25640 1910 25650 1980
rect 25850 1910 25860 1980
rect 25640 1860 25860 1910
rect 26140 2090 26360 2140
rect 26140 2020 26150 2090
rect 26350 2020 26360 2090
rect 26140 1980 26360 2020
rect 26140 1910 26150 1980
rect 26350 1910 26360 1980
rect 26140 1860 26360 1910
rect 0 1850 26500 1860
rect 0 1650 20 1850
rect 90 1650 410 1850
rect 480 1650 520 1850
rect 590 1650 910 1850
rect 980 1650 1020 1850
rect 1090 1650 1410 1850
rect 1480 1650 1520 1850
rect 1590 1650 1910 1850
rect 1980 1650 2020 1850
rect 2090 1650 2410 1850
rect 2480 1650 2520 1850
rect 2590 1650 2910 1850
rect 2980 1650 3020 1850
rect 3090 1650 3410 1850
rect 3480 1650 3520 1850
rect 3590 1650 3910 1850
rect 3980 1650 4020 1850
rect 4090 1650 4410 1850
rect 4480 1650 4520 1850
rect 4590 1650 4910 1850
rect 4980 1650 5020 1850
rect 5090 1650 5410 1850
rect 5480 1650 5520 1850
rect 5590 1650 5910 1850
rect 5980 1650 6020 1850
rect 6090 1650 6410 1850
rect 6480 1650 6520 1850
rect 6590 1650 6910 1850
rect 6980 1650 7020 1850
rect 7090 1650 7410 1850
rect 7480 1650 7520 1850
rect 7590 1650 7910 1850
rect 7980 1650 8020 1850
rect 8090 1650 8410 1850
rect 8480 1650 8520 1850
rect 8590 1650 8910 1850
rect 8980 1650 9020 1850
rect 9090 1650 9410 1850
rect 9480 1650 9520 1850
rect 9590 1650 9910 1850
rect 9980 1650 10020 1850
rect 10090 1650 10410 1850
rect 10480 1650 10520 1850
rect 10590 1650 10910 1850
rect 10980 1650 11020 1850
rect 11090 1650 11410 1850
rect 11480 1650 11520 1850
rect 11590 1650 11910 1850
rect 11980 1650 12020 1850
rect 12090 1650 12410 1850
rect 12480 1650 12520 1850
rect 12590 1650 12910 1850
rect 12980 1650 13020 1850
rect 13090 1650 13410 1850
rect 13480 1650 13520 1850
rect 13590 1650 13910 1850
rect 13980 1650 14020 1850
rect 14090 1650 14410 1850
rect 14480 1650 14520 1850
rect 14590 1650 14910 1850
rect 14980 1650 15020 1850
rect 15090 1650 15410 1850
rect 15480 1650 15520 1850
rect 15590 1650 15910 1850
rect 15980 1650 16020 1850
rect 16090 1650 16410 1850
rect 16480 1650 16520 1850
rect 16590 1650 16910 1850
rect 16980 1650 17020 1850
rect 17090 1650 17410 1850
rect 17480 1650 17520 1850
rect 17590 1650 17910 1850
rect 17980 1650 18020 1850
rect 18090 1650 18410 1850
rect 18480 1650 18520 1850
rect 18590 1650 18910 1850
rect 18980 1650 19020 1850
rect 19090 1650 19410 1850
rect 19480 1650 19520 1850
rect 19590 1650 19910 1850
rect 19980 1650 20020 1850
rect 20090 1650 20410 1850
rect 20480 1650 20520 1850
rect 20590 1650 20910 1850
rect 20980 1650 21020 1850
rect 21090 1650 21410 1850
rect 21480 1650 21520 1850
rect 21590 1650 21910 1850
rect 21980 1650 22020 1850
rect 22090 1650 22410 1850
rect 22480 1650 22520 1850
rect 22590 1650 22910 1850
rect 22980 1650 23020 1850
rect 23090 1650 23410 1850
rect 23480 1650 23520 1850
rect 23590 1650 23910 1850
rect 23980 1650 24020 1850
rect 24090 1650 24410 1850
rect 24480 1650 24520 1850
rect 24590 1650 24910 1850
rect 24980 1650 25020 1850
rect 25090 1650 25410 1850
rect 25480 1650 25520 1850
rect 25590 1650 25910 1850
rect 25980 1650 26020 1850
rect 26090 1650 26410 1850
rect 26480 1650 26500 1850
rect 0 1640 26500 1650
rect 140 1590 360 1640
rect 140 1520 150 1590
rect 350 1520 360 1590
rect 140 1480 360 1520
rect 140 1410 150 1480
rect 350 1410 360 1480
rect 140 1360 360 1410
rect 640 1590 860 1640
rect 640 1520 650 1590
rect 850 1520 860 1590
rect 640 1480 860 1520
rect 640 1410 650 1480
rect 850 1410 860 1480
rect 640 1360 860 1410
rect 1140 1590 1360 1640
rect 1140 1520 1150 1590
rect 1350 1520 1360 1590
rect 1140 1480 1360 1520
rect 1140 1410 1150 1480
rect 1350 1410 1360 1480
rect 1140 1360 1360 1410
rect 1640 1590 1860 1640
rect 1640 1520 1650 1590
rect 1850 1520 1860 1590
rect 1640 1480 1860 1520
rect 1640 1410 1650 1480
rect 1850 1410 1860 1480
rect 1640 1360 1860 1410
rect 2140 1590 2360 1640
rect 2140 1520 2150 1590
rect 2350 1520 2360 1590
rect 2140 1480 2360 1520
rect 2140 1410 2150 1480
rect 2350 1410 2360 1480
rect 2140 1360 2360 1410
rect 2640 1590 2860 1640
rect 2640 1520 2650 1590
rect 2850 1520 2860 1590
rect 2640 1480 2860 1520
rect 2640 1410 2650 1480
rect 2850 1410 2860 1480
rect 2640 1360 2860 1410
rect 3140 1590 3360 1640
rect 3140 1520 3150 1590
rect 3350 1520 3360 1590
rect 3140 1480 3360 1520
rect 3140 1410 3150 1480
rect 3350 1410 3360 1480
rect 3140 1360 3360 1410
rect 3640 1590 3860 1640
rect 3640 1520 3650 1590
rect 3850 1520 3860 1590
rect 3640 1480 3860 1520
rect 3640 1410 3650 1480
rect 3850 1410 3860 1480
rect 3640 1360 3860 1410
rect 4140 1590 4360 1640
rect 4140 1520 4150 1590
rect 4350 1520 4360 1590
rect 4140 1480 4360 1520
rect 4140 1410 4150 1480
rect 4350 1410 4360 1480
rect 4140 1360 4360 1410
rect 4640 1590 4860 1640
rect 4640 1520 4650 1590
rect 4850 1520 4860 1590
rect 4640 1480 4860 1520
rect 4640 1410 4650 1480
rect 4850 1410 4860 1480
rect 4640 1360 4860 1410
rect 5140 1590 5360 1640
rect 5140 1520 5150 1590
rect 5350 1520 5360 1590
rect 5140 1480 5360 1520
rect 5140 1410 5150 1480
rect 5350 1410 5360 1480
rect 5140 1360 5360 1410
rect 5640 1590 5860 1640
rect 5640 1520 5650 1590
rect 5850 1520 5860 1590
rect 5640 1480 5860 1520
rect 5640 1410 5650 1480
rect 5850 1410 5860 1480
rect 5640 1360 5860 1410
rect 6140 1590 6360 1640
rect 6140 1520 6150 1590
rect 6350 1520 6360 1590
rect 6140 1480 6360 1520
rect 6140 1410 6150 1480
rect 6350 1410 6360 1480
rect 6140 1360 6360 1410
rect 6640 1590 6860 1640
rect 6640 1520 6650 1590
rect 6850 1520 6860 1590
rect 6640 1480 6860 1520
rect 6640 1410 6650 1480
rect 6850 1410 6860 1480
rect 6640 1360 6860 1410
rect 7140 1590 7360 1640
rect 7140 1520 7150 1590
rect 7350 1520 7360 1590
rect 7140 1480 7360 1520
rect 7140 1410 7150 1480
rect 7350 1410 7360 1480
rect 7140 1360 7360 1410
rect 7640 1590 7860 1640
rect 7640 1520 7650 1590
rect 7850 1520 7860 1590
rect 7640 1480 7860 1520
rect 7640 1410 7650 1480
rect 7850 1410 7860 1480
rect 7640 1360 7860 1410
rect 8140 1590 8360 1640
rect 8140 1520 8150 1590
rect 8350 1520 8360 1590
rect 8140 1480 8360 1520
rect 8140 1410 8150 1480
rect 8350 1410 8360 1480
rect 8140 1360 8360 1410
rect 8640 1590 8860 1640
rect 8640 1520 8650 1590
rect 8850 1520 8860 1590
rect 8640 1480 8860 1520
rect 8640 1410 8650 1480
rect 8850 1410 8860 1480
rect 8640 1360 8860 1410
rect 9140 1590 9360 1640
rect 9140 1520 9150 1590
rect 9350 1520 9360 1590
rect 9140 1480 9360 1520
rect 9140 1410 9150 1480
rect 9350 1410 9360 1480
rect 9140 1360 9360 1410
rect 9640 1590 9860 1640
rect 9640 1520 9650 1590
rect 9850 1520 9860 1590
rect 9640 1480 9860 1520
rect 9640 1410 9650 1480
rect 9850 1410 9860 1480
rect 9640 1360 9860 1410
rect 10140 1590 10360 1640
rect 10140 1520 10150 1590
rect 10350 1520 10360 1590
rect 10140 1480 10360 1520
rect 10140 1410 10150 1480
rect 10350 1410 10360 1480
rect 10140 1360 10360 1410
rect 10640 1590 10860 1640
rect 10640 1520 10650 1590
rect 10850 1520 10860 1590
rect 10640 1480 10860 1520
rect 10640 1410 10650 1480
rect 10850 1410 10860 1480
rect 10640 1360 10860 1410
rect 11140 1590 11360 1640
rect 11140 1520 11150 1590
rect 11350 1520 11360 1590
rect 11140 1480 11360 1520
rect 11140 1410 11150 1480
rect 11350 1410 11360 1480
rect 11140 1360 11360 1410
rect 11640 1590 11860 1640
rect 11640 1520 11650 1590
rect 11850 1520 11860 1590
rect 11640 1480 11860 1520
rect 11640 1410 11650 1480
rect 11850 1410 11860 1480
rect 11640 1360 11860 1410
rect 12140 1590 12360 1640
rect 12140 1520 12150 1590
rect 12350 1520 12360 1590
rect 12140 1480 12360 1520
rect 12140 1410 12150 1480
rect 12350 1410 12360 1480
rect 12140 1360 12360 1410
rect 12640 1590 12860 1640
rect 12640 1520 12650 1590
rect 12850 1520 12860 1590
rect 12640 1480 12860 1520
rect 12640 1410 12650 1480
rect 12850 1410 12860 1480
rect 12640 1360 12860 1410
rect 13140 1590 13360 1640
rect 13140 1520 13150 1590
rect 13350 1520 13360 1590
rect 13140 1480 13360 1520
rect 13140 1410 13150 1480
rect 13350 1410 13360 1480
rect 13140 1360 13360 1410
rect 13640 1590 13860 1640
rect 13640 1520 13650 1590
rect 13850 1520 13860 1590
rect 13640 1480 13860 1520
rect 13640 1410 13650 1480
rect 13850 1410 13860 1480
rect 13640 1360 13860 1410
rect 14140 1590 14360 1640
rect 14140 1520 14150 1590
rect 14350 1520 14360 1590
rect 14140 1480 14360 1520
rect 14140 1410 14150 1480
rect 14350 1410 14360 1480
rect 14140 1360 14360 1410
rect 14640 1590 14860 1640
rect 14640 1520 14650 1590
rect 14850 1520 14860 1590
rect 14640 1480 14860 1520
rect 14640 1410 14650 1480
rect 14850 1410 14860 1480
rect 14640 1360 14860 1410
rect 15140 1590 15360 1640
rect 15140 1520 15150 1590
rect 15350 1520 15360 1590
rect 15140 1480 15360 1520
rect 15140 1410 15150 1480
rect 15350 1410 15360 1480
rect 15140 1360 15360 1410
rect 15640 1590 15860 1640
rect 15640 1520 15650 1590
rect 15850 1520 15860 1590
rect 15640 1480 15860 1520
rect 15640 1410 15650 1480
rect 15850 1410 15860 1480
rect 15640 1360 15860 1410
rect 16140 1590 16360 1640
rect 16140 1520 16150 1590
rect 16350 1520 16360 1590
rect 16140 1480 16360 1520
rect 16140 1410 16150 1480
rect 16350 1410 16360 1480
rect 16140 1360 16360 1410
rect 16640 1590 16860 1640
rect 16640 1520 16650 1590
rect 16850 1520 16860 1590
rect 16640 1480 16860 1520
rect 16640 1410 16650 1480
rect 16850 1410 16860 1480
rect 16640 1360 16860 1410
rect 17140 1590 17360 1640
rect 17140 1520 17150 1590
rect 17350 1520 17360 1590
rect 17140 1480 17360 1520
rect 17140 1410 17150 1480
rect 17350 1410 17360 1480
rect 17140 1360 17360 1410
rect 17640 1590 17860 1640
rect 17640 1520 17650 1590
rect 17850 1520 17860 1590
rect 17640 1480 17860 1520
rect 17640 1410 17650 1480
rect 17850 1410 17860 1480
rect 17640 1360 17860 1410
rect 18140 1590 18360 1640
rect 18140 1520 18150 1590
rect 18350 1520 18360 1590
rect 18140 1480 18360 1520
rect 18140 1410 18150 1480
rect 18350 1410 18360 1480
rect 18140 1360 18360 1410
rect 18640 1590 18860 1640
rect 18640 1520 18650 1590
rect 18850 1520 18860 1590
rect 18640 1480 18860 1520
rect 18640 1410 18650 1480
rect 18850 1410 18860 1480
rect 18640 1360 18860 1410
rect 19140 1590 19360 1640
rect 19140 1520 19150 1590
rect 19350 1520 19360 1590
rect 19140 1480 19360 1520
rect 19140 1410 19150 1480
rect 19350 1410 19360 1480
rect 19140 1360 19360 1410
rect 19640 1590 19860 1640
rect 19640 1520 19650 1590
rect 19850 1520 19860 1590
rect 19640 1480 19860 1520
rect 19640 1410 19650 1480
rect 19850 1410 19860 1480
rect 19640 1360 19860 1410
rect 20140 1590 20360 1640
rect 20140 1520 20150 1590
rect 20350 1520 20360 1590
rect 20140 1480 20360 1520
rect 20140 1410 20150 1480
rect 20350 1410 20360 1480
rect 20140 1360 20360 1410
rect 20640 1590 20860 1640
rect 20640 1520 20650 1590
rect 20850 1520 20860 1590
rect 20640 1480 20860 1520
rect 20640 1410 20650 1480
rect 20850 1410 20860 1480
rect 20640 1360 20860 1410
rect 21140 1590 21360 1640
rect 21140 1520 21150 1590
rect 21350 1520 21360 1590
rect 21140 1480 21360 1520
rect 21140 1410 21150 1480
rect 21350 1410 21360 1480
rect 21140 1360 21360 1410
rect 21640 1590 21860 1640
rect 21640 1520 21650 1590
rect 21850 1520 21860 1590
rect 21640 1480 21860 1520
rect 21640 1410 21650 1480
rect 21850 1410 21860 1480
rect 21640 1360 21860 1410
rect 22140 1590 22360 1640
rect 22140 1520 22150 1590
rect 22350 1520 22360 1590
rect 22140 1480 22360 1520
rect 22140 1410 22150 1480
rect 22350 1410 22360 1480
rect 22140 1360 22360 1410
rect 22640 1590 22860 1640
rect 22640 1520 22650 1590
rect 22850 1520 22860 1590
rect 22640 1480 22860 1520
rect 22640 1410 22650 1480
rect 22850 1410 22860 1480
rect 22640 1360 22860 1410
rect 23140 1590 23360 1640
rect 23140 1520 23150 1590
rect 23350 1520 23360 1590
rect 23140 1480 23360 1520
rect 23140 1410 23150 1480
rect 23350 1410 23360 1480
rect 23140 1360 23360 1410
rect 23640 1590 23860 1640
rect 23640 1520 23650 1590
rect 23850 1520 23860 1590
rect 23640 1480 23860 1520
rect 23640 1410 23650 1480
rect 23850 1410 23860 1480
rect 23640 1360 23860 1410
rect 24140 1590 24360 1640
rect 24140 1520 24150 1590
rect 24350 1520 24360 1590
rect 24140 1480 24360 1520
rect 24140 1410 24150 1480
rect 24350 1410 24360 1480
rect 24140 1360 24360 1410
rect 24640 1590 24860 1640
rect 24640 1520 24650 1590
rect 24850 1520 24860 1590
rect 24640 1480 24860 1520
rect 24640 1410 24650 1480
rect 24850 1410 24860 1480
rect 24640 1360 24860 1410
rect 25140 1590 25360 1640
rect 25140 1520 25150 1590
rect 25350 1520 25360 1590
rect 25140 1480 25360 1520
rect 25140 1410 25150 1480
rect 25350 1410 25360 1480
rect 25140 1360 25360 1410
rect 25640 1590 25860 1640
rect 25640 1520 25650 1590
rect 25850 1520 25860 1590
rect 25640 1480 25860 1520
rect 25640 1410 25650 1480
rect 25850 1410 25860 1480
rect 25640 1360 25860 1410
rect 26140 1590 26360 1640
rect 26140 1520 26150 1590
rect 26350 1520 26360 1590
rect 26140 1480 26360 1520
rect 26140 1410 26150 1480
rect 26350 1410 26360 1480
rect 26140 1360 26360 1410
rect 0 1350 26500 1360
rect 0 1150 20 1350
rect 90 1150 410 1350
rect 480 1150 520 1350
rect 590 1150 910 1350
rect 980 1150 1020 1350
rect 1090 1150 1410 1350
rect 1480 1150 1520 1350
rect 1590 1150 1910 1350
rect 1980 1150 2020 1350
rect 2090 1150 2410 1350
rect 2480 1150 2520 1350
rect 2590 1150 2910 1350
rect 2980 1150 3020 1350
rect 3090 1150 3410 1350
rect 3480 1150 3520 1350
rect 3590 1150 3910 1350
rect 3980 1150 4020 1350
rect 4090 1150 4410 1350
rect 4480 1150 4520 1350
rect 4590 1150 4910 1350
rect 4980 1150 5020 1350
rect 5090 1150 5410 1350
rect 5480 1150 5520 1350
rect 5590 1150 5910 1350
rect 5980 1150 6020 1350
rect 6090 1150 6410 1350
rect 6480 1150 6520 1350
rect 6590 1150 6910 1350
rect 6980 1150 7020 1350
rect 7090 1150 7410 1350
rect 7480 1150 7520 1350
rect 7590 1150 7910 1350
rect 7980 1150 8020 1350
rect 8090 1150 8410 1350
rect 8480 1150 8520 1350
rect 8590 1150 8910 1350
rect 8980 1150 9020 1350
rect 9090 1150 9410 1350
rect 9480 1150 9520 1350
rect 9590 1150 9910 1350
rect 9980 1150 10020 1350
rect 10090 1150 10410 1350
rect 10480 1150 10520 1350
rect 10590 1150 10910 1350
rect 10980 1150 11020 1350
rect 11090 1150 11410 1350
rect 11480 1150 11520 1350
rect 11590 1150 11910 1350
rect 11980 1150 12020 1350
rect 12090 1150 12410 1350
rect 12480 1150 12520 1350
rect 12590 1150 12910 1350
rect 12980 1150 13020 1350
rect 13090 1150 13410 1350
rect 13480 1150 13520 1350
rect 13590 1150 13910 1350
rect 13980 1150 14020 1350
rect 14090 1150 14410 1350
rect 14480 1150 14520 1350
rect 14590 1150 14910 1350
rect 14980 1150 15020 1350
rect 15090 1150 15410 1350
rect 15480 1150 15520 1350
rect 15590 1150 15910 1350
rect 15980 1150 16020 1350
rect 16090 1150 16410 1350
rect 16480 1150 16520 1350
rect 16590 1150 16910 1350
rect 16980 1150 17020 1350
rect 17090 1150 17410 1350
rect 17480 1150 17520 1350
rect 17590 1150 17910 1350
rect 17980 1150 18020 1350
rect 18090 1150 18410 1350
rect 18480 1150 18520 1350
rect 18590 1150 18910 1350
rect 18980 1150 19020 1350
rect 19090 1150 19410 1350
rect 19480 1150 19520 1350
rect 19590 1150 19910 1350
rect 19980 1150 20020 1350
rect 20090 1150 20410 1350
rect 20480 1150 20520 1350
rect 20590 1150 20910 1350
rect 20980 1150 21020 1350
rect 21090 1150 21410 1350
rect 21480 1150 21520 1350
rect 21590 1150 21910 1350
rect 21980 1150 22020 1350
rect 22090 1150 22410 1350
rect 22480 1150 22520 1350
rect 22590 1150 22910 1350
rect 22980 1150 23020 1350
rect 23090 1150 23410 1350
rect 23480 1150 23520 1350
rect 23590 1150 23910 1350
rect 23980 1150 24020 1350
rect 24090 1150 24410 1350
rect 24480 1150 24520 1350
rect 24590 1150 24910 1350
rect 24980 1150 25020 1350
rect 25090 1150 25410 1350
rect 25480 1150 25520 1350
rect 25590 1150 25910 1350
rect 25980 1150 26020 1350
rect 26090 1150 26410 1350
rect 26480 1150 26500 1350
rect 0 1140 26500 1150
rect 140 1090 360 1140
rect 140 1020 150 1090
rect 350 1020 360 1090
rect 140 1000 360 1020
rect 640 1090 860 1140
rect 640 1020 650 1090
rect 850 1020 860 1090
rect 640 1000 860 1020
rect 1140 1090 1360 1140
rect 1140 1020 1150 1090
rect 1350 1020 1360 1090
rect 1140 1000 1360 1020
rect 1640 1090 1860 1140
rect 1640 1020 1650 1090
rect 1850 1020 1860 1090
rect 1640 1000 1860 1020
rect 2140 1090 2360 1140
rect 2140 1020 2150 1090
rect 2350 1020 2360 1090
rect 2140 1000 2360 1020
rect 2640 1090 2860 1140
rect 2640 1020 2650 1090
rect 2850 1020 2860 1090
rect 2640 1000 2860 1020
rect 3140 1090 3360 1140
rect 3140 1020 3150 1090
rect 3350 1020 3360 1090
rect 3140 1000 3360 1020
rect 3640 1090 3860 1140
rect 3640 1020 3650 1090
rect 3850 1020 3860 1090
rect 3640 1000 3860 1020
rect 4140 1090 4360 1140
rect 4140 1020 4150 1090
rect 4350 1020 4360 1090
rect 4140 1000 4360 1020
rect 4640 1090 4860 1140
rect 4640 1020 4650 1090
rect 4850 1020 4860 1090
rect 4640 1000 4860 1020
rect 5140 1090 5360 1140
rect 5140 1020 5150 1090
rect 5350 1020 5360 1090
rect 5140 1000 5360 1020
rect 5640 1090 5860 1140
rect 5640 1020 5650 1090
rect 5850 1020 5860 1090
rect 5640 1000 5860 1020
rect 6140 1090 6360 1140
rect 6140 1020 6150 1090
rect 6350 1020 6360 1090
rect 6140 1000 6360 1020
rect 6640 1090 6860 1140
rect 6640 1020 6650 1090
rect 6850 1020 6860 1090
rect 6640 1000 6860 1020
rect 7140 1090 7360 1140
rect 7140 1020 7150 1090
rect 7350 1020 7360 1090
rect 7140 1000 7360 1020
rect 7640 1090 7860 1140
rect 7640 1020 7650 1090
rect 7850 1020 7860 1090
rect 7640 1000 7860 1020
rect 8140 1090 8360 1140
rect 8140 1020 8150 1090
rect 8350 1020 8360 1090
rect 8140 1000 8360 1020
rect 8640 1090 8860 1140
rect 8640 1020 8650 1090
rect 8850 1020 8860 1090
rect 8640 1000 8860 1020
rect 9140 1090 9360 1140
rect 9140 1020 9150 1090
rect 9350 1020 9360 1090
rect 9140 1000 9360 1020
rect 9640 1090 9860 1140
rect 9640 1020 9650 1090
rect 9850 1020 9860 1090
rect 9640 1000 9860 1020
rect 10140 1090 10360 1140
rect 10140 1020 10150 1090
rect 10350 1020 10360 1090
rect 10140 1000 10360 1020
rect 10640 1090 10860 1140
rect 10640 1020 10650 1090
rect 10850 1020 10860 1090
rect 10640 1000 10860 1020
rect 11140 1090 11360 1140
rect 11140 1020 11150 1090
rect 11350 1020 11360 1090
rect 11140 1000 11360 1020
rect 11640 1090 11860 1140
rect 11640 1020 11650 1090
rect 11850 1020 11860 1090
rect 11640 1000 11860 1020
rect 12140 1090 12360 1140
rect 12140 1020 12150 1090
rect 12350 1020 12360 1090
rect 12140 1000 12360 1020
rect 12640 1090 12860 1140
rect 12640 1020 12650 1090
rect 12850 1020 12860 1090
rect 12640 1000 12860 1020
rect 13140 1090 13360 1140
rect 13140 1020 13150 1090
rect 13350 1020 13360 1090
rect 13140 1000 13360 1020
rect 13640 1090 13860 1140
rect 13640 1020 13650 1090
rect 13850 1020 13860 1090
rect 13640 1000 13860 1020
rect 14140 1090 14360 1140
rect 14140 1020 14150 1090
rect 14350 1020 14360 1090
rect 14140 1000 14360 1020
rect 14640 1090 14860 1140
rect 14640 1020 14650 1090
rect 14850 1020 14860 1090
rect 14640 1000 14860 1020
rect 15140 1090 15360 1140
rect 15140 1020 15150 1090
rect 15350 1020 15360 1090
rect 15140 1000 15360 1020
rect 15640 1090 15860 1140
rect 15640 1020 15650 1090
rect 15850 1020 15860 1090
rect 15640 1000 15860 1020
rect 16140 1090 16360 1140
rect 16140 1020 16150 1090
rect 16350 1020 16360 1090
rect 16140 1000 16360 1020
rect 16640 1090 16860 1140
rect 16640 1020 16650 1090
rect 16850 1020 16860 1090
rect 16640 1000 16860 1020
rect 17140 1090 17360 1140
rect 17140 1020 17150 1090
rect 17350 1020 17360 1090
rect 17140 1000 17360 1020
rect 17640 1090 17860 1140
rect 17640 1020 17650 1090
rect 17850 1020 17860 1090
rect 17640 1000 17860 1020
rect 18140 1090 18360 1140
rect 18140 1020 18150 1090
rect 18350 1020 18360 1090
rect 18140 1000 18360 1020
rect 18640 1090 18860 1140
rect 18640 1020 18650 1090
rect 18850 1020 18860 1090
rect 18640 1000 18860 1020
rect 19140 1090 19360 1140
rect 19140 1020 19150 1090
rect 19350 1020 19360 1090
rect 19140 1000 19360 1020
rect 19640 1090 19860 1140
rect 19640 1020 19650 1090
rect 19850 1020 19860 1090
rect 19640 1000 19860 1020
rect 20140 1090 20360 1140
rect 20140 1020 20150 1090
rect 20350 1020 20360 1090
rect 20140 1000 20360 1020
rect 20640 1090 20860 1140
rect 20640 1020 20650 1090
rect 20850 1020 20860 1090
rect 20640 1000 20860 1020
rect 21140 1090 21360 1140
rect 21140 1020 21150 1090
rect 21350 1020 21360 1090
rect 21140 1000 21360 1020
rect 21640 1090 21860 1140
rect 21640 1020 21650 1090
rect 21850 1020 21860 1090
rect 21640 1000 21860 1020
rect 22140 1090 22360 1140
rect 22140 1020 22150 1090
rect 22350 1020 22360 1090
rect 22140 1000 22360 1020
rect 22640 1090 22860 1140
rect 22640 1020 22650 1090
rect 22850 1020 22860 1090
rect 22640 1000 22860 1020
rect 23140 1090 23360 1140
rect 23140 1020 23150 1090
rect 23350 1020 23360 1090
rect 23140 1000 23360 1020
rect 23640 1090 23860 1140
rect 23640 1020 23650 1090
rect 23850 1020 23860 1090
rect 23640 1000 23860 1020
rect 24140 1090 24360 1140
rect 24140 1020 24150 1090
rect 24350 1020 24360 1090
rect 24140 1000 24360 1020
rect 24640 1090 24860 1140
rect 24640 1020 24650 1090
rect 24850 1020 24860 1090
rect 24640 1000 24860 1020
rect 25140 1090 25360 1140
rect 25140 1020 25150 1090
rect 25350 1020 25360 1090
rect 25140 1000 25360 1020
rect 25640 1090 25860 1140
rect 25640 1020 25650 1090
rect 25850 1020 25860 1090
rect 25640 1000 25860 1020
rect 26140 1090 26360 1140
rect 26140 1020 26150 1090
rect 26350 1020 26360 1090
rect 26140 1000 26360 1020
<< via2 >>
rect -3290 40190 -3110 40450
rect 1540 46010 1552 46080
rect 1552 46010 6186 46080
rect 6186 46010 6200 46080
rect 1465 40585 1531 42345
rect 1623 43585 1689 45345
rect 1781 40585 1847 42345
rect 1939 43585 2005 45345
rect 2097 40585 2163 42345
rect 2255 43585 2321 45345
rect 2413 40585 2479 42345
rect 2571 43585 2637 45345
rect 2729 40585 2795 42345
rect 2887 43585 2953 45345
rect 3045 40585 3111 42345
rect 3203 43585 3269 45345
rect 3361 40585 3427 42345
rect 3519 43585 3585 45345
rect 3677 40585 3743 42345
rect 3835 43585 3901 45345
rect 3993 40585 4059 42345
rect 4151 43585 4217 45345
rect 4309 40585 4375 42345
rect 4467 43585 4533 45345
rect 4625 40585 4691 42345
rect 4783 43585 4849 45345
rect 4941 40585 5007 42345
rect 5099 43585 5165 45345
rect 5257 40585 5323 42345
rect 5415 43585 5481 45345
rect 5573 40585 5639 42345
rect 5731 43585 5797 45345
rect 5889 40585 5955 42345
rect 6047 43585 6113 45345
rect 6205 40585 6271 42345
rect 1540 39840 1552 39910
rect 1552 39840 6186 39910
rect 6186 39840 6190 39910
rect 7840 46010 7852 46080
rect 7852 46010 12486 46080
rect 12486 46010 12500 46080
rect 7765 40585 7831 42345
rect 7923 43585 7989 45345
rect 8081 40585 8147 42345
rect 8239 43585 8305 45345
rect 8397 40585 8463 42345
rect 8555 43585 8621 45345
rect 8713 40585 8779 42345
rect 8871 43585 8937 45345
rect 9029 40585 9095 42345
rect 9187 43585 9253 45345
rect 9345 40585 9411 42345
rect 9503 43585 9569 45345
rect 9661 40585 9727 42345
rect 9819 43585 9885 45345
rect 9977 40585 10043 42345
rect 10135 43585 10201 45345
rect 10293 40585 10359 42345
rect 10451 43585 10517 45345
rect 10609 40585 10675 42345
rect 10767 43585 10833 45345
rect 10925 40585 10991 42345
rect 11083 43585 11149 45345
rect 11241 40585 11307 42345
rect 11399 43585 11465 45345
rect 11557 40585 11623 42345
rect 11715 43585 11781 45345
rect 11873 40585 11939 42345
rect 12031 43585 12097 45345
rect 12189 40585 12255 42345
rect 12347 43585 12413 45345
rect 12505 40585 12571 42345
rect 7840 39840 7852 39910
rect 7852 39840 12486 39910
rect 12486 39840 12490 39910
rect 14140 46010 14152 46080
rect 14152 46010 18786 46080
rect 18786 46010 18800 46080
rect 14065 40585 14131 42345
rect 14223 43585 14289 45345
rect 14381 40585 14447 42345
rect 14539 43585 14605 45345
rect 14697 40585 14763 42345
rect 14855 43585 14921 45345
rect 15013 40585 15079 42345
rect 15171 43585 15237 45345
rect 15329 40585 15395 42345
rect 15487 43585 15553 45345
rect 15645 40585 15711 42345
rect 15803 43585 15869 45345
rect 15961 40585 16027 42345
rect 16119 43585 16185 45345
rect 16277 40585 16343 42345
rect 16435 43585 16501 45345
rect 16593 40585 16659 42345
rect 16751 43585 16817 45345
rect 16909 40585 16975 42345
rect 17067 43585 17133 45345
rect 17225 40585 17291 42345
rect 17383 43585 17449 45345
rect 17541 40585 17607 42345
rect 17699 43585 17765 45345
rect 17857 40585 17923 42345
rect 18015 43585 18081 45345
rect 18173 40585 18239 42345
rect 18331 43585 18397 45345
rect 18489 40585 18555 42345
rect 18647 43585 18713 45345
rect 18805 40585 18871 42345
rect 14140 39840 14152 39910
rect 14152 39840 18786 39910
rect 18786 39840 18790 39910
rect 20440 46010 20452 46080
rect 20452 46010 25086 46080
rect 25086 46010 25100 46080
rect 20365 40585 20431 42345
rect 20523 43585 20589 45345
rect 20681 40585 20747 42345
rect 20839 43585 20905 45345
rect 20997 40585 21063 42345
rect 21155 43585 21221 45345
rect 21313 40585 21379 42345
rect 21471 43585 21537 45345
rect 21629 40585 21695 42345
rect 21787 43585 21853 45345
rect 21945 40585 22011 42345
rect 22103 43585 22169 45345
rect 22261 40585 22327 42345
rect 22419 43585 22485 45345
rect 22577 40585 22643 42345
rect 22735 43585 22801 45345
rect 22893 40585 22959 42345
rect 23051 43585 23117 45345
rect 23209 40585 23275 42345
rect 23367 43585 23433 45345
rect 23525 40585 23591 42345
rect 23683 43585 23749 45345
rect 23841 40585 23907 42345
rect 23999 43585 24065 45345
rect 24157 40585 24223 42345
rect 24315 43585 24381 45345
rect 24473 40585 24539 42345
rect 24631 43585 24697 45345
rect 24789 40585 24855 42345
rect 24947 43585 25013 45345
rect 25105 40585 25171 42345
rect 20440 39840 20452 39910
rect 20452 39840 25086 39910
rect 25086 39840 25090 39910
rect 29910 40190 30090 40450
rect -3290 38690 -3110 38910
rect 1540 39010 1552 39080
rect 1552 39010 6186 39080
rect 6186 39010 6200 39080
rect 1465 33585 1531 35345
rect 1623 36585 1689 38345
rect 1781 33585 1847 35345
rect 1939 36585 2005 38345
rect 2097 33585 2163 35345
rect 2255 36585 2321 38345
rect 2413 33585 2479 35345
rect 2571 36585 2637 38345
rect 2729 33585 2795 35345
rect 2887 36585 2953 38345
rect 3045 33585 3111 35345
rect 3203 36585 3269 38345
rect 3361 33585 3427 35345
rect 3519 36585 3585 38345
rect 3677 33585 3743 35345
rect 3835 36585 3901 38345
rect 3993 33585 4059 35345
rect 4151 36585 4217 38345
rect 4309 33585 4375 35345
rect 4467 36585 4533 38345
rect 4625 33585 4691 35345
rect 4783 36585 4849 38345
rect 4941 33585 5007 35345
rect 5099 36585 5165 38345
rect 5257 33585 5323 35345
rect 5415 36585 5481 38345
rect 5573 33585 5639 35345
rect 5731 36585 5797 38345
rect 5889 33585 5955 35345
rect 6047 36585 6113 38345
rect 6205 33585 6271 35345
rect 1540 32840 1552 32910
rect 1552 32840 6186 32910
rect 6186 32840 6190 32910
rect 7840 39010 7852 39080
rect 7852 39010 12486 39080
rect 12486 39010 12500 39080
rect 7765 33585 7831 35345
rect 7923 36585 7989 38345
rect 8081 33585 8147 35345
rect 8239 36585 8305 38345
rect 8397 33585 8463 35345
rect 8555 36585 8621 38345
rect 8713 33585 8779 35345
rect 8871 36585 8937 38345
rect 9029 33585 9095 35345
rect 9187 36585 9253 38345
rect 9345 33585 9411 35345
rect 9503 36585 9569 38345
rect 9661 33585 9727 35345
rect 9819 36585 9885 38345
rect 9977 33585 10043 35345
rect 10135 36585 10201 38345
rect 10293 33585 10359 35345
rect 10451 36585 10517 38345
rect 10609 33585 10675 35345
rect 10767 36585 10833 38345
rect 10925 33585 10991 35345
rect 11083 36585 11149 38345
rect 11241 33585 11307 35345
rect 11399 36585 11465 38345
rect 11557 33585 11623 35345
rect 11715 36585 11781 38345
rect 11873 33585 11939 35345
rect 12031 36585 12097 38345
rect 12189 33585 12255 35345
rect 12347 36585 12413 38345
rect 12505 33585 12571 35345
rect 7840 32840 7852 32910
rect 7852 32840 12486 32910
rect 12486 32840 12490 32910
rect 14140 39010 14152 39080
rect 14152 39010 18786 39080
rect 18786 39010 18800 39080
rect 14065 33585 14131 35345
rect 14223 36585 14289 38345
rect 14381 33585 14447 35345
rect 14539 36585 14605 38345
rect 14697 33585 14763 35345
rect 14855 36585 14921 38345
rect 15013 33585 15079 35345
rect 15171 36585 15237 38345
rect 15329 33585 15395 35345
rect 15487 36585 15553 38345
rect 15645 33585 15711 35345
rect 15803 36585 15869 38345
rect 15961 33585 16027 35345
rect 16119 36585 16185 38345
rect 16277 33585 16343 35345
rect 16435 36585 16501 38345
rect 16593 33585 16659 35345
rect 16751 36585 16817 38345
rect 16909 33585 16975 35345
rect 17067 36585 17133 38345
rect 17225 33585 17291 35345
rect 17383 36585 17449 38345
rect 17541 33585 17607 35345
rect 17699 36585 17765 38345
rect 17857 33585 17923 35345
rect 18015 36585 18081 38345
rect 18173 33585 18239 35345
rect 18331 36585 18397 38345
rect 18489 33585 18555 35345
rect 18647 36585 18713 38345
rect 18805 33585 18871 35345
rect 14140 32840 14152 32910
rect 14152 32840 18786 32910
rect 18786 32840 18790 32910
rect 20440 39010 20452 39080
rect 20452 39010 25086 39080
rect 25086 39010 25100 39080
rect 20365 33585 20431 35345
rect 20523 36585 20589 38345
rect 20681 33585 20747 35345
rect 20839 36585 20905 38345
rect 20997 33585 21063 35345
rect 21155 36585 21221 38345
rect 21313 33585 21379 35345
rect 21471 36585 21537 38345
rect 21629 33585 21695 35345
rect 21787 36585 21853 38345
rect 21945 33585 22011 35345
rect 22103 36585 22169 38345
rect 22261 33585 22327 35345
rect 22419 36585 22485 38345
rect 22577 33585 22643 35345
rect 22735 36585 22801 38345
rect 22893 33585 22959 35345
rect 23051 36585 23117 38345
rect 23209 33585 23275 35345
rect 23367 36585 23433 38345
rect 23525 33585 23591 35345
rect 23683 36585 23749 38345
rect 23841 33585 23907 35345
rect 23999 36585 24065 38345
rect 24157 33585 24223 35345
rect 24315 36585 24381 38345
rect 24473 33585 24539 35345
rect 24631 36585 24697 38345
rect 24789 33585 24855 35345
rect 24947 36585 25013 38345
rect 25105 33585 25171 35345
rect 20440 32840 20452 32910
rect 20452 32840 25086 32910
rect 25086 32840 25090 32910
rect 29910 38690 30090 38910
rect -4290 27030 -4110 27250
rect -4290 25490 -4110 25710
rect 1540 30710 1552 30780
rect 1552 30710 6186 30780
rect 6186 30710 6200 30780
rect 1465 25285 1531 27045
rect 1623 28285 1689 30045
rect 1781 25285 1847 27045
rect 1939 28285 2005 30045
rect 2097 25285 2163 27045
rect 2255 28285 2321 30045
rect 2413 25285 2479 27045
rect 2571 28285 2637 30045
rect 2729 25285 2795 27045
rect 2887 28285 2953 30045
rect 3045 25285 3111 27045
rect 3203 28285 3269 30045
rect 3361 25285 3427 27045
rect 3519 28285 3585 30045
rect 3677 25285 3743 27045
rect 3835 28285 3901 30045
rect 3993 25285 4059 27045
rect 4151 28285 4217 30045
rect 4309 25285 4375 27045
rect 4467 28285 4533 30045
rect 4625 25285 4691 27045
rect 4783 28285 4849 30045
rect 4941 25285 5007 27045
rect 5099 28285 5165 30045
rect 5257 25285 5323 27045
rect 5415 28285 5481 30045
rect 5573 25285 5639 27045
rect 5731 28285 5797 30045
rect 5889 25285 5955 27045
rect 6047 28285 6113 30045
rect 6205 25285 6271 27045
rect 1540 24540 1552 24610
rect 1552 24540 6186 24610
rect 6186 24540 6190 24610
rect 7840 30710 7852 30780
rect 7852 30710 12486 30780
rect 12486 30710 12500 30780
rect 7765 25285 7831 27045
rect 7923 28285 7989 30045
rect 8081 25285 8147 27045
rect 8239 28285 8305 30045
rect 8397 25285 8463 27045
rect 8555 28285 8621 30045
rect 8713 25285 8779 27045
rect 8871 28285 8937 30045
rect 9029 25285 9095 27045
rect 9187 28285 9253 30045
rect 9345 25285 9411 27045
rect 9503 28285 9569 30045
rect 9661 25285 9727 27045
rect 9819 28285 9885 30045
rect 9977 25285 10043 27045
rect 10135 28285 10201 30045
rect 10293 25285 10359 27045
rect 10451 28285 10517 30045
rect 10609 25285 10675 27045
rect 10767 28285 10833 30045
rect 10925 25285 10991 27045
rect 11083 28285 11149 30045
rect 11241 25285 11307 27045
rect 11399 28285 11465 30045
rect 11557 25285 11623 27045
rect 11715 28285 11781 30045
rect 11873 25285 11939 27045
rect 12031 28285 12097 30045
rect 12189 25285 12255 27045
rect 12347 28285 12413 30045
rect 12505 25285 12571 27045
rect 7840 24540 7852 24610
rect 7852 24540 12486 24610
rect 12486 24540 12490 24610
rect 14140 30710 14152 30780
rect 14152 30710 18786 30780
rect 18786 30710 18800 30780
rect 14065 25285 14131 27045
rect 14223 28285 14289 30045
rect 14381 25285 14447 27045
rect 14539 28285 14605 30045
rect 14697 25285 14763 27045
rect 14855 28285 14921 30045
rect 15013 25285 15079 27045
rect 15171 28285 15237 30045
rect 15329 25285 15395 27045
rect 15487 28285 15553 30045
rect 15645 25285 15711 27045
rect 15803 28285 15869 30045
rect 15961 25285 16027 27045
rect 16119 28285 16185 30045
rect 16277 25285 16343 27045
rect 16435 28285 16501 30045
rect 16593 25285 16659 27045
rect 16751 28285 16817 30045
rect 16909 25285 16975 27045
rect 17067 28285 17133 30045
rect 17225 25285 17291 27045
rect 17383 28285 17449 30045
rect 17541 25285 17607 27045
rect 17699 28285 17765 30045
rect 17857 25285 17923 27045
rect 18015 28285 18081 30045
rect 18173 25285 18239 27045
rect 18331 28285 18397 30045
rect 18489 25285 18555 27045
rect 18647 28285 18713 30045
rect 18805 25285 18871 27045
rect 14140 24540 14152 24610
rect 14152 24540 18786 24610
rect 18786 24540 18790 24610
rect 20440 30710 20452 30780
rect 20452 30710 25086 30780
rect 25086 30710 25100 30780
rect 20365 25285 20431 27045
rect 20523 28285 20589 30045
rect 20681 25285 20747 27045
rect 20839 28285 20905 30045
rect 20997 25285 21063 27045
rect 21155 28285 21221 30045
rect 21313 25285 21379 27045
rect 21471 28285 21537 30045
rect 21629 25285 21695 27045
rect 21787 28285 21853 30045
rect 21945 25285 22011 27045
rect 22103 28285 22169 30045
rect 22261 25285 22327 27045
rect 22419 28285 22485 30045
rect 22577 25285 22643 27045
rect 22735 28285 22801 30045
rect 22893 25285 22959 27045
rect 23051 28285 23117 30045
rect 23209 25285 23275 27045
rect 23367 28285 23433 30045
rect 23525 25285 23591 27045
rect 23683 28285 23749 30045
rect 23841 25285 23907 27045
rect 23999 28285 24065 30045
rect 24157 25285 24223 27045
rect 24315 28285 24381 30045
rect 24473 25285 24539 27045
rect 24631 28285 24697 30045
rect 24789 25285 24855 27045
rect 24947 28285 25013 30045
rect 25105 25285 25171 27045
rect 20440 24540 20452 24610
rect 20452 24540 25086 24610
rect 25086 24540 25090 24610
rect 30910 27030 31090 27250
rect 30910 25490 31090 25710
rect 1540 23710 1552 23780
rect 1552 23710 6186 23780
rect 6186 23710 6200 23780
rect 1465 18285 1531 20045
rect 1623 21285 1689 23045
rect 1781 18285 1847 20045
rect 1939 21285 2005 23045
rect 2097 18285 2163 20045
rect 2255 21285 2321 23045
rect 2413 18285 2479 20045
rect 2571 21285 2637 23045
rect 2729 18285 2795 20045
rect 2887 21285 2953 23045
rect 3045 18285 3111 20045
rect 3203 21285 3269 23045
rect 3361 18285 3427 20045
rect 3519 21285 3585 23045
rect 3677 18285 3743 20045
rect 3835 21285 3901 23045
rect 3993 18285 4059 20045
rect 4151 21285 4217 23045
rect 4309 18285 4375 20045
rect 4467 21285 4533 23045
rect 4625 18285 4691 20045
rect 4783 21285 4849 23045
rect 4941 18285 5007 20045
rect 5099 21285 5165 23045
rect 5257 18285 5323 20045
rect 5415 21285 5481 23045
rect 5573 18285 5639 20045
rect 5731 21285 5797 23045
rect 5889 18285 5955 20045
rect 6047 21285 6113 23045
rect 6205 18285 6271 20045
rect 1540 17540 1552 17610
rect 1552 17540 6186 17610
rect 6186 17540 6190 17610
rect 7840 23710 7852 23780
rect 7852 23710 12486 23780
rect 12486 23710 12500 23780
rect 7765 18285 7831 20045
rect 7923 21285 7989 23045
rect 8081 18285 8147 20045
rect 8239 21285 8305 23045
rect 8397 18285 8463 20045
rect 8555 21285 8621 23045
rect 8713 18285 8779 20045
rect 8871 21285 8937 23045
rect 9029 18285 9095 20045
rect 9187 21285 9253 23045
rect 9345 18285 9411 20045
rect 9503 21285 9569 23045
rect 9661 18285 9727 20045
rect 9819 21285 9885 23045
rect 9977 18285 10043 20045
rect 10135 21285 10201 23045
rect 10293 18285 10359 20045
rect 10451 21285 10517 23045
rect 10609 18285 10675 20045
rect 10767 21285 10833 23045
rect 10925 18285 10991 20045
rect 11083 21285 11149 23045
rect 11241 18285 11307 20045
rect 11399 21285 11465 23045
rect 11557 18285 11623 20045
rect 11715 21285 11781 23045
rect 11873 18285 11939 20045
rect 12031 21285 12097 23045
rect 12189 18285 12255 20045
rect 12347 21285 12413 23045
rect 12505 18285 12571 20045
rect 7840 17540 7852 17610
rect 7852 17540 12486 17610
rect 12486 17540 12490 17610
rect 14140 23710 14152 23780
rect 14152 23710 18786 23780
rect 18786 23710 18800 23780
rect 14065 18285 14131 20045
rect 14223 21285 14289 23045
rect 14381 18285 14447 20045
rect 14539 21285 14605 23045
rect 14697 18285 14763 20045
rect 14855 21285 14921 23045
rect 15013 18285 15079 20045
rect 15171 21285 15237 23045
rect 15329 18285 15395 20045
rect 15487 21285 15553 23045
rect 15645 18285 15711 20045
rect 15803 21285 15869 23045
rect 15961 18285 16027 20045
rect 16119 21285 16185 23045
rect 16277 18285 16343 20045
rect 16435 21285 16501 23045
rect 16593 18285 16659 20045
rect 16751 21285 16817 23045
rect 16909 18285 16975 20045
rect 17067 21285 17133 23045
rect 17225 18285 17291 20045
rect 17383 21285 17449 23045
rect 17541 18285 17607 20045
rect 17699 21285 17765 23045
rect 17857 18285 17923 20045
rect 18015 21285 18081 23045
rect 18173 18285 18239 20045
rect 18331 21285 18397 23045
rect 18489 18285 18555 20045
rect 18647 21285 18713 23045
rect 18805 18285 18871 20045
rect 14140 17540 14152 17610
rect 14152 17540 18786 17610
rect 18786 17540 18790 17610
rect 20440 23710 20452 23780
rect 20452 23710 25086 23780
rect 25086 23710 25100 23780
rect 20365 18285 20431 20045
rect 20523 21285 20589 23045
rect 20681 18285 20747 20045
rect 20839 21285 20905 23045
rect 20997 18285 21063 20045
rect 21155 21285 21221 23045
rect 21313 18285 21379 20045
rect 21471 21285 21537 23045
rect 21629 18285 21695 20045
rect 21787 21285 21853 23045
rect 21945 18285 22011 20045
rect 22103 21285 22169 23045
rect 22261 18285 22327 20045
rect 22419 21285 22485 23045
rect 22577 18285 22643 20045
rect 22735 21285 22801 23045
rect 22893 18285 22959 20045
rect 23051 21285 23117 23045
rect 23209 18285 23275 20045
rect 23367 21285 23433 23045
rect 23525 18285 23591 20045
rect 23683 21285 23749 23045
rect 23841 18285 23907 20045
rect 23999 21285 24065 23045
rect 24157 18285 24223 20045
rect 24315 21285 24381 23045
rect 24473 18285 24539 20045
rect 24631 21285 24697 23045
rect 24789 18285 24855 20045
rect 24947 21285 25013 23045
rect 25105 18285 25171 20045
rect 20440 17540 20452 17610
rect 20452 17540 25086 17610
rect 25086 17540 25090 17610
rect -4290 13420 -4110 13900
rect -4290 12610 -4110 13090
rect 1540 15410 1552 15480
rect 1552 15410 6186 15480
rect 6186 15410 6200 15480
rect 1465 9985 1531 11745
rect 1623 12985 1689 14745
rect 1781 9985 1847 11745
rect 1939 12985 2005 14745
rect 2097 9985 2163 11745
rect 2255 12985 2321 14745
rect 2413 9985 2479 11745
rect 2571 12985 2637 14745
rect 2729 9985 2795 11745
rect 2887 12985 2953 14745
rect 3045 9985 3111 11745
rect 3203 12985 3269 14745
rect 3361 9985 3427 11745
rect 3519 12985 3585 14745
rect 3677 9985 3743 11745
rect 3835 12985 3901 14745
rect 3993 9985 4059 11745
rect 4151 12985 4217 14745
rect 4309 9985 4375 11745
rect 4467 12985 4533 14745
rect 4625 9985 4691 11745
rect 4783 12985 4849 14745
rect 4941 9985 5007 11745
rect 5099 12985 5165 14745
rect 5257 9985 5323 11745
rect 5415 12985 5481 14745
rect 5573 9985 5639 11745
rect 5731 12985 5797 14745
rect 5889 9985 5955 11745
rect 6047 12985 6113 14745
rect 6205 9985 6271 11745
rect 1540 9240 1552 9310
rect 1552 9240 6186 9310
rect 6186 9240 6190 9310
rect 7840 15410 7852 15480
rect 7852 15410 12486 15480
rect 12486 15410 12500 15480
rect 7765 9985 7831 11745
rect 7923 12985 7989 14745
rect 8081 9985 8147 11745
rect 8239 12985 8305 14745
rect 8397 9985 8463 11745
rect 8555 12985 8621 14745
rect 8713 9985 8779 11745
rect 8871 12985 8937 14745
rect 9029 9985 9095 11745
rect 9187 12985 9253 14745
rect 9345 9985 9411 11745
rect 9503 12985 9569 14745
rect 9661 9985 9727 11745
rect 9819 12985 9885 14745
rect 9977 9985 10043 11745
rect 10135 12985 10201 14745
rect 10293 9985 10359 11745
rect 10451 12985 10517 14745
rect 10609 9985 10675 11745
rect 10767 12985 10833 14745
rect 10925 9985 10991 11745
rect 11083 12985 11149 14745
rect 11241 9985 11307 11745
rect 11399 12985 11465 14745
rect 11557 9985 11623 11745
rect 11715 12985 11781 14745
rect 11873 9985 11939 11745
rect 12031 12985 12097 14745
rect 12189 9985 12255 11745
rect 12347 12985 12413 14745
rect 12505 9985 12571 11745
rect 7840 9240 7852 9310
rect 7852 9240 12486 9310
rect 12486 9240 12490 9310
rect 14140 15410 14152 15480
rect 14152 15410 18786 15480
rect 18786 15410 18800 15480
rect 14065 9985 14131 11745
rect 14223 12985 14289 14745
rect 14381 9985 14447 11745
rect 14539 12985 14605 14745
rect 14697 9985 14763 11745
rect 14855 12985 14921 14745
rect 15013 9985 15079 11745
rect 15171 12985 15237 14745
rect 15329 9985 15395 11745
rect 15487 12985 15553 14745
rect 15645 9985 15711 11745
rect 15803 12985 15869 14745
rect 15961 9985 16027 11745
rect 16119 12985 16185 14745
rect 16277 9985 16343 11745
rect 16435 12985 16501 14745
rect 16593 9985 16659 11745
rect 16751 12985 16817 14745
rect 16909 9985 16975 11745
rect 17067 12985 17133 14745
rect 17225 9985 17291 11745
rect 17383 12985 17449 14745
rect 17541 9985 17607 11745
rect 17699 12985 17765 14745
rect 17857 9985 17923 11745
rect 18015 12985 18081 14745
rect 18173 9985 18239 11745
rect 18331 12985 18397 14745
rect 18489 9985 18555 11745
rect 18647 12985 18713 14745
rect 18805 9985 18871 11745
rect 14140 9240 14152 9310
rect 14152 9240 18786 9310
rect 18786 9240 18790 9310
rect 20440 15410 20452 15480
rect 20452 15410 25086 15480
rect 25086 15410 25100 15480
rect 20365 9985 20431 11745
rect 20523 12985 20589 14745
rect 20681 9985 20747 11745
rect 20839 12985 20905 14745
rect 20997 9985 21063 11745
rect 21155 12985 21221 14745
rect 21313 9985 21379 11745
rect 21471 12985 21537 14745
rect 21629 9985 21695 11745
rect 21787 12985 21853 14745
rect 21945 9985 22011 11745
rect 22103 12985 22169 14745
rect 22261 9985 22327 11745
rect 22419 12985 22485 14745
rect 22577 9985 22643 11745
rect 22735 12985 22801 14745
rect 22893 9985 22959 11745
rect 23051 12985 23117 14745
rect 23209 9985 23275 11745
rect 23367 12985 23433 14745
rect 23525 9985 23591 11745
rect 23683 12985 23749 14745
rect 23841 9985 23907 11745
rect 23999 12985 24065 14745
rect 24157 9985 24223 11745
rect 24315 12985 24381 14745
rect 24473 9985 24539 11745
rect 24631 12985 24697 14745
rect 24789 9985 24855 11745
rect 24947 12985 25013 14745
rect 25105 9985 25171 11745
rect 20440 9240 20452 9310
rect 20452 9240 25086 9310
rect 25086 9240 25090 9310
rect 30910 13420 31090 13900
rect 30910 12610 31090 13090
rect 1540 8410 1552 8480
rect 1552 8410 6186 8480
rect 6186 8410 6200 8480
rect 1465 2985 1531 4745
rect 1623 5985 1689 7745
rect 1781 2985 1847 4745
rect 1939 5985 2005 7745
rect 2097 2985 2163 4745
rect 2255 5985 2321 7745
rect 2413 2985 2479 4745
rect 2571 5985 2637 7745
rect 2729 2985 2795 4745
rect 2887 5985 2953 7745
rect 3045 2985 3111 4745
rect 3203 5985 3269 7745
rect 3361 2985 3427 4745
rect 3519 5985 3585 7745
rect 3677 2985 3743 4745
rect 3835 5985 3901 7745
rect 3993 2985 4059 4745
rect 4151 5985 4217 7745
rect 4309 2985 4375 4745
rect 4467 5985 4533 7745
rect 4625 2985 4691 4745
rect 4783 5985 4849 7745
rect 4941 2985 5007 4745
rect 5099 5985 5165 7745
rect 5257 2985 5323 4745
rect 5415 5985 5481 7745
rect 5573 2985 5639 4745
rect 5731 5985 5797 7745
rect 5889 2985 5955 4745
rect 6047 5985 6113 7745
rect 6205 2985 6271 4745
rect 1540 2240 1552 2310
rect 1552 2240 6186 2310
rect 6186 2240 6190 2310
rect 7840 8410 7852 8480
rect 7852 8410 12486 8480
rect 12486 8410 12500 8480
rect 7765 2985 7831 4745
rect 7923 5985 7989 7745
rect 8081 2985 8147 4745
rect 8239 5985 8305 7745
rect 8397 2985 8463 4745
rect 8555 5985 8621 7745
rect 8713 2985 8779 4745
rect 8871 5985 8937 7745
rect 9029 2985 9095 4745
rect 9187 5985 9253 7745
rect 9345 2985 9411 4745
rect 9503 5985 9569 7745
rect 9661 2985 9727 4745
rect 9819 5985 9885 7745
rect 9977 2985 10043 4745
rect 10135 5985 10201 7745
rect 10293 2985 10359 4745
rect 10451 5985 10517 7745
rect 10609 2985 10675 4745
rect 10767 5985 10833 7745
rect 10925 2985 10991 4745
rect 11083 5985 11149 7745
rect 11241 2985 11307 4745
rect 11399 5985 11465 7745
rect 11557 2985 11623 4745
rect 11715 5985 11781 7745
rect 11873 2985 11939 4745
rect 12031 5985 12097 7745
rect 12189 2985 12255 4745
rect 12347 5985 12413 7745
rect 12505 2985 12571 4745
rect 7840 2240 7852 2310
rect 7852 2240 12486 2310
rect 12486 2240 12490 2310
rect 14140 8410 14152 8480
rect 14152 8410 18786 8480
rect 18786 8410 18800 8480
rect 14065 2985 14131 4745
rect 14223 5985 14289 7745
rect 14381 2985 14447 4745
rect 14539 5985 14605 7745
rect 14697 2985 14763 4745
rect 14855 5985 14921 7745
rect 15013 2985 15079 4745
rect 15171 5985 15237 7745
rect 15329 2985 15395 4745
rect 15487 5985 15553 7745
rect 15645 2985 15711 4745
rect 15803 5985 15869 7745
rect 15961 2985 16027 4745
rect 16119 5985 16185 7745
rect 16277 2985 16343 4745
rect 16435 5985 16501 7745
rect 16593 2985 16659 4745
rect 16751 5985 16817 7745
rect 16909 2985 16975 4745
rect 17067 5985 17133 7745
rect 17225 2985 17291 4745
rect 17383 5985 17449 7745
rect 17541 2985 17607 4745
rect 17699 5985 17765 7745
rect 17857 2985 17923 4745
rect 18015 5985 18081 7745
rect 18173 2985 18239 4745
rect 18331 5985 18397 7745
rect 18489 2985 18555 4745
rect 18647 5985 18713 7745
rect 18805 2985 18871 4745
rect 14140 2240 14152 2310
rect 14152 2240 18786 2310
rect 18786 2240 18790 2310
rect 20440 8410 20452 8480
rect 20452 8410 25086 8480
rect 25086 8410 25100 8480
rect 20365 2985 20431 4745
rect 20523 5985 20589 7745
rect 20681 2985 20747 4745
rect 20839 5985 20905 7745
rect 20997 2985 21063 4745
rect 21155 5985 21221 7745
rect 21313 2985 21379 4745
rect 21471 5985 21537 7745
rect 21629 2985 21695 4745
rect 21787 5985 21853 7745
rect 21945 2985 22011 4745
rect 22103 5985 22169 7745
rect 22261 2985 22327 4745
rect 22419 5985 22485 7745
rect 22577 2985 22643 4745
rect 22735 5985 22801 7745
rect 22893 2985 22959 4745
rect 23051 5985 23117 7745
rect 23209 2985 23275 4745
rect 23367 5985 23433 7745
rect 23525 2985 23591 4745
rect 23683 5985 23749 7745
rect 23841 2985 23907 4745
rect 23999 5985 24065 7745
rect 24157 2985 24223 4745
rect 24315 5985 24381 7745
rect 24473 2985 24539 4745
rect 24631 5985 24697 7745
rect 24789 2985 24855 4745
rect 24947 5985 25013 7745
rect 25105 2985 25171 4745
rect 20440 2240 20452 2310
rect 20452 2240 25086 2310
rect 25086 2240 25090 2310
<< metal3 >>
rect 1400 46080 6400 46200
rect 1400 46010 1540 46080
rect 6200 46010 6400 46080
rect 1400 46000 6400 46010
rect 7700 46080 12700 46200
rect 7700 46010 7840 46080
rect 12500 46010 12700 46080
rect 7700 46000 12700 46010
rect 14000 46080 19000 46200
rect 14000 46010 14140 46080
rect 18800 46010 19000 46080
rect 14000 46000 19000 46010
rect 20300 46080 25300 46200
rect 20300 46010 20440 46080
rect 25100 46010 25300 46080
rect 20300 46000 25300 46010
rect 1300 45400 6410 45500
rect 1300 43600 1400 45400
rect 2700 45345 6410 45400
rect 2700 43600 2887 45345
rect 1300 43585 1623 43600
rect 1689 43585 1939 43600
rect 2005 43585 2255 43600
rect 2321 43585 2571 43600
rect 2637 43585 2887 43600
rect 2953 43585 3203 45345
rect 3269 43585 3519 45345
rect 3585 43585 3835 45345
rect 3901 43585 4151 45345
rect 4217 43585 4467 45345
rect 4533 43585 4783 45345
rect 4849 43585 5099 45345
rect 5165 43585 5415 45345
rect 5481 43585 5731 45345
rect 5797 43585 6047 45345
rect 6113 43585 6410 45345
rect 1300 43500 6410 43585
rect 7600 45400 12710 45500
rect 7600 43600 7700 45400
rect 8900 45345 12710 45400
rect 7600 43585 7923 43600
rect 7989 43585 8239 43600
rect 8305 43585 8555 43600
rect 8621 43585 8871 43600
rect 8937 43585 9187 45345
rect 9253 43585 9503 45345
rect 9569 43585 9819 45345
rect 9885 43585 10135 45345
rect 10201 43585 10451 45345
rect 10517 43585 10767 45345
rect 10833 43585 11083 45345
rect 11149 43585 11399 45345
rect 11465 43585 11715 45345
rect 11781 43585 12031 45345
rect 12097 43585 12347 45345
rect 12413 43585 12710 45345
rect 7600 43500 12710 43585
rect 13900 45400 19010 45500
rect 13900 43600 14000 45400
rect 15300 45345 19010 45400
rect 15300 43600 15487 45345
rect 13900 43585 14223 43600
rect 14289 43585 14539 43600
rect 14605 43585 14855 43600
rect 14921 43585 15171 43600
rect 15237 43585 15487 43600
rect 15553 43585 15803 45345
rect 15869 43585 16119 45345
rect 16185 43585 16435 45345
rect 16501 43585 16751 45345
rect 16817 43585 17067 45345
rect 17133 43585 17383 45345
rect 17449 43585 17699 45345
rect 17765 43585 18015 45345
rect 18081 43585 18331 45345
rect 18397 43585 18647 45345
rect 18713 43585 19010 45345
rect 13900 43500 19010 43585
rect 20200 45400 25310 45500
rect 20200 43600 20300 45400
rect 21500 45345 25310 45400
rect 20200 43585 20523 43600
rect 20589 43585 20839 43600
rect 20905 43585 21155 43600
rect 21221 43585 21471 43600
rect 21537 43585 21787 45345
rect 21853 43585 22103 45345
rect 22169 43585 22419 45345
rect 22485 43585 22735 45345
rect 22801 43585 23051 45345
rect 23117 43585 23367 45345
rect 23433 43585 23683 45345
rect 23749 43585 23999 45345
rect 24065 43585 24315 45345
rect 24381 43585 24631 45345
rect 24697 43585 24947 45345
rect 25013 43585 25310 45345
rect 20200 43500 25310 43585
rect 1300 42400 6410 42500
rect 1300 40600 1400 42400
rect 2700 42345 6410 42400
rect 2700 40600 2729 42345
rect 1300 40585 1465 40600
rect 1531 40585 1781 40600
rect 1847 40585 2097 40600
rect 2163 40585 2413 40600
rect 2479 40585 2729 40600
rect 2795 40585 3045 42345
rect 3111 40585 3361 42345
rect 3427 40585 3677 42345
rect 3743 40585 3993 42345
rect 4059 40585 4309 42345
rect 4375 40585 4625 42345
rect 4691 40585 4941 42345
rect 5007 40585 5257 42345
rect 5323 40585 5573 42345
rect 5639 40585 5889 42345
rect 5955 40585 6205 42345
rect 6271 40585 6410 42345
rect 1300 40500 6410 40585
rect 7630 42400 12900 42500
rect 7630 42345 11500 42400
rect 7630 40585 7765 42345
rect 7831 40585 8081 42345
rect 8147 40585 8397 42345
rect 8463 40585 8713 42345
rect 8779 40585 9029 42345
rect 9095 40585 9345 42345
rect 9411 40585 9661 42345
rect 9727 40585 9977 42345
rect 10043 40585 10293 42345
rect 10359 40585 10609 42345
rect 10675 40585 10925 42345
rect 10991 40585 11241 42345
rect 11307 40600 11500 42345
rect 12800 40600 12900 42400
rect 11307 40585 11557 40600
rect 11623 40585 11873 40600
rect 11939 40585 12189 40600
rect 12255 40585 12505 40600
rect 12571 40585 12900 40600
rect 7630 40500 12900 40585
rect 13900 42400 19010 42500
rect 13900 40600 14000 42400
rect 15300 42345 19010 42400
rect 15300 40600 15329 42345
rect 13900 40585 14065 40600
rect 14131 40585 14381 40600
rect 14447 40585 14697 40600
rect 14763 40585 15013 40600
rect 15079 40585 15329 40600
rect 15395 40585 15645 42345
rect 15711 40585 15961 42345
rect 16027 40585 16277 42345
rect 16343 40585 16593 42345
rect 16659 40585 16909 42345
rect 16975 40585 17225 42345
rect 17291 40585 17541 42345
rect 17607 40585 17857 42345
rect 17923 40585 18173 42345
rect 18239 40585 18489 42345
rect 18555 40585 18805 42345
rect 18871 40585 19010 42345
rect 13900 40500 19010 40585
rect 20230 42400 25500 42500
rect 20230 42345 24100 42400
rect 20230 40585 20365 42345
rect 20431 40585 20681 42345
rect 20747 40585 20997 42345
rect 21063 40585 21313 42345
rect 21379 40585 21629 42345
rect 21695 40585 21945 42345
rect 22011 40585 22261 42345
rect 22327 40585 22577 42345
rect 22643 40585 22893 42345
rect 22959 40585 23209 42345
rect 23275 40585 23525 42345
rect 23591 40585 23841 42345
rect 23907 40600 24100 42345
rect 25400 40600 25500 42400
rect 23907 40585 24157 40600
rect 24223 40585 24473 40600
rect 24539 40585 24789 40600
rect 24855 40585 25105 40600
rect 25171 40585 25500 40600
rect 20230 40500 25500 40585
rect -3400 40480 -3000 40500
rect -3400 40410 -3380 40480
rect -3400 40190 -3390 40410
rect -3020 40410 -3000 40480
rect -3010 40190 -3000 40410
rect 29800 40480 30200 40500
rect 29800 40410 29820 40480
rect -3400 40180 -3000 40190
rect 3000 40100 4900 40200
rect 3000 40000 3200 40100
rect 1300 39910 3200 40000
rect 4700 40000 4900 40100
rect 15600 40100 17500 40200
rect 29800 40190 29810 40410
rect 30180 40410 30200 40480
rect 30190 40190 30200 40410
rect 29800 40180 30200 40190
rect 15600 40000 15800 40100
rect 4700 39910 7300 40000
rect 1300 39840 1540 39910
rect 6190 39880 7300 39910
rect 6190 39840 6920 39880
rect 1300 39800 3200 39840
rect 4700 39800 6920 39840
rect 1300 39720 6920 39800
rect 7280 39720 7300 39880
rect 1300 39700 7300 39720
rect 7500 39910 13600 40000
rect 7500 39840 7840 39910
rect 12490 39880 13600 39910
rect 12490 39840 13220 39880
rect 7500 39720 13220 39840
rect 13580 39720 13600 39880
rect 7500 39700 13600 39720
rect 13800 39910 15800 40000
rect 17300 40000 17500 40100
rect 17300 39910 19900 40000
rect 13800 39840 14140 39910
rect 18790 39880 19900 39910
rect 18790 39840 19520 39880
rect 13800 39800 15800 39840
rect 17300 39800 19520 39840
rect 13800 39720 19520 39800
rect 19880 39720 19900 39880
rect 13800 39700 19900 39720
rect 20100 39910 25300 40000
rect 20100 39840 20440 39910
rect 25090 39840 25300 39910
rect 20100 39700 25300 39840
rect 7500 39500 7800 39700
rect 9300 39600 11900 39700
rect 13800 39600 14000 39700
rect 20100 39600 20400 39700
rect 21900 39600 24500 39700
rect 6400 39300 7800 39500
rect 12700 39400 14000 39600
rect 19000 39400 20400 39600
rect 3000 39200 4900 39300
rect 6400 39200 6700 39300
rect 9300 39200 11900 39300
rect 12700 39200 13000 39400
rect 15600 39200 17500 39300
rect 19000 39200 19300 39400
rect 21900 39200 24500 39300
rect 1300 39080 3200 39200
rect 4700 39080 6700 39200
rect 1300 39010 1540 39080
rect 6200 39010 6700 39080
rect -3400 38910 -3000 38920
rect -3400 38690 -3390 38910
rect -3010 38690 -3000 38910
rect 1300 38900 3200 39010
rect 4700 38900 6700 39010
rect 6900 39180 13000 39200
rect 6900 39020 6920 39180
rect 7280 39080 13000 39180
rect 7280 39020 7840 39080
rect 6900 39010 7840 39020
rect 12500 39010 13000 39080
rect 6900 38900 13000 39010
rect 13200 39180 15800 39200
rect 13200 39020 13220 39180
rect 13580 39080 15800 39180
rect 17300 39080 19300 39200
rect 13580 39020 14140 39080
rect 13200 39010 14140 39020
rect 18800 39010 19300 39080
rect 13200 38900 15800 39010
rect 17300 38900 19300 39010
rect 19500 39180 25300 39200
rect 19500 39020 19520 39180
rect 19880 39080 25300 39180
rect 19880 39020 20440 39080
rect 19500 39010 20440 39020
rect 25100 39010 25300 39080
rect 19500 38900 25300 39010
rect 29800 38910 30200 38920
rect 3000 38800 4900 38900
rect 15600 38800 17500 38900
rect -3400 38680 -3000 38690
rect 29800 38690 29810 38910
rect 30190 38690 30200 38910
rect 29800 38680 30200 38690
rect 1330 38400 6410 38500
rect 1330 38345 3300 38400
rect 4600 38345 6410 38400
rect 1330 36585 1623 38345
rect 1689 36585 1939 38345
rect 2005 36585 2255 38345
rect 2321 36585 2571 38345
rect 2637 36585 2887 38345
rect 2953 36585 3203 38345
rect 3269 36600 3300 38345
rect 4600 36600 4783 38345
rect 3269 36585 3519 36600
rect 3585 36585 3835 36600
rect 3901 36585 4151 36600
rect 4217 36585 4467 36600
rect 4533 36585 4783 36600
rect 4849 36585 5099 38345
rect 5165 36585 5415 38345
rect 5481 36585 5731 38345
rect 5797 36585 6047 38345
rect 6113 36585 6410 38345
rect 1330 36500 6410 36585
rect 7600 38400 12710 38500
rect 7600 36600 7700 38400
rect 9000 38345 12710 38400
rect 9000 36600 9187 38345
rect 7600 36585 7923 36600
rect 7989 36585 8239 36600
rect 8305 36585 8555 36600
rect 8621 36585 8871 36600
rect 8937 36585 9187 36600
rect 9253 36585 9503 38345
rect 9569 36585 9819 38345
rect 9885 36585 10135 38345
rect 10201 36585 10451 38345
rect 10517 36585 10767 38345
rect 10833 36585 11083 38345
rect 11149 36585 11399 38345
rect 11465 36585 11715 38345
rect 11781 36585 12031 38345
rect 12097 36585 12347 38345
rect 12413 36585 12710 38345
rect 7600 36500 12710 36585
rect 13930 38400 19010 38500
rect 13930 38345 15900 38400
rect 17200 38345 19010 38400
rect 13930 36585 14223 38345
rect 14289 36585 14539 38345
rect 14605 36585 14855 38345
rect 14921 36585 15171 38345
rect 15237 36585 15487 38345
rect 15553 36585 15803 38345
rect 15869 36600 15900 38345
rect 17200 36600 17383 38345
rect 15869 36585 16119 36600
rect 16185 36585 16435 36600
rect 16501 36585 16751 36600
rect 16817 36585 17067 36600
rect 17133 36585 17383 36600
rect 17449 36585 17699 38345
rect 17765 36585 18015 38345
rect 18081 36585 18331 38345
rect 18397 36585 18647 38345
rect 18713 36585 19010 38345
rect 13930 36500 19010 36585
rect 20200 38400 25310 38500
rect 20200 36600 20300 38400
rect 21600 38345 25310 38400
rect 21600 36600 21787 38345
rect 20200 36585 20523 36600
rect 20589 36585 20839 36600
rect 20905 36585 21155 36600
rect 21221 36585 21471 36600
rect 21537 36585 21787 36600
rect 21853 36585 22103 38345
rect 22169 36585 22419 38345
rect 22485 36585 22735 38345
rect 22801 36585 23051 38345
rect 23117 36585 23367 38345
rect 23433 36585 23683 38345
rect 23749 36585 23999 38345
rect 24065 36585 24315 38345
rect 24381 36585 24631 38345
rect 24697 36585 24947 38345
rect 25013 36585 25310 38345
rect 20200 36500 25310 36585
rect 1330 35400 6600 35500
rect 1330 35345 5200 35400
rect 1330 33585 1465 35345
rect 1531 33585 1781 35345
rect 1847 33585 2097 35345
rect 2163 33585 2413 35345
rect 2479 33585 2729 35345
rect 2795 33585 3045 35345
rect 3111 33585 3361 35345
rect 3427 33585 3677 35345
rect 3743 33585 3993 35345
rect 4059 33585 4309 35345
rect 4375 33585 4625 35345
rect 4691 33585 4941 35345
rect 5007 33600 5200 35345
rect 6500 33600 6600 35400
rect 5007 33585 5257 33600
rect 5323 33585 5573 33600
rect 5639 33585 5889 33600
rect 5955 33585 6205 33600
rect 6271 33585 6600 33600
rect 1330 33500 6600 33585
rect 7630 35400 12710 35500
rect 7630 35345 9600 35400
rect 10900 35345 12710 35400
rect 7630 33585 7765 35345
rect 7831 33585 8081 35345
rect 8147 33585 8397 35345
rect 8463 33585 8713 35345
rect 8779 33585 9029 35345
rect 9095 33585 9345 35345
rect 9411 33600 9600 35345
rect 10900 33600 10925 35345
rect 9411 33585 9661 33600
rect 9727 33585 9977 33600
rect 10043 33585 10293 33600
rect 10359 33585 10609 33600
rect 10675 33585 10925 33600
rect 10991 33585 11241 35345
rect 11307 33585 11557 35345
rect 11623 33585 11873 35345
rect 11939 33585 12189 35345
rect 12255 33585 12505 35345
rect 12571 33585 12710 35345
rect 7630 33500 12710 33585
rect 13930 35400 19200 35500
rect 13930 35345 17800 35400
rect 13930 33585 14065 35345
rect 14131 33585 14381 35345
rect 14447 33585 14697 35345
rect 14763 33585 15013 35345
rect 15079 33585 15329 35345
rect 15395 33585 15645 35345
rect 15711 33585 15961 35345
rect 16027 33585 16277 35345
rect 16343 33585 16593 35345
rect 16659 33585 16909 35345
rect 16975 33585 17225 35345
rect 17291 33585 17541 35345
rect 17607 33600 17800 35345
rect 19100 33600 19200 35400
rect 17607 33585 17857 33600
rect 17923 33585 18173 33600
rect 18239 33585 18489 33600
rect 18555 33585 18805 33600
rect 18871 33585 19200 33600
rect 13930 33500 19200 33585
rect 20200 35400 25500 35500
rect 20200 35345 22200 35400
rect 23500 35345 25500 35400
rect 20200 33585 20365 35345
rect 20431 33585 20681 35345
rect 20747 33585 20997 35345
rect 21063 33585 21313 35345
rect 21379 33585 21629 35345
rect 21695 33585 21945 35345
rect 22011 33600 22200 35345
rect 23500 33600 23525 35345
rect 22011 33585 22261 33600
rect 22327 33585 22577 33600
rect 22643 33585 22893 33600
rect 22959 33585 23209 33600
rect 23275 33585 23525 33600
rect 23591 33585 23841 35345
rect 23907 33585 24157 35345
rect 24223 33585 24473 35345
rect 24539 33585 24789 35345
rect 24855 33585 25105 35345
rect 25171 33585 25500 35345
rect 20200 33500 25500 33585
rect 1400 32910 6400 32930
rect 1400 32840 1540 32910
rect 6190 32840 6400 32910
rect 1400 32730 6400 32840
rect 7700 32910 12700 32930
rect 7700 32840 7840 32910
rect 12490 32840 12700 32910
rect 7700 32730 12700 32840
rect 14000 32910 19000 32930
rect 14000 32840 14140 32910
rect 18790 32840 19000 32910
rect 14000 32730 19000 32840
rect 20300 32910 25300 32930
rect 20300 32840 20440 32910
rect 25090 32840 25300 32910
rect 20300 32730 25300 32840
rect -4400 31700 2800 31800
rect -4400 31100 1400 31700
rect 2700 31100 2800 31700
rect -4400 31000 2800 31100
rect 24000 31700 31200 31800
rect 24000 31100 24100 31700
rect 25400 31100 31200 31700
rect 24000 31000 31200 31100
rect -4400 27250 -3900 31000
rect 1400 30780 6400 30900
rect 1400 30710 1540 30780
rect 6200 30710 6400 30780
rect 1400 30700 6400 30710
rect 7700 30780 12700 30900
rect 7700 30710 7840 30780
rect 12500 30710 12700 30780
rect 7700 30700 12700 30710
rect 14000 30780 19000 30900
rect 14000 30710 14140 30780
rect 18800 30710 19000 30780
rect 14000 30700 19000 30710
rect 20300 30780 25300 30900
rect 20300 30710 20440 30780
rect 25100 30710 25300 30780
rect 20300 30700 25300 30710
rect 1300 30100 6410 30200
rect 1300 28300 1400 30100
rect 2700 30045 6410 30100
rect 2700 28300 2887 30045
rect 1300 28285 1623 28300
rect 1689 28285 1939 28300
rect 2005 28285 2255 28300
rect 2321 28285 2571 28300
rect 2637 28285 2887 28300
rect 2953 28285 3203 30045
rect 3269 28285 3519 30045
rect 3585 28285 3835 30045
rect 3901 28285 4151 30045
rect 4217 28285 4467 30045
rect 4533 28285 4783 30045
rect 4849 28285 5099 30045
rect 5165 28285 5415 30045
rect 5481 28285 5731 30045
rect 5797 28285 6047 30045
rect 6113 28285 6410 30045
rect 1300 28200 6410 28285
rect 7600 30100 12710 30200
rect 7600 28300 7700 30100
rect 8900 30045 12710 30100
rect 7600 28285 7923 28300
rect 7989 28285 8239 28300
rect 8305 28285 8555 28300
rect 8621 28285 8871 28300
rect 8937 28285 9187 30045
rect 9253 28285 9503 30045
rect 9569 28285 9819 30045
rect 9885 28285 10135 30045
rect 10201 28285 10451 30045
rect 10517 28285 10767 30045
rect 10833 28285 11083 30045
rect 11149 28285 11399 30045
rect 11465 28285 11715 30045
rect 11781 28285 12031 30045
rect 12097 28285 12347 30045
rect 12413 28285 12710 30045
rect 7600 28200 12710 28285
rect 13900 30100 19010 30200
rect 13900 28300 14000 30100
rect 15300 30045 19010 30100
rect 15300 28300 15487 30045
rect 13900 28285 14223 28300
rect 14289 28285 14539 28300
rect 14605 28285 14855 28300
rect 14921 28285 15171 28300
rect 15237 28285 15487 28300
rect 15553 28285 15803 30045
rect 15869 28285 16119 30045
rect 16185 28285 16435 30045
rect 16501 28285 16751 30045
rect 16817 28285 17067 30045
rect 17133 28285 17383 30045
rect 17449 28285 17699 30045
rect 17765 28285 18015 30045
rect 18081 28285 18331 30045
rect 18397 28285 18647 30045
rect 18713 28285 19010 30045
rect 13900 28200 19010 28285
rect 20200 30100 25310 30200
rect 20200 28300 20300 30100
rect 21500 30045 25310 30100
rect 20200 28285 20523 28300
rect 20589 28285 20839 28300
rect 20905 28285 21155 28300
rect 21221 28285 21471 28300
rect 21537 28285 21787 30045
rect 21853 28285 22103 30045
rect 22169 28285 22419 30045
rect 22485 28285 22735 30045
rect 22801 28285 23051 30045
rect 23117 28285 23367 30045
rect 23433 28285 23683 30045
rect 23749 28285 23999 30045
rect 24065 28285 24315 30045
rect 24381 28285 24631 30045
rect 24697 28285 24947 30045
rect 25013 28285 25310 30045
rect 20200 28200 25310 28285
rect -4400 27030 -4290 27250
rect -4110 27030 -3900 27250
rect 30700 27250 31200 31000
rect -4400 27000 -3900 27030
rect 1300 27100 6410 27200
rect -4400 25710 -4000 25720
rect -4400 25490 -4390 25710
rect -4010 25490 -4000 25710
rect -4400 25480 -4000 25490
rect 1300 25300 1400 27100
rect 2700 27045 6410 27100
rect 2700 25300 2729 27045
rect 1300 25285 1465 25300
rect 1531 25285 1781 25300
rect 1847 25285 2097 25300
rect 2163 25285 2413 25300
rect 2479 25285 2729 25300
rect 2795 25285 3045 27045
rect 3111 25285 3361 27045
rect 3427 25285 3677 27045
rect 3743 25285 3993 27045
rect 4059 25285 4309 27045
rect 4375 25285 4625 27045
rect 4691 25285 4941 27045
rect 5007 25285 5257 27045
rect 5323 25285 5573 27045
rect 5639 25285 5889 27045
rect 5955 25285 6205 27045
rect 6271 25285 6410 27045
rect 1300 25200 6410 25285
rect 7630 27100 12900 27200
rect 7630 27045 11500 27100
rect 7630 25285 7765 27045
rect 7831 25285 8081 27045
rect 8147 25285 8397 27045
rect 8463 25285 8713 27045
rect 8779 25285 9029 27045
rect 9095 25285 9345 27045
rect 9411 25285 9661 27045
rect 9727 25285 9977 27045
rect 10043 25285 10293 27045
rect 10359 25285 10609 27045
rect 10675 25285 10925 27045
rect 10991 25285 11241 27045
rect 11307 25300 11500 27045
rect 12800 25300 12900 27100
rect 11307 25285 11557 25300
rect 11623 25285 11873 25300
rect 11939 25285 12189 25300
rect 12255 25285 12505 25300
rect 12571 25285 12900 25300
rect 7630 25200 12900 25285
rect 13900 27100 19010 27200
rect 13900 25300 14000 27100
rect 15300 27045 19010 27100
rect 15300 25300 15329 27045
rect 13900 25285 14065 25300
rect 14131 25285 14381 25300
rect 14447 25285 14697 25300
rect 14763 25285 15013 25300
rect 15079 25285 15329 25300
rect 15395 25285 15645 27045
rect 15711 25285 15961 27045
rect 16027 25285 16277 27045
rect 16343 25285 16593 27045
rect 16659 25285 16909 27045
rect 16975 25285 17225 27045
rect 17291 25285 17541 27045
rect 17607 25285 17857 27045
rect 17923 25285 18173 27045
rect 18239 25285 18489 27045
rect 18555 25285 18805 27045
rect 18871 25285 19010 27045
rect 13900 25200 19010 25285
rect 20230 27100 25500 27200
rect 20230 27045 24100 27100
rect 20230 25285 20365 27045
rect 20431 25285 20681 27045
rect 20747 25285 20997 27045
rect 21063 25285 21313 27045
rect 21379 25285 21629 27045
rect 21695 25285 21945 27045
rect 22011 25285 22261 27045
rect 22327 25285 22577 27045
rect 22643 25285 22893 27045
rect 22959 25285 23209 27045
rect 23275 25285 23525 27045
rect 23591 25285 23841 27045
rect 23907 25300 24100 27045
rect 25400 25300 25500 27100
rect 30700 27030 30910 27250
rect 31090 27030 31200 27250
rect 30700 27000 31200 27030
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25480 31200 25490
rect 23907 25285 24157 25300
rect 24223 25285 24473 25300
rect 24539 25285 24789 25300
rect 24855 25285 25105 25300
rect 25171 25285 25500 25300
rect 20230 25200 25500 25285
rect 3000 24800 4900 24900
rect 3000 24700 3200 24800
rect 1300 24610 3200 24700
rect 4700 24700 4900 24800
rect 15600 24800 17500 24900
rect 15600 24700 15800 24800
rect 4700 24610 7300 24700
rect 1300 24540 1540 24610
rect 6190 24580 7300 24610
rect 6190 24540 6920 24580
rect 1300 24500 3200 24540
rect 4700 24500 6920 24540
rect 1300 24420 6920 24500
rect 7280 24420 7300 24580
rect 1300 24400 7300 24420
rect 7500 24610 13600 24700
rect 7500 24540 7840 24610
rect 12490 24580 13600 24610
rect 12490 24540 13220 24580
rect 7500 24420 13220 24540
rect 13580 24420 13600 24580
rect 7500 24400 13600 24420
rect 13800 24610 15800 24700
rect 17300 24700 17500 24800
rect 17300 24610 19900 24700
rect 13800 24540 14140 24610
rect 18790 24580 19900 24610
rect 18790 24540 19520 24580
rect 13800 24500 15800 24540
rect 17300 24500 19520 24540
rect 13800 24420 19520 24500
rect 19880 24420 19900 24580
rect 13800 24400 19900 24420
rect 20100 24610 25300 24700
rect 20100 24540 20440 24610
rect 25090 24540 25300 24610
rect 20100 24400 25300 24540
rect 7500 24200 7800 24400
rect 9300 24300 11900 24400
rect 13800 24300 14000 24400
rect 20100 24300 20400 24400
rect 21900 24300 24500 24400
rect 6400 24000 7800 24200
rect 12700 24100 14000 24300
rect 19000 24100 20400 24300
rect 3000 23900 4900 24000
rect 6400 23900 6700 24000
rect 9300 23900 11900 24000
rect 12700 23900 13000 24100
rect 15600 23900 17500 24000
rect 19000 23900 19300 24100
rect 21900 23900 24500 24000
rect 1300 23780 3200 23900
rect 4700 23780 6700 23900
rect 1300 23710 1540 23780
rect 6200 23710 6700 23780
rect 1300 23600 3200 23710
rect 4700 23600 6700 23710
rect 6900 23880 13000 23900
rect 6900 23720 6920 23880
rect 7280 23780 13000 23880
rect 7280 23720 7840 23780
rect 6900 23710 7840 23720
rect 12500 23710 13000 23780
rect 6900 23600 13000 23710
rect 13200 23880 15800 23900
rect 13200 23720 13220 23880
rect 13580 23780 15800 23880
rect 17300 23780 19300 23900
rect 13580 23720 14140 23780
rect 13200 23710 14140 23720
rect 18800 23710 19300 23780
rect 13200 23600 15800 23710
rect 17300 23600 19300 23710
rect 19500 23880 25300 23900
rect 19500 23720 19520 23880
rect 19880 23780 25300 23880
rect 19880 23720 20440 23780
rect 19500 23710 20440 23720
rect 25100 23710 25300 23780
rect 19500 23600 25300 23710
rect 3000 23500 4900 23600
rect 15600 23500 17500 23600
rect 1330 23100 6410 23200
rect 1330 23045 3300 23100
rect 4600 23045 6410 23100
rect 1330 21285 1623 23045
rect 1689 21285 1939 23045
rect 2005 21285 2255 23045
rect 2321 21285 2571 23045
rect 2637 21285 2887 23045
rect 2953 21285 3203 23045
rect 3269 21300 3300 23045
rect 4600 21300 4783 23045
rect 3269 21285 3519 21300
rect 3585 21285 3835 21300
rect 3901 21285 4151 21300
rect 4217 21285 4467 21300
rect 4533 21285 4783 21300
rect 4849 21285 5099 23045
rect 5165 21285 5415 23045
rect 5481 21285 5731 23045
rect 5797 21285 6047 23045
rect 6113 21285 6410 23045
rect 1330 21200 6410 21285
rect 7600 23100 12710 23200
rect 7600 21300 7700 23100
rect 9000 23045 12710 23100
rect 9000 21300 9187 23045
rect 7600 21285 7923 21300
rect 7989 21285 8239 21300
rect 8305 21285 8555 21300
rect 8621 21285 8871 21300
rect 8937 21285 9187 21300
rect 9253 21285 9503 23045
rect 9569 21285 9819 23045
rect 9885 21285 10135 23045
rect 10201 21285 10451 23045
rect 10517 21285 10767 23045
rect 10833 21285 11083 23045
rect 11149 21285 11399 23045
rect 11465 21285 11715 23045
rect 11781 21285 12031 23045
rect 12097 21285 12347 23045
rect 12413 21285 12710 23045
rect 7600 21200 12710 21285
rect 13930 23100 19010 23200
rect 13930 23045 15900 23100
rect 17200 23045 19010 23100
rect 13930 21285 14223 23045
rect 14289 21285 14539 23045
rect 14605 21285 14855 23045
rect 14921 21285 15171 23045
rect 15237 21285 15487 23045
rect 15553 21285 15803 23045
rect 15869 21300 15900 23045
rect 17200 21300 17383 23045
rect 15869 21285 16119 21300
rect 16185 21285 16435 21300
rect 16501 21285 16751 21300
rect 16817 21285 17067 21300
rect 17133 21285 17383 21300
rect 17449 21285 17699 23045
rect 17765 21285 18015 23045
rect 18081 21285 18331 23045
rect 18397 21285 18647 23045
rect 18713 21285 19010 23045
rect 13930 21200 19010 21285
rect 20200 23100 25310 23200
rect 20200 21300 20300 23100
rect 21600 23045 25310 23100
rect 21600 21300 21787 23045
rect 20200 21285 20523 21300
rect 20589 21285 20839 21300
rect 20905 21285 21155 21300
rect 21221 21285 21471 21300
rect 21537 21285 21787 21300
rect 21853 21285 22103 23045
rect 22169 21285 22419 23045
rect 22485 21285 22735 23045
rect 22801 21285 23051 23045
rect 23117 21285 23367 23045
rect 23433 21285 23683 23045
rect 23749 21285 23999 23045
rect 24065 21285 24315 23045
rect 24381 21285 24631 23045
rect 24697 21285 24947 23045
rect 25013 21285 25310 23045
rect 20200 21200 25310 21285
rect 1330 20100 6600 20200
rect 1330 20045 5200 20100
rect 1330 18285 1465 20045
rect 1531 18285 1781 20045
rect 1847 18285 2097 20045
rect 2163 18285 2413 20045
rect 2479 18285 2729 20045
rect 2795 18285 3045 20045
rect 3111 18285 3361 20045
rect 3427 18285 3677 20045
rect 3743 18285 3993 20045
rect 4059 18285 4309 20045
rect 4375 18285 4625 20045
rect 4691 18285 4941 20045
rect 5007 18300 5200 20045
rect 6500 18300 6600 20100
rect 5007 18285 5257 18300
rect 5323 18285 5573 18300
rect 5639 18285 5889 18300
rect 5955 18285 6205 18300
rect 6271 18285 6600 18300
rect 1330 18200 6600 18285
rect 7630 20100 12710 20200
rect 7630 20045 9600 20100
rect 10900 20045 12710 20100
rect 7630 18285 7765 20045
rect 7831 18285 8081 20045
rect 8147 18285 8397 20045
rect 8463 18285 8713 20045
rect 8779 18285 9029 20045
rect 9095 18285 9345 20045
rect 9411 18300 9600 20045
rect 10900 18300 10925 20045
rect 9411 18285 9661 18300
rect 9727 18285 9977 18300
rect 10043 18285 10293 18300
rect 10359 18285 10609 18300
rect 10675 18285 10925 18300
rect 10991 18285 11241 20045
rect 11307 18285 11557 20045
rect 11623 18285 11873 20045
rect 11939 18285 12189 20045
rect 12255 18285 12505 20045
rect 12571 18285 12710 20045
rect 7630 18200 12710 18285
rect 13930 20100 19200 20200
rect 13930 20045 17800 20100
rect 13930 18285 14065 20045
rect 14131 18285 14381 20045
rect 14447 18285 14697 20045
rect 14763 18285 15013 20045
rect 15079 18285 15329 20045
rect 15395 18285 15645 20045
rect 15711 18285 15961 20045
rect 16027 18285 16277 20045
rect 16343 18285 16593 20045
rect 16659 18285 16909 20045
rect 16975 18285 17225 20045
rect 17291 18285 17541 20045
rect 17607 18300 17800 20045
rect 19100 18300 19200 20100
rect 17607 18285 17857 18300
rect 17923 18285 18173 18300
rect 18239 18285 18489 18300
rect 18555 18285 18805 18300
rect 18871 18285 19200 18300
rect 13930 18200 19200 18285
rect 20200 20100 25500 20200
rect 20200 20045 22200 20100
rect 23500 20045 25500 20100
rect 20200 18285 20365 20045
rect 20431 18285 20681 20045
rect 20747 18285 20997 20045
rect 21063 18285 21313 20045
rect 21379 18285 21629 20045
rect 21695 18285 21945 20045
rect 22011 18300 22200 20045
rect 23500 18300 23525 20045
rect 22011 18285 22261 18300
rect 22327 18285 22577 18300
rect 22643 18285 22893 18300
rect 22959 18285 23209 18300
rect 23275 18285 23525 18300
rect 23591 18285 23841 20045
rect 23907 18285 24157 20045
rect 24223 18285 24473 20045
rect 24539 18285 24789 20045
rect 24855 18285 25105 20045
rect 25171 18285 25500 20045
rect 20200 18200 25500 18285
rect 1400 17610 6400 17630
rect 1400 17540 1540 17610
rect 6190 17540 6400 17610
rect 1400 17430 6400 17540
rect 7700 17610 12700 17630
rect 7700 17540 7840 17610
rect 12490 17540 12700 17610
rect 7700 17430 12700 17540
rect 14000 17610 19000 17630
rect 14000 17540 14140 17610
rect 18790 17540 19000 17610
rect 14000 17430 19000 17540
rect 20300 17610 25300 17630
rect 20300 17540 20440 17610
rect 25090 17540 25300 17610
rect 20300 17430 25300 17540
rect 1400 15480 6400 15600
rect 1400 15410 1540 15480
rect 6200 15410 6400 15480
rect 1400 15400 6400 15410
rect 7700 15480 12700 15600
rect 7700 15410 7840 15480
rect 12500 15410 12700 15480
rect 7700 15400 12700 15410
rect 14000 15480 19000 15600
rect 14000 15410 14140 15480
rect 18800 15410 19000 15480
rect 14000 15400 19000 15410
rect 20300 15480 25300 15600
rect 20300 15410 20440 15480
rect 25100 15410 25300 15480
rect 20300 15400 25300 15410
rect 1300 14800 6410 14900
rect -4400 14000 -4000 14010
rect -4400 13420 -4390 14000
rect -4010 13420 -4000 14000
rect -4400 13410 -4000 13420
rect -4400 13090 -4000 13100
rect -4400 12510 -4390 13090
rect -4010 12510 -4000 13090
rect 1300 13000 1400 14800
rect 2700 14745 6410 14800
rect 2700 13000 2887 14745
rect 1300 12985 1623 13000
rect 1689 12985 1939 13000
rect 2005 12985 2255 13000
rect 2321 12985 2571 13000
rect 2637 12985 2887 13000
rect 2953 12985 3203 14745
rect 3269 12985 3519 14745
rect 3585 12985 3835 14745
rect 3901 12985 4151 14745
rect 4217 12985 4467 14745
rect 4533 12985 4783 14745
rect 4849 12985 5099 14745
rect 5165 12985 5415 14745
rect 5481 12985 5731 14745
rect 5797 12985 6047 14745
rect 6113 12985 6410 14745
rect 1300 12900 6410 12985
rect 7600 14800 12710 14900
rect 7600 13000 7700 14800
rect 8900 14745 12710 14800
rect 7600 12985 7923 13000
rect 7989 12985 8239 13000
rect 8305 12985 8555 13000
rect 8621 12985 8871 13000
rect 8937 12985 9187 14745
rect 9253 12985 9503 14745
rect 9569 12985 9819 14745
rect 9885 12985 10135 14745
rect 10201 12985 10451 14745
rect 10517 12985 10767 14745
rect 10833 12985 11083 14745
rect 11149 12985 11399 14745
rect 11465 12985 11715 14745
rect 11781 12985 12031 14745
rect 12097 12985 12347 14745
rect 12413 12985 12710 14745
rect 7600 12900 12710 12985
rect 13900 14800 19010 14900
rect 13900 13000 14000 14800
rect 15300 14745 19010 14800
rect 15300 13000 15487 14745
rect 13900 12985 14223 13000
rect 14289 12985 14539 13000
rect 14605 12985 14855 13000
rect 14921 12985 15171 13000
rect 15237 12985 15487 13000
rect 15553 12985 15803 14745
rect 15869 12985 16119 14745
rect 16185 12985 16435 14745
rect 16501 12985 16751 14745
rect 16817 12985 17067 14745
rect 17133 12985 17383 14745
rect 17449 12985 17699 14745
rect 17765 12985 18015 14745
rect 18081 12985 18331 14745
rect 18397 12985 18647 14745
rect 18713 12985 19010 14745
rect 13900 12900 19010 12985
rect 20200 14800 25310 14900
rect 20200 13000 20300 14800
rect 21500 14745 25310 14800
rect 20200 12985 20523 13000
rect 20589 12985 20839 13000
rect 20905 12985 21155 13000
rect 21221 12985 21471 13000
rect 21537 12985 21787 14745
rect 21853 12985 22103 14745
rect 22169 12985 22419 14745
rect 22485 12985 22735 14745
rect 22801 12985 23051 14745
rect 23117 12985 23367 14745
rect 23433 12985 23683 14745
rect 23749 12985 23999 14745
rect 24065 12985 24315 14745
rect 24381 12985 24631 14745
rect 24697 12985 24947 14745
rect 25013 12985 25310 14745
rect 30800 14000 31200 14010
rect 30800 13420 30810 14000
rect 31190 13420 31200 14000
rect 30800 13410 31200 13420
rect 20200 12900 25310 12985
rect 30800 13090 31200 13100
rect -4400 12500 -4000 12510
rect 30800 12510 30810 13090
rect 31190 12510 31200 13090
rect 30800 12500 31200 12510
rect 1300 11800 6410 11900
rect 1300 10000 1400 11800
rect 2700 11745 6410 11800
rect 2700 10000 2729 11745
rect 1300 9985 1465 10000
rect 1531 9985 1781 10000
rect 1847 9985 2097 10000
rect 2163 9985 2413 10000
rect 2479 9985 2729 10000
rect 2795 9985 3045 11745
rect 3111 9985 3361 11745
rect 3427 9985 3677 11745
rect 3743 9985 3993 11745
rect 4059 9985 4309 11745
rect 4375 9985 4625 11745
rect 4691 9985 4941 11745
rect 5007 9985 5257 11745
rect 5323 9985 5573 11745
rect 5639 9985 5889 11745
rect 5955 9985 6205 11745
rect 6271 9985 6410 11745
rect 1300 9900 6410 9985
rect 7630 11800 12900 11900
rect 7630 11745 11500 11800
rect 7630 9985 7765 11745
rect 7831 9985 8081 11745
rect 8147 9985 8397 11745
rect 8463 9985 8713 11745
rect 8779 9985 9029 11745
rect 9095 9985 9345 11745
rect 9411 9985 9661 11745
rect 9727 9985 9977 11745
rect 10043 9985 10293 11745
rect 10359 9985 10609 11745
rect 10675 9985 10925 11745
rect 10991 9985 11241 11745
rect 11307 10000 11500 11745
rect 12800 10000 12900 11800
rect 11307 9985 11557 10000
rect 11623 9985 11873 10000
rect 11939 9985 12189 10000
rect 12255 9985 12505 10000
rect 12571 9985 12900 10000
rect 7630 9900 12900 9985
rect 13900 11800 19010 11900
rect 13900 10000 14000 11800
rect 15300 11745 19010 11800
rect 15300 10000 15329 11745
rect 13900 9985 14065 10000
rect 14131 9985 14381 10000
rect 14447 9985 14697 10000
rect 14763 9985 15013 10000
rect 15079 9985 15329 10000
rect 15395 9985 15645 11745
rect 15711 9985 15961 11745
rect 16027 9985 16277 11745
rect 16343 9985 16593 11745
rect 16659 9985 16909 11745
rect 16975 9985 17225 11745
rect 17291 9985 17541 11745
rect 17607 9985 17857 11745
rect 17923 9985 18173 11745
rect 18239 9985 18489 11745
rect 18555 9985 18805 11745
rect 18871 9985 19010 11745
rect 13900 9900 19010 9985
rect 20230 11800 25500 11900
rect 20230 11745 24100 11800
rect 20230 9985 20365 11745
rect 20431 9985 20681 11745
rect 20747 9985 20997 11745
rect 21063 9985 21313 11745
rect 21379 9985 21629 11745
rect 21695 9985 21945 11745
rect 22011 9985 22261 11745
rect 22327 9985 22577 11745
rect 22643 9985 22893 11745
rect 22959 9985 23209 11745
rect 23275 9985 23525 11745
rect 23591 9985 23841 11745
rect 23907 10000 24100 11745
rect 25400 10000 25500 11800
rect 23907 9985 24157 10000
rect 24223 9985 24473 10000
rect 24539 9985 24789 10000
rect 24855 9985 25105 10000
rect 25171 9985 25500 10000
rect 20230 9900 25500 9985
rect 3000 9500 4900 9600
rect 3000 9400 3200 9500
rect 1300 9310 3200 9400
rect 4700 9400 4900 9500
rect 15600 9500 17500 9600
rect 15600 9400 15800 9500
rect 4700 9310 7300 9400
rect 1300 9240 1540 9310
rect 6190 9280 7300 9310
rect 6190 9240 6920 9280
rect 1300 9200 3200 9240
rect 4700 9200 6920 9240
rect 1300 9120 6920 9200
rect 7280 9120 7300 9280
rect 1300 9100 7300 9120
rect 7500 9310 13600 9400
rect 7500 9240 7840 9310
rect 12490 9280 13600 9310
rect 12490 9240 13220 9280
rect 7500 9120 13220 9240
rect 13580 9120 13600 9280
rect 7500 9100 13600 9120
rect 13800 9310 15800 9400
rect 17300 9400 17500 9500
rect 17300 9310 19900 9400
rect 13800 9240 14140 9310
rect 18790 9280 19900 9310
rect 18790 9240 19520 9280
rect 13800 9200 15800 9240
rect 17300 9200 19520 9240
rect 13800 9120 19520 9200
rect 19880 9120 19900 9280
rect 13800 9100 19900 9120
rect 20100 9310 25300 9400
rect 20100 9240 20440 9310
rect 25090 9240 25300 9310
rect 20100 9100 25300 9240
rect 7500 8900 7800 9100
rect 9300 9000 11900 9100
rect 13800 9000 14000 9100
rect 20100 9000 20400 9100
rect 21900 9000 24500 9100
rect 6400 8700 7800 8900
rect 12700 8800 14000 9000
rect 19000 8800 20400 9000
rect 3000 8600 4900 8700
rect 6400 8600 6700 8700
rect 9300 8600 11900 8700
rect 12700 8600 13000 8800
rect 15600 8600 17500 8700
rect 19000 8600 19300 8800
rect 21900 8600 24500 8700
rect 1300 8480 3200 8600
rect 4700 8480 6700 8600
rect 1300 8410 1540 8480
rect 6200 8410 6700 8480
rect 1300 8300 3200 8410
rect 4700 8300 6700 8410
rect 6900 8580 13000 8600
rect 6900 8420 6920 8580
rect 7280 8480 13000 8580
rect 7280 8420 7840 8480
rect 6900 8410 7840 8420
rect 12500 8410 13000 8480
rect 6900 8300 13000 8410
rect 13200 8580 15800 8600
rect 13200 8420 13220 8580
rect 13580 8480 15800 8580
rect 17300 8480 19300 8600
rect 13580 8420 14140 8480
rect 13200 8410 14140 8420
rect 18800 8410 19300 8480
rect 13200 8300 15800 8410
rect 17300 8300 19300 8410
rect 19500 8580 25300 8600
rect 19500 8420 19520 8580
rect 19880 8480 25300 8580
rect 19880 8420 20440 8480
rect 19500 8410 20440 8420
rect 25100 8410 25300 8480
rect 19500 8300 25300 8410
rect 3000 8200 4900 8300
rect 15600 8200 17500 8300
rect 1330 7800 6410 7900
rect 1330 7745 3300 7800
rect 4600 7745 6410 7800
rect 1330 5985 1623 7745
rect 1689 5985 1939 7745
rect 2005 5985 2255 7745
rect 2321 5985 2571 7745
rect 2637 5985 2887 7745
rect 2953 5985 3203 7745
rect 3269 6000 3300 7745
rect 4600 6000 4783 7745
rect 3269 5985 3519 6000
rect 3585 5985 3835 6000
rect 3901 5985 4151 6000
rect 4217 5985 4467 6000
rect 4533 5985 4783 6000
rect 4849 5985 5099 7745
rect 5165 5985 5415 7745
rect 5481 5985 5731 7745
rect 5797 5985 6047 7745
rect 6113 5985 6410 7745
rect 1330 5900 6410 5985
rect 7600 7800 12710 7900
rect 7600 6000 7700 7800
rect 9000 7745 12710 7800
rect 9000 6000 9187 7745
rect 7600 5985 7923 6000
rect 7989 5985 8239 6000
rect 8305 5985 8555 6000
rect 8621 5985 8871 6000
rect 8937 5985 9187 6000
rect 9253 5985 9503 7745
rect 9569 5985 9819 7745
rect 9885 5985 10135 7745
rect 10201 5985 10451 7745
rect 10517 5985 10767 7745
rect 10833 5985 11083 7745
rect 11149 5985 11399 7745
rect 11465 5985 11715 7745
rect 11781 5985 12031 7745
rect 12097 5985 12347 7745
rect 12413 5985 12710 7745
rect 7600 5900 12710 5985
rect 13930 7800 19010 7900
rect 13930 7745 15900 7800
rect 17200 7745 19010 7800
rect 13930 5985 14223 7745
rect 14289 5985 14539 7745
rect 14605 5985 14855 7745
rect 14921 5985 15171 7745
rect 15237 5985 15487 7745
rect 15553 5985 15803 7745
rect 15869 6000 15900 7745
rect 17200 6000 17383 7745
rect 15869 5985 16119 6000
rect 16185 5985 16435 6000
rect 16501 5985 16751 6000
rect 16817 5985 17067 6000
rect 17133 5985 17383 6000
rect 17449 5985 17699 7745
rect 17765 5985 18015 7745
rect 18081 5985 18331 7745
rect 18397 5985 18647 7745
rect 18713 5985 19010 7745
rect 13930 5900 19010 5985
rect 20200 7800 25310 7900
rect 20200 6000 20300 7800
rect 21600 7745 25310 7800
rect 21600 6000 21787 7745
rect 20200 5985 20523 6000
rect 20589 5985 20839 6000
rect 20905 5985 21155 6000
rect 21221 5985 21471 6000
rect 21537 5985 21787 6000
rect 21853 5985 22103 7745
rect 22169 5985 22419 7745
rect 22485 5985 22735 7745
rect 22801 5985 23051 7745
rect 23117 5985 23367 7745
rect 23433 5985 23683 7745
rect 23749 5985 23999 7745
rect 24065 5985 24315 7745
rect 24381 5985 24631 7745
rect 24697 5985 24947 7745
rect 25013 5985 25310 7745
rect 20200 5900 25310 5985
rect 1330 4800 6600 4900
rect 1330 4745 5200 4800
rect 1330 2985 1465 4745
rect 1531 2985 1781 4745
rect 1847 2985 2097 4745
rect 2163 2985 2413 4745
rect 2479 2985 2729 4745
rect 2795 2985 3045 4745
rect 3111 2985 3361 4745
rect 3427 2985 3677 4745
rect 3743 2985 3993 4745
rect 4059 2985 4309 4745
rect 4375 2985 4625 4745
rect 4691 2985 4941 4745
rect 5007 3000 5200 4745
rect 6500 3000 6600 4800
rect 5007 2985 5257 3000
rect 5323 2985 5573 3000
rect 5639 2985 5889 3000
rect 5955 2985 6205 3000
rect 6271 2985 6600 3000
rect 1330 2900 6600 2985
rect 7630 4800 12710 4900
rect 7630 4745 9600 4800
rect 10900 4745 12710 4800
rect 7630 2985 7765 4745
rect 7831 2985 8081 4745
rect 8147 2985 8397 4745
rect 8463 2985 8713 4745
rect 8779 2985 9029 4745
rect 9095 2985 9345 4745
rect 9411 3000 9600 4745
rect 10900 3000 10925 4745
rect 9411 2985 9661 3000
rect 9727 2985 9977 3000
rect 10043 2985 10293 3000
rect 10359 2985 10609 3000
rect 10675 2985 10925 3000
rect 10991 2985 11241 4745
rect 11307 2985 11557 4745
rect 11623 2985 11873 4745
rect 11939 2985 12189 4745
rect 12255 2985 12505 4745
rect 12571 2985 12710 4745
rect 7630 2900 12710 2985
rect 13930 4800 19200 4900
rect 13930 4745 17800 4800
rect 13930 2985 14065 4745
rect 14131 2985 14381 4745
rect 14447 2985 14697 4745
rect 14763 2985 15013 4745
rect 15079 2985 15329 4745
rect 15395 2985 15645 4745
rect 15711 2985 15961 4745
rect 16027 2985 16277 4745
rect 16343 2985 16593 4745
rect 16659 2985 16909 4745
rect 16975 2985 17225 4745
rect 17291 2985 17541 4745
rect 17607 3000 17800 4745
rect 19100 3000 19200 4800
rect 17607 2985 17857 3000
rect 17923 2985 18173 3000
rect 18239 2985 18489 3000
rect 18555 2985 18805 3000
rect 18871 2985 19200 3000
rect 13930 2900 19200 2985
rect 20200 4800 25500 4900
rect 20200 4745 22200 4800
rect 23500 4745 25500 4800
rect 20200 2985 20365 4745
rect 20431 2985 20681 4745
rect 20747 2985 20997 4745
rect 21063 2985 21313 4745
rect 21379 2985 21629 4745
rect 21695 2985 21945 4745
rect 22011 3000 22200 4745
rect 23500 3000 23525 4745
rect 22011 2985 22261 3000
rect 22327 2985 22577 3000
rect 22643 2985 22893 3000
rect 22959 2985 23209 3000
rect 23275 2985 23525 3000
rect 23591 2985 23841 4745
rect 23907 2985 24157 4745
rect 24223 2985 24473 4745
rect 24539 2985 24789 4745
rect 24855 2985 25105 4745
rect 25171 2985 25500 4745
rect 20200 2900 25500 2985
rect 1400 2310 6400 2330
rect 1400 2240 1540 2310
rect 6190 2240 6400 2310
rect 1400 2130 6400 2240
rect 7700 2310 12700 2330
rect 7700 2240 7840 2310
rect 12490 2240 12700 2310
rect 7700 2130 12700 2240
rect 14000 2310 19000 2330
rect 14000 2240 14140 2310
rect 18790 2240 19000 2310
rect 14000 2130 19000 2240
rect 20300 2310 25300 2330
rect 20300 2240 20440 2310
rect 25090 2240 25300 2310
rect 20300 2130 25300 2240
<< via3 >>
rect 1400 45345 2700 45400
rect 1400 43600 1623 45345
rect 1623 43600 1689 45345
rect 1689 43600 1939 45345
rect 1939 43600 2005 45345
rect 2005 43600 2255 45345
rect 2255 43600 2321 45345
rect 2321 43600 2571 45345
rect 2571 43600 2637 45345
rect 2637 43600 2700 45345
rect 7700 45345 8900 45400
rect 7700 43600 7923 45345
rect 7923 43600 7989 45345
rect 7989 43600 8239 45345
rect 8239 43600 8305 45345
rect 8305 43600 8555 45345
rect 8555 43600 8621 45345
rect 8621 43600 8871 45345
rect 8871 43600 8900 45345
rect 14000 45345 15300 45400
rect 14000 43600 14223 45345
rect 14223 43600 14289 45345
rect 14289 43600 14539 45345
rect 14539 43600 14605 45345
rect 14605 43600 14855 45345
rect 14855 43600 14921 45345
rect 14921 43600 15171 45345
rect 15171 43600 15237 45345
rect 15237 43600 15300 45345
rect 20300 45345 21500 45400
rect 20300 43600 20523 45345
rect 20523 43600 20589 45345
rect 20589 43600 20839 45345
rect 20839 43600 20905 45345
rect 20905 43600 21155 45345
rect 21155 43600 21221 45345
rect 21221 43600 21471 45345
rect 21471 43600 21500 45345
rect 1400 42345 2700 42400
rect 1400 40600 1465 42345
rect 1465 40600 1531 42345
rect 1531 40600 1781 42345
rect 1781 40600 1847 42345
rect 1847 40600 2097 42345
rect 2097 40600 2163 42345
rect 2163 40600 2413 42345
rect 2413 40600 2479 42345
rect 2479 40600 2700 42345
rect 11500 42345 12800 42400
rect 11500 40600 11557 42345
rect 11557 40600 11623 42345
rect 11623 40600 11873 42345
rect 11873 40600 11939 42345
rect 11939 40600 12189 42345
rect 12189 40600 12255 42345
rect 12255 40600 12505 42345
rect 12505 40600 12571 42345
rect 12571 40600 12800 42345
rect 14000 42345 15300 42400
rect 14000 40600 14065 42345
rect 14065 40600 14131 42345
rect 14131 40600 14381 42345
rect 14381 40600 14447 42345
rect 14447 40600 14697 42345
rect 14697 40600 14763 42345
rect 14763 40600 15013 42345
rect 15013 40600 15079 42345
rect 15079 40600 15300 42345
rect 24100 42345 25400 42400
rect 24100 40600 24157 42345
rect 24157 40600 24223 42345
rect 24223 40600 24473 42345
rect 24473 40600 24539 42345
rect 24539 40600 24789 42345
rect 24789 40600 24855 42345
rect 24855 40600 25105 42345
rect 25105 40600 25171 42345
rect 25171 40600 25400 42345
rect -3380 40450 -3020 40480
rect -3380 40410 -3290 40450
rect -3390 40190 -3290 40410
rect -3290 40190 -3110 40450
rect -3110 40410 -3020 40450
rect -3110 40190 -3010 40410
rect 29820 40450 30180 40480
rect 29820 40410 29910 40450
rect 3200 39910 4700 40100
rect 29810 40190 29910 40410
rect 29910 40190 30090 40450
rect 30090 40410 30180 40450
rect 30090 40190 30190 40410
rect 3200 39840 4700 39910
rect 3200 39800 4700 39840
rect 6920 39720 7280 39880
rect 13220 39720 13580 39880
rect 15800 39910 17300 40100
rect 15800 39840 17300 39910
rect 15800 39800 17300 39840
rect 19520 39720 19880 39880
rect 3200 39080 4700 39200
rect 3200 39010 4700 39080
rect -3390 38690 -3290 38910
rect -3290 38690 -3110 38910
rect -3110 38690 -3010 38910
rect 3200 38900 4700 39010
rect 6920 39020 7280 39180
rect 13220 39020 13580 39180
rect 15800 39080 17300 39200
rect 15800 39010 17300 39080
rect 15800 38900 17300 39010
rect 19520 39020 19880 39180
rect 29810 38690 29910 38910
rect 29910 38690 30090 38910
rect 30090 38690 30190 38910
rect 3300 38345 4600 38400
rect 3300 36600 3519 38345
rect 3519 36600 3585 38345
rect 3585 36600 3835 38345
rect 3835 36600 3901 38345
rect 3901 36600 4151 38345
rect 4151 36600 4217 38345
rect 4217 36600 4467 38345
rect 4467 36600 4533 38345
rect 4533 36600 4600 38345
rect 7700 38345 9000 38400
rect 7700 36600 7923 38345
rect 7923 36600 7989 38345
rect 7989 36600 8239 38345
rect 8239 36600 8305 38345
rect 8305 36600 8555 38345
rect 8555 36600 8621 38345
rect 8621 36600 8871 38345
rect 8871 36600 8937 38345
rect 8937 36600 9000 38345
rect 15900 38345 17200 38400
rect 15900 36600 16119 38345
rect 16119 36600 16185 38345
rect 16185 36600 16435 38345
rect 16435 36600 16501 38345
rect 16501 36600 16751 38345
rect 16751 36600 16817 38345
rect 16817 36600 17067 38345
rect 17067 36600 17133 38345
rect 17133 36600 17200 38345
rect 20300 38345 21600 38400
rect 20300 36600 20523 38345
rect 20523 36600 20589 38345
rect 20589 36600 20839 38345
rect 20839 36600 20905 38345
rect 20905 36600 21155 38345
rect 21155 36600 21221 38345
rect 21221 36600 21471 38345
rect 21471 36600 21537 38345
rect 21537 36600 21600 38345
rect 5200 35345 6500 35400
rect 5200 33600 5257 35345
rect 5257 33600 5323 35345
rect 5323 33600 5573 35345
rect 5573 33600 5639 35345
rect 5639 33600 5889 35345
rect 5889 33600 5955 35345
rect 5955 33600 6205 35345
rect 6205 33600 6271 35345
rect 6271 33600 6500 35345
rect 9600 35345 10900 35400
rect 9600 33600 9661 35345
rect 9661 33600 9727 35345
rect 9727 33600 9977 35345
rect 9977 33600 10043 35345
rect 10043 33600 10293 35345
rect 10293 33600 10359 35345
rect 10359 33600 10609 35345
rect 10609 33600 10675 35345
rect 10675 33600 10900 35345
rect 17800 35345 19100 35400
rect 17800 33600 17857 35345
rect 17857 33600 17923 35345
rect 17923 33600 18173 35345
rect 18173 33600 18239 35345
rect 18239 33600 18489 35345
rect 18489 33600 18555 35345
rect 18555 33600 18805 35345
rect 18805 33600 18871 35345
rect 18871 33600 19100 35345
rect 22200 35345 23500 35400
rect 22200 33600 22261 35345
rect 22261 33600 22327 35345
rect 22327 33600 22577 35345
rect 22577 33600 22643 35345
rect 22643 33600 22893 35345
rect 22893 33600 22959 35345
rect 22959 33600 23209 35345
rect 23209 33600 23275 35345
rect 23275 33600 23500 35345
rect 1400 31100 2700 31700
rect 24100 31100 25400 31700
rect 1400 30045 2700 30100
rect 1400 28300 1623 30045
rect 1623 28300 1689 30045
rect 1689 28300 1939 30045
rect 1939 28300 2005 30045
rect 2005 28300 2255 30045
rect 2255 28300 2321 30045
rect 2321 28300 2571 30045
rect 2571 28300 2637 30045
rect 2637 28300 2700 30045
rect 7700 30045 8900 30100
rect 7700 28300 7923 30045
rect 7923 28300 7989 30045
rect 7989 28300 8239 30045
rect 8239 28300 8305 30045
rect 8305 28300 8555 30045
rect 8555 28300 8621 30045
rect 8621 28300 8871 30045
rect 8871 28300 8900 30045
rect 14000 30045 15300 30100
rect 14000 28300 14223 30045
rect 14223 28300 14289 30045
rect 14289 28300 14539 30045
rect 14539 28300 14605 30045
rect 14605 28300 14855 30045
rect 14855 28300 14921 30045
rect 14921 28300 15171 30045
rect 15171 28300 15237 30045
rect 15237 28300 15300 30045
rect 20300 30045 21500 30100
rect 20300 28300 20523 30045
rect 20523 28300 20589 30045
rect 20589 28300 20839 30045
rect 20839 28300 20905 30045
rect 20905 28300 21155 30045
rect 21155 28300 21221 30045
rect 21221 28300 21471 30045
rect 21471 28300 21500 30045
rect -4390 25490 -4290 25710
rect -4290 25490 -4110 25710
rect -4110 25490 -4010 25710
rect 1400 27045 2700 27100
rect 1400 25300 1465 27045
rect 1465 25300 1531 27045
rect 1531 25300 1781 27045
rect 1781 25300 1847 27045
rect 1847 25300 2097 27045
rect 2097 25300 2163 27045
rect 2163 25300 2413 27045
rect 2413 25300 2479 27045
rect 2479 25300 2700 27045
rect 11500 27045 12800 27100
rect 11500 25300 11557 27045
rect 11557 25300 11623 27045
rect 11623 25300 11873 27045
rect 11873 25300 11939 27045
rect 11939 25300 12189 27045
rect 12189 25300 12255 27045
rect 12255 25300 12505 27045
rect 12505 25300 12571 27045
rect 12571 25300 12800 27045
rect 14000 27045 15300 27100
rect 14000 25300 14065 27045
rect 14065 25300 14131 27045
rect 14131 25300 14381 27045
rect 14381 25300 14447 27045
rect 14447 25300 14697 27045
rect 14697 25300 14763 27045
rect 14763 25300 15013 27045
rect 15013 25300 15079 27045
rect 15079 25300 15300 27045
rect 24100 27045 25400 27100
rect 24100 25300 24157 27045
rect 24157 25300 24223 27045
rect 24223 25300 24473 27045
rect 24473 25300 24539 27045
rect 24539 25300 24789 27045
rect 24789 25300 24855 27045
rect 24855 25300 25105 27045
rect 25105 25300 25171 27045
rect 25171 25300 25400 27045
rect 30810 25490 30910 25710
rect 30910 25490 31090 25710
rect 31090 25490 31190 25710
rect 3200 24610 4700 24800
rect 3200 24540 4700 24610
rect 3200 24500 4700 24540
rect 6920 24420 7280 24580
rect 13220 24420 13580 24580
rect 15800 24610 17300 24800
rect 15800 24540 17300 24610
rect 15800 24500 17300 24540
rect 19520 24420 19880 24580
rect 3200 23780 4700 23900
rect 3200 23710 4700 23780
rect 3200 23600 4700 23710
rect 6920 23720 7280 23880
rect 13220 23720 13580 23880
rect 15800 23780 17300 23900
rect 15800 23710 17300 23780
rect 15800 23600 17300 23710
rect 19520 23720 19880 23880
rect 3300 23045 4600 23100
rect 3300 21300 3519 23045
rect 3519 21300 3585 23045
rect 3585 21300 3835 23045
rect 3835 21300 3901 23045
rect 3901 21300 4151 23045
rect 4151 21300 4217 23045
rect 4217 21300 4467 23045
rect 4467 21300 4533 23045
rect 4533 21300 4600 23045
rect 7700 23045 9000 23100
rect 7700 21300 7923 23045
rect 7923 21300 7989 23045
rect 7989 21300 8239 23045
rect 8239 21300 8305 23045
rect 8305 21300 8555 23045
rect 8555 21300 8621 23045
rect 8621 21300 8871 23045
rect 8871 21300 8937 23045
rect 8937 21300 9000 23045
rect 15900 23045 17200 23100
rect 15900 21300 16119 23045
rect 16119 21300 16185 23045
rect 16185 21300 16435 23045
rect 16435 21300 16501 23045
rect 16501 21300 16751 23045
rect 16751 21300 16817 23045
rect 16817 21300 17067 23045
rect 17067 21300 17133 23045
rect 17133 21300 17200 23045
rect 20300 23045 21600 23100
rect 20300 21300 20523 23045
rect 20523 21300 20589 23045
rect 20589 21300 20839 23045
rect 20839 21300 20905 23045
rect 20905 21300 21155 23045
rect 21155 21300 21221 23045
rect 21221 21300 21471 23045
rect 21471 21300 21537 23045
rect 21537 21300 21600 23045
rect 5200 20045 6500 20100
rect 5200 18300 5257 20045
rect 5257 18300 5323 20045
rect 5323 18300 5573 20045
rect 5573 18300 5639 20045
rect 5639 18300 5889 20045
rect 5889 18300 5955 20045
rect 5955 18300 6205 20045
rect 6205 18300 6271 20045
rect 6271 18300 6500 20045
rect 9600 20045 10900 20100
rect 9600 18300 9661 20045
rect 9661 18300 9727 20045
rect 9727 18300 9977 20045
rect 9977 18300 10043 20045
rect 10043 18300 10293 20045
rect 10293 18300 10359 20045
rect 10359 18300 10609 20045
rect 10609 18300 10675 20045
rect 10675 18300 10900 20045
rect 17800 20045 19100 20100
rect 17800 18300 17857 20045
rect 17857 18300 17923 20045
rect 17923 18300 18173 20045
rect 18173 18300 18239 20045
rect 18239 18300 18489 20045
rect 18489 18300 18555 20045
rect 18555 18300 18805 20045
rect 18805 18300 18871 20045
rect 18871 18300 19100 20045
rect 22200 20045 23500 20100
rect 22200 18300 22261 20045
rect 22261 18300 22327 20045
rect 22327 18300 22577 20045
rect 22577 18300 22643 20045
rect 22643 18300 22893 20045
rect 22893 18300 22959 20045
rect 22959 18300 23209 20045
rect 23209 18300 23275 20045
rect 23275 18300 23500 20045
rect -4390 13900 -4010 14000
rect -4390 13420 -4290 13900
rect -4290 13420 -4110 13900
rect -4110 13420 -4010 13900
rect -4390 12610 -4290 13090
rect -4290 12610 -4110 13090
rect -4110 12610 -4010 13090
rect -4390 12510 -4010 12610
rect 1400 14745 2700 14800
rect 1400 13000 1623 14745
rect 1623 13000 1689 14745
rect 1689 13000 1939 14745
rect 1939 13000 2005 14745
rect 2005 13000 2255 14745
rect 2255 13000 2321 14745
rect 2321 13000 2571 14745
rect 2571 13000 2637 14745
rect 2637 13000 2700 14745
rect 7700 14745 8900 14800
rect 7700 13000 7923 14745
rect 7923 13000 7989 14745
rect 7989 13000 8239 14745
rect 8239 13000 8305 14745
rect 8305 13000 8555 14745
rect 8555 13000 8621 14745
rect 8621 13000 8871 14745
rect 8871 13000 8900 14745
rect 14000 14745 15300 14800
rect 14000 13000 14223 14745
rect 14223 13000 14289 14745
rect 14289 13000 14539 14745
rect 14539 13000 14605 14745
rect 14605 13000 14855 14745
rect 14855 13000 14921 14745
rect 14921 13000 15171 14745
rect 15171 13000 15237 14745
rect 15237 13000 15300 14745
rect 20300 14745 21500 14800
rect 20300 13000 20523 14745
rect 20523 13000 20589 14745
rect 20589 13000 20839 14745
rect 20839 13000 20905 14745
rect 20905 13000 21155 14745
rect 21155 13000 21221 14745
rect 21221 13000 21471 14745
rect 21471 13000 21500 14745
rect 30810 13900 31190 14000
rect 30810 13420 30910 13900
rect 30910 13420 31090 13900
rect 31090 13420 31190 13900
rect 30810 12610 30910 13090
rect 30910 12610 31090 13090
rect 31090 12610 31190 13090
rect 30810 12510 31190 12610
rect 1400 11745 2700 11800
rect 1400 10000 1465 11745
rect 1465 10000 1531 11745
rect 1531 10000 1781 11745
rect 1781 10000 1847 11745
rect 1847 10000 2097 11745
rect 2097 10000 2163 11745
rect 2163 10000 2413 11745
rect 2413 10000 2479 11745
rect 2479 10000 2700 11745
rect 11500 11745 12800 11800
rect 11500 10000 11557 11745
rect 11557 10000 11623 11745
rect 11623 10000 11873 11745
rect 11873 10000 11939 11745
rect 11939 10000 12189 11745
rect 12189 10000 12255 11745
rect 12255 10000 12505 11745
rect 12505 10000 12571 11745
rect 12571 10000 12800 11745
rect 14000 11745 15300 11800
rect 14000 10000 14065 11745
rect 14065 10000 14131 11745
rect 14131 10000 14381 11745
rect 14381 10000 14447 11745
rect 14447 10000 14697 11745
rect 14697 10000 14763 11745
rect 14763 10000 15013 11745
rect 15013 10000 15079 11745
rect 15079 10000 15300 11745
rect 24100 11745 25400 11800
rect 24100 10000 24157 11745
rect 24157 10000 24223 11745
rect 24223 10000 24473 11745
rect 24473 10000 24539 11745
rect 24539 10000 24789 11745
rect 24789 10000 24855 11745
rect 24855 10000 25105 11745
rect 25105 10000 25171 11745
rect 25171 10000 25400 11745
rect 3200 9310 4700 9500
rect 3200 9240 4700 9310
rect 3200 9200 4700 9240
rect 6920 9120 7280 9280
rect 13220 9120 13580 9280
rect 15800 9310 17300 9500
rect 15800 9240 17300 9310
rect 15800 9200 17300 9240
rect 19520 9120 19880 9280
rect 3200 8480 4700 8600
rect 3200 8410 4700 8480
rect 3200 8300 4700 8410
rect 6920 8420 7280 8580
rect 13220 8420 13580 8580
rect 15800 8480 17300 8600
rect 15800 8410 17300 8480
rect 15800 8300 17300 8410
rect 19520 8420 19880 8580
rect 3300 7745 4600 7800
rect 3300 6000 3519 7745
rect 3519 6000 3585 7745
rect 3585 6000 3835 7745
rect 3835 6000 3901 7745
rect 3901 6000 4151 7745
rect 4151 6000 4217 7745
rect 4217 6000 4467 7745
rect 4467 6000 4533 7745
rect 4533 6000 4600 7745
rect 7700 7745 9000 7800
rect 7700 6000 7923 7745
rect 7923 6000 7989 7745
rect 7989 6000 8239 7745
rect 8239 6000 8305 7745
rect 8305 6000 8555 7745
rect 8555 6000 8621 7745
rect 8621 6000 8871 7745
rect 8871 6000 8937 7745
rect 8937 6000 9000 7745
rect 15900 7745 17200 7800
rect 15900 6000 16119 7745
rect 16119 6000 16185 7745
rect 16185 6000 16435 7745
rect 16435 6000 16501 7745
rect 16501 6000 16751 7745
rect 16751 6000 16817 7745
rect 16817 6000 17067 7745
rect 17067 6000 17133 7745
rect 17133 6000 17200 7745
rect 20300 7745 21600 7800
rect 20300 6000 20523 7745
rect 20523 6000 20589 7745
rect 20589 6000 20839 7745
rect 20839 6000 20905 7745
rect 20905 6000 21155 7745
rect 21155 6000 21221 7745
rect 21221 6000 21471 7745
rect 21471 6000 21537 7745
rect 21537 6000 21600 7745
rect 5200 4745 6500 4800
rect 5200 3000 5257 4745
rect 5257 3000 5323 4745
rect 5323 3000 5573 4745
rect 5573 3000 5639 4745
rect 5639 3000 5889 4745
rect 5889 3000 5955 4745
rect 5955 3000 6205 4745
rect 6205 3000 6271 4745
rect 6271 3000 6500 4745
rect 9600 4745 10900 4800
rect 9600 3000 9661 4745
rect 9661 3000 9727 4745
rect 9727 3000 9977 4745
rect 9977 3000 10043 4745
rect 10043 3000 10293 4745
rect 10293 3000 10359 4745
rect 10359 3000 10609 4745
rect 10609 3000 10675 4745
rect 10675 3000 10900 4745
rect 17800 4745 19100 4800
rect 17800 3000 17857 4745
rect 17857 3000 17923 4745
rect 17923 3000 18173 4745
rect 18173 3000 18239 4745
rect 18239 3000 18489 4745
rect 18489 3000 18555 4745
rect 18555 3000 18805 4745
rect 18805 3000 18871 4745
rect 18871 3000 19100 4745
rect 22200 4745 23500 4800
rect 22200 3000 22261 4745
rect 22261 3000 22327 4745
rect 22327 3000 22577 4745
rect 22577 3000 22643 4745
rect 22643 3000 22893 4745
rect 22893 3000 22959 4745
rect 22959 3000 23209 4745
rect 23209 3000 23275 4745
rect 23275 3000 23500 4745
<< metal4 >>
rect 1300 48000 2800 48100
rect 1300 46800 1400 48000
rect 2700 46800 2800 48000
rect -3400 40800 800 46000
rect 1300 45400 2800 46800
rect 9500 48000 11000 48100
rect 9500 46800 9600 48000
rect 10900 46800 11000 48000
rect 1300 43600 1400 45400
rect 2700 43600 2800 45400
rect 1300 43500 2800 43600
rect 5100 46200 6600 46300
rect 5100 45000 5200 46200
rect 6500 45000 6600 46200
rect -3400 40480 -3000 40500
rect -3400 40410 -3380 40480
rect -3400 40190 -3390 40410
rect -3020 40410 -3000 40480
rect -3010 40190 -3000 40410
rect -3400 40100 -3000 40190
rect -1000 39100 800 40800
rect -3440 38960 -3000 39000
rect -3440 38700 -3400 38960
rect -3020 38910 -3000 38960
rect -3010 38700 -3000 38910
rect -3440 38690 -3390 38700
rect -3010 38690 -1600 38700
rect -3440 38660 -1600 38690
rect -3400 38600 -1600 38660
rect -3400 37600 -3300 38600
rect -1700 37600 -1600 38600
rect -3400 37500 -1600 37600
rect -4400 25710 -4000 25720
rect -4400 25490 -4390 25710
rect -4010 25490 -4000 25710
rect -4400 25450 -4370 25490
rect -4030 25450 -4000 25490
rect -4400 25430 -4000 25450
rect -3400 24900 -1600 37100
rect -6400 14300 -1600 24900
rect -1000 25500 -600 39100
rect 700 25500 800 39100
rect 1300 42400 2800 42500
rect 1300 40600 1400 42400
rect 2700 40600 2800 42400
rect 1300 33100 2800 40600
rect 3100 40100 4800 40200
rect 3100 39800 3200 40100
rect 4700 39800 4800 40100
rect 3100 39700 4800 39800
rect 3100 39200 4800 39300
rect 3100 38900 3200 39200
rect 4700 38900 4800 39200
rect 3100 38800 4800 38900
rect 1300 31900 1400 33100
rect 2700 31900 2800 33100
rect 1300 31700 2800 31900
rect 1300 31100 1400 31700
rect 2700 31100 2800 31700
rect 1300 30100 2800 31100
rect 1300 28300 1400 30100
rect 2700 28300 2800 30100
rect 3200 38400 4700 38500
rect 3200 36600 3300 38400
rect 4600 36600 4700 38400
rect 3200 30900 4700 36600
rect 5100 35400 6600 45000
rect 7600 46200 9100 46300
rect 7600 43600 7700 46200
rect 9000 45000 9100 46200
rect 8900 43600 9100 45000
rect 7600 43500 9100 43600
rect 6900 39880 7300 39900
rect 6900 39720 6920 39880
rect 7280 39720 7300 39880
rect 6900 39180 7300 39720
rect 6900 39020 6920 39180
rect 7280 39020 7300 39180
rect 6900 39000 7300 39020
rect 5100 33600 5200 35400
rect 6500 33600 6600 35400
rect 5100 33500 6600 33600
rect 7600 38400 9100 38500
rect 7600 36600 7700 38400
rect 9000 36600 9100 38400
rect 7600 33100 9100 36600
rect 9500 35400 11000 46800
rect 13900 48000 15400 48100
rect 13900 46800 14000 48000
rect 15300 46800 15400 48000
rect 13900 45400 15400 46800
rect 22100 48000 23600 48100
rect 22100 46800 22200 48000
rect 23500 46800 23600 48000
rect 13900 43600 14000 45400
rect 15300 43600 15400 45400
rect 13900 43500 15400 43600
rect 17700 46200 19200 46300
rect 17700 45000 17800 46200
rect 19100 45000 19200 46200
rect 9500 33600 9600 35400
rect 10900 33600 11000 35400
rect 9500 33500 11000 33600
rect 11400 42400 12900 42500
rect 11400 40600 11500 42400
rect 12800 40600 12900 42400
rect 7600 31900 7700 33100
rect 9000 31900 9100 33100
rect 7600 31800 9100 31900
rect 9500 33100 11000 33200
rect 9500 31900 9600 33100
rect 10900 31900 11000 33100
rect 3200 29700 3300 30900
rect 4600 29700 4700 30900
rect 3200 29600 4700 29700
rect 5100 30900 6600 31000
rect 5100 29700 5200 30900
rect 6500 29700 6600 30900
rect 1300 28200 2800 28300
rect -1000 23200 800 25500
rect -1000 18500 -600 23200
rect 700 18500 800 23200
rect -1000 17800 800 18500
rect -1000 16600 -900 17800
rect 700 16600 800 17800
rect -1000 16500 800 16600
rect 1300 27100 2800 27200
rect 1300 25300 1400 27100
rect 2700 25300 2800 27100
rect 1300 17800 2800 25300
rect 3100 24800 4800 24900
rect 3100 24500 3200 24800
rect 4700 24500 4800 24800
rect 3100 24400 4800 24500
rect 3100 23900 4800 24000
rect 3100 23600 3200 23900
rect 4700 23600 4800 23900
rect 3100 23500 4800 23600
rect 1300 16600 1400 17800
rect 2700 16600 2800 17800
rect -4400 14000 -4000 14010
rect -4400 13420 -4390 14000
rect -4010 13420 -4000 14000
rect -4400 13410 -4000 13420
rect -3400 13900 -1600 14300
rect 1300 14800 2800 16600
rect -3400 13100 800 13900
rect -4400 13090 800 13100
rect -4400 12510 -4390 13090
rect -4010 12510 800 13090
rect 1300 13000 1400 14800
rect 2700 13000 2800 14800
rect 3200 23100 4700 23200
rect 3200 21300 3300 23100
rect 4600 21300 4700 23100
rect 3200 15600 4700 21300
rect 5100 20100 6600 29700
rect 7600 30900 9100 31000
rect 7600 28300 7700 30900
rect 9000 29700 9100 30900
rect 8900 28300 9100 29700
rect 7600 28200 9100 28300
rect 6900 24580 7300 24600
rect 6900 24420 6920 24580
rect 7280 24420 7300 24580
rect 6900 23880 7300 24420
rect 6900 23720 6920 23880
rect 7280 23720 7300 23880
rect 6900 23700 7300 23720
rect 5100 18300 5200 20100
rect 6500 18300 6600 20100
rect 5100 18200 6600 18300
rect 7600 23100 9100 23200
rect 7600 21300 7700 23100
rect 9000 21300 9100 23100
rect 7600 17800 9100 21300
rect 9500 20100 11000 31900
rect 11400 30900 12900 40600
rect 13900 42400 15400 42500
rect 13900 40600 14000 42400
rect 15300 40600 15400 42400
rect 13200 39880 13600 39900
rect 13200 39720 13220 39880
rect 13580 39720 13600 39880
rect 13200 39180 13600 39720
rect 13200 39020 13220 39180
rect 13580 39020 13600 39180
rect 13200 39000 13600 39020
rect 11400 29700 11500 30900
rect 12800 29700 12900 30900
rect 11400 29600 12900 29700
rect 13900 33100 15400 40600
rect 15700 40100 17400 40200
rect 15700 39800 15800 40100
rect 17300 39800 17400 40100
rect 15700 39700 17400 39800
rect 15700 39200 17400 39300
rect 15700 38900 15800 39200
rect 17300 38900 17400 39200
rect 15700 38800 17400 38900
rect 13900 31900 14000 33100
rect 15300 31900 15400 33100
rect 13900 30100 15400 31900
rect 13900 28300 14000 30100
rect 15300 28300 15400 30100
rect 15800 38400 17300 38500
rect 15800 36600 15900 38400
rect 17200 36600 17300 38400
rect 15800 30900 17300 36600
rect 17700 35400 19200 45000
rect 20200 46200 21700 46300
rect 20200 43600 20300 46200
rect 21600 45000 21700 46200
rect 21500 43600 21700 45000
rect 20200 43500 21700 43600
rect 19500 39880 19900 39900
rect 19500 39720 19520 39880
rect 19880 39720 19900 39880
rect 19500 39180 19900 39720
rect 19500 39020 19520 39180
rect 19880 39020 19900 39180
rect 19500 39000 19900 39020
rect 17700 33600 17800 35400
rect 19100 33600 19200 35400
rect 17700 33500 19200 33600
rect 20200 38400 21700 38500
rect 20200 36600 20300 38400
rect 21600 36600 21700 38400
rect 20200 33100 21700 36600
rect 22100 35400 23600 46800
rect 22100 33600 22200 35400
rect 23500 33600 23600 35400
rect 22100 33500 23600 33600
rect 24000 42400 25500 42500
rect 24000 40600 24100 42400
rect 25400 40600 25500 42400
rect 20200 31900 20300 33100
rect 21600 31900 21700 33100
rect 20200 31800 21700 31900
rect 22100 33100 23600 33200
rect 22100 31900 22200 33100
rect 23500 31900 23600 33100
rect 15800 29700 15900 30900
rect 17200 29700 17300 30900
rect 15800 29600 17300 29700
rect 17700 30900 19200 31000
rect 17700 29700 17800 30900
rect 19100 29700 19200 30900
rect 13900 28200 15400 28300
rect 9500 18300 9600 20100
rect 10900 18300 11000 20100
rect 9500 18200 11000 18300
rect 11400 27100 12900 27200
rect 11400 25300 11500 27100
rect 12800 25300 12900 27100
rect 7600 16600 7700 17800
rect 9000 16600 9100 17800
rect 7600 16500 9100 16600
rect 9500 17800 11000 17900
rect 9500 16600 9600 17800
rect 10900 16600 11000 17800
rect 3200 14400 3300 15600
rect 4600 14400 4700 15600
rect 3200 14300 4700 14400
rect 5100 15600 6600 15700
rect 5100 14400 5200 15600
rect 6500 14400 6600 15600
rect 1300 12900 2800 13000
rect -4400 12500 800 12510
rect -3400 12100 800 12500
rect -3400 11100 -600 12100
rect -1000 8000 -600 11100
rect 700 10100 800 12100
rect 200 10000 800 10100
rect 1300 11800 2800 11900
rect 1300 10000 1400 11800
rect 2700 10000 2800 11800
rect 200 8000 300 10000
rect -1000 7900 300 8000
rect -1000 7400 800 7900
rect -7200 3600 800 7400
rect 1300 3600 2800 10000
rect 3100 9500 4800 9600
rect 3100 9200 3200 9500
rect 4700 9200 4800 9500
rect 3100 9100 4800 9200
rect 3100 8600 4800 8700
rect 3100 8300 3200 8600
rect 4700 8300 4800 8600
rect 3100 8200 4800 8300
rect -7200 3500 2800 3600
rect -7200 2300 1400 3500
rect 2700 2300 2800 3500
rect -7200 1200 2800 2300
rect -7200 400 -7100 1200
rect 2600 400 2800 1200
rect 3200 7800 4700 7900
rect 3200 6000 3300 7800
rect 4600 6000 4700 7800
rect 3200 1700 4700 6000
rect 5100 4800 6600 14400
rect 7600 15600 9100 15700
rect 7600 13000 7700 15600
rect 9000 14400 9100 15600
rect 8900 13000 9100 14400
rect 7600 12900 9100 13000
rect 6900 9280 7300 9300
rect 6900 9120 6920 9280
rect 7280 9120 7300 9280
rect 6900 8580 7300 9120
rect 6900 8420 6920 8580
rect 7280 8420 7300 8580
rect 6900 8400 7300 8420
rect 5100 3000 5200 4800
rect 6500 3000 6600 4800
rect 5100 2900 6600 3000
rect 7600 7800 9100 7900
rect 7600 6000 7700 7800
rect 9000 6000 9100 7800
rect 7600 3500 9100 6000
rect 7600 2300 7700 3500
rect 9000 2300 9100 3500
rect 9500 4800 11000 16600
rect 11400 15600 12900 25300
rect 13900 27100 15400 27200
rect 13900 25300 14000 27100
rect 15300 25300 15400 27100
rect 13200 24580 13600 24600
rect 13200 24420 13220 24580
rect 13580 24420 13600 24580
rect 13200 23880 13600 24420
rect 13200 23720 13220 23880
rect 13580 23720 13600 23880
rect 13200 23700 13600 23720
rect 11400 14400 11500 15600
rect 12800 14400 12900 15600
rect 11400 14300 12900 14400
rect 13900 17800 15400 25300
rect 15700 24800 17400 24900
rect 15700 24500 15800 24800
rect 17300 24500 17400 24800
rect 15700 24400 17400 24500
rect 15700 23900 17400 24000
rect 15700 23600 15800 23900
rect 17300 23600 17400 23900
rect 15700 23500 17400 23600
rect 13900 16600 14000 17800
rect 15300 16600 15400 17800
rect 13900 14800 15400 16600
rect 13900 13000 14000 14800
rect 15300 13000 15400 14800
rect 15800 23100 17300 23200
rect 15800 21300 15900 23100
rect 17200 21300 17300 23100
rect 15800 15600 17300 21300
rect 17700 20100 19200 29700
rect 20200 30900 21700 31000
rect 20200 28300 20300 30900
rect 21600 29700 21700 30900
rect 21500 28300 21700 29700
rect 20200 28200 21700 28300
rect 19500 24580 19900 24600
rect 19500 24420 19520 24580
rect 19880 24420 19900 24580
rect 19500 23880 19900 24420
rect 19500 23720 19520 23880
rect 19880 23720 19900 23880
rect 19500 23700 19900 23720
rect 17700 18300 17800 20100
rect 19100 18300 19200 20100
rect 17700 18200 19200 18300
rect 20200 23100 21700 23200
rect 20200 21300 20300 23100
rect 21600 21300 21700 23100
rect 20200 17800 21700 21300
rect 22100 20100 23600 31900
rect 24000 31700 25500 40600
rect 24000 31100 24100 31700
rect 25400 31100 25500 31700
rect 24000 30900 25500 31100
rect 24000 29700 24100 30900
rect 25400 29700 25500 30900
rect 24000 29600 25500 29700
rect 26000 40800 30200 46000
rect 26000 40700 27800 40800
rect 26000 39900 26100 40700
rect 27700 39900 27800 40700
rect 29800 40480 30200 40500
rect 29800 40410 29820 40480
rect 29800 40190 29810 40410
rect 30180 40410 30200 40480
rect 30190 40190 30200 40410
rect 29800 40100 30200 40190
rect 26000 38100 27800 39900
rect 29700 38960 30200 39000
rect 29700 38910 29820 38960
rect 30180 38910 30200 38960
rect 29700 38700 29810 38910
rect 22100 18300 22200 20100
rect 23500 18300 23600 20100
rect 22100 18200 23600 18300
rect 24000 27100 25500 27200
rect 24000 25300 24100 27100
rect 25400 25300 25500 27100
rect 20200 16600 20300 17800
rect 21600 16600 21700 17800
rect 20200 16500 21700 16600
rect 22100 17800 23600 17900
rect 22100 16600 22200 17800
rect 23500 16600 23600 17800
rect 15800 14400 15900 15600
rect 17200 14400 17300 15600
rect 15800 14300 17300 14400
rect 17700 15600 19200 15700
rect 17700 14400 17800 15600
rect 19100 14400 19200 15600
rect 13900 12900 15400 13000
rect 9500 3000 9600 4800
rect 10900 3000 11000 4800
rect 9500 2900 11000 3000
rect 11400 11800 12900 11900
rect 11400 10000 11500 11800
rect 12800 10000 12900 11800
rect 7600 2200 9100 2300
rect 3200 500 3300 1700
rect 4600 500 4700 1700
rect 3200 400 4700 500
rect 11400 1700 12900 10000
rect 13900 11800 15400 11900
rect 13900 10000 14000 11800
rect 15300 10000 15400 11800
rect 13200 9280 13600 9300
rect 13200 9120 13220 9280
rect 13580 9120 13600 9280
rect 13200 8580 13600 9120
rect 13200 8420 13220 8580
rect 13580 8420 13600 8580
rect 13200 8400 13600 8420
rect 13900 3500 15400 10000
rect 15700 9500 17400 9600
rect 15700 9200 15800 9500
rect 17300 9200 17400 9500
rect 15700 9100 17400 9200
rect 15700 8600 17400 8700
rect 15700 8300 15800 8600
rect 17300 8300 17400 8600
rect 15700 8200 17400 8300
rect 13900 2300 14000 3500
rect 15300 2300 15400 3500
rect 13900 2200 15400 2300
rect 15800 7800 17300 7900
rect 15800 6000 15900 7800
rect 17200 6000 17300 7800
rect 11400 500 11500 1700
rect 12800 500 12900 1700
rect 11400 400 12900 500
rect 15800 1700 17300 6000
rect 17700 4800 19200 14400
rect 20200 15600 21700 15700
rect 20200 13000 20300 15600
rect 21600 14400 21700 15600
rect 21500 13000 21700 14400
rect 20200 12900 21700 13000
rect 19500 9280 19900 9300
rect 19500 9120 19520 9280
rect 19880 9120 19900 9280
rect 19500 8580 19900 9120
rect 19500 8420 19520 8580
rect 19880 8420 19900 8580
rect 19500 8400 19900 8420
rect 17700 3000 17800 4800
rect 19100 3000 19200 4800
rect 17700 2900 19200 3000
rect 20200 7800 21700 7900
rect 20200 6000 20300 7800
rect 21600 6000 21700 7800
rect 20200 3500 21700 6000
rect 20200 2300 20300 3500
rect 21600 2300 21700 3500
rect 22100 4800 23600 16600
rect 24000 15600 25500 25300
rect 26000 25500 26100 38100
rect 27400 25500 27800 38100
rect 28400 38690 29810 38700
rect 30190 38690 30200 38910
rect 28400 38600 30200 38690
rect 28400 37600 28500 38600
rect 30100 37600 30200 38600
rect 28400 37500 30200 37600
rect 26000 23200 27800 25500
rect 26000 18500 26100 23200
rect 27400 18500 27800 23200
rect 26000 17800 27800 18500
rect 26000 16600 26100 17800
rect 27700 16600 27800 17800
rect 26000 16500 27800 16600
rect 28400 24900 30200 37100
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25450 30830 25490
rect 31170 25450 31200 25490
rect 30800 25430 31200 25450
rect 24000 14400 24100 15600
rect 25400 14400 25500 15600
rect 24000 14300 25500 14400
rect 28400 14300 33200 24900
rect 28400 13900 30200 14300
rect 26000 13100 30200 13900
rect 30800 14000 31200 14010
rect 30800 13420 30810 14000
rect 31190 13420 31200 14000
rect 30800 13410 31200 13420
rect 26000 13090 31200 13100
rect 26000 12510 30810 13090
rect 31190 12510 31200 13090
rect 26000 12500 31200 12510
rect 26000 12100 30200 12500
rect 22100 3000 22200 4800
rect 23500 3000 23600 4800
rect 22100 2900 23600 3000
rect 24000 11800 25500 11900
rect 24000 10000 24100 11800
rect 25400 10000 25500 11800
rect 26000 10100 26100 12100
rect 27400 11100 30200 12100
rect 26000 10000 26600 10100
rect 24000 3600 25500 10000
rect 26500 8000 26600 10000
rect 27400 8000 27800 11100
rect 26500 7900 27800 8000
rect 26000 7400 27800 7900
rect 26000 3600 34000 7400
rect 20200 2200 21700 2300
rect 15800 500 15900 1700
rect 17200 500 17300 1700
rect 15800 400 17300 500
rect 24000 1700 34000 3600
rect 24000 500 24100 1700
rect 25400 1200 34000 1700
rect 25400 500 25600 1200
rect 24000 400 25600 500
rect 33900 400 34000 1200
rect -7200 200 2800 400
rect 25500 200 34000 400
<< via4 >>
rect 1400 46800 2700 48000
rect 9600 46800 10900 48000
rect 5200 45000 6500 46200
rect -3370 40210 -3030 40450
rect -3400 38910 -3020 38960
rect -3400 38700 -3390 38910
rect -3390 38700 -3020 38910
rect -3300 37600 -1700 38600
rect -4370 25490 -4030 25690
rect -4370 25450 -4030 25490
rect -600 25500 700 39100
rect 3200 39800 4700 40100
rect 3200 38900 4700 39200
rect 1400 31900 2700 33100
rect 7700 45400 9000 46200
rect 7700 45000 8900 45400
rect 8900 45000 9000 45400
rect 14000 46800 15300 48000
rect 22200 46800 23500 48000
rect 17800 45000 19100 46200
rect 7700 31900 9000 33100
rect 9600 31900 10900 33100
rect 3300 29700 4600 30900
rect 5200 29700 6500 30900
rect -600 18500 700 23200
rect -900 16600 700 17800
rect 3200 24500 4700 24800
rect 3200 23600 4700 23900
rect 1400 16600 2700 17800
rect -4370 13440 -4030 13980
rect 7700 30100 9000 30900
rect 7700 29700 8900 30100
rect 8900 29700 9000 30100
rect 11500 29700 12800 30900
rect 15800 39800 17300 40100
rect 15800 38900 17300 39200
rect 14000 31900 15300 33100
rect 20300 45400 21600 46200
rect 20300 45000 21500 45400
rect 21500 45000 21600 45400
rect 20300 31900 21600 33100
rect 22200 31900 23500 33100
rect 15900 29700 17200 30900
rect 17800 29700 19100 30900
rect 7700 16600 9000 17800
rect 9600 16600 10900 17800
rect 3300 14400 4600 15600
rect 5200 14400 6500 15600
rect -600 10100 700 12100
rect -600 8000 200 10100
rect 3200 9200 4700 9500
rect 3200 8300 4700 8600
rect 1400 2300 2700 3500
rect -7100 400 2600 1200
rect 7700 14800 9000 15600
rect 7700 14400 8900 14800
rect 8900 14400 9000 14800
rect 7700 2300 9000 3500
rect 11500 14400 12800 15600
rect 15800 24500 17300 24800
rect 15800 23600 17300 23900
rect 14000 16600 15300 17800
rect 20300 30100 21600 30900
rect 20300 29700 21500 30100
rect 21500 29700 21600 30100
rect 24100 29700 25400 30900
rect 26100 39900 27700 40700
rect 29830 40210 30170 40450
rect 29820 38910 30180 38960
rect 29820 38720 30180 38910
rect 20300 16600 21600 17800
rect 22200 16600 23500 17800
rect 15900 14400 17200 15600
rect 17800 14400 19100 15600
rect 3300 500 4600 1700
rect 15800 9200 17300 9500
rect 15800 8300 17300 8600
rect 14000 2300 15300 3500
rect 11500 500 12800 1700
rect 20300 14800 21600 15600
rect 20300 14400 21500 14800
rect 21500 14400 21600 14800
rect 20300 2300 21600 3500
rect 26100 25500 27400 38100
rect 28500 37600 30100 38600
rect 26100 18500 27400 23200
rect 26100 16600 27700 17800
rect 30830 25490 31170 25690
rect 30830 25450 31170 25490
rect 24100 14400 25400 15600
rect 30830 13440 31170 13980
rect 26100 10100 27400 12100
rect 26600 8000 27400 10100
rect 15900 500 17200 1700
rect 24100 500 25400 1700
rect 25600 400 33900 1200
<< mimcap2 >>
rect -3300 45800 700 45900
rect -3300 41000 -3200 45800
rect 600 41000 700 45800
rect -3300 40900 700 41000
rect 26100 45800 30100 45900
rect 26100 41000 26200 45800
rect 30000 41000 30100 45800
rect 26100 40900 30100 41000
rect -3300 36900 -1700 37000
rect -3300 26700 -3200 36900
rect -1800 26700 -1700 36900
rect -3300 26600 -1700 26700
rect 28500 36900 30100 37000
rect 28500 26700 28600 36900
rect 30000 26700 30100 36900
rect 28500 26600 30100 26700
rect -6300 24700 -1700 24800
rect -6300 14500 -6200 24700
rect -1800 14500 -1700 24700
rect -6300 14400 -1700 14500
rect 28500 24700 33100 24800
rect 28500 14500 28600 24700
rect 33000 14500 33100 24700
rect 28500 14400 33100 14500
rect -7100 7200 700 7300
rect -7100 2400 -7000 7200
rect 600 2400 700 7200
rect -7100 2300 700 2400
rect 26100 7200 33900 7300
rect 26100 2400 26200 7200
rect 33800 2400 33900 7200
rect 26100 2300 33900 2400
<< mimcap2contact >>
rect -3200 41000 600 45800
rect 26200 41000 30000 45800
rect -3200 26700 -1800 36900
rect 28600 26700 30000 36900
rect -6200 14500 -1800 24700
rect 28600 14500 33000 24700
rect -7000 2400 600 7200
rect 26200 2400 33800 7200
<< metal5 >>
rect 1300 48100 2800 48500
rect 1300 48000 23600 48100
rect 1300 47600 1400 48000
rect -600 46800 1400 47600
rect 2700 46800 9600 48000
rect 10900 46800 14000 48000
rect 15300 46800 22200 48000
rect 23500 46800 23600 48000
rect -600 46700 23600 46800
rect 24000 47600 25500 48500
rect 24000 46700 27400 47600
rect -600 46000 800 46700
rect 24000 46300 25500 46700
rect -3400 45800 800 46000
rect -3400 41000 -3200 45800
rect 600 41000 800 45800
rect 5100 46200 25500 46300
rect 5100 45000 5200 46200
rect 6500 45000 7700 46200
rect 9000 45000 17800 46200
rect 19100 45000 20300 46200
rect 21600 45000 25500 46200
rect 5100 44900 25500 45000
rect 26000 46000 27400 46700
rect 26000 45800 30200 46000
rect -3400 40800 800 41000
rect 26000 41000 26200 45800
rect 30000 41000 30200 45800
rect 26000 40800 30200 41000
rect -3400 40450 -3000 40800
rect -3400 40210 -3370 40450
rect -3030 40210 -3000 40450
rect -3400 40100 -3000 40210
rect 26000 40700 27800 40800
rect -2400 40100 25400 40200
rect -2500 40000 3200 40100
rect -2600 39900 3200 40000
rect -2700 39800 3200 39900
rect 4700 39800 15800 40100
rect 17300 39800 25400 40100
rect 26000 39900 26100 40700
rect 27700 39900 27800 40700
rect 29800 40450 30200 40800
rect 29800 40210 29830 40450
rect 30170 40210 30200 40450
rect 29800 40100 30200 40210
rect 26000 39800 27800 39900
rect -2800 39700 25400 39800
rect -2900 39600 -1400 39700
rect -3000 39500 -1500 39600
rect -3000 39000 -1600 39500
rect 1200 39200 29200 39300
rect -3440 38960 -1600 39000
rect -3440 38700 -3400 38960
rect -3020 38700 -1600 38960
rect -3440 38660 -1600 38700
rect -3400 38600 -1600 38660
rect -3400 37600 -3300 38600
rect -1700 37600 -1600 38600
rect -3400 36900 -1600 37600
rect -3400 26700 -3200 36900
rect -1800 26700 -1600 36900
rect -3400 26500 -1600 26700
rect -700 39100 800 39200
rect -4400 25690 -4000 25720
rect -4400 25450 -4370 25690
rect -4030 25450 -4000 25690
rect -4400 24900 -4000 25450
rect -700 25500 -600 39100
rect 700 25500 800 39100
rect 1200 38900 3200 39200
rect 4700 38900 15800 39200
rect 17300 39100 29300 39200
rect 17300 39000 29400 39100
rect 17300 38960 30220 39000
rect 17300 38900 29820 38960
rect 1200 38800 29820 38900
rect 28200 38720 29820 38800
rect 30180 38720 30220 38960
rect 28200 38700 30220 38720
rect 28300 38660 30220 38700
rect 28300 38600 30200 38660
rect 26000 38100 27500 38200
rect 1300 33100 25500 33200
rect 1300 31900 1400 33100
rect 2700 31900 7700 33100
rect 9000 31900 9600 33100
rect 10900 31900 14000 33100
rect 15300 31900 20300 33100
rect 21600 31900 22200 33100
rect 23500 31900 25500 33100
rect 1300 31800 25500 31900
rect 1300 30900 25500 31000
rect 1300 29700 3300 30900
rect 4600 29700 5200 30900
rect 6500 29700 7700 30900
rect 9000 29700 11500 30900
rect 12800 29700 15900 30900
rect 17200 29700 17800 30900
rect 19100 29700 20300 30900
rect 21600 29700 24100 30900
rect 25400 29700 25500 30900
rect 1300 29600 25500 29700
rect -700 25400 800 25500
rect 26000 25500 26100 38100
rect 27400 25500 27500 38100
rect 28400 37600 28500 38600
rect 30100 37600 30200 38600
rect 28400 36900 30200 37600
rect 28400 26700 28600 36900
rect 30000 26700 30200 36900
rect 28400 26500 30200 26700
rect 26000 25400 27500 25500
rect 30800 25690 31200 25720
rect 30800 25450 30830 25690
rect 31170 25450 31200 25690
rect 30800 24900 31200 25450
rect -6400 24800 33200 24900
rect -6400 24700 3200 24800
rect -6400 14500 -6200 24700
rect -1800 24500 3200 24700
rect 4700 24500 15800 24800
rect 17300 24700 33200 24800
rect 17300 24500 28600 24700
rect -1800 24400 28600 24500
rect -1800 24000 2100 24400
rect 24700 24000 28600 24400
rect -1800 23900 28600 24000
rect -1800 23800 3200 23900
rect -1800 14500 -1600 23800
rect 1200 23600 3200 23800
rect 4700 23600 15800 23900
rect 17300 23800 28600 23900
rect 17300 23600 25400 23800
rect 1200 23500 25400 23600
rect -700 23200 800 23300
rect -700 18500 -600 23200
rect 700 18500 800 23200
rect -700 18400 800 18500
rect 26000 23200 27500 23300
rect 26000 18500 26100 23200
rect 27400 18500 27500 23200
rect 26000 18400 27500 18500
rect -6400 14300 -1600 14500
rect -1200 17800 28000 17900
rect -1200 16600 -900 17800
rect 700 16600 1400 17800
rect 2700 16600 7700 17800
rect 9000 16600 9600 17800
rect 10900 16600 14000 17800
rect 15300 16600 20300 17800
rect 21600 16600 22200 17800
rect 23500 16600 26100 17800
rect 27700 16600 28000 17800
rect -1200 16500 28000 16600
rect -4400 13980 -4000 14300
rect -4400 13440 -4370 13980
rect -4030 13440 -4000 13980
rect -1200 13900 0 16500
rect 1300 15600 25500 15700
rect 1300 14400 3300 15600
rect 4600 14400 5200 15600
rect 6500 14400 7700 15600
rect 9000 14400 11500 15600
rect 12800 14400 15900 15600
rect 17200 14400 17800 15600
rect 19100 14400 20300 15600
rect 21600 14400 24100 15600
rect 25400 14400 25500 15600
rect 1300 14300 25500 14400
rect -4400 13410 -4000 13440
rect -3400 12600 0 13900
rect 26800 13900 28000 16500
rect 28400 14500 28600 23800
rect 33000 14500 33200 24700
rect 28400 14300 33200 14500
rect 30800 13980 31200 14300
rect 26800 12600 30200 13900
rect 30800 13440 30830 13980
rect 31170 13440 31200 13980
rect 30800 13410 31200 13440
rect -3400 7400 -1600 12600
rect -700 12100 800 12200
rect -700 8000 -600 12100
rect 700 10100 800 12100
rect 200 10000 800 10100
rect 26000 12100 27500 12200
rect 26000 10100 26100 12100
rect 26000 10000 26600 10100
rect 200 8000 300 10000
rect 700 9500 25400 9600
rect 700 9200 3200 9500
rect 4700 9200 15800 9500
rect 17300 9200 25400 9500
rect 700 9100 25400 9200
rect 1200 8600 25900 8700
rect 1200 8300 3200 8600
rect 4700 8300 15800 8600
rect 17300 8300 25900 8600
rect 1200 8200 25900 8300
rect -700 7900 300 8000
rect 26500 8000 26600 10000
rect 27400 8000 27500 12100
rect 26500 7900 27500 8000
rect 28400 7400 30200 12600
rect -7200 7200 800 7400
rect -7200 2400 -7000 7200
rect 600 2400 800 7200
rect 26000 7200 34000 7400
rect -7200 2200 800 2400
rect 1300 3500 21700 3600
rect 1300 2300 1400 3500
rect 2700 2300 7700 3500
rect 9000 2300 14000 3500
rect 15300 2300 20300 3500
rect 21600 2300 21700 3500
rect 1300 2200 21700 2300
rect 26000 2400 26200 7200
rect 33800 2400 34000 7200
rect 26000 2200 34000 2400
rect 1300 1400 2800 2200
rect -7200 1200 2800 1400
rect -7200 400 -7100 1200
rect 2600 400 2800 1200
rect 3200 1700 25500 1800
rect 3200 500 3300 1700
rect 4600 500 11500 1700
rect 12800 500 15900 1700
rect 17200 500 24100 1700
rect 25400 1400 25500 1700
rect 25400 1200 34000 1400
rect 25400 500 25600 1200
rect 3200 400 25600 500
rect 33900 400 34000 1200
rect -7200 200 2800 400
rect 1300 0 2800 200
rect 24000 200 34000 400
rect 24000 0 25500 200
<< comment >>
rect 1300 46400 1400 46600
rect 5100 46500 5300 46600
rect 7600 46500 7800 46600
rect 9500 46500 9600 46700
rect 1300 46300 1500 46400
rect 5100 46312 5200 46500
rect 7600 46312 7700 46500
rect 9500 46400 9700 46500
rect 14000 46400 14100 46600
rect 17700 46500 17900 46600
rect 20200 46500 20400 46600
rect 22100 46500 22200 46700
rect 14000 46300 14200 46400
rect 17700 46312 17800 46500
rect 20200 46312 20300 46500
rect 22100 46400 22300 46500
rect 200 46100 300 46200
rect 100 45900 200 46100
rect 300 45900 400 46000
rect 100 45800 400 45900
rect 300 45700 400 45800
rect 1300 32500 1400 32700
rect 3200 32600 3400 32700
rect 1300 32400 1500 32500
rect 3200 32412 3300 32600
rect 7600 32500 7700 32700
rect 11400 32600 11600 32700
rect 7600 32400 7800 32500
rect 11400 32412 11500 32600
rect 13900 32500 14000 32700
rect 15800 32600 16000 32700
rect 13900 32400 14100 32500
rect 15800 32412 15900 32600
rect 20200 32500 20300 32700
rect 24000 32600 24200 32700
rect 20200 32400 20400 32500
rect 24000 32412 24100 32600
rect 0 31400 300 31500
rect 200 31300 300 31400
rect 100 31200 300 31300
rect 200 31100 300 31200
rect 0 31000 300 31100
rect 1300 31100 1400 31300
rect 5100 31200 5300 31300
rect 7600 31200 7800 31300
rect 9500 31200 9600 31400
rect 1300 31000 1500 31100
rect 5100 31012 5200 31200
rect 7600 31012 7700 31200
rect 9500 31100 9700 31200
rect 14000 31100 14100 31300
rect 17700 31200 17900 31300
rect 20200 31200 20400 31300
rect 22100 31200 22200 31400
rect 14000 31000 14200 31100
rect 17700 31012 17800 31200
rect 20200 31012 20300 31200
rect 22100 31100 22300 31200
rect 1300 17200 1400 17400
rect 3200 17300 3400 17400
rect 1300 17100 1500 17200
rect 3200 17112 3300 17300
rect 7600 17200 7700 17400
rect 11400 17300 11600 17400
rect 7600 17100 7800 17200
rect 11400 17112 11500 17300
rect 13900 17200 14000 17400
rect 15800 17300 16000 17400
rect 13900 17100 14100 17200
rect 15800 17112 15900 17300
rect 20200 17200 20300 17400
rect 24000 17300 24200 17400
rect 20200 17100 20400 17200
rect 24000 17112 24100 17300
rect 1300 15800 1400 16000
rect 5100 15900 5300 16000
rect 7600 15900 7800 16000
rect 9500 15900 9600 16100
rect 1300 15700 1500 15800
rect 5100 15712 5200 15900
rect 7600 15712 7700 15900
rect 9500 15800 9700 15900
rect 14000 15800 14100 16000
rect 17700 15900 17900 16000
rect 20200 15900 20400 16000
rect 22100 15900 22200 16100
rect 14000 15700 14200 15800
rect 17700 15712 17800 15900
rect 20200 15712 20300 15900
rect 22100 15800 22300 15900
rect 100 15600 400 15700
rect 300 15500 400 15600
rect 200 15400 400 15500
rect 100 15300 200 15400
rect 100 15200 400 15300
rect 1300 1900 1400 2100
rect 3200 2000 3400 2100
rect 1300 1800 1500 1900
rect 3200 1812 3300 2000
rect 7600 1900 7700 2100
rect 11400 2000 11600 2100
rect 7600 1800 7800 1900
rect 11400 1812 11500 2000
rect 13900 1900 14000 2100
rect 15800 2000 16000 2100
rect 13900 1800 14100 1900
rect 15800 1812 15900 2000
rect 20200 1900 20300 2100
rect 24000 2000 24200 2100
rect 20200 1800 20400 1900
rect 24000 1812 24100 2000
rect 400 800 500 900
rect 300 700 500 800
rect 400 500 500 700
rect 300 400 600 500
<< res0p35 >>
rect -4236 13096 -4162 13420
<< labels >>
rlabel metal5 1300 48100 2800 48500 1 VDN
rlabel metal5 900 39700 1200 40200 1 VGN
rlabel metal3 800 31000 1000 31800 1 N2
rlabel metal5 900 16500 1200 17900 1 N
rlabel metal5 700 9100 1000 9600 1 VINN
rlabel metal5 1300 0 2800 400 1 VSS
rlabel metal5 800 23800 1000 24800 1 MIDGATE
rlabel metal5 24000 48300 25500 48500 1 VDP
rlabel metal3 25600 31100 25900 31700 1 P2
rlabel metal5 25600 16500 25900 17900 1 P
rlabel metal5 24000 0 25500 200 1 VSSH
rlabel metal5 25700 38800 25900 39300 1 VGP
rlabel metal5 25700 8200 25900 8700 1 VINP
rlabel metal1 -3920 13900 -3540 14000 1 SUB
rlabel metal5 1300 0 2800 400 1 cascode_1_0/SD1L
rlabel metal5 24000 0 25500 400 1 cascode_1_0/SD1R
rlabel metal5 1300 14300 1600 15700 1 cascode_1_0/SD2R
rlabel metal5 1300 16500 1600 17900 1 cascode_1_0/SD2L
rlabel metal5 1300 29600 1600 31000 1 cascode_1_0/SD3R
rlabel metal5 1300 31800 1600 33200 1 cascode_1_0/SD3L
rlabel metal5 1300 48100 2800 48500 1 cascode_1_0/SD4L
rlabel metal5 24000 48100 25500 48500 1 cascode_1_0/SD4R
rlabel metal5 1200 9100 1300 9600 1 cascode_1_0/G12L
rlabel metal5 1200 8200 1300 8700 1 cascode_1_0/G12R
rlabel metal5 1200 23500 1300 24000 1 cascode_1_0/G23R
rlabel metal5 1200 24400 1300 24900 1 cascode_1_0/G23L
rlabel metal5 1200 38800 1300 39300 1 cascode_1_0/G34R
rlabel metal5 1200 39700 1300 40200 1 cascode_1_0/G34L
rlabel metal5 1200 39700 1300 40200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/GL
rlabel metal5 1200 38800 1300 39300 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/GR
rlabel metal2 13930 39120 14000 39180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/SUB
rlabel metal2 1330 39120 1400 39180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SUB
rlabel metal3 1440 39000 1500 39200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/G
rlabel metal3 1520 36510 1560 38470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD1
rlabel metal3 1490 33510 1530 35470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_7/SD2
rlabel metal2 7630 39120 7700 39180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SUB
rlabel metal3 7740 39000 7800 39200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/G
rlabel metal3 7820 36510 7860 38470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD1
rlabel metal3 7790 33510 7830 35470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_6/SD2
rlabel metal2 13930 39120 14000 39180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_5/SUB
rlabel metal3 14040 39000 14100 39200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_5/G
rlabel metal3 14120 36510 14160 38470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_5/SD1
rlabel metal3 14090 33510 14130 35470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_5/SD2
rlabel metal2 20230 39120 20300 39180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SUB
rlabel metal3 20340 39000 20400 39200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/G
rlabel metal3 20420 36510 20460 38470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD1
rlabel metal3 20390 33510 20430 35470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_4/SD2
rlabel metal2 20230 46120 20300 46180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_3/SUB
rlabel metal3 20340 46000 20400 46200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_3/G
rlabel metal3 20420 43510 20460 45470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_3/SD1
rlabel metal3 20390 40510 20430 42470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_3/SD2
rlabel metal2 13930 46120 14000 46180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SUB
rlabel metal3 14040 46000 14100 46200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/G
rlabel metal3 14120 43510 14160 45470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD1
rlabel metal3 14090 40510 14130 42470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_2/SD2
rlabel metal2 7630 46120 7700 46180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/SUB
rlabel metal3 7740 46000 7800 46200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/G
rlabel metal3 7820 43510 7860 45470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/SD1
rlabel metal3 7790 40510 7830 42470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_1/SD2
rlabel metal2 1330 46120 1400 46180 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SUB
rlabel metal3 1440 46000 1500 46200 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/G
rlabel metal3 1520 43510 1560 45470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD1
rlabel metal3 1490 40510 1530 42470 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_2/NMOS_30_0p5_30_1_0/SD2
rlabel metal5 1200 24400 1300 24900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/GL
rlabel metal5 1200 23500 1300 24000 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/GR
rlabel metal2 13930 23820 14000 23880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/SUB
rlabel metal2 1330 23820 1400 23880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SUB
rlabel metal3 1440 23700 1500 23900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/G
rlabel metal3 1520 21210 1560 23170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD1
rlabel metal3 1490 18210 1530 20170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_7/SD2
rlabel metal2 7630 23820 7700 23880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_6/SUB
rlabel metal3 7740 23700 7800 23900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_6/G
rlabel metal3 7820 21210 7860 23170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_6/SD1
rlabel metal3 7790 18210 7830 20170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_6/SD2
rlabel metal2 13930 23820 14000 23880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/SUB
rlabel metal3 14040 23700 14100 23900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/G
rlabel metal3 14120 21210 14160 23170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/SD1
rlabel metal3 14090 18210 14130 20170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_5/SD2
rlabel metal2 20230 23820 20300 23880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_4/SUB
rlabel metal3 20340 23700 20400 23900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_4/G
rlabel metal3 20420 21210 20460 23170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_4/SD1
rlabel metal3 20390 18210 20430 20170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_4/SD2
rlabel metal2 20230 30820 20300 30880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SUB
rlabel metal3 20340 30700 20400 30900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/G
rlabel metal3 20420 28210 20460 30170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD1
rlabel metal3 20390 25210 20430 27170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_3/SD2
rlabel metal2 13930 30820 14000 30880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SUB
rlabel metal3 14040 30700 14100 30900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/G
rlabel metal3 14120 28210 14160 30170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD1
rlabel metal3 14090 25210 14130 27170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_2/SD2
rlabel metal2 7630 30820 7700 30880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SUB
rlabel metal3 7740 30700 7800 30900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/G
rlabel metal3 7820 28210 7860 30170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD1
rlabel metal3 7790 25210 7830 27170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_1/SD2
rlabel metal2 1330 30820 1400 30880 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SUB
rlabel metal3 1440 30700 1500 30900 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/G
rlabel metal3 1520 28210 1560 30170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD1
rlabel metal3 1490 25210 1530 27170 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_1/NMOS_30_0p5_30_1_0/SD2
rlabel metal5 1200 9100 1300 9600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/GL
rlabel metal5 1200 8200 1300 8700 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/GR
rlabel metal2 13930 8520 14000 8580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/SUB
rlabel metal2 1330 8520 1400 8580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SUB
rlabel metal3 1440 8400 1500 8600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/G
rlabel metal3 1520 5910 1560 7870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD1
rlabel metal3 1490 2910 1530 4870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_7/SD2
rlabel metal2 7630 8520 7700 8580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SUB
rlabel metal3 7740 8400 7800 8600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/G
rlabel metal3 7820 5910 7860 7870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD1
rlabel metal3 7790 2910 7830 4870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_6/SD2
rlabel metal2 13930 8520 14000 8580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SUB
rlabel metal3 14040 8400 14100 8600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/G
rlabel metal3 14120 5910 14160 7870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD1
rlabel metal3 14090 2910 14130 4870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_5/SD2
rlabel metal2 20230 8520 20300 8580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SUB
rlabel metal3 20340 8400 20400 8600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/G
rlabel metal3 20420 5910 20460 7870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD1
rlabel metal3 20390 2910 20430 4870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_4/SD2
rlabel metal2 20230 15520 20300 15580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SUB
rlabel metal3 20340 15400 20400 15600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/G
rlabel metal3 20420 12910 20460 14870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD1
rlabel metal3 20390 9910 20430 11870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_3/SD2
rlabel metal2 13930 15520 14000 15580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SUB
rlabel metal3 14040 15400 14100 15600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/G
rlabel metal3 14120 12910 14160 14870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD1
rlabel metal3 14090 9910 14130 11870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_2/SD2
rlabel metal2 7630 15520 7700 15580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SUB
rlabel metal3 7740 15400 7800 15600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/G
rlabel metal3 7820 12910 7860 14870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD1
rlabel metal3 7790 9910 7830 11870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_1/SD2
rlabel metal2 1330 15520 1400 15580 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SUB
rlabel metal3 1440 15400 1500 15600 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/G
rlabel metal3 1520 12910 1560 14870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD1
rlabel metal3 1490 9910 1530 11870 1 cascode_1_0/NMOS_30_0p5_30_diff4x_2s_0/NMOS_30_0p5_30_1_0/SD2
<< end >>
