magic
tech sky130B
timestamp 1662579390
<< nwell >>
rect -569 -518 569 518
<< pwell >>
rect -638 518 638 587
rect -638 -518 -569 518
rect 569 -518 638 518
rect -638 -587 638 -518
<< psubdiff >>
rect -620 552 -572 569
rect 572 552 620 569
rect -620 521 -603 552
rect 603 521 620 552
rect -620 -552 -603 -521
rect 603 -552 620 -521
rect -620 -569 -572 -552
rect 572 -569 620 -552
<< nsubdiff >>
rect -551 483 -503 500
rect 503 483 551 500
rect -551 452 -534 483
rect 534 452 551 483
rect -551 315 -534 346
rect 534 315 551 346
rect -551 298 -503 315
rect 503 298 551 315
rect -551 217 -503 234
rect 503 217 551 234
rect -551 186 -534 217
rect 534 186 551 217
rect -551 49 -534 80
rect 534 49 551 80
rect -551 32 -503 49
rect 503 32 551 49
rect -551 -49 -503 -32
rect 503 -49 551 -32
rect -551 -80 -534 -49
rect 534 -80 551 -49
rect -551 -217 -534 -186
rect 534 -217 551 -186
rect -551 -234 -503 -217
rect 503 -234 551 -217
rect -551 -315 -503 -298
rect 503 -315 551 -298
rect -551 -346 -534 -315
rect 534 -346 551 -315
rect -551 -483 -534 -452
rect 534 -483 551 -452
rect -551 -500 -503 -483
rect 503 -500 551 -483
<< psubdiffcont >>
rect -572 552 572 569
rect -620 -521 -603 521
rect 603 -521 620 521
rect -572 -569 572 -552
<< nsubdiffcont >>
rect -503 483 503 500
rect -551 346 -534 452
rect 534 346 551 452
rect -503 298 503 315
rect -503 217 503 234
rect -551 80 -534 186
rect 534 80 551 186
rect -503 32 503 49
rect -503 -49 503 -32
rect -551 -186 -534 -80
rect 534 -186 551 -80
rect -503 -234 503 -217
rect -503 -315 503 -298
rect -551 -452 -534 -346
rect 534 -452 551 -346
rect -503 -500 503 -483
<< pdiode >>
rect -500 443 500 449
rect -500 355 -494 443
rect 494 355 500 443
rect -500 349 500 355
rect -500 177 500 183
rect -500 89 -494 177
rect 494 89 500 177
rect -500 83 500 89
rect -500 -89 500 -83
rect -500 -177 -494 -89
rect 494 -177 500 -89
rect -500 -183 500 -177
rect -500 -355 500 -349
rect -500 -443 -494 -355
rect 494 -443 500 -355
rect -500 -449 500 -443
<< pdiodec >>
rect -494 355 494 443
rect -494 89 494 177
rect -494 -177 494 -89
rect -494 -443 494 -355
<< locali >>
rect -620 552 -572 569
rect 572 552 620 569
rect -620 521 -603 552
rect 603 521 620 552
rect -551 483 -503 500
rect 503 483 551 500
rect -551 452 -534 483
rect 534 452 551 483
rect -502 355 -494 443
rect 494 355 502 443
rect -551 315 -534 346
rect 534 315 551 346
rect -551 298 -503 315
rect 503 298 551 315
rect -551 217 -503 234
rect 503 217 551 234
rect -551 186 -534 217
rect 534 186 551 217
rect -502 89 -494 177
rect 494 89 502 177
rect -551 49 -534 80
rect 534 49 551 80
rect -551 32 -503 49
rect 503 32 551 49
rect -551 -49 -503 -32
rect 503 -49 551 -32
rect -551 -80 -534 -49
rect 534 -80 551 -49
rect -502 -177 -494 -89
rect 494 -177 502 -89
rect -551 -217 -534 -186
rect 534 -217 551 -186
rect -551 -234 -503 -217
rect 503 -234 551 -217
rect -551 -315 -503 -298
rect 503 -315 551 -298
rect -551 -346 -534 -315
rect 534 -346 551 -315
rect -502 -443 -494 -355
rect 494 -443 502 -355
rect -551 -483 -534 -452
rect 534 -483 551 -452
rect -551 -500 -503 -483
rect 503 -500 551 -483
rect -620 -552 -603 -521
rect 603 -552 620 -521
rect -620 -569 -572 -552
rect 572 -569 620 -552
<< viali >>
rect -494 355 494 443
rect -494 89 494 177
rect -494 -177 494 -89
rect -494 -443 494 -355
<< metal1 >>
rect -500 443 500 446
rect -500 355 -494 443
rect 494 355 500 443
rect -500 352 500 355
rect -500 177 500 180
rect -500 89 -494 177
rect 494 89 500 177
rect -500 86 500 89
rect -500 -89 500 -86
rect -500 -177 -494 -89
rect 494 -177 500 -89
rect -500 -180 500 -177
rect -500 -355 500 -352
rect -500 -443 -494 -355
rect 494 -443 500 -355
rect -500 -446 500 -443
<< properties >>
string FIXED_BBOX -542 306 542 491
string gencell sky130_fd_pr__diode_pd2nw_05v5
string library sky130
string parameters w 10 l 1 area 10.0 peri 22.0 nx 1 ny 4 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
