magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< locali >>
rect 4182 25143 4216 25177
rect 558 24964 624 24998
rect 558 24772 624 24806
rect 4182 24593 4216 24627
rect 4182 24353 4216 24387
rect 558 24174 624 24208
rect 558 23982 624 24016
rect 4182 23803 4216 23837
rect 4182 23563 4216 23597
rect 558 23384 624 23418
rect 558 23192 624 23226
rect 4182 23013 4216 23047
rect 4182 22773 4216 22807
rect 558 22594 624 22628
rect 558 22402 624 22436
rect 4182 22223 4216 22257
rect 4182 21983 4216 22017
rect 558 21804 624 21838
rect 558 21612 624 21646
rect 4182 21433 4216 21467
rect 4182 21193 4216 21227
rect 558 21014 624 21048
rect 558 20822 624 20856
rect 4182 20643 4216 20677
rect 4182 20403 4216 20437
rect 558 20224 624 20258
rect 558 20032 624 20066
rect 4182 19853 4216 19887
rect 4182 19613 4216 19647
rect 558 19434 624 19468
rect 558 19242 624 19276
rect 4182 19063 4216 19097
rect 4182 18823 4216 18857
rect 558 18644 624 18678
rect 558 18452 624 18486
rect 4182 18273 4216 18307
rect 4182 18033 4216 18067
rect 558 17854 624 17888
rect 558 17662 624 17696
rect 4182 17483 4216 17517
rect 4182 17243 4216 17277
rect 558 17064 624 17098
rect 558 16872 624 16906
rect 4182 16693 4216 16727
rect 4182 16453 4216 16487
rect 558 16274 624 16308
rect 558 16082 624 16116
rect 4182 15903 4216 15937
rect 4182 15663 4216 15697
rect 558 15484 624 15518
rect 558 15292 624 15326
rect 4182 15113 4216 15147
rect 4182 14873 4216 14907
rect 558 14694 624 14728
rect 558 14502 624 14536
rect 4182 14323 4216 14357
rect 4182 14083 4216 14117
rect 558 13904 624 13938
rect 558 13712 624 13746
rect 4182 13533 4216 13567
rect 4182 13293 4216 13327
rect 558 13114 624 13148
rect 558 12922 624 12956
rect 4182 12743 4216 12777
rect 4182 12503 4216 12537
rect 558 12324 624 12358
rect 558 12132 624 12166
rect 4182 11953 4216 11987
rect 4182 11713 4216 11747
rect 558 11534 624 11568
rect 558 11342 624 11376
rect 4182 11163 4216 11197
rect 4182 10923 4216 10957
rect 558 10744 624 10778
rect 558 10552 624 10586
rect 4182 10373 4216 10407
rect 4182 10133 4216 10167
rect 558 9954 624 9988
rect 558 9762 624 9796
rect 4182 9583 4216 9617
rect 4182 9343 4216 9377
rect 558 9164 624 9198
rect 558 8972 624 9006
rect 4182 8793 4216 8827
rect 4182 8553 4216 8587
rect 558 8374 624 8408
rect 558 8182 624 8216
rect 4182 8003 4216 8037
rect 4182 7763 4216 7797
rect 558 7584 624 7618
rect 558 7392 624 7426
rect 4182 7213 4216 7247
rect 4182 6973 4216 7007
rect 558 6794 624 6828
rect 558 6602 624 6636
rect 4182 6423 4216 6457
rect 4182 6183 4216 6217
rect 558 6004 624 6038
rect 558 5812 624 5846
rect 4182 5633 4216 5667
rect 4182 5393 4216 5427
rect 558 5214 624 5248
rect 558 5022 624 5056
rect 4182 4843 4216 4877
rect 4182 4603 4216 4637
rect 558 4424 624 4458
rect 558 4232 624 4266
rect 4182 4053 4216 4087
rect 4182 3813 4216 3847
rect 558 3634 624 3668
rect 558 3442 624 3476
rect 4182 3263 4216 3297
rect 4182 3023 4216 3057
rect 558 2844 624 2878
rect 558 2652 624 2686
rect 4182 2473 4216 2507
rect 4182 2233 4216 2267
rect 558 2054 624 2088
rect 558 1862 624 1896
rect 4182 1683 4216 1717
rect 4182 1443 4216 1477
rect 558 1264 624 1298
rect 558 1072 624 1106
rect 4182 893 4216 927
rect 4182 653 4216 687
rect 558 474 624 508
rect 558 282 624 316
rect 4182 103 4216 137
<< metal1 >>
rect 559 25063 623 25115
rect 726 25068 790 25120
rect 1151 25069 1215 25121
rect 1994 25056 2058 25108
rect 3442 25056 3506 25108
rect 559 24655 623 24707
rect 726 24650 790 24702
rect 1151 24649 1215 24701
rect 1994 24662 2058 24714
rect 3442 24662 3506 24714
rect 559 24273 623 24325
rect 726 24278 790 24330
rect 1151 24279 1215 24331
rect 1994 24266 2058 24318
rect 3442 24266 3506 24318
rect 559 23865 623 23917
rect 726 23860 790 23912
rect 1151 23859 1215 23911
rect 1994 23872 2058 23924
rect 3442 23872 3506 23924
rect 559 23483 623 23535
rect 726 23488 790 23540
rect 1151 23489 1215 23541
rect 1994 23476 2058 23528
rect 3442 23476 3506 23528
rect 559 23075 623 23127
rect 726 23070 790 23122
rect 1151 23069 1215 23121
rect 1994 23082 2058 23134
rect 3442 23082 3506 23134
rect 559 22693 623 22745
rect 726 22698 790 22750
rect 1151 22699 1215 22751
rect 1994 22686 2058 22738
rect 3442 22686 3506 22738
rect 559 22285 623 22337
rect 726 22280 790 22332
rect 1151 22279 1215 22331
rect 1994 22292 2058 22344
rect 3442 22292 3506 22344
rect 559 21903 623 21955
rect 726 21908 790 21960
rect 1151 21909 1215 21961
rect 1994 21896 2058 21948
rect 3442 21896 3506 21948
rect 559 21495 623 21547
rect 726 21490 790 21542
rect 1151 21489 1215 21541
rect 1994 21502 2058 21554
rect 3442 21502 3506 21554
rect 559 21113 623 21165
rect 726 21118 790 21170
rect 1151 21119 1215 21171
rect 1994 21106 2058 21158
rect 3442 21106 3506 21158
rect 559 20705 623 20757
rect 726 20700 790 20752
rect 1151 20699 1215 20751
rect 1994 20712 2058 20764
rect 3442 20712 3506 20764
rect 559 20323 623 20375
rect 726 20328 790 20380
rect 1151 20329 1215 20381
rect 1994 20316 2058 20368
rect 3442 20316 3506 20368
rect 559 19915 623 19967
rect 726 19910 790 19962
rect 1151 19909 1215 19961
rect 1994 19922 2058 19974
rect 3442 19922 3506 19974
rect 559 19533 623 19585
rect 726 19538 790 19590
rect 1151 19539 1215 19591
rect 1994 19526 2058 19578
rect 3442 19526 3506 19578
rect 559 19125 623 19177
rect 726 19120 790 19172
rect 1151 19119 1215 19171
rect 1994 19132 2058 19184
rect 3442 19132 3506 19184
rect 559 18743 623 18795
rect 726 18748 790 18800
rect 1151 18749 1215 18801
rect 1994 18736 2058 18788
rect 3442 18736 3506 18788
rect 559 18335 623 18387
rect 726 18330 790 18382
rect 1151 18329 1215 18381
rect 1994 18342 2058 18394
rect 3442 18342 3506 18394
rect 559 17953 623 18005
rect 726 17958 790 18010
rect 1151 17959 1215 18011
rect 1994 17946 2058 17998
rect 3442 17946 3506 17998
rect 559 17545 623 17597
rect 726 17540 790 17592
rect 1151 17539 1215 17591
rect 1994 17552 2058 17604
rect 3442 17552 3506 17604
rect 559 17163 623 17215
rect 726 17168 790 17220
rect 1151 17169 1215 17221
rect 1994 17156 2058 17208
rect 3442 17156 3506 17208
rect 559 16755 623 16807
rect 726 16750 790 16802
rect 1151 16749 1215 16801
rect 1994 16762 2058 16814
rect 3442 16762 3506 16814
rect 559 16373 623 16425
rect 726 16378 790 16430
rect 1151 16379 1215 16431
rect 1994 16366 2058 16418
rect 3442 16366 3506 16418
rect 559 15965 623 16017
rect 726 15960 790 16012
rect 1151 15959 1215 16011
rect 1994 15972 2058 16024
rect 3442 15972 3506 16024
rect 559 15583 623 15635
rect 726 15588 790 15640
rect 1151 15589 1215 15641
rect 1994 15576 2058 15628
rect 3442 15576 3506 15628
rect 559 15175 623 15227
rect 726 15170 790 15222
rect 1151 15169 1215 15221
rect 1994 15182 2058 15234
rect 3442 15182 3506 15234
rect 559 14793 623 14845
rect 726 14798 790 14850
rect 1151 14799 1215 14851
rect 1994 14786 2058 14838
rect 3442 14786 3506 14838
rect 559 14385 623 14437
rect 726 14380 790 14432
rect 1151 14379 1215 14431
rect 1994 14392 2058 14444
rect 3442 14392 3506 14444
rect 559 14003 623 14055
rect 726 14008 790 14060
rect 1151 14009 1215 14061
rect 1994 13996 2058 14048
rect 3442 13996 3506 14048
rect 559 13595 623 13647
rect 726 13590 790 13642
rect 1151 13589 1215 13641
rect 1994 13602 2058 13654
rect 3442 13602 3506 13654
rect 559 13213 623 13265
rect 726 13218 790 13270
rect 1151 13219 1215 13271
rect 1994 13206 2058 13258
rect 3442 13206 3506 13258
rect 559 12805 623 12857
rect 726 12800 790 12852
rect 1151 12799 1215 12851
rect 1994 12812 2058 12864
rect 3442 12812 3506 12864
rect 559 12423 623 12475
rect 726 12428 790 12480
rect 1151 12429 1215 12481
rect 1994 12416 2058 12468
rect 3442 12416 3506 12468
rect 559 12015 623 12067
rect 726 12010 790 12062
rect 1151 12009 1215 12061
rect 1994 12022 2058 12074
rect 3442 12022 3506 12074
rect 559 11633 623 11685
rect 726 11638 790 11690
rect 1151 11639 1215 11691
rect 1994 11626 2058 11678
rect 3442 11626 3506 11678
rect 559 11225 623 11277
rect 726 11220 790 11272
rect 1151 11219 1215 11271
rect 1994 11232 2058 11284
rect 3442 11232 3506 11284
rect 559 10843 623 10895
rect 726 10848 790 10900
rect 1151 10849 1215 10901
rect 1994 10836 2058 10888
rect 3442 10836 3506 10888
rect 559 10435 623 10487
rect 726 10430 790 10482
rect 1151 10429 1215 10481
rect 1994 10442 2058 10494
rect 3442 10442 3506 10494
rect 559 10053 623 10105
rect 726 10058 790 10110
rect 1151 10059 1215 10111
rect 1994 10046 2058 10098
rect 3442 10046 3506 10098
rect 559 9645 623 9697
rect 726 9640 790 9692
rect 1151 9639 1215 9691
rect 1994 9652 2058 9704
rect 3442 9652 3506 9704
rect 559 9263 623 9315
rect 726 9268 790 9320
rect 1151 9269 1215 9321
rect 1994 9256 2058 9308
rect 3442 9256 3506 9308
rect 559 8855 623 8907
rect 726 8850 790 8902
rect 1151 8849 1215 8901
rect 1994 8862 2058 8914
rect 3442 8862 3506 8914
rect 559 8473 623 8525
rect 726 8478 790 8530
rect 1151 8479 1215 8531
rect 1994 8466 2058 8518
rect 3442 8466 3506 8518
rect 559 8065 623 8117
rect 726 8060 790 8112
rect 1151 8059 1215 8111
rect 1994 8072 2058 8124
rect 3442 8072 3506 8124
rect 559 7683 623 7735
rect 726 7688 790 7740
rect 1151 7689 1215 7741
rect 1994 7676 2058 7728
rect 3442 7676 3506 7728
rect 559 7275 623 7327
rect 726 7270 790 7322
rect 1151 7269 1215 7321
rect 1994 7282 2058 7334
rect 3442 7282 3506 7334
rect 559 6893 623 6945
rect 726 6898 790 6950
rect 1151 6899 1215 6951
rect 1994 6886 2058 6938
rect 3442 6886 3506 6938
rect 559 6485 623 6537
rect 726 6480 790 6532
rect 1151 6479 1215 6531
rect 1994 6492 2058 6544
rect 3442 6492 3506 6544
rect 559 6103 623 6155
rect 726 6108 790 6160
rect 1151 6109 1215 6161
rect 1994 6096 2058 6148
rect 3442 6096 3506 6148
rect 559 5695 623 5747
rect 726 5690 790 5742
rect 1151 5689 1215 5741
rect 1994 5702 2058 5754
rect 3442 5702 3506 5754
rect 559 5313 623 5365
rect 726 5318 790 5370
rect 1151 5319 1215 5371
rect 1994 5306 2058 5358
rect 3442 5306 3506 5358
rect 559 4905 623 4957
rect 726 4900 790 4952
rect 1151 4899 1215 4951
rect 1994 4912 2058 4964
rect 3442 4912 3506 4964
rect 559 4523 623 4575
rect 726 4528 790 4580
rect 1151 4529 1215 4581
rect 1994 4516 2058 4568
rect 3442 4516 3506 4568
rect 559 4115 623 4167
rect 726 4110 790 4162
rect 1151 4109 1215 4161
rect 1994 4122 2058 4174
rect 3442 4122 3506 4174
rect 559 3733 623 3785
rect 726 3738 790 3790
rect 1151 3739 1215 3791
rect 1994 3726 2058 3778
rect 3442 3726 3506 3778
rect 559 3325 623 3377
rect 726 3320 790 3372
rect 1151 3319 1215 3371
rect 1994 3332 2058 3384
rect 3442 3332 3506 3384
rect 559 2943 623 2995
rect 726 2948 790 3000
rect 1151 2949 1215 3001
rect 1994 2936 2058 2988
rect 3442 2936 3506 2988
rect 559 2535 623 2587
rect 726 2530 790 2582
rect 1151 2529 1215 2581
rect 1994 2542 2058 2594
rect 3442 2542 3506 2594
rect 559 2153 623 2205
rect 726 2158 790 2210
rect 1151 2159 1215 2211
rect 1994 2146 2058 2198
rect 3442 2146 3506 2198
rect 559 1745 623 1797
rect 726 1740 790 1792
rect 1151 1739 1215 1791
rect 1994 1752 2058 1804
rect 3442 1752 3506 1804
rect 559 1363 623 1415
rect 726 1368 790 1420
rect 1151 1369 1215 1421
rect 1994 1356 2058 1408
rect 3442 1356 3506 1408
rect 559 955 623 1007
rect 726 950 790 1002
rect 1151 949 1215 1001
rect 1994 962 2058 1014
rect 3442 962 3506 1014
rect 559 573 623 625
rect 726 578 790 630
rect 1151 579 1215 631
rect 1994 566 2058 618
rect 3442 566 3506 618
rect 559 165 623 217
rect 726 160 790 212
rect 1151 159 1215 211
rect 1994 172 2058 224
rect 3442 172 3506 224
<< metal2 >>
rect 577 0 605 25280
rect 730 25070 786 25118
rect 1155 25071 1211 25119
rect 1998 25058 2054 25106
rect 3446 25058 3502 25106
rect 730 24652 786 24700
rect 1155 24651 1211 24699
rect 1998 24663 2054 24711
rect 3446 24663 3502 24711
rect 730 24280 786 24328
rect 1155 24281 1211 24329
rect 1998 24268 2054 24316
rect 3446 24268 3502 24316
rect 730 23862 786 23910
rect 1155 23861 1211 23909
rect 1998 23873 2054 23921
rect 3446 23873 3502 23921
rect 730 23490 786 23538
rect 1155 23491 1211 23539
rect 1998 23478 2054 23526
rect 3446 23478 3502 23526
rect 730 23072 786 23120
rect 1155 23071 1211 23119
rect 1998 23083 2054 23131
rect 3446 23083 3502 23131
rect 730 22700 786 22748
rect 1155 22701 1211 22749
rect 1998 22688 2054 22736
rect 3446 22688 3502 22736
rect 730 22282 786 22330
rect 1155 22281 1211 22329
rect 1998 22293 2054 22341
rect 3446 22293 3502 22341
rect 730 21910 786 21958
rect 1155 21911 1211 21959
rect 1998 21898 2054 21946
rect 3446 21898 3502 21946
rect 730 21492 786 21540
rect 1155 21491 1211 21539
rect 1998 21503 2054 21551
rect 3446 21503 3502 21551
rect 730 21120 786 21168
rect 1155 21121 1211 21169
rect 1998 21108 2054 21156
rect 3446 21108 3502 21156
rect 730 20702 786 20750
rect 1155 20701 1211 20749
rect 1998 20713 2054 20761
rect 3446 20713 3502 20761
rect 730 20330 786 20378
rect 1155 20331 1211 20379
rect 1998 20318 2054 20366
rect 3446 20318 3502 20366
rect 730 19912 786 19960
rect 1155 19911 1211 19959
rect 1998 19923 2054 19971
rect 3446 19923 3502 19971
rect 730 19540 786 19588
rect 1155 19541 1211 19589
rect 1998 19528 2054 19576
rect 3446 19528 3502 19576
rect 730 19122 786 19170
rect 1155 19121 1211 19169
rect 1998 19133 2054 19181
rect 3446 19133 3502 19181
rect 730 18750 786 18798
rect 1155 18751 1211 18799
rect 1998 18738 2054 18786
rect 3446 18738 3502 18786
rect 730 18332 786 18380
rect 1155 18331 1211 18379
rect 1998 18343 2054 18391
rect 3446 18343 3502 18391
rect 730 17960 786 18008
rect 1155 17961 1211 18009
rect 1998 17948 2054 17996
rect 3446 17948 3502 17996
rect 730 17542 786 17590
rect 1155 17541 1211 17589
rect 1998 17553 2054 17601
rect 3446 17553 3502 17601
rect 730 17170 786 17218
rect 1155 17171 1211 17219
rect 1998 17158 2054 17206
rect 3446 17158 3502 17206
rect 730 16752 786 16800
rect 1155 16751 1211 16799
rect 1998 16763 2054 16811
rect 3446 16763 3502 16811
rect 730 16380 786 16428
rect 1155 16381 1211 16429
rect 1998 16368 2054 16416
rect 3446 16368 3502 16416
rect 730 15962 786 16010
rect 1155 15961 1211 16009
rect 1998 15973 2054 16021
rect 3446 15973 3502 16021
rect 730 15590 786 15638
rect 1155 15591 1211 15639
rect 1998 15578 2054 15626
rect 3446 15578 3502 15626
rect 730 15172 786 15220
rect 1155 15171 1211 15219
rect 1998 15183 2054 15231
rect 3446 15183 3502 15231
rect 730 14800 786 14848
rect 1155 14801 1211 14849
rect 1998 14788 2054 14836
rect 3446 14788 3502 14836
rect 730 14382 786 14430
rect 1155 14381 1211 14429
rect 1998 14393 2054 14441
rect 3446 14393 3502 14441
rect 730 14010 786 14058
rect 1155 14011 1211 14059
rect 1998 13998 2054 14046
rect 3446 13998 3502 14046
rect 730 13592 786 13640
rect 1155 13591 1211 13639
rect 1998 13603 2054 13651
rect 3446 13603 3502 13651
rect 730 13220 786 13268
rect 1155 13221 1211 13269
rect 1998 13208 2054 13256
rect 3446 13208 3502 13256
rect 730 12802 786 12850
rect 1155 12801 1211 12849
rect 1998 12813 2054 12861
rect 3446 12813 3502 12861
rect 730 12430 786 12478
rect 1155 12431 1211 12479
rect 1998 12418 2054 12466
rect 3446 12418 3502 12466
rect 730 12012 786 12060
rect 1155 12011 1211 12059
rect 1998 12023 2054 12071
rect 3446 12023 3502 12071
rect 730 11640 786 11688
rect 1155 11641 1211 11689
rect 1998 11628 2054 11676
rect 3446 11628 3502 11676
rect 730 11222 786 11270
rect 1155 11221 1211 11269
rect 1998 11233 2054 11281
rect 3446 11233 3502 11281
rect 730 10850 786 10898
rect 1155 10851 1211 10899
rect 1998 10838 2054 10886
rect 3446 10838 3502 10886
rect 730 10432 786 10480
rect 1155 10431 1211 10479
rect 1998 10443 2054 10491
rect 3446 10443 3502 10491
rect 730 10060 786 10108
rect 1155 10061 1211 10109
rect 1998 10048 2054 10096
rect 3446 10048 3502 10096
rect 730 9642 786 9690
rect 1155 9641 1211 9689
rect 1998 9653 2054 9701
rect 3446 9653 3502 9701
rect 730 9270 786 9318
rect 1155 9271 1211 9319
rect 1998 9258 2054 9306
rect 3446 9258 3502 9306
rect 730 8852 786 8900
rect 1155 8851 1211 8899
rect 1998 8863 2054 8911
rect 3446 8863 3502 8911
rect 730 8480 786 8528
rect 1155 8481 1211 8529
rect 1998 8468 2054 8516
rect 3446 8468 3502 8516
rect 730 8062 786 8110
rect 1155 8061 1211 8109
rect 1998 8073 2054 8121
rect 3446 8073 3502 8121
rect 730 7690 786 7738
rect 1155 7691 1211 7739
rect 1998 7678 2054 7726
rect 3446 7678 3502 7726
rect 730 7272 786 7320
rect 1155 7271 1211 7319
rect 1998 7283 2054 7331
rect 3446 7283 3502 7331
rect 730 6900 786 6948
rect 1155 6901 1211 6949
rect 1998 6888 2054 6936
rect 3446 6888 3502 6936
rect 730 6482 786 6530
rect 1155 6481 1211 6529
rect 1998 6493 2054 6541
rect 3446 6493 3502 6541
rect 730 6110 786 6158
rect 1155 6111 1211 6159
rect 1998 6098 2054 6146
rect 3446 6098 3502 6146
rect 730 5692 786 5740
rect 1155 5691 1211 5739
rect 1998 5703 2054 5751
rect 3446 5703 3502 5751
rect 730 5320 786 5368
rect 1155 5321 1211 5369
rect 1998 5308 2054 5356
rect 3446 5308 3502 5356
rect 730 4902 786 4950
rect 1155 4901 1211 4949
rect 1998 4913 2054 4961
rect 3446 4913 3502 4961
rect 730 4530 786 4578
rect 1155 4531 1211 4579
rect 1998 4518 2054 4566
rect 3446 4518 3502 4566
rect 730 4112 786 4160
rect 1155 4111 1211 4159
rect 1998 4123 2054 4171
rect 3446 4123 3502 4171
rect 730 3740 786 3788
rect 1155 3741 1211 3789
rect 1998 3728 2054 3776
rect 3446 3728 3502 3776
rect 730 3322 786 3370
rect 1155 3321 1211 3369
rect 1998 3333 2054 3381
rect 3446 3333 3502 3381
rect 730 2950 786 2998
rect 1155 2951 1211 2999
rect 1998 2938 2054 2986
rect 3446 2938 3502 2986
rect 730 2532 786 2580
rect 1155 2531 1211 2579
rect 1998 2543 2054 2591
rect 3446 2543 3502 2591
rect 730 2160 786 2208
rect 1155 2161 1211 2209
rect 1998 2148 2054 2196
rect 3446 2148 3502 2196
rect 730 1742 786 1790
rect 1155 1741 1211 1789
rect 1998 1753 2054 1801
rect 3446 1753 3502 1801
rect 730 1370 786 1418
rect 1155 1371 1211 1419
rect 1998 1358 2054 1406
rect 3446 1358 3502 1406
rect 730 952 786 1000
rect 1155 951 1211 999
rect 1998 963 2054 1011
rect 3446 963 3502 1011
rect 730 580 786 628
rect 1155 581 1211 629
rect 1998 568 2054 616
rect 3446 568 3502 616
rect 730 162 786 210
rect 1155 161 1211 209
rect 1998 173 2054 221
rect 3446 173 3502 221
<< metal3 >>
rect 683 25062 833 25126
rect 1108 25063 1258 25127
rect 1951 25050 2101 25114
rect 3399 25050 3549 25114
rect 683 24644 833 24708
rect 1108 24643 1258 24707
rect 1951 24656 2101 24720
rect 3399 24656 3549 24720
rect 683 24272 833 24336
rect 1108 24273 1258 24337
rect 1951 24260 2101 24324
rect 3399 24260 3549 24324
rect 683 23854 833 23918
rect 1108 23853 1258 23917
rect 1951 23866 2101 23930
rect 3399 23866 3549 23930
rect 683 23482 833 23546
rect 1108 23483 1258 23547
rect 1951 23470 2101 23534
rect 3399 23470 3549 23534
rect 683 23064 833 23128
rect 1108 23063 1258 23127
rect 1951 23076 2101 23140
rect 3399 23076 3549 23140
rect 683 22692 833 22756
rect 1108 22693 1258 22757
rect 1951 22680 2101 22744
rect 3399 22680 3549 22744
rect 683 22274 833 22338
rect 1108 22273 1258 22337
rect 1951 22286 2101 22350
rect 3399 22286 3549 22350
rect 683 21902 833 21966
rect 1108 21903 1258 21967
rect 1951 21890 2101 21954
rect 3399 21890 3549 21954
rect 683 21484 833 21548
rect 1108 21483 1258 21547
rect 1951 21496 2101 21560
rect 3399 21496 3549 21560
rect 683 21112 833 21176
rect 1108 21113 1258 21177
rect 1951 21100 2101 21164
rect 3399 21100 3549 21164
rect 683 20694 833 20758
rect 1108 20693 1258 20757
rect 1951 20706 2101 20770
rect 3399 20706 3549 20770
rect 683 20322 833 20386
rect 1108 20323 1258 20387
rect 1951 20310 2101 20374
rect 3399 20310 3549 20374
rect 683 19904 833 19968
rect 1108 19903 1258 19967
rect 1951 19916 2101 19980
rect 3399 19916 3549 19980
rect 683 19532 833 19596
rect 1108 19533 1258 19597
rect 1951 19520 2101 19584
rect 3399 19520 3549 19584
rect 683 19114 833 19178
rect 1108 19113 1258 19177
rect 1951 19126 2101 19190
rect 3399 19126 3549 19190
rect 683 18742 833 18806
rect 1108 18743 1258 18807
rect 1951 18730 2101 18794
rect 3399 18730 3549 18794
rect 683 18324 833 18388
rect 1108 18323 1258 18387
rect 1951 18336 2101 18400
rect 3399 18336 3549 18400
rect 683 17952 833 18016
rect 1108 17953 1258 18017
rect 1951 17940 2101 18004
rect 3399 17940 3549 18004
rect 683 17534 833 17598
rect 1108 17533 1258 17597
rect 1951 17546 2101 17610
rect 3399 17546 3549 17610
rect 683 17162 833 17226
rect 1108 17163 1258 17227
rect 1951 17150 2101 17214
rect 3399 17150 3549 17214
rect 683 16744 833 16808
rect 1108 16743 1258 16807
rect 1951 16756 2101 16820
rect 3399 16756 3549 16820
rect 683 16372 833 16436
rect 1108 16373 1258 16437
rect 1951 16360 2101 16424
rect 3399 16360 3549 16424
rect 683 15954 833 16018
rect 1108 15953 1258 16017
rect 1951 15966 2101 16030
rect 3399 15966 3549 16030
rect 683 15582 833 15646
rect 1108 15583 1258 15647
rect 1951 15570 2101 15634
rect 3399 15570 3549 15634
rect 683 15164 833 15228
rect 1108 15163 1258 15227
rect 1951 15176 2101 15240
rect 3399 15176 3549 15240
rect 683 14792 833 14856
rect 1108 14793 1258 14857
rect 1951 14780 2101 14844
rect 3399 14780 3549 14844
rect 683 14374 833 14438
rect 1108 14373 1258 14437
rect 1951 14386 2101 14450
rect 3399 14386 3549 14450
rect 683 14002 833 14066
rect 1108 14003 1258 14067
rect 1951 13990 2101 14054
rect 3399 13990 3549 14054
rect 683 13584 833 13648
rect 1108 13583 1258 13647
rect 1951 13596 2101 13660
rect 3399 13596 3549 13660
rect 683 13212 833 13276
rect 1108 13213 1258 13277
rect 1951 13200 2101 13264
rect 3399 13200 3549 13264
rect 683 12794 833 12858
rect 1108 12793 1258 12857
rect 1951 12806 2101 12870
rect 3399 12806 3549 12870
rect 683 12422 833 12486
rect 1108 12423 1258 12487
rect 1951 12410 2101 12474
rect 3399 12410 3549 12474
rect 683 12004 833 12068
rect 1108 12003 1258 12067
rect 1951 12016 2101 12080
rect 3399 12016 3549 12080
rect 683 11632 833 11696
rect 1108 11633 1258 11697
rect 1951 11620 2101 11684
rect 3399 11620 3549 11684
rect 683 11214 833 11278
rect 1108 11213 1258 11277
rect 1951 11226 2101 11290
rect 3399 11226 3549 11290
rect 683 10842 833 10906
rect 1108 10843 1258 10907
rect 1951 10830 2101 10894
rect 3399 10830 3549 10894
rect 683 10424 833 10488
rect 1108 10423 1258 10487
rect 1951 10436 2101 10500
rect 3399 10436 3549 10500
rect 683 10052 833 10116
rect 1108 10053 1258 10117
rect 1951 10040 2101 10104
rect 3399 10040 3549 10104
rect 683 9634 833 9698
rect 1108 9633 1258 9697
rect 1951 9646 2101 9710
rect 3399 9646 3549 9710
rect 683 9262 833 9326
rect 1108 9263 1258 9327
rect 1951 9250 2101 9314
rect 3399 9250 3549 9314
rect 683 8844 833 8908
rect 1108 8843 1258 8907
rect 1951 8856 2101 8920
rect 3399 8856 3549 8920
rect 683 8472 833 8536
rect 1108 8473 1258 8537
rect 1951 8460 2101 8524
rect 3399 8460 3549 8524
rect 683 8054 833 8118
rect 1108 8053 1258 8117
rect 1951 8066 2101 8130
rect 3399 8066 3549 8130
rect 683 7682 833 7746
rect 1108 7683 1258 7747
rect 1951 7670 2101 7734
rect 3399 7670 3549 7734
rect 683 7264 833 7328
rect 1108 7263 1258 7327
rect 1951 7276 2101 7340
rect 3399 7276 3549 7340
rect 683 6892 833 6956
rect 1108 6893 1258 6957
rect 1951 6880 2101 6944
rect 3399 6880 3549 6944
rect 683 6474 833 6538
rect 1108 6473 1258 6537
rect 1951 6486 2101 6550
rect 3399 6486 3549 6550
rect 683 6102 833 6166
rect 1108 6103 1258 6167
rect 1951 6090 2101 6154
rect 3399 6090 3549 6154
rect 683 5684 833 5748
rect 1108 5683 1258 5747
rect 1951 5696 2101 5760
rect 3399 5696 3549 5760
rect 683 5312 833 5376
rect 1108 5313 1258 5377
rect 1951 5300 2101 5364
rect 3399 5300 3549 5364
rect 683 4894 833 4958
rect 1108 4893 1258 4957
rect 1951 4906 2101 4970
rect 3399 4906 3549 4970
rect 683 4522 833 4586
rect 1108 4523 1258 4587
rect 1951 4510 2101 4574
rect 3399 4510 3549 4574
rect 683 4104 833 4168
rect 1108 4103 1258 4167
rect 1951 4116 2101 4180
rect 3399 4116 3549 4180
rect 683 3732 833 3796
rect 1108 3733 1258 3797
rect 1951 3720 2101 3784
rect 3399 3720 3549 3784
rect 683 3314 833 3378
rect 1108 3313 1258 3377
rect 1951 3326 2101 3390
rect 3399 3326 3549 3390
rect 683 2942 833 3006
rect 1108 2943 1258 3007
rect 1951 2930 2101 2994
rect 3399 2930 3549 2994
rect 683 2524 833 2588
rect 1108 2523 1258 2587
rect 1951 2536 2101 2600
rect 3399 2536 3549 2600
rect 683 2152 833 2216
rect 1108 2153 1258 2217
rect 1951 2140 2101 2204
rect 3399 2140 3549 2204
rect 683 1734 833 1798
rect 1108 1733 1258 1797
rect 1951 1746 2101 1810
rect 3399 1746 3549 1810
rect 683 1362 833 1426
rect 1108 1363 1258 1427
rect 1951 1350 2101 1414
rect 3399 1350 3549 1414
rect 683 944 833 1008
rect 1108 943 1258 1007
rect 1951 956 2101 1020
rect 3399 956 3549 1020
rect 683 572 833 636
rect 1108 573 1258 637
rect 1951 560 2101 624
rect 3399 560 3549 624
rect 683 154 833 218
rect 1108 153 1258 217
rect 1951 166 2101 230
rect 3399 166 3549 230
<< metal4 >>
rect 725 -63 791 25343
rect 1150 -65 1216 25345
rect 1993 -33 2059 25313
rect 3441 -33 3507 25313
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 562 0 1 25056
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 562 0 1 24648
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_2
timestamp 1661296025
transform 1 0 562 0 1 24266
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_3
timestamp 1661296025
transform 1 0 562 0 1 23858
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_4
timestamp 1661296025
transform 1 0 562 0 1 23476
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_5
timestamp 1661296025
transform 1 0 562 0 1 23068
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_6
timestamp 1661296025
transform 1 0 562 0 1 22686
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_7
timestamp 1661296025
transform 1 0 562 0 1 22278
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_8
timestamp 1661296025
transform 1 0 562 0 1 21896
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_9
timestamp 1661296025
transform 1 0 562 0 1 21488
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_10
timestamp 1661296025
transform 1 0 562 0 1 21106
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_11
timestamp 1661296025
transform 1 0 562 0 1 20698
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_12
timestamp 1661296025
transform 1 0 562 0 1 20316
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_13
timestamp 1661296025
transform 1 0 562 0 1 19908
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_14
timestamp 1661296025
transform 1 0 562 0 1 19526
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_15
timestamp 1661296025
transform 1 0 562 0 1 19118
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_16
timestamp 1661296025
transform 1 0 562 0 1 18736
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_17
timestamp 1661296025
transform 1 0 562 0 1 18328
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_18
timestamp 1661296025
transform 1 0 562 0 1 17946
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_19
timestamp 1661296025
transform 1 0 562 0 1 17538
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_20
timestamp 1661296025
transform 1 0 562 0 1 17156
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_21
timestamp 1661296025
transform 1 0 562 0 1 16748
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_22
timestamp 1661296025
transform 1 0 562 0 1 16366
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_23
timestamp 1661296025
transform 1 0 562 0 1 15958
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_24
timestamp 1661296025
transform 1 0 562 0 1 15576
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_25
timestamp 1661296025
transform 1 0 562 0 1 15168
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_26
timestamp 1661296025
transform 1 0 562 0 1 14786
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_27
timestamp 1661296025
transform 1 0 562 0 1 14378
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_28
timestamp 1661296025
transform 1 0 562 0 1 13996
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_29
timestamp 1661296025
transform 1 0 562 0 1 13588
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_30
timestamp 1661296025
transform 1 0 562 0 1 13206
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_31
timestamp 1661296025
transform 1 0 562 0 1 12798
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_32
timestamp 1661296025
transform 1 0 562 0 1 12416
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_33
timestamp 1661296025
transform 1 0 562 0 1 12008
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_34
timestamp 1661296025
transform 1 0 562 0 1 11626
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_35
timestamp 1661296025
transform 1 0 562 0 1 11218
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_36
timestamp 1661296025
transform 1 0 562 0 1 10836
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_37
timestamp 1661296025
transform 1 0 562 0 1 10428
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_38
timestamp 1661296025
transform 1 0 562 0 1 10046
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_39
timestamp 1661296025
transform 1 0 562 0 1 9638
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_40
timestamp 1661296025
transform 1 0 562 0 1 9256
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_41
timestamp 1661296025
transform 1 0 562 0 1 8848
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_42
timestamp 1661296025
transform 1 0 562 0 1 8466
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_43
timestamp 1661296025
transform 1 0 562 0 1 8058
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_44
timestamp 1661296025
transform 1 0 562 0 1 7676
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_45
timestamp 1661296025
transform 1 0 562 0 1 7268
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_46
timestamp 1661296025
transform 1 0 562 0 1 6886
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_47
timestamp 1661296025
transform 1 0 562 0 1 6478
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_48
timestamp 1661296025
transform 1 0 562 0 1 6096
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_49
timestamp 1661296025
transform 1 0 562 0 1 5688
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_50
timestamp 1661296025
transform 1 0 562 0 1 5306
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_51
timestamp 1661296025
transform 1 0 562 0 1 4898
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_52
timestamp 1661296025
transform 1 0 562 0 1 4516
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_53
timestamp 1661296025
transform 1 0 562 0 1 4108
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_54
timestamp 1661296025
transform 1 0 562 0 1 3726
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_55
timestamp 1661296025
transform 1 0 562 0 1 3318
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_56
timestamp 1661296025
transform 1 0 562 0 1 2936
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_57
timestamp 1661296025
transform 1 0 562 0 1 2528
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_58
timestamp 1661296025
transform 1 0 562 0 1 2146
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_59
timestamp 1661296025
transform 1 0 562 0 1 1738
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_60
timestamp 1661296025
transform 1 0 562 0 1 1356
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_61
timestamp 1661296025
transform 1 0 562 0 1 948
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_62
timestamp 1661296025
transform 1 0 562 0 1 566
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_63
timestamp 1661296025
transform 1 0 562 0 1 158
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_0
timestamp 1661296025
transform 1 0 726 0 1 25062
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_1
timestamp 1661296025
transform 1 0 726 0 1 24644
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_2
timestamp 1661296025
transform 1 0 726 0 1 24272
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_3
timestamp 1661296025
transform 1 0 726 0 1 23854
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_4
timestamp 1661296025
transform 1 0 726 0 1 23482
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_5
timestamp 1661296025
transform 1 0 726 0 1 23064
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_6
timestamp 1661296025
transform 1 0 726 0 1 22692
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_7
timestamp 1661296025
transform 1 0 726 0 1 22274
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_8
timestamp 1661296025
transform 1 0 726 0 1 21902
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_9
timestamp 1661296025
transform 1 0 726 0 1 21484
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_10
timestamp 1661296025
transform 1 0 726 0 1 21112
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_11
timestamp 1661296025
transform 1 0 726 0 1 20694
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_12
timestamp 1661296025
transform 1 0 726 0 1 20322
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_13
timestamp 1661296025
transform 1 0 726 0 1 19904
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_14
timestamp 1661296025
transform 1 0 726 0 1 19532
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_15
timestamp 1661296025
transform 1 0 726 0 1 19114
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_16
timestamp 1661296025
transform 1 0 726 0 1 18742
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_17
timestamp 1661296025
transform 1 0 726 0 1 18324
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_18
timestamp 1661296025
transform 1 0 726 0 1 17952
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_19
timestamp 1661296025
transform 1 0 726 0 1 17534
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_20
timestamp 1661296025
transform 1 0 726 0 1 17162
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_21
timestamp 1661296025
transform 1 0 726 0 1 16744
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_22
timestamp 1661296025
transform 1 0 726 0 1 16372
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_23
timestamp 1661296025
transform 1 0 726 0 1 15954
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_24
timestamp 1661296025
transform 1 0 726 0 1 15582
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_25
timestamp 1661296025
transform 1 0 726 0 1 15164
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_26
timestamp 1661296025
transform 1 0 726 0 1 14792
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_27
timestamp 1661296025
transform 1 0 726 0 1 14374
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_28
timestamp 1661296025
transform 1 0 726 0 1 14002
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_29
timestamp 1661296025
transform 1 0 726 0 1 13584
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_30
timestamp 1661296025
transform 1 0 726 0 1 13212
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_31
timestamp 1661296025
transform 1 0 726 0 1 12794
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_32
timestamp 1661296025
transform 1 0 726 0 1 12422
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_33
timestamp 1661296025
transform 1 0 726 0 1 12004
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_34
timestamp 1661296025
transform 1 0 726 0 1 11632
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_35
timestamp 1661296025
transform 1 0 726 0 1 11214
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_36
timestamp 1661296025
transform 1 0 726 0 1 10842
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_37
timestamp 1661296025
transform 1 0 726 0 1 10424
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_38
timestamp 1661296025
transform 1 0 726 0 1 10052
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_39
timestamp 1661296025
transform 1 0 726 0 1 9634
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_40
timestamp 1661296025
transform 1 0 726 0 1 9262
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_41
timestamp 1661296025
transform 1 0 726 0 1 8844
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_42
timestamp 1661296025
transform 1 0 726 0 1 8472
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_43
timestamp 1661296025
transform 1 0 726 0 1 8054
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_44
timestamp 1661296025
transform 1 0 726 0 1 7682
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_45
timestamp 1661296025
transform 1 0 726 0 1 7264
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_46
timestamp 1661296025
transform 1 0 726 0 1 6892
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_47
timestamp 1661296025
transform 1 0 726 0 1 6474
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_48
timestamp 1661296025
transform 1 0 726 0 1 6102
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_49
timestamp 1661296025
transform 1 0 726 0 1 5684
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_50
timestamp 1661296025
transform 1 0 726 0 1 5312
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_51
timestamp 1661296025
transform 1 0 726 0 1 4894
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_52
timestamp 1661296025
transform 1 0 726 0 1 4522
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_53
timestamp 1661296025
transform 1 0 726 0 1 4104
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_54
timestamp 1661296025
transform 1 0 726 0 1 3732
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_55
timestamp 1661296025
transform 1 0 726 0 1 3314
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_56
timestamp 1661296025
transform 1 0 726 0 1 2942
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_57
timestamp 1661296025
transform 1 0 726 0 1 2524
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_58
timestamp 1661296025
transform 1 0 726 0 1 2152
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_59
timestamp 1661296025
transform 1 0 726 0 1 1734
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_60
timestamp 1661296025
transform 1 0 726 0 1 1362
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_61
timestamp 1661296025
transform 1 0 726 0 1 944
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_62
timestamp 1661296025
transform 1 0 726 0 1 572
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_63
timestamp 1661296025
transform 1 0 726 0 1 154
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_64
timestamp 1661296025
transform 1 0 1994 0 1 25050
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_65
timestamp 1661296025
transform 1 0 1994 0 1 24656
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_66
timestamp 1661296025
transform 1 0 1994 0 1 24260
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_67
timestamp 1661296025
transform 1 0 1994 0 1 23866
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_68
timestamp 1661296025
transform 1 0 1994 0 1 23470
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_69
timestamp 1661296025
transform 1 0 1994 0 1 23076
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_70
timestamp 1661296025
transform 1 0 1994 0 1 22680
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_71
timestamp 1661296025
transform 1 0 1994 0 1 22286
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_72
timestamp 1661296025
transform 1 0 1994 0 1 21890
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_73
timestamp 1661296025
transform 1 0 1994 0 1 21496
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_74
timestamp 1661296025
transform 1 0 1994 0 1 21100
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_75
timestamp 1661296025
transform 1 0 1994 0 1 20706
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_76
timestamp 1661296025
transform 1 0 1994 0 1 20310
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_77
timestamp 1661296025
transform 1 0 1994 0 1 19916
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_78
timestamp 1661296025
transform 1 0 1994 0 1 19520
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_79
timestamp 1661296025
transform 1 0 1994 0 1 19126
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_80
timestamp 1661296025
transform 1 0 1994 0 1 18730
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_81
timestamp 1661296025
transform 1 0 1994 0 1 18336
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_82
timestamp 1661296025
transform 1 0 1994 0 1 17940
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_83
timestamp 1661296025
transform 1 0 1994 0 1 17546
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_84
timestamp 1661296025
transform 1 0 1994 0 1 17150
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_85
timestamp 1661296025
transform 1 0 1994 0 1 16756
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_86
timestamp 1661296025
transform 1 0 1994 0 1 16360
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_87
timestamp 1661296025
transform 1 0 1994 0 1 15966
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_88
timestamp 1661296025
transform 1 0 1994 0 1 15570
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_89
timestamp 1661296025
transform 1 0 1994 0 1 15176
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_90
timestamp 1661296025
transform 1 0 1994 0 1 14780
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_91
timestamp 1661296025
transform 1 0 1994 0 1 14386
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_92
timestamp 1661296025
transform 1 0 1994 0 1 13990
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_93
timestamp 1661296025
transform 1 0 1994 0 1 13596
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_94
timestamp 1661296025
transform 1 0 1994 0 1 13200
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_95
timestamp 1661296025
transform 1 0 1994 0 1 12806
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_96
timestamp 1661296025
transform 1 0 1994 0 1 12410
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_97
timestamp 1661296025
transform 1 0 1994 0 1 12016
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_98
timestamp 1661296025
transform 1 0 1994 0 1 11620
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_99
timestamp 1661296025
transform 1 0 1994 0 1 11226
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_100
timestamp 1661296025
transform 1 0 1994 0 1 10830
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_101
timestamp 1661296025
transform 1 0 1994 0 1 10436
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_102
timestamp 1661296025
transform 1 0 1994 0 1 10040
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_103
timestamp 1661296025
transform 1 0 1994 0 1 9646
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_104
timestamp 1661296025
transform 1 0 1994 0 1 9250
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_105
timestamp 1661296025
transform 1 0 1994 0 1 8856
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_106
timestamp 1661296025
transform 1 0 1994 0 1 8460
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_107
timestamp 1661296025
transform 1 0 1994 0 1 8066
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_108
timestamp 1661296025
transform 1 0 1994 0 1 7670
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_109
timestamp 1661296025
transform 1 0 1994 0 1 7276
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_110
timestamp 1661296025
transform 1 0 1994 0 1 6880
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_111
timestamp 1661296025
transform 1 0 1994 0 1 6486
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_112
timestamp 1661296025
transform 1 0 1994 0 1 6090
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_113
timestamp 1661296025
transform 1 0 1994 0 1 5696
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_114
timestamp 1661296025
transform 1 0 1994 0 1 5300
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_115
timestamp 1661296025
transform 1 0 1994 0 1 4906
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_116
timestamp 1661296025
transform 1 0 1994 0 1 4510
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_117
timestamp 1661296025
transform 1 0 1994 0 1 4116
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_118
timestamp 1661296025
transform 1 0 1994 0 1 3720
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_119
timestamp 1661296025
transform 1 0 1994 0 1 3326
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_120
timestamp 1661296025
transform 1 0 1994 0 1 2930
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_121
timestamp 1661296025
transform 1 0 1994 0 1 2536
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_122
timestamp 1661296025
transform 1 0 1994 0 1 2140
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_123
timestamp 1661296025
transform 1 0 1994 0 1 1746
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_124
timestamp 1661296025
transform 1 0 1994 0 1 1350
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_125
timestamp 1661296025
transform 1 0 1994 0 1 956
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_126
timestamp 1661296025
transform 1 0 1994 0 1 560
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_127
timestamp 1661296025
transform 1 0 1994 0 1 166
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_128
timestamp 1661296025
transform 1 0 3442 0 1 25050
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_129
timestamp 1661296025
transform 1 0 3442 0 1 24656
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_130
timestamp 1661296025
transform 1 0 3442 0 1 24260
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_131
timestamp 1661296025
transform 1 0 3442 0 1 23866
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_132
timestamp 1661296025
transform 1 0 3442 0 1 23470
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_133
timestamp 1661296025
transform 1 0 3442 0 1 23076
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_134
timestamp 1661296025
transform 1 0 3442 0 1 22680
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_135
timestamp 1661296025
transform 1 0 3442 0 1 22286
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_136
timestamp 1661296025
transform 1 0 3442 0 1 21890
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_137
timestamp 1661296025
transform 1 0 3442 0 1 21496
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_138
timestamp 1661296025
transform 1 0 3442 0 1 21100
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_139
timestamp 1661296025
transform 1 0 3442 0 1 20706
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_140
timestamp 1661296025
transform 1 0 3442 0 1 20310
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_141
timestamp 1661296025
transform 1 0 3442 0 1 19916
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_142
timestamp 1661296025
transform 1 0 3442 0 1 19520
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_143
timestamp 1661296025
transform 1 0 3442 0 1 19126
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_144
timestamp 1661296025
transform 1 0 3442 0 1 18730
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_145
timestamp 1661296025
transform 1 0 3442 0 1 18336
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_146
timestamp 1661296025
transform 1 0 3442 0 1 17940
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_147
timestamp 1661296025
transform 1 0 3442 0 1 17546
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_148
timestamp 1661296025
transform 1 0 3442 0 1 17150
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_149
timestamp 1661296025
transform 1 0 3442 0 1 16756
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_150
timestamp 1661296025
transform 1 0 3442 0 1 16360
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_151
timestamp 1661296025
transform 1 0 3442 0 1 15966
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_152
timestamp 1661296025
transform 1 0 3442 0 1 15570
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_153
timestamp 1661296025
transform 1 0 3442 0 1 15176
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_154
timestamp 1661296025
transform 1 0 3442 0 1 14780
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_155
timestamp 1661296025
transform 1 0 3442 0 1 14386
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_156
timestamp 1661296025
transform 1 0 3442 0 1 13990
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_157
timestamp 1661296025
transform 1 0 3442 0 1 13596
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_158
timestamp 1661296025
transform 1 0 3442 0 1 13200
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_159
timestamp 1661296025
transform 1 0 3442 0 1 12806
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_160
timestamp 1661296025
transform 1 0 3442 0 1 12410
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_161
timestamp 1661296025
transform 1 0 3442 0 1 12016
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_162
timestamp 1661296025
transform 1 0 3442 0 1 11620
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_163
timestamp 1661296025
transform 1 0 3442 0 1 11226
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_164
timestamp 1661296025
transform 1 0 3442 0 1 10830
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_165
timestamp 1661296025
transform 1 0 3442 0 1 10436
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_166
timestamp 1661296025
transform 1 0 3442 0 1 10040
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_167
timestamp 1661296025
transform 1 0 3442 0 1 9646
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_168
timestamp 1661296025
transform 1 0 3442 0 1 9250
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_169
timestamp 1661296025
transform 1 0 3442 0 1 8856
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_170
timestamp 1661296025
transform 1 0 3442 0 1 8460
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_171
timestamp 1661296025
transform 1 0 3442 0 1 8066
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_172
timestamp 1661296025
transform 1 0 3442 0 1 7670
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_173
timestamp 1661296025
transform 1 0 3442 0 1 7276
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_174
timestamp 1661296025
transform 1 0 3442 0 1 6880
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_175
timestamp 1661296025
transform 1 0 3442 0 1 6486
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_176
timestamp 1661296025
transform 1 0 3442 0 1 6090
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_177
timestamp 1661296025
transform 1 0 3442 0 1 5696
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_178
timestamp 1661296025
transform 1 0 3442 0 1 5300
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_179
timestamp 1661296025
transform 1 0 3442 0 1 4906
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_180
timestamp 1661296025
transform 1 0 3442 0 1 4510
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_181
timestamp 1661296025
transform 1 0 3442 0 1 4116
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_182
timestamp 1661296025
transform 1 0 3442 0 1 3720
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_183
timestamp 1661296025
transform 1 0 3442 0 1 3326
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_184
timestamp 1661296025
transform 1 0 3442 0 1 2930
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_185
timestamp 1661296025
transform 1 0 3442 0 1 2536
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_186
timestamp 1661296025
transform 1 0 3442 0 1 2140
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_187
timestamp 1661296025
transform 1 0 3442 0 1 1746
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_188
timestamp 1661296025
transform 1 0 3442 0 1 1350
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_189
timestamp 1661296025
transform 1 0 3442 0 1 956
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_190
timestamp 1661296025
transform 1 0 3442 0 1 560
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_191
timestamp 1661296025
transform 1 0 3442 0 1 166
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_192
timestamp 1661296025
transform 1 0 1151 0 1 25063
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_193
timestamp 1661296025
transform 1 0 1151 0 1 24643
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_194
timestamp 1661296025
transform 1 0 1151 0 1 24273
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_195
timestamp 1661296025
transform 1 0 1151 0 1 23853
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_196
timestamp 1661296025
transform 1 0 1151 0 1 23483
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_197
timestamp 1661296025
transform 1 0 1151 0 1 23063
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_198
timestamp 1661296025
transform 1 0 1151 0 1 22693
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_199
timestamp 1661296025
transform 1 0 1151 0 1 22273
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_200
timestamp 1661296025
transform 1 0 1151 0 1 21903
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_201
timestamp 1661296025
transform 1 0 1151 0 1 21483
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_202
timestamp 1661296025
transform 1 0 1151 0 1 21113
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_203
timestamp 1661296025
transform 1 0 1151 0 1 20693
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_204
timestamp 1661296025
transform 1 0 1151 0 1 20323
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_205
timestamp 1661296025
transform 1 0 1151 0 1 19903
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_206
timestamp 1661296025
transform 1 0 1151 0 1 19533
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_207
timestamp 1661296025
transform 1 0 1151 0 1 19113
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_208
timestamp 1661296025
transform 1 0 1151 0 1 18743
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_209
timestamp 1661296025
transform 1 0 1151 0 1 18323
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_210
timestamp 1661296025
transform 1 0 1151 0 1 17953
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_211
timestamp 1661296025
transform 1 0 1151 0 1 17533
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_212
timestamp 1661296025
transform 1 0 1151 0 1 17163
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_213
timestamp 1661296025
transform 1 0 1151 0 1 16743
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_214
timestamp 1661296025
transform 1 0 1151 0 1 16373
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_215
timestamp 1661296025
transform 1 0 1151 0 1 15953
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_216
timestamp 1661296025
transform 1 0 1151 0 1 15583
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_217
timestamp 1661296025
transform 1 0 1151 0 1 15163
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_218
timestamp 1661296025
transform 1 0 1151 0 1 14793
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_219
timestamp 1661296025
transform 1 0 1151 0 1 14373
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_220
timestamp 1661296025
transform 1 0 1151 0 1 14003
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_221
timestamp 1661296025
transform 1 0 1151 0 1 13583
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_222
timestamp 1661296025
transform 1 0 1151 0 1 13213
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_223
timestamp 1661296025
transform 1 0 1151 0 1 12793
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_224
timestamp 1661296025
transform 1 0 1151 0 1 12423
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_225
timestamp 1661296025
transform 1 0 1151 0 1 12003
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_226
timestamp 1661296025
transform 1 0 1151 0 1 11633
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_227
timestamp 1661296025
transform 1 0 1151 0 1 11213
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_228
timestamp 1661296025
transform 1 0 1151 0 1 10843
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_229
timestamp 1661296025
transform 1 0 1151 0 1 10423
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_230
timestamp 1661296025
transform 1 0 1151 0 1 10053
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_231
timestamp 1661296025
transform 1 0 1151 0 1 9633
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_232
timestamp 1661296025
transform 1 0 1151 0 1 9263
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_233
timestamp 1661296025
transform 1 0 1151 0 1 8843
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_234
timestamp 1661296025
transform 1 0 1151 0 1 8473
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_235
timestamp 1661296025
transform 1 0 1151 0 1 8053
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_236
timestamp 1661296025
transform 1 0 1151 0 1 7683
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_237
timestamp 1661296025
transform 1 0 1151 0 1 7263
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_238
timestamp 1661296025
transform 1 0 1151 0 1 6893
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_239
timestamp 1661296025
transform 1 0 1151 0 1 6473
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_240
timestamp 1661296025
transform 1 0 1151 0 1 6103
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_241
timestamp 1661296025
transform 1 0 1151 0 1 5683
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_242
timestamp 1661296025
transform 1 0 1151 0 1 5313
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_243
timestamp 1661296025
transform 1 0 1151 0 1 4893
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_244
timestamp 1661296025
transform 1 0 1151 0 1 4523
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_245
timestamp 1661296025
transform 1 0 1151 0 1 4103
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_246
timestamp 1661296025
transform 1 0 1151 0 1 3733
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_247
timestamp 1661296025
transform 1 0 1151 0 1 3313
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_248
timestamp 1661296025
transform 1 0 1151 0 1 2943
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_249
timestamp 1661296025
transform 1 0 1151 0 1 2523
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_250
timestamp 1661296025
transform 1 0 1151 0 1 2153
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_251
timestamp 1661296025
transform 1 0 1151 0 1 1733
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_252
timestamp 1661296025
transform 1 0 1151 0 1 1363
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_253
timestamp 1661296025
transform 1 0 1151 0 1 943
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_254
timestamp 1661296025
transform 1 0 1151 0 1 573
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_255
timestamp 1661296025
transform 1 0 1151 0 1 153
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_256
timestamp 1661296025
transform 1 0 559 0 1 25057
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_257
timestamp 1661296025
transform 1 0 559 0 1 24649
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_258
timestamp 1661296025
transform 1 0 559 0 1 24267
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_259
timestamp 1661296025
transform 1 0 559 0 1 23859
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_260
timestamp 1661296025
transform 1 0 559 0 1 23477
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_261
timestamp 1661296025
transform 1 0 559 0 1 23069
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_262
timestamp 1661296025
transform 1 0 559 0 1 22687
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_263
timestamp 1661296025
transform 1 0 559 0 1 22279
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_264
timestamp 1661296025
transform 1 0 559 0 1 21897
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_265
timestamp 1661296025
transform 1 0 559 0 1 21489
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_266
timestamp 1661296025
transform 1 0 559 0 1 21107
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_267
timestamp 1661296025
transform 1 0 559 0 1 20699
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_268
timestamp 1661296025
transform 1 0 559 0 1 20317
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_269
timestamp 1661296025
transform 1 0 559 0 1 19909
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_270
timestamp 1661296025
transform 1 0 559 0 1 19527
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_271
timestamp 1661296025
transform 1 0 559 0 1 19119
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_272
timestamp 1661296025
transform 1 0 559 0 1 18737
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_273
timestamp 1661296025
transform 1 0 559 0 1 18329
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_274
timestamp 1661296025
transform 1 0 559 0 1 17947
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_275
timestamp 1661296025
transform 1 0 559 0 1 17539
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_276
timestamp 1661296025
transform 1 0 559 0 1 17157
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_277
timestamp 1661296025
transform 1 0 559 0 1 16749
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_278
timestamp 1661296025
transform 1 0 559 0 1 16367
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_279
timestamp 1661296025
transform 1 0 559 0 1 15959
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_280
timestamp 1661296025
transform 1 0 559 0 1 15577
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_281
timestamp 1661296025
transform 1 0 559 0 1 15169
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_282
timestamp 1661296025
transform 1 0 559 0 1 14787
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_283
timestamp 1661296025
transform 1 0 559 0 1 14379
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_284
timestamp 1661296025
transform 1 0 559 0 1 13997
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_285
timestamp 1661296025
transform 1 0 559 0 1 13589
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_286
timestamp 1661296025
transform 1 0 559 0 1 13207
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_287
timestamp 1661296025
transform 1 0 559 0 1 12799
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_288
timestamp 1661296025
transform 1 0 559 0 1 12417
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_289
timestamp 1661296025
transform 1 0 559 0 1 12009
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_290
timestamp 1661296025
transform 1 0 559 0 1 11627
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_291
timestamp 1661296025
transform 1 0 559 0 1 11219
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_292
timestamp 1661296025
transform 1 0 559 0 1 10837
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_293
timestamp 1661296025
transform 1 0 559 0 1 10429
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_294
timestamp 1661296025
transform 1 0 559 0 1 10047
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_295
timestamp 1661296025
transform 1 0 559 0 1 9639
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_296
timestamp 1661296025
transform 1 0 559 0 1 9257
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_297
timestamp 1661296025
transform 1 0 559 0 1 8849
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_298
timestamp 1661296025
transform 1 0 559 0 1 8467
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_299
timestamp 1661296025
transform 1 0 559 0 1 8059
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_300
timestamp 1661296025
transform 1 0 559 0 1 7677
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_301
timestamp 1661296025
transform 1 0 559 0 1 7269
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_302
timestamp 1661296025
transform 1 0 559 0 1 6887
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_303
timestamp 1661296025
transform 1 0 559 0 1 6479
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_304
timestamp 1661296025
transform 1 0 559 0 1 6097
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_305
timestamp 1661296025
transform 1 0 559 0 1 5689
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_306
timestamp 1661296025
transform 1 0 559 0 1 5307
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_307
timestamp 1661296025
transform 1 0 559 0 1 4899
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_308
timestamp 1661296025
transform 1 0 559 0 1 4517
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_309
timestamp 1661296025
transform 1 0 559 0 1 4109
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_310
timestamp 1661296025
transform 1 0 559 0 1 3727
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_311
timestamp 1661296025
transform 1 0 559 0 1 3319
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_312
timestamp 1661296025
transform 1 0 559 0 1 2937
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_313
timestamp 1661296025
transform 1 0 559 0 1 2529
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_314
timestamp 1661296025
transform 1 0 559 0 1 2147
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_315
timestamp 1661296025
transform 1 0 559 0 1 1739
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_316
timestamp 1661296025
transform 1 0 559 0 1 1357
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_317
timestamp 1661296025
transform 1 0 559 0 1 949
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_318
timestamp 1661296025
transform 1 0 559 0 1 567
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_319
timestamp 1661296025
transform 1 0 559 0 1 159
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_0
timestamp 1661296025
transform 1 0 725 0 1 25057
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_1
timestamp 1661296025
transform 1 0 725 0 1 24639
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_2
timestamp 1661296025
transform 1 0 725 0 1 24267
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_3
timestamp 1661296025
transform 1 0 725 0 1 23849
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_4
timestamp 1661296025
transform 1 0 725 0 1 23477
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_5
timestamp 1661296025
transform 1 0 725 0 1 23059
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_6
timestamp 1661296025
transform 1 0 725 0 1 22687
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_7
timestamp 1661296025
transform 1 0 725 0 1 22269
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_8
timestamp 1661296025
transform 1 0 725 0 1 21897
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_9
timestamp 1661296025
transform 1 0 725 0 1 21479
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_10
timestamp 1661296025
transform 1 0 725 0 1 21107
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_11
timestamp 1661296025
transform 1 0 725 0 1 20689
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_12
timestamp 1661296025
transform 1 0 725 0 1 20317
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_13
timestamp 1661296025
transform 1 0 725 0 1 19899
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_14
timestamp 1661296025
transform 1 0 725 0 1 19527
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_15
timestamp 1661296025
transform 1 0 725 0 1 19109
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_16
timestamp 1661296025
transform 1 0 725 0 1 18737
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_17
timestamp 1661296025
transform 1 0 725 0 1 18319
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_18
timestamp 1661296025
transform 1 0 725 0 1 17947
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_19
timestamp 1661296025
transform 1 0 725 0 1 17529
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_20
timestamp 1661296025
transform 1 0 725 0 1 17157
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_21
timestamp 1661296025
transform 1 0 725 0 1 16739
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_22
timestamp 1661296025
transform 1 0 725 0 1 16367
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_23
timestamp 1661296025
transform 1 0 725 0 1 15949
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_24
timestamp 1661296025
transform 1 0 725 0 1 15577
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_25
timestamp 1661296025
transform 1 0 725 0 1 15159
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_26
timestamp 1661296025
transform 1 0 725 0 1 14787
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_27
timestamp 1661296025
transform 1 0 725 0 1 14369
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_28
timestamp 1661296025
transform 1 0 725 0 1 13997
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_29
timestamp 1661296025
transform 1 0 725 0 1 13579
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_30
timestamp 1661296025
transform 1 0 725 0 1 13207
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_31
timestamp 1661296025
transform 1 0 725 0 1 12789
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_32
timestamp 1661296025
transform 1 0 725 0 1 12417
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_33
timestamp 1661296025
transform 1 0 725 0 1 11999
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_34
timestamp 1661296025
transform 1 0 725 0 1 11627
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_35
timestamp 1661296025
transform 1 0 725 0 1 11209
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_36
timestamp 1661296025
transform 1 0 725 0 1 10837
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_37
timestamp 1661296025
transform 1 0 725 0 1 10419
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_38
timestamp 1661296025
transform 1 0 725 0 1 10047
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_39
timestamp 1661296025
transform 1 0 725 0 1 9629
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_40
timestamp 1661296025
transform 1 0 725 0 1 9257
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_41
timestamp 1661296025
transform 1 0 725 0 1 8839
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_42
timestamp 1661296025
transform 1 0 725 0 1 8467
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_43
timestamp 1661296025
transform 1 0 725 0 1 8049
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_44
timestamp 1661296025
transform 1 0 725 0 1 7677
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_45
timestamp 1661296025
transform 1 0 725 0 1 7259
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_46
timestamp 1661296025
transform 1 0 725 0 1 6887
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_47
timestamp 1661296025
transform 1 0 725 0 1 6469
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_48
timestamp 1661296025
transform 1 0 725 0 1 6097
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_49
timestamp 1661296025
transform 1 0 725 0 1 5679
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_50
timestamp 1661296025
transform 1 0 725 0 1 5307
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_51
timestamp 1661296025
transform 1 0 725 0 1 4889
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_52
timestamp 1661296025
transform 1 0 725 0 1 4517
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_53
timestamp 1661296025
transform 1 0 725 0 1 4099
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_54
timestamp 1661296025
transform 1 0 725 0 1 3727
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_55
timestamp 1661296025
transform 1 0 725 0 1 3309
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_56
timestamp 1661296025
transform 1 0 725 0 1 2937
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_57
timestamp 1661296025
transform 1 0 725 0 1 2519
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_58
timestamp 1661296025
transform 1 0 725 0 1 2147
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_59
timestamp 1661296025
transform 1 0 725 0 1 1729
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_60
timestamp 1661296025
transform 1 0 725 0 1 1357
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_61
timestamp 1661296025
transform 1 0 725 0 1 939
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_62
timestamp 1661296025
transform 1 0 725 0 1 567
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_63
timestamp 1661296025
transform 1 0 725 0 1 149
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_64
timestamp 1661296025
transform 1 0 1993 0 1 25046
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_65
timestamp 1661296025
transform 1 0 1993 0 1 24650
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_66
timestamp 1661296025
transform 1 0 1993 0 1 24256
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_67
timestamp 1661296025
transform 1 0 1993 0 1 23860
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_68
timestamp 1661296025
transform 1 0 1993 0 1 23466
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_69
timestamp 1661296025
transform 1 0 1993 0 1 23070
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_70
timestamp 1661296025
transform 1 0 1993 0 1 22676
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_71
timestamp 1661296025
transform 1 0 1993 0 1 22280
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_72
timestamp 1661296025
transform 1 0 1993 0 1 21886
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_73
timestamp 1661296025
transform 1 0 1993 0 1 21490
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_74
timestamp 1661296025
transform 1 0 1993 0 1 21096
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_75
timestamp 1661296025
transform 1 0 1993 0 1 20700
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_76
timestamp 1661296025
transform 1 0 1993 0 1 20306
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_77
timestamp 1661296025
transform 1 0 1993 0 1 19910
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_78
timestamp 1661296025
transform 1 0 1993 0 1 19516
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_79
timestamp 1661296025
transform 1 0 1993 0 1 19120
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_80
timestamp 1661296025
transform 1 0 1993 0 1 18726
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_81
timestamp 1661296025
transform 1 0 1993 0 1 18330
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_82
timestamp 1661296025
transform 1 0 1993 0 1 17936
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_83
timestamp 1661296025
transform 1 0 1993 0 1 17540
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_84
timestamp 1661296025
transform 1 0 1993 0 1 17146
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_85
timestamp 1661296025
transform 1 0 1993 0 1 16750
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_86
timestamp 1661296025
transform 1 0 1993 0 1 16356
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_87
timestamp 1661296025
transform 1 0 1993 0 1 15960
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_88
timestamp 1661296025
transform 1 0 1993 0 1 15566
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_89
timestamp 1661296025
transform 1 0 1993 0 1 15170
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_90
timestamp 1661296025
transform 1 0 1993 0 1 14776
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_91
timestamp 1661296025
transform 1 0 1993 0 1 14380
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_92
timestamp 1661296025
transform 1 0 1993 0 1 13986
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_93
timestamp 1661296025
transform 1 0 1993 0 1 13590
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_94
timestamp 1661296025
transform 1 0 1993 0 1 13196
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_95
timestamp 1661296025
transform 1 0 1993 0 1 12800
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_96
timestamp 1661296025
transform 1 0 1993 0 1 12406
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_97
timestamp 1661296025
transform 1 0 1993 0 1 12010
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_98
timestamp 1661296025
transform 1 0 1993 0 1 11616
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_99
timestamp 1661296025
transform 1 0 1993 0 1 11220
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_100
timestamp 1661296025
transform 1 0 1993 0 1 10826
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_101
timestamp 1661296025
transform 1 0 1993 0 1 10430
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_102
timestamp 1661296025
transform 1 0 1993 0 1 10036
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_103
timestamp 1661296025
transform 1 0 1993 0 1 9640
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_104
timestamp 1661296025
transform 1 0 1993 0 1 9246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_105
timestamp 1661296025
transform 1 0 1993 0 1 8850
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_106
timestamp 1661296025
transform 1 0 1993 0 1 8456
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_107
timestamp 1661296025
transform 1 0 1993 0 1 8060
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_108
timestamp 1661296025
transform 1 0 1993 0 1 7666
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_109
timestamp 1661296025
transform 1 0 1993 0 1 7270
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_110
timestamp 1661296025
transform 1 0 1993 0 1 6876
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_111
timestamp 1661296025
transform 1 0 1993 0 1 6480
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_112
timestamp 1661296025
transform 1 0 1993 0 1 6086
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_113
timestamp 1661296025
transform 1 0 1993 0 1 5690
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_114
timestamp 1661296025
transform 1 0 1993 0 1 5296
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_115
timestamp 1661296025
transform 1 0 1993 0 1 4900
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_116
timestamp 1661296025
transform 1 0 1993 0 1 4506
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_117
timestamp 1661296025
transform 1 0 1993 0 1 4110
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_118
timestamp 1661296025
transform 1 0 1993 0 1 3716
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_119
timestamp 1661296025
transform 1 0 1993 0 1 3320
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_120
timestamp 1661296025
transform 1 0 1993 0 1 2926
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_121
timestamp 1661296025
transform 1 0 1993 0 1 2530
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_122
timestamp 1661296025
transform 1 0 1993 0 1 2136
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_123
timestamp 1661296025
transform 1 0 1993 0 1 1740
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_124
timestamp 1661296025
transform 1 0 1993 0 1 1346
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_125
timestamp 1661296025
transform 1 0 1993 0 1 950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_126
timestamp 1661296025
transform 1 0 1993 0 1 556
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_127
timestamp 1661296025
transform 1 0 1993 0 1 160
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_128
timestamp 1661296025
transform 1 0 3441 0 1 25046
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_129
timestamp 1661296025
transform 1 0 3441 0 1 24650
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_130
timestamp 1661296025
transform 1 0 3441 0 1 24256
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_131
timestamp 1661296025
transform 1 0 3441 0 1 23860
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_132
timestamp 1661296025
transform 1 0 3441 0 1 23466
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_133
timestamp 1661296025
transform 1 0 3441 0 1 23070
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_134
timestamp 1661296025
transform 1 0 3441 0 1 22676
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_135
timestamp 1661296025
transform 1 0 3441 0 1 22280
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_136
timestamp 1661296025
transform 1 0 3441 0 1 21886
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_137
timestamp 1661296025
transform 1 0 3441 0 1 21490
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_138
timestamp 1661296025
transform 1 0 3441 0 1 21096
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_139
timestamp 1661296025
transform 1 0 3441 0 1 20700
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_140
timestamp 1661296025
transform 1 0 3441 0 1 20306
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_141
timestamp 1661296025
transform 1 0 3441 0 1 19910
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_142
timestamp 1661296025
transform 1 0 3441 0 1 19516
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_143
timestamp 1661296025
transform 1 0 3441 0 1 19120
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_144
timestamp 1661296025
transform 1 0 3441 0 1 18726
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_145
timestamp 1661296025
transform 1 0 3441 0 1 18330
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_146
timestamp 1661296025
transform 1 0 3441 0 1 17936
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_147
timestamp 1661296025
transform 1 0 3441 0 1 17540
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_148
timestamp 1661296025
transform 1 0 3441 0 1 17146
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_149
timestamp 1661296025
transform 1 0 3441 0 1 16750
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_150
timestamp 1661296025
transform 1 0 3441 0 1 16356
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_151
timestamp 1661296025
transform 1 0 3441 0 1 15960
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_152
timestamp 1661296025
transform 1 0 3441 0 1 15566
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_153
timestamp 1661296025
transform 1 0 3441 0 1 15170
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_154
timestamp 1661296025
transform 1 0 3441 0 1 14776
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_155
timestamp 1661296025
transform 1 0 3441 0 1 14380
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_156
timestamp 1661296025
transform 1 0 3441 0 1 13986
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_157
timestamp 1661296025
transform 1 0 3441 0 1 13590
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_158
timestamp 1661296025
transform 1 0 3441 0 1 13196
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_159
timestamp 1661296025
transform 1 0 3441 0 1 12800
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_160
timestamp 1661296025
transform 1 0 3441 0 1 12406
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_161
timestamp 1661296025
transform 1 0 3441 0 1 12010
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_162
timestamp 1661296025
transform 1 0 3441 0 1 11616
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_163
timestamp 1661296025
transform 1 0 3441 0 1 11220
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_164
timestamp 1661296025
transform 1 0 3441 0 1 10826
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_165
timestamp 1661296025
transform 1 0 3441 0 1 10430
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_166
timestamp 1661296025
transform 1 0 3441 0 1 10036
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_167
timestamp 1661296025
transform 1 0 3441 0 1 9640
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_168
timestamp 1661296025
transform 1 0 3441 0 1 9246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_169
timestamp 1661296025
transform 1 0 3441 0 1 8850
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_170
timestamp 1661296025
transform 1 0 3441 0 1 8456
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_171
timestamp 1661296025
transform 1 0 3441 0 1 8060
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_172
timestamp 1661296025
transform 1 0 3441 0 1 7666
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_173
timestamp 1661296025
transform 1 0 3441 0 1 7270
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_174
timestamp 1661296025
transform 1 0 3441 0 1 6876
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_175
timestamp 1661296025
transform 1 0 3441 0 1 6480
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_176
timestamp 1661296025
transform 1 0 3441 0 1 6086
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_177
timestamp 1661296025
transform 1 0 3441 0 1 5690
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_178
timestamp 1661296025
transform 1 0 3441 0 1 5296
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_179
timestamp 1661296025
transform 1 0 3441 0 1 4900
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_180
timestamp 1661296025
transform 1 0 3441 0 1 4506
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_181
timestamp 1661296025
transform 1 0 3441 0 1 4110
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_182
timestamp 1661296025
transform 1 0 3441 0 1 3716
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_183
timestamp 1661296025
transform 1 0 3441 0 1 3320
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_184
timestamp 1661296025
transform 1 0 3441 0 1 2926
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_185
timestamp 1661296025
transform 1 0 3441 0 1 2530
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_186
timestamp 1661296025
transform 1 0 3441 0 1 2136
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_187
timestamp 1661296025
transform 1 0 3441 0 1 1740
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_188
timestamp 1661296025
transform 1 0 3441 0 1 1346
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_189
timestamp 1661296025
transform 1 0 3441 0 1 950
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_190
timestamp 1661296025
transform 1 0 3441 0 1 556
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_191
timestamp 1661296025
transform 1 0 3441 0 1 160
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_192
timestamp 1661296025
transform 1 0 1150 0 1 25058
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_193
timestamp 1661296025
transform 1 0 1150 0 1 24638
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_194
timestamp 1661296025
transform 1 0 1150 0 1 24268
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_195
timestamp 1661296025
transform 1 0 1150 0 1 23848
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_196
timestamp 1661296025
transform 1 0 1150 0 1 23478
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_197
timestamp 1661296025
transform 1 0 1150 0 1 23058
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_198
timestamp 1661296025
transform 1 0 1150 0 1 22688
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_199
timestamp 1661296025
transform 1 0 1150 0 1 22268
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_200
timestamp 1661296025
transform 1 0 1150 0 1 21898
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_201
timestamp 1661296025
transform 1 0 1150 0 1 21478
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_202
timestamp 1661296025
transform 1 0 1150 0 1 21108
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_203
timestamp 1661296025
transform 1 0 1150 0 1 20688
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_204
timestamp 1661296025
transform 1 0 1150 0 1 20318
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_205
timestamp 1661296025
transform 1 0 1150 0 1 19898
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_206
timestamp 1661296025
transform 1 0 1150 0 1 19528
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_207
timestamp 1661296025
transform 1 0 1150 0 1 19108
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_208
timestamp 1661296025
transform 1 0 1150 0 1 18738
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_209
timestamp 1661296025
transform 1 0 1150 0 1 18318
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_210
timestamp 1661296025
transform 1 0 1150 0 1 17948
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_211
timestamp 1661296025
transform 1 0 1150 0 1 17528
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_212
timestamp 1661296025
transform 1 0 1150 0 1 17158
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_213
timestamp 1661296025
transform 1 0 1150 0 1 16738
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_214
timestamp 1661296025
transform 1 0 1150 0 1 16368
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_215
timestamp 1661296025
transform 1 0 1150 0 1 15948
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_216
timestamp 1661296025
transform 1 0 1150 0 1 15578
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_217
timestamp 1661296025
transform 1 0 1150 0 1 15158
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_218
timestamp 1661296025
transform 1 0 1150 0 1 14788
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_219
timestamp 1661296025
transform 1 0 1150 0 1 14368
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_220
timestamp 1661296025
transform 1 0 1150 0 1 13998
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_221
timestamp 1661296025
transform 1 0 1150 0 1 13578
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_222
timestamp 1661296025
transform 1 0 1150 0 1 13208
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_223
timestamp 1661296025
transform 1 0 1150 0 1 12788
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_224
timestamp 1661296025
transform 1 0 1150 0 1 12418
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_225
timestamp 1661296025
transform 1 0 1150 0 1 11998
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_226
timestamp 1661296025
transform 1 0 1150 0 1 11628
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_227
timestamp 1661296025
transform 1 0 1150 0 1 11208
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_228
timestamp 1661296025
transform 1 0 1150 0 1 10838
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_229
timestamp 1661296025
transform 1 0 1150 0 1 10418
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_230
timestamp 1661296025
transform 1 0 1150 0 1 10048
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_231
timestamp 1661296025
transform 1 0 1150 0 1 9628
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_232
timestamp 1661296025
transform 1 0 1150 0 1 9258
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_233
timestamp 1661296025
transform 1 0 1150 0 1 8838
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_234
timestamp 1661296025
transform 1 0 1150 0 1 8468
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_235
timestamp 1661296025
transform 1 0 1150 0 1 8048
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_236
timestamp 1661296025
transform 1 0 1150 0 1 7678
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_237
timestamp 1661296025
transform 1 0 1150 0 1 7258
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_238
timestamp 1661296025
transform 1 0 1150 0 1 6888
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_239
timestamp 1661296025
transform 1 0 1150 0 1 6468
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_240
timestamp 1661296025
transform 1 0 1150 0 1 6098
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_241
timestamp 1661296025
transform 1 0 1150 0 1 5678
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_242
timestamp 1661296025
transform 1 0 1150 0 1 5308
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_243
timestamp 1661296025
transform 1 0 1150 0 1 4888
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_244
timestamp 1661296025
transform 1 0 1150 0 1 4518
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_245
timestamp 1661296025
transform 1 0 1150 0 1 4098
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_246
timestamp 1661296025
transform 1 0 1150 0 1 3728
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_247
timestamp 1661296025
transform 1 0 1150 0 1 3308
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_248
timestamp 1661296025
transform 1 0 1150 0 1 2938
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_249
timestamp 1661296025
transform 1 0 1150 0 1 2518
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_250
timestamp 1661296025
transform 1 0 1150 0 1 2148
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_251
timestamp 1661296025
transform 1 0 1150 0 1 1728
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_252
timestamp 1661296025
transform 1 0 1150 0 1 1358
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_253
timestamp 1661296025
transform 1 0 1150 0 1 938
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_254
timestamp 1661296025
transform 1 0 1150 0 1 568
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_255
timestamp 1661296025
transform 1 0 1150 0 1 148
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_0
timestamp 1661296025
transform 1 0 720 0 1 25061
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_1
timestamp 1661296025
transform 1 0 720 0 1 24643
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_2
timestamp 1661296025
transform 1 0 720 0 1 24271
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_3
timestamp 1661296025
transform 1 0 720 0 1 23853
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_4
timestamp 1661296025
transform 1 0 720 0 1 23481
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_5
timestamp 1661296025
transform 1 0 720 0 1 23063
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_6
timestamp 1661296025
transform 1 0 720 0 1 22691
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_7
timestamp 1661296025
transform 1 0 720 0 1 22273
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_8
timestamp 1661296025
transform 1 0 720 0 1 21901
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_9
timestamp 1661296025
transform 1 0 720 0 1 21483
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_10
timestamp 1661296025
transform 1 0 720 0 1 21111
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_11
timestamp 1661296025
transform 1 0 720 0 1 20693
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_12
timestamp 1661296025
transform 1 0 720 0 1 20321
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_13
timestamp 1661296025
transform 1 0 720 0 1 19903
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_14
timestamp 1661296025
transform 1 0 720 0 1 19531
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_15
timestamp 1661296025
transform 1 0 720 0 1 19113
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_16
timestamp 1661296025
transform 1 0 720 0 1 18741
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_17
timestamp 1661296025
transform 1 0 720 0 1 18323
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_18
timestamp 1661296025
transform 1 0 720 0 1 17951
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_19
timestamp 1661296025
transform 1 0 720 0 1 17533
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_20
timestamp 1661296025
transform 1 0 720 0 1 17161
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_21
timestamp 1661296025
transform 1 0 720 0 1 16743
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_22
timestamp 1661296025
transform 1 0 720 0 1 16371
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_23
timestamp 1661296025
transform 1 0 720 0 1 15953
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_24
timestamp 1661296025
transform 1 0 720 0 1 15581
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_25
timestamp 1661296025
transform 1 0 720 0 1 15163
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_26
timestamp 1661296025
transform 1 0 720 0 1 14791
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_27
timestamp 1661296025
transform 1 0 720 0 1 14373
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_28
timestamp 1661296025
transform 1 0 720 0 1 14001
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_29
timestamp 1661296025
transform 1 0 720 0 1 13583
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_30
timestamp 1661296025
transform 1 0 720 0 1 13211
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_31
timestamp 1661296025
transform 1 0 720 0 1 12793
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_32
timestamp 1661296025
transform 1 0 720 0 1 12421
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_33
timestamp 1661296025
transform 1 0 720 0 1 12003
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_34
timestamp 1661296025
transform 1 0 720 0 1 11631
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_35
timestamp 1661296025
transform 1 0 720 0 1 11213
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_36
timestamp 1661296025
transform 1 0 720 0 1 10841
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_37
timestamp 1661296025
transform 1 0 720 0 1 10423
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_38
timestamp 1661296025
transform 1 0 720 0 1 10051
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_39
timestamp 1661296025
transform 1 0 720 0 1 9633
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_40
timestamp 1661296025
transform 1 0 720 0 1 9261
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_41
timestamp 1661296025
transform 1 0 720 0 1 8843
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_42
timestamp 1661296025
transform 1 0 720 0 1 8471
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_43
timestamp 1661296025
transform 1 0 720 0 1 8053
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_44
timestamp 1661296025
transform 1 0 720 0 1 7681
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_45
timestamp 1661296025
transform 1 0 720 0 1 7263
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_46
timestamp 1661296025
transform 1 0 720 0 1 6891
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_47
timestamp 1661296025
transform 1 0 720 0 1 6473
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_48
timestamp 1661296025
transform 1 0 720 0 1 6101
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_49
timestamp 1661296025
transform 1 0 720 0 1 5683
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_50
timestamp 1661296025
transform 1 0 720 0 1 5311
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_51
timestamp 1661296025
transform 1 0 720 0 1 4893
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_52
timestamp 1661296025
transform 1 0 720 0 1 4521
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_53
timestamp 1661296025
transform 1 0 720 0 1 4103
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_54
timestamp 1661296025
transform 1 0 720 0 1 3731
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_55
timestamp 1661296025
transform 1 0 720 0 1 3313
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_56
timestamp 1661296025
transform 1 0 720 0 1 2941
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_57
timestamp 1661296025
transform 1 0 720 0 1 2523
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_58
timestamp 1661296025
transform 1 0 720 0 1 2151
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_59
timestamp 1661296025
transform 1 0 720 0 1 1733
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_60
timestamp 1661296025
transform 1 0 720 0 1 1361
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_61
timestamp 1661296025
transform 1 0 720 0 1 943
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_62
timestamp 1661296025
transform 1 0 720 0 1 571
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_63
timestamp 1661296025
transform 1 0 720 0 1 153
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_64
timestamp 1661296025
transform 1 0 1988 0 1 25050
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_65
timestamp 1661296025
transform 1 0 1988 0 1 24654
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_66
timestamp 1661296025
transform 1 0 1988 0 1 24260
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_67
timestamp 1661296025
transform 1 0 1988 0 1 23864
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_68
timestamp 1661296025
transform 1 0 1988 0 1 23470
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_69
timestamp 1661296025
transform 1 0 1988 0 1 23074
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_70
timestamp 1661296025
transform 1 0 1988 0 1 22680
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_71
timestamp 1661296025
transform 1 0 1988 0 1 22284
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_72
timestamp 1661296025
transform 1 0 1988 0 1 21890
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_73
timestamp 1661296025
transform 1 0 1988 0 1 21494
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_74
timestamp 1661296025
transform 1 0 1988 0 1 21100
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_75
timestamp 1661296025
transform 1 0 1988 0 1 20704
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_76
timestamp 1661296025
transform 1 0 1988 0 1 20310
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_77
timestamp 1661296025
transform 1 0 1988 0 1 19914
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_78
timestamp 1661296025
transform 1 0 1988 0 1 19520
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_79
timestamp 1661296025
transform 1 0 1988 0 1 19124
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_80
timestamp 1661296025
transform 1 0 1988 0 1 18730
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_81
timestamp 1661296025
transform 1 0 1988 0 1 18334
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_82
timestamp 1661296025
transform 1 0 1988 0 1 17940
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_83
timestamp 1661296025
transform 1 0 1988 0 1 17544
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_84
timestamp 1661296025
transform 1 0 1988 0 1 17150
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_85
timestamp 1661296025
transform 1 0 1988 0 1 16754
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_86
timestamp 1661296025
transform 1 0 1988 0 1 16360
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_87
timestamp 1661296025
transform 1 0 1988 0 1 15964
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_88
timestamp 1661296025
transform 1 0 1988 0 1 15570
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_89
timestamp 1661296025
transform 1 0 1988 0 1 15174
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_90
timestamp 1661296025
transform 1 0 1988 0 1 14780
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_91
timestamp 1661296025
transform 1 0 1988 0 1 14384
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_92
timestamp 1661296025
transform 1 0 1988 0 1 13990
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_93
timestamp 1661296025
transform 1 0 1988 0 1 13594
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_94
timestamp 1661296025
transform 1 0 1988 0 1 13200
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_95
timestamp 1661296025
transform 1 0 1988 0 1 12804
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_96
timestamp 1661296025
transform 1 0 1988 0 1 12410
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_97
timestamp 1661296025
transform 1 0 1988 0 1 12014
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_98
timestamp 1661296025
transform 1 0 1988 0 1 11620
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_99
timestamp 1661296025
transform 1 0 1988 0 1 11224
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_100
timestamp 1661296025
transform 1 0 1988 0 1 10830
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_101
timestamp 1661296025
transform 1 0 1988 0 1 10434
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_102
timestamp 1661296025
transform 1 0 1988 0 1 10040
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_103
timestamp 1661296025
transform 1 0 1988 0 1 9644
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_104
timestamp 1661296025
transform 1 0 1988 0 1 9250
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_105
timestamp 1661296025
transform 1 0 1988 0 1 8854
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_106
timestamp 1661296025
transform 1 0 1988 0 1 8460
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_107
timestamp 1661296025
transform 1 0 1988 0 1 8064
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_108
timestamp 1661296025
transform 1 0 1988 0 1 7670
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_109
timestamp 1661296025
transform 1 0 1988 0 1 7274
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_110
timestamp 1661296025
transform 1 0 1988 0 1 6880
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_111
timestamp 1661296025
transform 1 0 1988 0 1 6484
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_112
timestamp 1661296025
transform 1 0 1988 0 1 6090
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_113
timestamp 1661296025
transform 1 0 1988 0 1 5694
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_114
timestamp 1661296025
transform 1 0 1988 0 1 5300
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_115
timestamp 1661296025
transform 1 0 1988 0 1 4904
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_116
timestamp 1661296025
transform 1 0 1988 0 1 4510
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_117
timestamp 1661296025
transform 1 0 1988 0 1 4114
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_118
timestamp 1661296025
transform 1 0 1988 0 1 3720
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_119
timestamp 1661296025
transform 1 0 1988 0 1 3324
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_120
timestamp 1661296025
transform 1 0 1988 0 1 2930
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_121
timestamp 1661296025
transform 1 0 1988 0 1 2534
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_122
timestamp 1661296025
transform 1 0 1988 0 1 2140
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_123
timestamp 1661296025
transform 1 0 1988 0 1 1744
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_124
timestamp 1661296025
transform 1 0 1988 0 1 1350
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_125
timestamp 1661296025
transform 1 0 1988 0 1 954
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_126
timestamp 1661296025
transform 1 0 1988 0 1 560
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_127
timestamp 1661296025
transform 1 0 1988 0 1 164
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_128
timestamp 1661296025
transform 1 0 3436 0 1 25050
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_129
timestamp 1661296025
transform 1 0 3436 0 1 24654
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_130
timestamp 1661296025
transform 1 0 3436 0 1 24260
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_131
timestamp 1661296025
transform 1 0 3436 0 1 23864
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_132
timestamp 1661296025
transform 1 0 3436 0 1 23470
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_133
timestamp 1661296025
transform 1 0 3436 0 1 23074
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_134
timestamp 1661296025
transform 1 0 3436 0 1 22680
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_135
timestamp 1661296025
transform 1 0 3436 0 1 22284
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_136
timestamp 1661296025
transform 1 0 3436 0 1 21890
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_137
timestamp 1661296025
transform 1 0 3436 0 1 21494
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_138
timestamp 1661296025
transform 1 0 3436 0 1 21100
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_139
timestamp 1661296025
transform 1 0 3436 0 1 20704
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_140
timestamp 1661296025
transform 1 0 3436 0 1 20310
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_141
timestamp 1661296025
transform 1 0 3436 0 1 19914
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_142
timestamp 1661296025
transform 1 0 3436 0 1 19520
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_143
timestamp 1661296025
transform 1 0 3436 0 1 19124
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_144
timestamp 1661296025
transform 1 0 3436 0 1 18730
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_145
timestamp 1661296025
transform 1 0 3436 0 1 18334
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_146
timestamp 1661296025
transform 1 0 3436 0 1 17940
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_147
timestamp 1661296025
transform 1 0 3436 0 1 17544
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_148
timestamp 1661296025
transform 1 0 3436 0 1 17150
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_149
timestamp 1661296025
transform 1 0 3436 0 1 16754
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_150
timestamp 1661296025
transform 1 0 3436 0 1 16360
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_151
timestamp 1661296025
transform 1 0 3436 0 1 15964
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_152
timestamp 1661296025
transform 1 0 3436 0 1 15570
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_153
timestamp 1661296025
transform 1 0 3436 0 1 15174
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_154
timestamp 1661296025
transform 1 0 3436 0 1 14780
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_155
timestamp 1661296025
transform 1 0 3436 0 1 14384
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_156
timestamp 1661296025
transform 1 0 3436 0 1 13990
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_157
timestamp 1661296025
transform 1 0 3436 0 1 13594
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_158
timestamp 1661296025
transform 1 0 3436 0 1 13200
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_159
timestamp 1661296025
transform 1 0 3436 0 1 12804
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_160
timestamp 1661296025
transform 1 0 3436 0 1 12410
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_161
timestamp 1661296025
transform 1 0 3436 0 1 12014
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_162
timestamp 1661296025
transform 1 0 3436 0 1 11620
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_163
timestamp 1661296025
transform 1 0 3436 0 1 11224
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_164
timestamp 1661296025
transform 1 0 3436 0 1 10830
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_165
timestamp 1661296025
transform 1 0 3436 0 1 10434
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_166
timestamp 1661296025
transform 1 0 3436 0 1 10040
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_167
timestamp 1661296025
transform 1 0 3436 0 1 9644
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_168
timestamp 1661296025
transform 1 0 3436 0 1 9250
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_169
timestamp 1661296025
transform 1 0 3436 0 1 8854
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_170
timestamp 1661296025
transform 1 0 3436 0 1 8460
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_171
timestamp 1661296025
transform 1 0 3436 0 1 8064
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_172
timestamp 1661296025
transform 1 0 3436 0 1 7670
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_173
timestamp 1661296025
transform 1 0 3436 0 1 7274
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_174
timestamp 1661296025
transform 1 0 3436 0 1 6880
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_175
timestamp 1661296025
transform 1 0 3436 0 1 6484
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_176
timestamp 1661296025
transform 1 0 3436 0 1 6090
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_177
timestamp 1661296025
transform 1 0 3436 0 1 5694
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_178
timestamp 1661296025
transform 1 0 3436 0 1 5300
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_179
timestamp 1661296025
transform 1 0 3436 0 1 4904
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_180
timestamp 1661296025
transform 1 0 3436 0 1 4510
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_181
timestamp 1661296025
transform 1 0 3436 0 1 4114
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_182
timestamp 1661296025
transform 1 0 3436 0 1 3720
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_183
timestamp 1661296025
transform 1 0 3436 0 1 3324
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_184
timestamp 1661296025
transform 1 0 3436 0 1 2930
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_185
timestamp 1661296025
transform 1 0 3436 0 1 2534
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_186
timestamp 1661296025
transform 1 0 3436 0 1 2140
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_187
timestamp 1661296025
transform 1 0 3436 0 1 1744
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_188
timestamp 1661296025
transform 1 0 3436 0 1 1350
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_189
timestamp 1661296025
transform 1 0 3436 0 1 954
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_190
timestamp 1661296025
transform 1 0 3436 0 1 560
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_191
timestamp 1661296025
transform 1 0 3436 0 1 164
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_192
timestamp 1661296025
transform 1 0 1145 0 1 25062
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_193
timestamp 1661296025
transform 1 0 1145 0 1 24642
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_194
timestamp 1661296025
transform 1 0 1145 0 1 24272
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_195
timestamp 1661296025
transform 1 0 1145 0 1 23852
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_196
timestamp 1661296025
transform 1 0 1145 0 1 23482
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_197
timestamp 1661296025
transform 1 0 1145 0 1 23062
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_198
timestamp 1661296025
transform 1 0 1145 0 1 22692
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_199
timestamp 1661296025
transform 1 0 1145 0 1 22272
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_200
timestamp 1661296025
transform 1 0 1145 0 1 21902
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_201
timestamp 1661296025
transform 1 0 1145 0 1 21482
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_202
timestamp 1661296025
transform 1 0 1145 0 1 21112
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_203
timestamp 1661296025
transform 1 0 1145 0 1 20692
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_204
timestamp 1661296025
transform 1 0 1145 0 1 20322
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_205
timestamp 1661296025
transform 1 0 1145 0 1 19902
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_206
timestamp 1661296025
transform 1 0 1145 0 1 19532
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_207
timestamp 1661296025
transform 1 0 1145 0 1 19112
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_208
timestamp 1661296025
transform 1 0 1145 0 1 18742
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_209
timestamp 1661296025
transform 1 0 1145 0 1 18322
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_210
timestamp 1661296025
transform 1 0 1145 0 1 17952
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_211
timestamp 1661296025
transform 1 0 1145 0 1 17532
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_212
timestamp 1661296025
transform 1 0 1145 0 1 17162
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_213
timestamp 1661296025
transform 1 0 1145 0 1 16742
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_214
timestamp 1661296025
transform 1 0 1145 0 1 16372
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_215
timestamp 1661296025
transform 1 0 1145 0 1 15952
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_216
timestamp 1661296025
transform 1 0 1145 0 1 15582
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_217
timestamp 1661296025
transform 1 0 1145 0 1 15162
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_218
timestamp 1661296025
transform 1 0 1145 0 1 14792
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_219
timestamp 1661296025
transform 1 0 1145 0 1 14372
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_220
timestamp 1661296025
transform 1 0 1145 0 1 14002
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_221
timestamp 1661296025
transform 1 0 1145 0 1 13582
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_222
timestamp 1661296025
transform 1 0 1145 0 1 13212
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_223
timestamp 1661296025
transform 1 0 1145 0 1 12792
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_224
timestamp 1661296025
transform 1 0 1145 0 1 12422
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_225
timestamp 1661296025
transform 1 0 1145 0 1 12002
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_226
timestamp 1661296025
transform 1 0 1145 0 1 11632
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_227
timestamp 1661296025
transform 1 0 1145 0 1 11212
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_228
timestamp 1661296025
transform 1 0 1145 0 1 10842
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_229
timestamp 1661296025
transform 1 0 1145 0 1 10422
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_230
timestamp 1661296025
transform 1 0 1145 0 1 10052
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_231
timestamp 1661296025
transform 1 0 1145 0 1 9632
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_232
timestamp 1661296025
transform 1 0 1145 0 1 9262
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_233
timestamp 1661296025
transform 1 0 1145 0 1 8842
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_234
timestamp 1661296025
transform 1 0 1145 0 1 8472
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_235
timestamp 1661296025
transform 1 0 1145 0 1 8052
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_236
timestamp 1661296025
transform 1 0 1145 0 1 7682
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_237
timestamp 1661296025
transform 1 0 1145 0 1 7262
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_238
timestamp 1661296025
transform 1 0 1145 0 1 6892
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_239
timestamp 1661296025
transform 1 0 1145 0 1 6472
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_240
timestamp 1661296025
transform 1 0 1145 0 1 6102
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_241
timestamp 1661296025
transform 1 0 1145 0 1 5682
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_242
timestamp 1661296025
transform 1 0 1145 0 1 5312
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_243
timestamp 1661296025
transform 1 0 1145 0 1 4892
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_244
timestamp 1661296025
transform 1 0 1145 0 1 4522
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_245
timestamp 1661296025
transform 1 0 1145 0 1 4102
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_246
timestamp 1661296025
transform 1 0 1145 0 1 3732
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_247
timestamp 1661296025
transform 1 0 1145 0 1 3312
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_248
timestamp 1661296025
transform 1 0 1145 0 1 2942
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_249
timestamp 1661296025
transform 1 0 1145 0 1 2522
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_250
timestamp 1661296025
transform 1 0 1145 0 1 2152
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_251
timestamp 1661296025
transform 1 0 1145 0 1 1732
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_252
timestamp 1661296025
transform 1 0 1145 0 1 1362
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_253
timestamp 1661296025
transform 1 0 1145 0 1 942
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_254
timestamp 1661296025
transform 1 0 1145 0 1 572
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_contact_22  sky130_sram_1r1w_24x128_8_contact_22_255
timestamp 1661296025
transform 1 0 1145 0 1 152
box 0 0 76 66
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_0
timestamp 1661296025
transform 1 0 488 0 -1 25280
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_1
timestamp 1661296025
transform 1 0 488 0 1 24490
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_2
timestamp 1661296025
transform 1 0 488 0 -1 24490
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_3
timestamp 1661296025
transform 1 0 488 0 1 23700
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_4
timestamp 1661296025
transform 1 0 488 0 -1 23700
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_5
timestamp 1661296025
transform 1 0 488 0 1 22910
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_6
timestamp 1661296025
transform 1 0 488 0 -1 22910
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_7
timestamp 1661296025
transform 1 0 488 0 1 22120
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_8
timestamp 1661296025
transform 1 0 488 0 -1 22120
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_9
timestamp 1661296025
transform 1 0 488 0 1 21330
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_10
timestamp 1661296025
transform 1 0 488 0 -1 21330
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_11
timestamp 1661296025
transform 1 0 488 0 1 20540
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_12
timestamp 1661296025
transform 1 0 488 0 -1 20540
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_13
timestamp 1661296025
transform 1 0 488 0 1 19750
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_14
timestamp 1661296025
transform 1 0 488 0 -1 19750
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_15
timestamp 1661296025
transform 1 0 488 0 1 18960
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_16
timestamp 1661296025
transform 1 0 488 0 -1 18960
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_17
timestamp 1661296025
transform 1 0 488 0 1 18170
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_18
timestamp 1661296025
transform 1 0 488 0 -1 18170
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_19
timestamp 1661296025
transform 1 0 488 0 1 17380
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_20
timestamp 1661296025
transform 1 0 488 0 -1 17380
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_21
timestamp 1661296025
transform 1 0 488 0 1 16590
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_22
timestamp 1661296025
transform 1 0 488 0 -1 16590
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_23
timestamp 1661296025
transform 1 0 488 0 1 15800
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_24
timestamp 1661296025
transform 1 0 488 0 -1 15800
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_25
timestamp 1661296025
transform 1 0 488 0 1 15010
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_26
timestamp 1661296025
transform 1 0 488 0 -1 15010
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_27
timestamp 1661296025
transform 1 0 488 0 1 14220
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_28
timestamp 1661296025
transform 1 0 488 0 -1 14220
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_29
timestamp 1661296025
transform 1 0 488 0 1 13430
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_30
timestamp 1661296025
transform 1 0 488 0 -1 13430
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_31
timestamp 1661296025
transform 1 0 488 0 1 12640
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_32
timestamp 1661296025
transform 1 0 488 0 -1 12640
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_33
timestamp 1661296025
transform 1 0 488 0 1 11850
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_34
timestamp 1661296025
transform 1 0 488 0 -1 11850
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_35
timestamp 1661296025
transform 1 0 488 0 1 11060
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_36
timestamp 1661296025
transform 1 0 488 0 -1 11060
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_37
timestamp 1661296025
transform 1 0 488 0 1 10270
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_38
timestamp 1661296025
transform 1 0 488 0 -1 10270
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_39
timestamp 1661296025
transform 1 0 488 0 1 9480
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_40
timestamp 1661296025
transform 1 0 488 0 -1 9480
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_41
timestamp 1661296025
transform 1 0 488 0 1 8690
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_42
timestamp 1661296025
transform 1 0 488 0 -1 8690
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_43
timestamp 1661296025
transform 1 0 488 0 1 7900
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_44
timestamp 1661296025
transform 1 0 488 0 -1 7900
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_45
timestamp 1661296025
transform 1 0 488 0 1 7110
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_46
timestamp 1661296025
transform 1 0 488 0 -1 7110
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_47
timestamp 1661296025
transform 1 0 488 0 1 6320
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_48
timestamp 1661296025
transform 1 0 488 0 -1 6320
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_49
timestamp 1661296025
transform 1 0 488 0 1 5530
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_50
timestamp 1661296025
transform 1 0 488 0 -1 5530
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_51
timestamp 1661296025
transform 1 0 488 0 1 4740
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_52
timestamp 1661296025
transform 1 0 488 0 -1 4740
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_53
timestamp 1661296025
transform 1 0 488 0 1 3950
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_54
timestamp 1661296025
transform 1 0 488 0 -1 3950
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_55
timestamp 1661296025
transform 1 0 488 0 1 3160
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_56
timestamp 1661296025
transform 1 0 488 0 -1 3160
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_57
timestamp 1661296025
transform 1 0 488 0 1 2370
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_58
timestamp 1661296025
transform 1 0 488 0 -1 2370
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_59
timestamp 1661296025
transform 1 0 488 0 1 1580
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_60
timestamp 1661296025
transform 1 0 488 0 -1 1580
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_61
timestamp 1661296025
transform 1 0 488 0 1 790
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_62
timestamp 1661296025
transform 1 0 488 0 -1 790
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_wordline_driver  sky130_sram_1r1w_24x128_8_wordline_driver_63
timestamp 1661296025
transform 1 0 488 0 1 0
box 70 -56 3740 490
<< labels >>
rlabel metal2 s 577 0 605 25280 4 en
port 1 nsew
rlabel locali s 591 299 591 299 4 in_0
port 2 nsew
rlabel locali s 4199 120 4199 120 4 wl_0
port 3 nsew
rlabel locali s 591 491 591 491 4 in_1
port 4 nsew
rlabel locali s 4199 670 4199 670 4 wl_1
port 5 nsew
rlabel locali s 591 1089 591 1089 4 in_2
port 6 nsew
rlabel locali s 4199 910 4199 910 4 wl_2
port 7 nsew
rlabel locali s 591 1281 591 1281 4 in_3
port 8 nsew
rlabel locali s 4199 1460 4199 1460 4 wl_3
port 9 nsew
rlabel locali s 591 1879 591 1879 4 in_4
port 10 nsew
rlabel locali s 4199 1700 4199 1700 4 wl_4
port 11 nsew
rlabel locali s 591 2071 591 2071 4 in_5
port 12 nsew
rlabel locali s 4199 2250 4199 2250 4 wl_5
port 13 nsew
rlabel locali s 591 2669 591 2669 4 in_6
port 14 nsew
rlabel locali s 4199 2490 4199 2490 4 wl_6
port 15 nsew
rlabel locali s 591 2861 591 2861 4 in_7
port 16 nsew
rlabel locali s 4199 3040 4199 3040 4 wl_7
port 17 nsew
rlabel locali s 591 3459 591 3459 4 in_8
port 18 nsew
rlabel locali s 4199 3280 4199 3280 4 wl_8
port 19 nsew
rlabel locali s 591 3651 591 3651 4 in_9
port 20 nsew
rlabel locali s 4199 3830 4199 3830 4 wl_9
port 21 nsew
rlabel locali s 591 4249 591 4249 4 in_10
port 22 nsew
rlabel locali s 4199 4070 4199 4070 4 wl_10
port 23 nsew
rlabel locali s 591 4441 591 4441 4 in_11
port 24 nsew
rlabel locali s 4199 4620 4199 4620 4 wl_11
port 25 nsew
rlabel locali s 591 5039 591 5039 4 in_12
port 26 nsew
rlabel locali s 4199 4860 4199 4860 4 wl_12
port 27 nsew
rlabel locali s 591 5231 591 5231 4 in_13
port 28 nsew
rlabel locali s 4199 5410 4199 5410 4 wl_13
port 29 nsew
rlabel locali s 591 5829 591 5829 4 in_14
port 30 nsew
rlabel locali s 4199 5650 4199 5650 4 wl_14
port 31 nsew
rlabel locali s 591 6021 591 6021 4 in_15
port 32 nsew
rlabel locali s 4199 6200 4199 6200 4 wl_15
port 33 nsew
rlabel locali s 591 6619 591 6619 4 in_16
port 34 nsew
rlabel locali s 4199 6440 4199 6440 4 wl_16
port 35 nsew
rlabel locali s 591 6811 591 6811 4 in_17
port 36 nsew
rlabel locali s 4199 6990 4199 6990 4 wl_17
port 37 nsew
rlabel locali s 591 7409 591 7409 4 in_18
port 38 nsew
rlabel locali s 4199 7230 4199 7230 4 wl_18
port 39 nsew
rlabel locali s 591 7601 591 7601 4 in_19
port 40 nsew
rlabel locali s 4199 7780 4199 7780 4 wl_19
port 41 nsew
rlabel locali s 591 8199 591 8199 4 in_20
port 42 nsew
rlabel locali s 4199 8020 4199 8020 4 wl_20
port 43 nsew
rlabel locali s 591 8391 591 8391 4 in_21
port 44 nsew
rlabel locali s 4199 8570 4199 8570 4 wl_21
port 45 nsew
rlabel locali s 591 8989 591 8989 4 in_22
port 46 nsew
rlabel locali s 4199 8810 4199 8810 4 wl_22
port 47 nsew
rlabel locali s 591 9181 591 9181 4 in_23
port 48 nsew
rlabel locali s 4199 9360 4199 9360 4 wl_23
port 49 nsew
rlabel locali s 591 9779 591 9779 4 in_24
port 50 nsew
rlabel locali s 4199 9600 4199 9600 4 wl_24
port 51 nsew
rlabel locali s 591 9971 591 9971 4 in_25
port 52 nsew
rlabel locali s 4199 10150 4199 10150 4 wl_25
port 53 nsew
rlabel locali s 591 10569 591 10569 4 in_26
port 54 nsew
rlabel locali s 4199 10390 4199 10390 4 wl_26
port 55 nsew
rlabel locali s 591 10761 591 10761 4 in_27
port 56 nsew
rlabel locali s 4199 10940 4199 10940 4 wl_27
port 57 nsew
rlabel locali s 591 11359 591 11359 4 in_28
port 58 nsew
rlabel locali s 4199 11180 4199 11180 4 wl_28
port 59 nsew
rlabel locali s 591 11551 591 11551 4 in_29
port 60 nsew
rlabel locali s 4199 11730 4199 11730 4 wl_29
port 61 nsew
rlabel locali s 591 12149 591 12149 4 in_30
port 62 nsew
rlabel locali s 4199 11970 4199 11970 4 wl_30
port 63 nsew
rlabel locali s 591 12341 591 12341 4 in_31
port 64 nsew
rlabel locali s 4199 12520 4199 12520 4 wl_31
port 65 nsew
rlabel locali s 591 12939 591 12939 4 in_32
port 66 nsew
rlabel locali s 4199 12760 4199 12760 4 wl_32
port 67 nsew
rlabel locali s 591 13131 591 13131 4 in_33
port 68 nsew
rlabel locali s 4199 13310 4199 13310 4 wl_33
port 69 nsew
rlabel locali s 591 13729 591 13729 4 in_34
port 70 nsew
rlabel locali s 4199 13550 4199 13550 4 wl_34
port 71 nsew
rlabel locali s 591 13921 591 13921 4 in_35
port 72 nsew
rlabel locali s 4199 14100 4199 14100 4 wl_35
port 73 nsew
rlabel locali s 591 14519 591 14519 4 in_36
port 74 nsew
rlabel locali s 4199 14340 4199 14340 4 wl_36
port 75 nsew
rlabel locali s 591 14711 591 14711 4 in_37
port 76 nsew
rlabel locali s 4199 14890 4199 14890 4 wl_37
port 77 nsew
rlabel locali s 591 15309 591 15309 4 in_38
port 78 nsew
rlabel locali s 4199 15130 4199 15130 4 wl_38
port 79 nsew
rlabel locali s 591 15501 591 15501 4 in_39
port 80 nsew
rlabel locali s 4199 15680 4199 15680 4 wl_39
port 81 nsew
rlabel locali s 591 16099 591 16099 4 in_40
port 82 nsew
rlabel locali s 4199 15920 4199 15920 4 wl_40
port 83 nsew
rlabel locali s 591 16291 591 16291 4 in_41
port 84 nsew
rlabel locali s 4199 16470 4199 16470 4 wl_41
port 85 nsew
rlabel locali s 591 16889 591 16889 4 in_42
port 86 nsew
rlabel locali s 4199 16710 4199 16710 4 wl_42
port 87 nsew
rlabel locali s 591 17081 591 17081 4 in_43
port 88 nsew
rlabel locali s 4199 17260 4199 17260 4 wl_43
port 89 nsew
rlabel locali s 591 17679 591 17679 4 in_44
port 90 nsew
rlabel locali s 4199 17500 4199 17500 4 wl_44
port 91 nsew
rlabel locali s 591 17871 591 17871 4 in_45
port 92 nsew
rlabel locali s 4199 18050 4199 18050 4 wl_45
port 93 nsew
rlabel locali s 591 18469 591 18469 4 in_46
port 94 nsew
rlabel locali s 4199 18290 4199 18290 4 wl_46
port 95 nsew
rlabel locali s 591 18661 591 18661 4 in_47
port 96 nsew
rlabel locali s 4199 18840 4199 18840 4 wl_47
port 97 nsew
rlabel locali s 591 19259 591 19259 4 in_48
port 98 nsew
rlabel locali s 4199 19080 4199 19080 4 wl_48
port 99 nsew
rlabel locali s 591 19451 591 19451 4 in_49
port 100 nsew
rlabel locali s 4199 19630 4199 19630 4 wl_49
port 101 nsew
rlabel locali s 591 20049 591 20049 4 in_50
port 102 nsew
rlabel locali s 4199 19870 4199 19870 4 wl_50
port 103 nsew
rlabel locali s 591 20241 591 20241 4 in_51
port 104 nsew
rlabel locali s 4199 20420 4199 20420 4 wl_51
port 105 nsew
rlabel locali s 591 20839 591 20839 4 in_52
port 106 nsew
rlabel locali s 4199 20660 4199 20660 4 wl_52
port 107 nsew
rlabel locali s 591 21031 591 21031 4 in_53
port 108 nsew
rlabel locali s 4199 21210 4199 21210 4 wl_53
port 109 nsew
rlabel locali s 591 21629 591 21629 4 in_54
port 110 nsew
rlabel locali s 4199 21450 4199 21450 4 wl_54
port 111 nsew
rlabel locali s 591 21821 591 21821 4 in_55
port 112 nsew
rlabel locali s 4199 22000 4199 22000 4 wl_55
port 113 nsew
rlabel locali s 591 22419 591 22419 4 in_56
port 114 nsew
rlabel locali s 4199 22240 4199 22240 4 wl_56
port 115 nsew
rlabel locali s 591 22611 591 22611 4 in_57
port 116 nsew
rlabel locali s 4199 22790 4199 22790 4 wl_57
port 117 nsew
rlabel locali s 591 23209 591 23209 4 in_58
port 118 nsew
rlabel locali s 4199 23030 4199 23030 4 wl_58
port 119 nsew
rlabel locali s 591 23401 591 23401 4 in_59
port 120 nsew
rlabel locali s 4199 23580 4199 23580 4 wl_59
port 121 nsew
rlabel locali s 591 23999 591 23999 4 in_60
port 122 nsew
rlabel locali s 4199 23820 4199 23820 4 wl_60
port 123 nsew
rlabel locali s 591 24191 591 24191 4 in_61
port 124 nsew
rlabel locali s 4199 24370 4199 24370 4 wl_61
port 125 nsew
rlabel locali s 591 24789 591 24789 4 in_62
port 126 nsew
rlabel locali s 4199 24610 4199 24610 4 wl_62
port 127 nsew
rlabel locali s 591 24981 591 24981 4 in_63
port 128 nsew
rlabel locali s 4199 25160 4199 25160 4 wl_63
port 129 nsew
rlabel metal4 s 1150 -65 1216 25345 4 vdd
port 130 nsew
rlabel metal4 s 3441 -33 3507 25313 4 vdd
port 130 nsew
rlabel metal4 s 1993 -33 2059 25313 4 gnd
port 131 nsew
rlabel metal4 s 725 -63 791 25343 4 gnd
port 131 nsew
<< properties >>
string FIXED_BBOX 0 0 4246 25280
<< end >>
