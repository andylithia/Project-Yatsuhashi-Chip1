magic
tech sky130B
timestamp 1659754370
<< metal1 >>
rect 13 685 43 720
<< metal2 >>
rect 0 341 10 577
rect 0 80 10 316
<< metal3 >>
rect 200 300 1041 350
use nfet_3x_2  nfet_3x_2_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/LNA
timestamp 1659754370
transform 1 0 0 0 1 30
box 0 -30 646 690
use nfet_3x_2  nfet_3x_2_1
timestamp 1659754370
transform 1 0 591 0 1 30
box 0 -30 646 690
<< labels >>
rlabel metal2 0 341 10 577 1 D
rlabel metal2 0 80 10 316 1 S
rlabel metal1 13 685 43 720 1 B
rlabel metal3 200 300 1041 350 1 G
<< end >>
