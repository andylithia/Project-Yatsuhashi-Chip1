** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/gmid_test/nmos_test.sch
**.subckt nmos_test
XM1 vds vgs GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W * 0.29' as='int((nf+2)/2) * W * 0.29'
+ pd='2*int((nf+1)/2) * (W + 0.29)' ps='2*int((nf+2)/2) * (W + 0.29)' nrd='0.29 / W / nf' nrs='0.29 / W / nf'
+ sa=0 sb=0 sd=0 mult=1 m=1
VGS vgs GND 0.9
VDD vds GND 1
**** begin user architecture code


.param L=0.15
.param W=1
.param NF=1
.op
.control
save @m.xm1.msky130_fd_pr__nfet_01v8[gm]
save @m.xm1.msky130_fd_pr__nfet_01v8[id]
save @m.xm1.msky130_fd_pr__nfet_01v8[gds]
save @m.xm1.msky130_fd_pr__nfet_01v8[cgs]
save @m.xm1.msky130_fd_pr__nfet_01v8[cgb]
save @m.xm1.msky130_fd_pr__nfet_01v8[cgd]
save @m.xm1.msky130_fd_pr__nfet_01v8[vth]

let w_start = 1
let w_stop  = 10
let delta_w = 1

let l_start = 0.15
let l_stop  = 1.5
let delta_l = 0.15


let w_test = w_start
while w_test le w_stop
 let l_test = l_start
 while l_test le l_stop
  alter @m.xm1.msky130_fd_pr__nfet_01v8[w] = w_test
  alter @m.xm1.msky130_fd_pr__nfet_01v8[l] = l_test
  op
  DC VGS 0 1.8 0.01
  * plot @m.xm1.msky130_fd_pr__nfet_01v8[id]
  * plot @m.xm1.msky130_fd_pr__nfet_01v8[vth]
  set filetype=ascii
  write ./gmid_test/data_L{$&l_test}_W{$&w_test}.raw
  let l_test = l_test + delta_l
 end
 let w_test = w_test + delta_w
end
.endc


.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
**** end user architecture code
**.ends
.GLOBAL GND
.end
