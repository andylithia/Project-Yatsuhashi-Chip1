magic
tech sky130B
magscale 1 2
timestamp 1660275428
<< dnwell >>
rect 4200 -4100 10500 900
<< nwell >>
rect 4120 694 10580 980
rect 4120 -3894 4406 694
rect 10294 -3894 10580 694
rect 4120 -4180 10580 -3894
<< nsubdiff >>
rect 4157 923 10543 943
rect 4157 889 4237 923
rect 10463 889 10543 923
rect 4157 869 10543 889
rect 4157 863 4231 869
rect 4157 -4063 4177 863
rect 4211 -4063 4231 863
rect 4157 -4069 4231 -4063
rect 10469 863 10543 869
rect 10469 -4063 10489 863
rect 10523 -4063 10543 863
rect 10469 -4069 10543 -4063
rect 4157 -4089 10543 -4069
rect 4157 -4123 4237 -4089
rect 10463 -4123 10543 -4089
rect 4157 -4143 10543 -4123
<< nsubdiffcont >>
rect 4237 889 10463 923
rect 4177 -4063 4211 863
rect 10489 -4063 10523 863
rect 4237 -4123 10463 -4089
<< locali >>
rect 4177 920 4237 923
rect 10463 920 10523 923
rect 4177 863 4180 920
rect 10520 863 10523 920
rect 4177 -4120 4180 -4063
rect 10520 -4120 10523 -4063
rect 4177 -4123 4237 -4120
rect 10463 -4123 10523 -4120
<< viali >>
rect 4180 889 4237 920
rect 4237 889 10463 920
rect 10463 889 10520 920
rect 4180 880 10520 889
rect 4180 863 4220 880
rect 4180 -4063 4211 863
rect 4211 -4063 4220 863
rect 10480 863 10520 880
rect 4660 500 9900 560
rect 4630 -3650 4670 460
rect 9950 -3650 9990 460
rect 4720 -3730 9900 -3690
rect 4180 -4080 4220 -4063
rect 10480 -4063 10489 863
rect 10489 -4063 10520 863
rect 10480 -4080 10520 -4063
rect 4180 -4089 10520 -4080
rect 4180 -4120 4237 -4089
rect 4237 -4120 10463 -4089
rect 10463 -4120 10520 -4089
<< metal1 >>
rect 4160 920 4280 940
rect 10420 920 10540 940
rect 4160 -4120 4180 920
rect 4220 820 4280 880
rect 10420 860 10480 880
rect 10440 820 10480 860
rect 4620 480 4660 580
rect 9880 560 10010 580
rect 9900 500 10010 560
rect 9880 480 10010 500
rect 4620 460 4690 480
rect 4620 -3650 4630 460
rect 4670 -3650 4690 460
rect 9940 460 10010 480
rect 4810 370 4820 430
rect 5060 370 5070 430
rect 5130 370 5140 430
rect 5380 370 5390 430
rect 5450 370 5460 430
rect 5700 370 5710 430
rect 5760 370 5770 430
rect 6010 370 6020 430
rect 6080 370 6090 430
rect 6330 370 6340 430
rect 6390 370 6400 430
rect 6640 370 6650 430
rect 6710 370 6720 430
rect 6960 370 6970 430
rect 7030 370 7040 430
rect 7280 370 7290 430
rect 7340 370 7350 430
rect 7590 370 7600 430
rect 7660 370 7670 430
rect 7910 370 7920 430
rect 7970 370 7980 430
rect 8220 370 8230 430
rect 8290 370 8300 430
rect 8540 370 8550 430
rect 8610 370 8620 430
rect 8860 370 8870 430
rect 8920 370 8930 430
rect 9170 370 9180 430
rect 9240 370 9250 430
rect 9490 370 9500 430
rect 9550 370 9560 430
rect 9800 370 9810 430
rect 4755 310 4810 340
rect 4755 -460 4810 -430
rect 4913 310 4968 340
rect 4913 -460 4968 -430
rect 5071 310 5126 340
rect 5071 -460 5126 -430
rect 5229 310 5284 340
rect 5229 -460 5284 -430
rect 5387 310 5442 340
rect 5387 -460 5442 -430
rect 5545 310 5600 340
rect 5545 -460 5600 -430
rect 5703 310 5758 340
rect 5703 -460 5758 -430
rect 5861 310 5916 340
rect 5861 -460 5916 -430
rect 6019 310 6074 340
rect 6019 -460 6074 -430
rect 6177 310 6232 340
rect 6177 -460 6232 -430
rect 6335 310 6390 340
rect 6335 -460 6390 -430
rect 6493 310 6548 340
rect 6493 -460 6548 -430
rect 6651 310 6706 340
rect 6651 -460 6706 -430
rect 6809 310 6864 340
rect 6809 -460 6864 -430
rect 6967 310 7022 340
rect 6967 -460 7022 -430
rect 7125 310 7180 340
rect 7125 -460 7180 -430
rect 7283 310 7338 340
rect 7283 -460 7338 -430
rect 7441 310 7496 340
rect 7441 -460 7496 -430
rect 7599 310 7654 340
rect 7599 -460 7654 -430
rect 7757 310 7812 340
rect 7757 -460 7812 -430
rect 7915 310 7970 340
rect 7915 -460 7970 -430
rect 8073 310 8128 340
rect 8073 -460 8128 -430
rect 8231 310 8286 340
rect 8231 -460 8286 -430
rect 8389 310 8444 340
rect 8389 -460 8444 -430
rect 8547 310 8602 340
rect 8547 -460 8602 -430
rect 8705 310 8760 340
rect 8705 -460 8760 -430
rect 8863 310 8918 340
rect 8863 -460 8918 -430
rect 9021 310 9076 340
rect 9021 -460 9076 -430
rect 9179 310 9234 340
rect 9179 -460 9234 -430
rect 9337 310 9392 340
rect 9337 -460 9392 -430
rect 9495 310 9550 340
rect 9495 -460 9550 -430
rect 9653 310 9708 340
rect 9653 -460 9708 -430
rect 9811 310 9866 340
rect 9811 -460 9866 -430
rect 4810 -560 4820 -500
rect 5060 -560 5070 -500
rect 5130 -560 5140 -500
rect 5380 -560 5390 -500
rect 5450 -515 5460 -500
rect 5449 -560 5460 -515
rect 5700 -560 5710 -500
rect 5760 -560 5770 -500
rect 6010 -560 6020 -500
rect 6080 -560 6090 -500
rect 6330 -560 6340 -500
rect 6390 -560 6400 -500
rect 6640 -560 6650 -500
rect 6710 -560 6720 -500
rect 6960 -560 6970 -500
rect 7030 -515 7040 -500
rect 7029 -560 7040 -515
rect 7280 -560 7290 -500
rect 7340 -560 7350 -500
rect 7590 -560 7600 -500
rect 7660 -560 7670 -500
rect 7910 -560 7920 -500
rect 7970 -560 7980 -500
rect 8220 -560 8230 -500
rect 8290 -560 8300 -500
rect 8540 -560 8550 -500
rect 8610 -515 8620 -500
rect 8609 -560 8620 -515
rect 8860 -560 8870 -500
rect 8920 -560 8930 -500
rect 9170 -560 9180 -500
rect 9240 -560 9250 -500
rect 9490 -560 9500 -500
rect 9550 -560 9560 -500
rect 9800 -560 9810 -500
rect 4817 -561 4909 -560
rect 4975 -561 5067 -560
rect 5133 -561 5225 -560
rect 5291 -561 5383 -560
rect 5449 -561 5541 -560
rect 5607 -561 5699 -560
rect 5765 -561 5857 -560
rect 5923 -561 6015 -560
rect 6081 -561 6173 -560
rect 6239 -561 6331 -560
rect 6397 -561 6489 -560
rect 6555 -561 6647 -560
rect 6713 -561 6805 -560
rect 6871 -561 6963 -560
rect 7029 -561 7121 -560
rect 7187 -561 7279 -560
rect 7345 -561 7437 -560
rect 7503 -561 7595 -560
rect 7661 -561 7753 -560
rect 7819 -561 7911 -560
rect 7977 -561 8069 -560
rect 8135 -561 8227 -560
rect 8293 -561 8385 -560
rect 8451 -561 8543 -560
rect 8609 -561 8701 -560
rect 8767 -561 8859 -560
rect 8925 -561 9017 -560
rect 9083 -561 9175 -560
rect 9241 -561 9333 -560
rect 9399 -561 9491 -560
rect 9557 -561 9649 -560
rect 9715 -561 9807 -560
rect 4810 -649 4820 -589
rect 5060 -590 5070 -589
rect 5130 -590 5140 -589
rect 5060 -649 5140 -590
rect 5380 -590 5390 -589
rect 5450 -590 5460 -589
rect 5380 -649 5460 -590
rect 5700 -590 5710 -589
rect 5760 -590 5770 -589
rect 5700 -649 5770 -590
rect 6010 -590 6020 -589
rect 6080 -590 6090 -589
rect 6010 -649 6090 -590
rect 6330 -590 6340 -589
rect 6390 -590 6400 -589
rect 6330 -649 6400 -590
rect 6640 -590 6650 -589
rect 6710 -590 6720 -589
rect 6640 -649 6720 -590
rect 6960 -590 6970 -589
rect 7030 -590 7040 -589
rect 6960 -649 7040 -590
rect 7280 -649 7290 -589
rect 7340 -649 7350 -589
rect 7590 -649 7600 -589
rect 7660 -649 7670 -589
rect 7910 -649 7920 -589
rect 7970 -649 7980 -589
rect 8220 -649 8230 -589
rect 8290 -649 8300 -589
rect 8540 -649 8550 -589
rect 8610 -604 8620 -589
rect 8609 -649 8620 -604
rect 8860 -649 8870 -589
rect 8920 -649 8930 -589
rect 9170 -649 9180 -589
rect 9240 -649 9250 -589
rect 9490 -649 9500 -589
rect 9550 -649 9560 -589
rect 9800 -649 9810 -589
rect 4810 -650 7290 -649
rect 7345 -650 7437 -649
rect 7503 -650 7595 -649
rect 7661 -650 7753 -649
rect 7819 -650 7911 -649
rect 7977 -650 8069 -649
rect 8135 -650 8227 -649
rect 8293 -650 8385 -649
rect 8451 -650 8543 -649
rect 8609 -650 8701 -649
rect 8767 -650 8859 -649
rect 8925 -650 9017 -649
rect 9083 -650 9175 -649
rect 9241 -650 9333 -649
rect 9399 -650 9491 -649
rect 9557 -650 9649 -649
rect 9715 -650 9807 -649
rect 4755 -708 4810 -678
rect 4755 -1478 4810 -1448
rect 4913 -708 4968 -678
rect 4913 -1478 4968 -1448
rect 5071 -708 5126 -678
rect 5071 -1478 5126 -1448
rect 5229 -708 5284 -678
rect 5229 -1478 5284 -1448
rect 5387 -708 5442 -678
rect 5387 -1478 5442 -1448
rect 5545 -708 5600 -678
rect 5545 -1478 5600 -1448
rect 5703 -708 5758 -678
rect 5703 -1478 5758 -1448
rect 5861 -708 5916 -678
rect 5861 -1478 5916 -1448
rect 6019 -708 6074 -678
rect 6019 -1478 6074 -1448
rect 6177 -708 6232 -678
rect 6177 -1478 6232 -1448
rect 6335 -708 6390 -678
rect 6335 -1478 6390 -1448
rect 6493 -708 6548 -678
rect 6493 -1478 6548 -1448
rect 6651 -708 6706 -678
rect 6651 -1478 6706 -1448
rect 6809 -708 6864 -678
rect 6809 -1478 6864 -1448
rect 6967 -708 7022 -678
rect 6967 -1478 7022 -1448
rect 7125 -708 7180 -678
rect 7125 -1478 7180 -1448
rect 7283 -708 7338 -678
rect 7283 -1478 7338 -1448
rect 7441 -708 7496 -678
rect 7441 -1478 7496 -1448
rect 7599 -708 7654 -678
rect 7599 -1478 7654 -1448
rect 7757 -708 7812 -678
rect 7757 -1478 7812 -1448
rect 7915 -708 7970 -678
rect 7915 -1478 7970 -1448
rect 8073 -708 8128 -678
rect 8073 -1478 8128 -1448
rect 8231 -708 8286 -678
rect 8231 -1478 8286 -1448
rect 8389 -708 8444 -678
rect 8389 -1478 8444 -1448
rect 8547 -708 8602 -678
rect 8547 -1478 8602 -1448
rect 8705 -708 8760 -678
rect 8705 -1478 8760 -1448
rect 8863 -708 8918 -678
rect 8863 -1478 8918 -1448
rect 9021 -708 9076 -678
rect 9021 -1478 9076 -1448
rect 9179 -708 9234 -678
rect 9179 -1478 9234 -1448
rect 9337 -708 9392 -678
rect 9337 -1478 9392 -1448
rect 9495 -708 9550 -678
rect 9495 -1478 9550 -1448
rect 9653 -708 9708 -678
rect 9653 -1478 9708 -1448
rect 9811 -708 9866 -678
rect 9811 -1478 9866 -1448
rect 4810 -1570 4820 -1510
rect 5060 -1570 5070 -1510
rect 5130 -1570 5140 -1510
rect 5380 -1570 5390 -1510
rect 5450 -1525 5460 -1510
rect 5449 -1570 5460 -1525
rect 5700 -1570 5710 -1510
rect 5760 -1570 5770 -1510
rect 6010 -1570 6020 -1510
rect 6080 -1570 6090 -1510
rect 6330 -1570 6340 -1510
rect 6390 -1570 6400 -1510
rect 6640 -1570 6650 -1510
rect 6710 -1570 6720 -1510
rect 6960 -1570 6970 -1510
rect 7030 -1525 7040 -1510
rect 7029 -1570 7040 -1525
rect 7280 -1570 7290 -1510
rect 7340 -1570 7350 -1510
rect 7590 -1570 7600 -1510
rect 7660 -1570 7670 -1510
rect 7910 -1570 7920 -1510
rect 7970 -1570 7980 -1510
rect 8220 -1570 8230 -1510
rect 8290 -1570 8300 -1510
rect 8540 -1570 8550 -1510
rect 8610 -1525 8620 -1510
rect 8609 -1570 8620 -1525
rect 8860 -1570 8870 -1510
rect 8920 -1570 8930 -1510
rect 9170 -1570 9180 -1510
rect 9240 -1570 9250 -1510
rect 9490 -1570 9500 -1510
rect 9550 -1570 9560 -1510
rect 9800 -1570 9810 -1510
rect 4817 -1571 4909 -1570
rect 4975 -1571 5067 -1570
rect 5133 -1571 5225 -1570
rect 5291 -1571 5383 -1570
rect 5449 -1571 5541 -1570
rect 5607 -1571 5699 -1570
rect 5765 -1571 5857 -1570
rect 5923 -1571 6015 -1570
rect 6081 -1571 6173 -1570
rect 6239 -1571 6331 -1570
rect 6397 -1571 6489 -1570
rect 6555 -1571 6647 -1570
rect 6713 -1571 6805 -1570
rect 6871 -1571 6963 -1570
rect 7029 -1571 7121 -1570
rect 7187 -1571 7279 -1570
rect 7345 -1571 7437 -1570
rect 7503 -1571 7595 -1570
rect 7661 -1571 7753 -1570
rect 7819 -1571 7911 -1570
rect 7977 -1571 8069 -1570
rect 8135 -1571 8227 -1570
rect 8293 -1571 8385 -1570
rect 8451 -1571 8543 -1570
rect 8609 -1571 8701 -1570
rect 8767 -1571 8859 -1570
rect 8925 -1571 9017 -1570
rect 9083 -1571 9175 -1570
rect 9241 -1571 9333 -1570
rect 9399 -1571 9491 -1570
rect 9557 -1571 9649 -1570
rect 9715 -1571 9807 -1570
rect 4810 -1667 4820 -1607
rect 5060 -1667 5070 -1607
rect 5130 -1667 5140 -1607
rect 5380 -1667 5390 -1607
rect 5450 -1622 5460 -1607
rect 5449 -1667 5460 -1622
rect 5700 -1667 5710 -1607
rect 5760 -1667 5770 -1607
rect 6010 -1667 6020 -1607
rect 6080 -1667 6090 -1607
rect 6330 -1667 6340 -1607
rect 6390 -1667 6400 -1607
rect 6640 -1667 6650 -1607
rect 6710 -1667 6720 -1607
rect 6960 -1667 6970 -1607
rect 7030 -1622 7040 -1607
rect 7029 -1667 7040 -1622
rect 7280 -1667 7290 -1607
rect 7340 -1667 7350 -1607
rect 7590 -1667 7600 -1607
rect 7660 -1667 7670 -1607
rect 7910 -1667 7920 -1607
rect 7970 -1667 7980 -1607
rect 8220 -1667 8230 -1607
rect 8290 -1667 8300 -1607
rect 8540 -1667 8550 -1607
rect 8610 -1622 8620 -1607
rect 8609 -1667 8620 -1622
rect 8860 -1667 8870 -1607
rect 8920 -1667 8930 -1607
rect 9170 -1667 9180 -1607
rect 9240 -1667 9250 -1607
rect 9490 -1667 9500 -1607
rect 9550 -1667 9560 -1607
rect 9800 -1667 9810 -1607
rect 4817 -1668 4909 -1667
rect 4975 -1668 5067 -1667
rect 5133 -1668 5225 -1667
rect 5291 -1668 5383 -1667
rect 5449 -1668 5541 -1667
rect 5607 -1668 5699 -1667
rect 5765 -1668 5857 -1667
rect 5923 -1668 6015 -1667
rect 6081 -1668 6173 -1667
rect 6239 -1668 6331 -1667
rect 6397 -1668 6489 -1667
rect 6555 -1668 6647 -1667
rect 6713 -1668 6805 -1667
rect 6871 -1668 6963 -1667
rect 7029 -1668 7121 -1667
rect 7187 -1668 7279 -1667
rect 7345 -1668 7437 -1667
rect 7503 -1668 7595 -1667
rect 7661 -1668 7753 -1667
rect 7819 -1668 7911 -1667
rect 7977 -1668 8069 -1667
rect 8135 -1668 8227 -1667
rect 8293 -1668 8385 -1667
rect 8451 -1668 8543 -1667
rect 8609 -1668 8701 -1667
rect 8767 -1668 8859 -1667
rect 8925 -1668 9017 -1667
rect 9083 -1668 9175 -1667
rect 9241 -1668 9333 -1667
rect 9399 -1668 9491 -1667
rect 9557 -1668 9649 -1667
rect 9715 -1668 9807 -1667
rect 4755 -1726 4810 -1696
rect 4755 -2496 4810 -2466
rect 4913 -1726 4968 -1696
rect 4913 -2496 4968 -2466
rect 5071 -1726 5126 -1696
rect 5071 -2496 5126 -2466
rect 5229 -1726 5284 -1696
rect 5229 -2496 5284 -2466
rect 5387 -1726 5442 -1696
rect 5387 -2496 5442 -2466
rect 5545 -1726 5600 -1696
rect 5545 -2496 5600 -2466
rect 5703 -1726 5758 -1696
rect 5703 -2496 5758 -2466
rect 5861 -1726 5916 -1696
rect 5861 -2496 5916 -2466
rect 6019 -1726 6074 -1696
rect 6019 -2496 6074 -2466
rect 6177 -1726 6232 -1696
rect 6177 -2496 6232 -2466
rect 6335 -1726 6390 -1696
rect 6335 -2496 6390 -2466
rect 6493 -1726 6548 -1696
rect 6493 -2496 6548 -2466
rect 6651 -1726 6706 -1696
rect 6651 -2496 6706 -2466
rect 6809 -1726 6864 -1696
rect 6809 -2496 6864 -2466
rect 6967 -1726 7022 -1696
rect 6967 -2496 7022 -2466
rect 7125 -1726 7180 -1696
rect 7125 -2496 7180 -2466
rect 7283 -1726 7338 -1696
rect 7283 -2496 7338 -2466
rect 7441 -1726 7496 -1696
rect 7441 -2496 7496 -2466
rect 7599 -1726 7654 -1696
rect 7599 -2496 7654 -2466
rect 7757 -1726 7812 -1696
rect 7757 -2496 7812 -2466
rect 7915 -1726 7970 -1696
rect 7915 -2496 7970 -2466
rect 8073 -1726 8128 -1696
rect 8073 -2496 8128 -2466
rect 8231 -1726 8286 -1696
rect 8231 -2496 8286 -2466
rect 8389 -1726 8444 -1696
rect 8389 -2496 8444 -2466
rect 8547 -1726 8602 -1696
rect 8547 -2496 8602 -2466
rect 8705 -1726 8760 -1696
rect 8705 -2496 8760 -2466
rect 8863 -1726 8918 -1696
rect 8863 -2496 8918 -2466
rect 9021 -1726 9076 -1696
rect 9021 -2496 9076 -2466
rect 9179 -1726 9234 -1696
rect 9179 -2496 9234 -2466
rect 9337 -1726 9392 -1696
rect 9337 -2496 9392 -2466
rect 9495 -1726 9550 -1696
rect 9495 -2496 9550 -2466
rect 9653 -1726 9708 -1696
rect 9653 -2496 9708 -2466
rect 9811 -1726 9866 -1696
rect 9811 -2496 9866 -2466
rect 4810 -2590 4820 -2530
rect 5060 -2590 5070 -2530
rect 5130 -2590 5140 -2530
rect 5380 -2590 5390 -2530
rect 5450 -2545 5460 -2530
rect 5449 -2590 5460 -2545
rect 5700 -2590 5710 -2530
rect 5760 -2590 5770 -2530
rect 6010 -2590 6020 -2530
rect 6080 -2590 6090 -2530
rect 6330 -2590 6340 -2530
rect 6390 -2590 6400 -2530
rect 6640 -2590 6650 -2530
rect 6710 -2590 6720 -2530
rect 6960 -2590 6970 -2530
rect 7030 -2545 7040 -2530
rect 7029 -2590 7040 -2545
rect 7280 -2590 7290 -2530
rect 7340 -2590 7350 -2530
rect 7590 -2590 7600 -2530
rect 7660 -2590 7670 -2530
rect 7910 -2590 7920 -2530
rect 7970 -2590 7980 -2530
rect 8220 -2590 8230 -2530
rect 8290 -2590 8300 -2530
rect 8540 -2590 8550 -2530
rect 8610 -2545 8620 -2530
rect 8609 -2590 8620 -2545
rect 8860 -2590 8870 -2530
rect 8920 -2590 8930 -2530
rect 9170 -2590 9180 -2530
rect 9240 -2590 9250 -2530
rect 9490 -2590 9500 -2530
rect 9550 -2590 9560 -2530
rect 9800 -2590 9810 -2530
rect 4817 -2591 4909 -2590
rect 4975 -2591 5067 -2590
rect 5133 -2591 5225 -2590
rect 5291 -2591 5383 -2590
rect 5449 -2591 5541 -2590
rect 5607 -2591 5699 -2590
rect 5765 -2591 5857 -2590
rect 5923 -2591 6015 -2590
rect 6081 -2591 6173 -2590
rect 6239 -2591 6331 -2590
rect 6397 -2591 6489 -2590
rect 6555 -2591 6647 -2590
rect 6713 -2591 6805 -2590
rect 6871 -2591 6963 -2590
rect 7029 -2591 7121 -2590
rect 7187 -2591 7279 -2590
rect 7345 -2591 7437 -2590
rect 7503 -2591 7595 -2590
rect 7661 -2591 7753 -2590
rect 7819 -2591 7911 -2590
rect 7977 -2591 8069 -2590
rect 8135 -2591 8227 -2590
rect 8293 -2591 8385 -2590
rect 8451 -2591 8543 -2590
rect 8609 -2591 8701 -2590
rect 8767 -2591 8859 -2590
rect 8925 -2591 9017 -2590
rect 9083 -2591 9175 -2590
rect 9241 -2591 9333 -2590
rect 9399 -2591 9491 -2590
rect 9557 -2591 9649 -2590
rect 9715 -2591 9807 -2590
rect 4810 -2684 4820 -2624
rect 5060 -2684 5070 -2624
rect 5130 -2684 5140 -2624
rect 5380 -2684 5390 -2624
rect 5450 -2639 5460 -2624
rect 5449 -2684 5460 -2639
rect 5700 -2684 5710 -2624
rect 5760 -2684 5770 -2624
rect 6010 -2684 6020 -2624
rect 6080 -2684 6090 -2624
rect 6330 -2684 6340 -2624
rect 6390 -2684 6400 -2624
rect 6640 -2684 6650 -2624
rect 6710 -2684 6720 -2624
rect 6960 -2684 6970 -2624
rect 7030 -2639 7040 -2624
rect 7029 -2684 7040 -2639
rect 7280 -2684 7290 -2624
rect 7340 -2684 7350 -2624
rect 7590 -2684 7600 -2624
rect 7660 -2684 7670 -2624
rect 7910 -2684 7920 -2624
rect 7970 -2684 7980 -2624
rect 8220 -2684 8230 -2624
rect 8290 -2684 8300 -2624
rect 8540 -2684 8550 -2624
rect 8610 -2639 8620 -2624
rect 8609 -2684 8620 -2639
rect 8860 -2684 8870 -2624
rect 8920 -2684 8930 -2624
rect 9170 -2684 9180 -2624
rect 9240 -2684 9250 -2624
rect 9490 -2684 9500 -2624
rect 9550 -2684 9560 -2624
rect 9800 -2684 9810 -2624
rect 4817 -2685 4909 -2684
rect 4975 -2685 5067 -2684
rect 5133 -2685 5225 -2684
rect 5291 -2685 5383 -2684
rect 5449 -2685 5541 -2684
rect 5607 -2685 5699 -2684
rect 5765 -2685 5857 -2684
rect 5923 -2685 6015 -2684
rect 6081 -2685 6173 -2684
rect 6239 -2685 6331 -2684
rect 6397 -2685 6489 -2684
rect 6555 -2685 6647 -2684
rect 6713 -2685 6805 -2684
rect 6871 -2685 6963 -2684
rect 7029 -2685 7121 -2684
rect 7187 -2685 7279 -2684
rect 7345 -2685 7437 -2684
rect 7503 -2685 7595 -2684
rect 7661 -2685 7753 -2684
rect 7819 -2685 7911 -2684
rect 7977 -2685 8069 -2684
rect 8135 -2685 8227 -2684
rect 8293 -2685 8385 -2684
rect 8451 -2685 8543 -2684
rect 8609 -2685 8701 -2684
rect 8767 -2685 8859 -2684
rect 8925 -2685 9017 -2684
rect 9083 -2685 9175 -2684
rect 9241 -2685 9333 -2684
rect 9399 -2685 9491 -2684
rect 9557 -2685 9649 -2684
rect 9715 -2685 9807 -2684
rect 4755 -2744 4810 -2714
rect 4755 -3514 4810 -3484
rect 4913 -2744 4968 -2714
rect 4913 -3514 4968 -3484
rect 5071 -2744 5126 -2714
rect 5071 -3514 5126 -3484
rect 5229 -2744 5284 -2714
rect 5229 -3514 5284 -3484
rect 5387 -2744 5442 -2714
rect 5387 -3514 5442 -3484
rect 5545 -2744 5600 -2714
rect 5545 -3514 5600 -3484
rect 5703 -2744 5758 -2714
rect 5703 -3514 5758 -3484
rect 5861 -2744 5916 -2714
rect 5861 -3514 5916 -3484
rect 6019 -2744 6074 -2714
rect 6019 -3514 6074 -3484
rect 6177 -2744 6232 -2714
rect 6177 -3514 6232 -3484
rect 6335 -2744 6390 -2714
rect 6335 -3514 6390 -3484
rect 6493 -2744 6548 -2714
rect 6493 -3514 6548 -3484
rect 6651 -2744 6706 -2714
rect 6651 -3514 6706 -3484
rect 6809 -2744 6864 -2714
rect 6809 -3514 6864 -3484
rect 6967 -2744 7022 -2714
rect 6967 -3514 7022 -3484
rect 7125 -2744 7180 -2714
rect 7125 -3514 7180 -3484
rect 7283 -2744 7338 -2714
rect 7283 -3514 7338 -3484
rect 7441 -2744 7496 -2714
rect 7441 -3514 7496 -3484
rect 7599 -2744 7654 -2714
rect 7599 -3514 7654 -3484
rect 7757 -2744 7812 -2714
rect 7757 -3514 7812 -3484
rect 7915 -2744 7970 -2714
rect 7915 -3514 7970 -3484
rect 8073 -2744 8128 -2714
rect 8073 -3514 8128 -3484
rect 8231 -2744 8286 -2714
rect 8231 -3514 8286 -3484
rect 8389 -2744 8444 -2714
rect 8389 -3514 8444 -3484
rect 8547 -2744 8602 -2714
rect 8547 -3514 8602 -3484
rect 8705 -2744 8760 -2714
rect 8705 -3514 8760 -3484
rect 8863 -2744 8918 -2714
rect 8863 -3514 8918 -3484
rect 9021 -2744 9076 -2714
rect 9021 -3514 9076 -3484
rect 9179 -2744 9234 -2714
rect 9179 -3514 9234 -3484
rect 9337 -2744 9392 -2714
rect 9337 -3514 9392 -3484
rect 9495 -2744 9550 -2714
rect 9495 -3514 9550 -3484
rect 9653 -2744 9708 -2714
rect 9653 -3514 9708 -3484
rect 9811 -2744 9866 -2714
rect 9811 -3514 9866 -3484
rect 4810 -3610 4820 -3550
rect 5060 -3610 5070 -3550
rect 5130 -3610 5140 -3550
rect 5380 -3610 5390 -3550
rect 5450 -3565 5460 -3550
rect 5449 -3610 5460 -3565
rect 5700 -3610 5710 -3550
rect 5760 -3610 5770 -3550
rect 6010 -3610 6020 -3550
rect 6080 -3610 6090 -3550
rect 6330 -3610 6340 -3550
rect 6390 -3610 6400 -3550
rect 6640 -3610 6650 -3550
rect 6710 -3610 6720 -3550
rect 6960 -3610 6970 -3550
rect 7030 -3565 7040 -3550
rect 7029 -3610 7040 -3565
rect 7280 -3610 7290 -3550
rect 7340 -3610 7350 -3550
rect 7590 -3610 7600 -3550
rect 7660 -3610 7670 -3550
rect 7910 -3610 7920 -3550
rect 7970 -3610 7980 -3550
rect 8220 -3610 8230 -3550
rect 8290 -3610 8300 -3550
rect 8540 -3610 8550 -3550
rect 8610 -3565 8620 -3550
rect 8609 -3610 8620 -3565
rect 8860 -3610 8870 -3550
rect 8920 -3610 8930 -3550
rect 9170 -3610 9180 -3550
rect 9240 -3610 9250 -3550
rect 9490 -3610 9500 -3550
rect 9550 -3610 9560 -3550
rect 9800 -3610 9810 -3550
rect 4817 -3611 4909 -3610
rect 4975 -3611 5067 -3610
rect 5133 -3611 5225 -3610
rect 5291 -3611 5383 -3610
rect 5449 -3611 5541 -3610
rect 5607 -3611 5699 -3610
rect 5765 -3611 5857 -3610
rect 5923 -3611 6015 -3610
rect 6081 -3611 6173 -3610
rect 6239 -3611 6331 -3610
rect 6397 -3611 6489 -3610
rect 6555 -3611 6647 -3610
rect 6713 -3611 6805 -3610
rect 6871 -3611 6963 -3610
rect 7029 -3611 7121 -3610
rect 7187 -3611 7279 -3610
rect 7345 -3611 7437 -3610
rect 7503 -3611 7595 -3610
rect 7661 -3611 7753 -3610
rect 7819 -3611 7911 -3610
rect 7977 -3611 8069 -3610
rect 8135 -3611 8227 -3610
rect 8293 -3611 8385 -3610
rect 8451 -3611 8543 -3610
rect 8609 -3611 8701 -3610
rect 8767 -3611 8859 -3610
rect 8925 -3611 9017 -3610
rect 9083 -3611 9175 -3610
rect 9241 -3611 9333 -3610
rect 9399 -3611 9491 -3610
rect 9557 -3611 9649 -3610
rect 9715 -3611 9807 -3610
rect 4620 -3680 4690 -3650
rect 9940 -3650 9950 460
rect 9990 -3650 10010 460
rect 9940 -3680 10010 -3650
rect 4620 -3690 10010 -3680
rect 4620 -3730 4720 -3690
rect 9900 -3730 10010 -3690
rect 4620 -3740 10010 -3730
rect 4220 -4060 4280 -4020
rect 10440 -4060 10480 -4020
rect 4220 -4080 4380 -4060
rect 10420 -4080 10480 -4060
rect 10520 -4120 10540 920
rect 4160 -4140 4380 -4120
rect 10420 -4140 10540 -4120
<< via1 >>
rect 4280 920 10420 940
rect 4280 880 10420 920
rect 4280 860 10420 880
rect 4200 -4020 4220 820
rect 4220 -4020 4280 820
rect 4660 560 9880 580
rect 4660 500 9880 560
rect 4660 480 9880 500
rect 4820 370 5060 430
rect 5140 370 5380 430
rect 5460 370 5700 430
rect 5770 370 6010 430
rect 6090 370 6330 430
rect 6400 370 6640 430
rect 6720 370 6960 430
rect 7040 370 7280 430
rect 7350 370 7590 430
rect 7670 370 7910 430
rect 7980 370 8220 430
rect 8300 370 8540 430
rect 8620 370 8860 430
rect 8930 370 9170 430
rect 9250 370 9490 430
rect 9560 370 9800 430
rect 4755 -430 4810 310
rect 4913 -430 4968 310
rect 5071 -430 5126 310
rect 5229 -430 5284 310
rect 5387 -430 5442 310
rect 5545 -430 5600 310
rect 5703 -430 5758 310
rect 5861 -430 5916 310
rect 6019 -430 6074 310
rect 6177 -430 6232 310
rect 6335 -430 6390 310
rect 6493 -430 6548 310
rect 6651 -430 6706 310
rect 6809 -430 6864 310
rect 6967 -430 7022 310
rect 7125 -430 7180 310
rect 7283 -430 7338 310
rect 7441 -430 7496 310
rect 7599 -430 7654 310
rect 7757 -430 7812 310
rect 7915 -430 7970 310
rect 8073 -430 8128 310
rect 8231 -430 8286 310
rect 8389 -430 8444 310
rect 8547 -430 8602 310
rect 8705 -430 8760 310
rect 8863 -430 8918 310
rect 9021 -430 9076 310
rect 9179 -430 9234 310
rect 9337 -430 9392 310
rect 9495 -430 9550 310
rect 9653 -430 9708 310
rect 9811 -430 9866 310
rect 4820 -560 5060 -500
rect 5140 -560 5380 -500
rect 5460 -560 5700 -500
rect 5770 -560 6010 -500
rect 6090 -560 6330 -500
rect 6400 -560 6640 -500
rect 6720 -560 6960 -500
rect 7040 -560 7280 -500
rect 7350 -560 7590 -500
rect 7670 -560 7910 -500
rect 7980 -560 8220 -500
rect 8300 -560 8540 -500
rect 8620 -560 8860 -500
rect 8930 -560 9170 -500
rect 9250 -560 9490 -500
rect 9560 -560 9800 -500
rect 4820 -649 5060 -589
rect 5140 -649 5380 -589
rect 5460 -649 5700 -589
rect 5770 -649 6010 -589
rect 6090 -649 6330 -589
rect 6400 -649 6640 -589
rect 6720 -649 6960 -589
rect 7040 -649 7280 -589
rect 7350 -649 7590 -589
rect 7670 -649 7910 -589
rect 7980 -649 8220 -589
rect 8300 -649 8540 -589
rect 8620 -649 8860 -589
rect 8930 -649 9170 -589
rect 9250 -649 9490 -589
rect 9560 -649 9800 -589
rect 4755 -1448 4810 -708
rect 4913 -1448 4968 -708
rect 5071 -1448 5126 -708
rect 5229 -1448 5284 -708
rect 5387 -1448 5442 -708
rect 5545 -1448 5600 -708
rect 5703 -1448 5758 -708
rect 5861 -1448 5916 -708
rect 6019 -1448 6074 -708
rect 6177 -1448 6232 -708
rect 6335 -1448 6390 -708
rect 6493 -1448 6548 -708
rect 6651 -1448 6706 -708
rect 6809 -1448 6864 -708
rect 6967 -1448 7022 -708
rect 7125 -1448 7180 -708
rect 7283 -1448 7338 -708
rect 7441 -1448 7496 -708
rect 7599 -1448 7654 -708
rect 7757 -1448 7812 -708
rect 7915 -1448 7970 -708
rect 8073 -1448 8128 -708
rect 8231 -1448 8286 -708
rect 8389 -1448 8444 -708
rect 8547 -1448 8602 -708
rect 8705 -1448 8760 -708
rect 8863 -1448 8918 -708
rect 9021 -1448 9076 -708
rect 9179 -1448 9234 -708
rect 9337 -1448 9392 -708
rect 9495 -1448 9550 -708
rect 9653 -1448 9708 -708
rect 9811 -1448 9866 -708
rect 4820 -1570 5060 -1510
rect 5140 -1570 5380 -1510
rect 5460 -1570 5700 -1510
rect 5770 -1570 6010 -1510
rect 6090 -1570 6330 -1510
rect 6400 -1570 6640 -1510
rect 6720 -1570 6960 -1510
rect 7040 -1570 7280 -1510
rect 7350 -1570 7590 -1510
rect 7670 -1570 7910 -1510
rect 7980 -1570 8220 -1510
rect 8300 -1570 8540 -1510
rect 8620 -1570 8860 -1510
rect 8930 -1570 9170 -1510
rect 9250 -1570 9490 -1510
rect 9560 -1570 9800 -1510
rect 4820 -1667 5060 -1607
rect 5140 -1667 5380 -1607
rect 5460 -1667 5700 -1607
rect 5770 -1667 6010 -1607
rect 6090 -1667 6330 -1607
rect 6400 -1667 6640 -1607
rect 6720 -1667 6960 -1607
rect 7040 -1667 7280 -1607
rect 7350 -1667 7590 -1607
rect 7670 -1667 7910 -1607
rect 7980 -1667 8220 -1607
rect 8300 -1667 8540 -1607
rect 8620 -1667 8860 -1607
rect 8930 -1667 9170 -1607
rect 9250 -1667 9490 -1607
rect 9560 -1667 9800 -1607
rect 4755 -2466 4810 -1726
rect 4913 -2466 4968 -1726
rect 5071 -2466 5126 -1726
rect 5229 -2466 5284 -1726
rect 5387 -2466 5442 -1726
rect 5545 -2466 5600 -1726
rect 5703 -2466 5758 -1726
rect 5861 -2466 5916 -1726
rect 6019 -2466 6074 -1726
rect 6177 -2466 6232 -1726
rect 6335 -2466 6390 -1726
rect 6493 -2466 6548 -1726
rect 6651 -2466 6706 -1726
rect 6809 -2466 6864 -1726
rect 6967 -2466 7022 -1726
rect 7125 -2466 7180 -1726
rect 7283 -2466 7338 -1726
rect 7441 -2466 7496 -1726
rect 7599 -2466 7654 -1726
rect 7757 -2466 7812 -1726
rect 7915 -2466 7970 -1726
rect 8073 -2466 8128 -1726
rect 8231 -2466 8286 -1726
rect 8389 -2466 8444 -1726
rect 8547 -2466 8602 -1726
rect 8705 -2466 8760 -1726
rect 8863 -2466 8918 -1726
rect 9021 -2466 9076 -1726
rect 9179 -2466 9234 -1726
rect 9337 -2466 9392 -1726
rect 9495 -2466 9550 -1726
rect 9653 -2466 9708 -1726
rect 9811 -2466 9866 -1726
rect 4820 -2590 5060 -2530
rect 5140 -2590 5380 -2530
rect 5460 -2590 5700 -2530
rect 5770 -2590 6010 -2530
rect 6090 -2590 6330 -2530
rect 6400 -2590 6640 -2530
rect 6720 -2590 6960 -2530
rect 7040 -2590 7280 -2530
rect 7350 -2590 7590 -2530
rect 7670 -2590 7910 -2530
rect 7980 -2590 8220 -2530
rect 8300 -2590 8540 -2530
rect 8620 -2590 8860 -2530
rect 8930 -2590 9170 -2530
rect 9250 -2590 9490 -2530
rect 9560 -2590 9800 -2530
rect 4820 -2684 5060 -2624
rect 5140 -2684 5380 -2624
rect 5460 -2684 5700 -2624
rect 5770 -2684 6010 -2624
rect 6090 -2684 6330 -2624
rect 6400 -2684 6640 -2624
rect 6720 -2684 6960 -2624
rect 7040 -2684 7280 -2624
rect 7350 -2684 7590 -2624
rect 7670 -2684 7910 -2624
rect 7980 -2684 8220 -2624
rect 8300 -2684 8540 -2624
rect 8620 -2684 8860 -2624
rect 8930 -2684 9170 -2624
rect 9250 -2684 9490 -2624
rect 9560 -2684 9800 -2624
rect 4755 -3484 4810 -2744
rect 4913 -3484 4968 -2744
rect 5071 -3484 5126 -2744
rect 5229 -3484 5284 -2744
rect 5387 -3484 5442 -2744
rect 5545 -3484 5600 -2744
rect 5703 -3484 5758 -2744
rect 5861 -3484 5916 -2744
rect 6019 -3484 6074 -2744
rect 6177 -3484 6232 -2744
rect 6335 -3484 6390 -2744
rect 6493 -3484 6548 -2744
rect 6651 -3484 6706 -2744
rect 6809 -3484 6864 -2744
rect 6967 -3484 7022 -2744
rect 7125 -3484 7180 -2744
rect 7283 -3484 7338 -2744
rect 7441 -3484 7496 -2744
rect 7599 -3484 7654 -2744
rect 7757 -3484 7812 -2744
rect 7915 -3484 7970 -2744
rect 8073 -3484 8128 -2744
rect 8231 -3484 8286 -2744
rect 8389 -3484 8444 -2744
rect 8547 -3484 8602 -2744
rect 8705 -3484 8760 -2744
rect 8863 -3484 8918 -2744
rect 9021 -3484 9076 -2744
rect 9179 -3484 9234 -2744
rect 9337 -3484 9392 -2744
rect 9495 -3484 9550 -2744
rect 9653 -3484 9708 -2744
rect 9811 -3484 9866 -2744
rect 4820 -3610 5060 -3550
rect 5140 -3610 5380 -3550
rect 5460 -3610 5700 -3550
rect 5770 -3610 6010 -3550
rect 6090 -3610 6330 -3550
rect 6400 -3610 6640 -3550
rect 6720 -3610 6960 -3550
rect 7040 -3610 7280 -3550
rect 7350 -3610 7590 -3550
rect 7670 -3610 7910 -3550
rect 7980 -3610 8220 -3550
rect 8300 -3610 8540 -3550
rect 8620 -3610 8860 -3550
rect 8930 -3610 9170 -3550
rect 9250 -3610 9490 -3550
rect 9560 -3610 9800 -3550
rect 10440 -4020 10480 820
rect 10480 -4020 10520 820
rect 4380 -4080 10420 -4060
rect 4380 -4120 10420 -4080
rect 4380 -4140 10420 -4120
<< metal2 >>
rect 4200 820 4280 940
rect 10420 860 10520 940
rect 10440 820 10520 860
rect 4640 640 9920 660
rect 4640 480 4660 640
rect 9880 480 9920 640
rect 4470 430 4820 450
rect 9820 430 10160 450
rect 4470 -3610 4480 430
rect 4560 370 4820 430
rect 5060 370 5140 430
rect 5380 370 5460 430
rect 5700 370 5770 430
rect 6010 370 6090 430
rect 6330 370 6400 430
rect 6640 370 6720 430
rect 6960 370 7040 430
rect 7280 370 7290 430
rect 7340 370 7350 430
rect 7590 370 7670 430
rect 7910 370 7980 430
rect 8220 370 8300 430
rect 8540 370 8620 430
rect 8860 370 8930 430
rect 9170 370 9250 430
rect 9490 370 9560 430
rect 9800 370 10070 430
rect 4560 -500 4570 370
rect 4755 310 4815 340
rect 4811 -430 4815 310
rect 4755 -460 4815 -430
rect 4913 310 4973 340
rect 4969 -430 4973 310
rect 4913 -460 4973 -430
rect 5071 310 5131 340
rect 5127 -430 5131 310
rect 5071 -460 5131 -430
rect 5229 310 5289 340
rect 5285 -430 5289 310
rect 5229 -460 5289 -430
rect 5387 310 5447 340
rect 5443 -430 5447 310
rect 5387 -460 5447 -430
rect 5545 310 5605 340
rect 5601 -430 5605 310
rect 5545 -460 5605 -430
rect 5703 310 5763 340
rect 5759 -430 5763 310
rect 5703 -460 5763 -430
rect 5861 310 5921 340
rect 5917 -430 5921 310
rect 5861 -460 5921 -430
rect 6019 310 6079 340
rect 6075 -430 6079 310
rect 6019 -460 6079 -430
rect 6177 310 6237 340
rect 6233 -430 6237 310
rect 6177 -460 6237 -430
rect 6335 310 6395 340
rect 6391 -430 6395 310
rect 6335 -460 6395 -430
rect 6493 310 6553 340
rect 6549 -430 6553 310
rect 6493 -460 6553 -430
rect 6651 310 6711 340
rect 6707 -430 6711 310
rect 6651 -460 6711 -430
rect 6809 310 6869 340
rect 6865 -430 6869 310
rect 6809 -460 6869 -430
rect 6967 310 7027 340
rect 7023 -430 7027 310
rect 6967 -460 7027 -430
rect 7125 310 7185 340
rect 7181 -430 7185 310
rect 7125 -460 7185 -430
rect 7283 310 7343 340
rect 7339 -430 7343 310
rect 7283 -460 7343 -430
rect 7441 310 7501 340
rect 7497 -430 7501 310
rect 7441 -460 7501 -430
rect 7599 310 7659 340
rect 7655 -430 7659 310
rect 7599 -460 7659 -430
rect 7757 310 7817 340
rect 7813 -430 7817 310
rect 7757 -460 7817 -430
rect 7915 310 7975 340
rect 7971 -430 7975 310
rect 7915 -460 7975 -430
rect 8073 310 8133 340
rect 8129 -430 8133 310
rect 8073 -460 8133 -430
rect 8231 310 8291 340
rect 8287 -430 8291 310
rect 8231 -460 8291 -430
rect 8389 310 8449 340
rect 8445 -430 8449 310
rect 8389 -460 8449 -430
rect 8547 310 8607 340
rect 8603 -430 8607 310
rect 8547 -460 8607 -430
rect 8705 310 8765 340
rect 8761 -430 8765 310
rect 8705 -460 8765 -430
rect 8863 310 8923 340
rect 8919 -430 8923 310
rect 8863 -460 8923 -430
rect 9021 310 9081 340
rect 9077 -430 9081 310
rect 9021 -460 9081 -430
rect 9179 310 9239 340
rect 9235 -430 9239 310
rect 9179 -460 9239 -430
rect 9337 310 9397 340
rect 9393 -430 9397 310
rect 9337 -460 9397 -430
rect 9495 310 9555 340
rect 9551 -430 9555 310
rect 9495 -460 9555 -430
rect 9653 310 9713 340
rect 9709 -430 9713 310
rect 9653 -460 9713 -430
rect 9811 310 9871 340
rect 9867 -430 9871 310
rect 9811 -460 9871 -430
rect 10060 -500 10070 370
rect 4560 -560 4820 -500
rect 5060 -560 5140 -500
rect 5380 -560 5460 -500
rect 5700 -560 5770 -500
rect 6010 -560 6090 -500
rect 6330 -560 6400 -500
rect 6640 -560 6720 -500
rect 6960 -560 7040 -500
rect 7280 -560 7290 -500
rect 4560 -589 7290 -560
rect 4560 -649 4820 -589
rect 5060 -611 5140 -589
rect 5060 -649 5070 -611
rect 5130 -649 5140 -611
rect 5380 -611 5460 -589
rect 5380 -649 5390 -611
rect 5450 -649 5460 -611
rect 5700 -611 5770 -589
rect 5700 -649 5710 -611
rect 5760 -649 5770 -611
rect 6010 -611 6090 -589
rect 6010 -649 6020 -611
rect 6080 -649 6090 -611
rect 6330 -611 6400 -589
rect 6330 -649 6340 -611
rect 6390 -649 6400 -611
rect 6640 -611 6720 -589
rect 6640 -649 6650 -611
rect 6710 -649 6720 -611
rect 6960 -611 7040 -589
rect 6960 -649 6970 -611
rect 7030 -649 7040 -611
rect 7280 -649 7290 -589
rect 7340 -560 7350 -500
rect 7590 -560 7670 -500
rect 7910 -560 7980 -500
rect 8220 -560 8300 -500
rect 8540 -560 8620 -500
rect 8860 -560 8930 -500
rect 9170 -560 9250 -500
rect 9490 -560 9560 -500
rect 9800 -560 10070 -500
rect 7340 -589 10070 -560
rect 7340 -649 7350 -589
rect 7590 -649 7670 -589
rect 7910 -649 7980 -589
rect 8220 -649 8300 -589
rect 8540 -649 8620 -589
rect 8860 -649 8930 -589
rect 9170 -649 9250 -589
rect 9490 -649 9560 -589
rect 9800 -649 10070 -589
rect 4560 -650 4810 -649
rect 7340 -650 10070 -649
rect 4560 -1510 4570 -650
rect 4755 -708 4815 -678
rect 4811 -1448 4815 -708
rect 4755 -1478 4815 -1448
rect 4913 -708 4973 -678
rect 4969 -1448 4973 -708
rect 4913 -1478 4973 -1448
rect 5071 -708 5131 -678
rect 5127 -1448 5131 -708
rect 5071 -1478 5131 -1448
rect 5229 -708 5289 -678
rect 5285 -1448 5289 -708
rect 5229 -1478 5289 -1448
rect 5387 -708 5447 -678
rect 5443 -1448 5447 -708
rect 5387 -1478 5447 -1448
rect 5545 -708 5605 -678
rect 5601 -1448 5605 -708
rect 5545 -1478 5605 -1448
rect 5703 -708 5763 -678
rect 5759 -1448 5763 -708
rect 5703 -1478 5763 -1448
rect 5861 -708 5921 -678
rect 5917 -1448 5921 -708
rect 5861 -1478 5921 -1448
rect 6019 -708 6079 -678
rect 6075 -1448 6079 -708
rect 6019 -1478 6079 -1448
rect 6177 -708 6237 -678
rect 6233 -1448 6237 -708
rect 6177 -1478 6237 -1448
rect 6335 -708 6395 -678
rect 6391 -1448 6395 -708
rect 6335 -1478 6395 -1448
rect 6493 -708 6553 -678
rect 6549 -1448 6553 -708
rect 6493 -1478 6553 -1448
rect 6651 -708 6711 -678
rect 6707 -1448 6711 -708
rect 6651 -1478 6711 -1448
rect 6809 -708 6869 -678
rect 6865 -1448 6869 -708
rect 6809 -1478 6869 -1448
rect 6967 -708 7027 -678
rect 7023 -1448 7027 -708
rect 6967 -1478 7027 -1448
rect 7125 -708 7185 -678
rect 7181 -1448 7185 -708
rect 7125 -1478 7185 -1448
rect 7283 -708 7343 -678
rect 7339 -1448 7343 -708
rect 7283 -1478 7343 -1448
rect 7441 -708 7501 -678
rect 7497 -1448 7501 -708
rect 7441 -1478 7501 -1448
rect 7599 -708 7659 -678
rect 7655 -1448 7659 -708
rect 7599 -1478 7659 -1448
rect 7757 -708 7817 -678
rect 7813 -1448 7817 -708
rect 7757 -1478 7817 -1448
rect 7915 -708 7975 -678
rect 7971 -1448 7975 -708
rect 7915 -1478 7975 -1448
rect 8073 -708 8133 -678
rect 8129 -1448 8133 -708
rect 8073 -1478 8133 -1448
rect 8231 -708 8291 -678
rect 8287 -1448 8291 -708
rect 8231 -1478 8291 -1448
rect 8389 -708 8449 -678
rect 8445 -1448 8449 -708
rect 8389 -1478 8449 -1448
rect 8547 -708 8607 -678
rect 8603 -1448 8607 -708
rect 8547 -1478 8607 -1448
rect 8705 -708 8765 -678
rect 8761 -1448 8765 -708
rect 8705 -1478 8765 -1448
rect 8863 -708 8923 -678
rect 8919 -1448 8923 -708
rect 8863 -1478 8923 -1448
rect 9021 -708 9081 -678
rect 9077 -1448 9081 -708
rect 9021 -1478 9081 -1448
rect 9179 -708 9239 -678
rect 9235 -1448 9239 -708
rect 9179 -1478 9239 -1448
rect 9337 -708 9397 -678
rect 9393 -1448 9397 -708
rect 9337 -1478 9397 -1448
rect 9495 -708 9555 -678
rect 9551 -1448 9555 -708
rect 9495 -1478 9555 -1448
rect 9653 -708 9713 -678
rect 9709 -1448 9713 -708
rect 9653 -1478 9713 -1448
rect 9811 -708 9871 -678
rect 9867 -1448 9871 -708
rect 9811 -1478 9871 -1448
rect 10060 -1510 10070 -650
rect 4560 -1570 4820 -1510
rect 5060 -1570 5140 -1510
rect 5380 -1570 5460 -1510
rect 5700 -1570 5770 -1510
rect 6010 -1570 6090 -1510
rect 6330 -1570 6400 -1510
rect 6640 -1570 6720 -1510
rect 6960 -1570 7040 -1510
rect 7280 -1570 7290 -1510
rect 4560 -1607 7290 -1570
rect 4560 -1660 4820 -1607
rect 4560 -2530 4570 -1660
rect 4810 -1667 4820 -1660
rect 5060 -1667 5140 -1607
rect 5380 -1667 5460 -1607
rect 5700 -1667 5770 -1607
rect 6010 -1667 6090 -1607
rect 6330 -1667 6400 -1607
rect 6640 -1667 6720 -1607
rect 6960 -1667 7040 -1607
rect 7280 -1667 7290 -1607
rect 7340 -1570 7350 -1510
rect 7590 -1570 7670 -1510
rect 7910 -1570 7980 -1510
rect 8220 -1570 8300 -1510
rect 8540 -1570 8620 -1510
rect 8860 -1570 8930 -1510
rect 9170 -1570 9250 -1510
rect 9490 -1570 9560 -1510
rect 9800 -1570 10070 -1510
rect 7340 -1607 10070 -1570
rect 7340 -1667 7350 -1607
rect 7590 -1667 7670 -1607
rect 7910 -1667 7980 -1607
rect 8220 -1667 8300 -1607
rect 8540 -1667 8620 -1607
rect 8860 -1667 8930 -1607
rect 9170 -1667 9250 -1607
rect 9490 -1667 9560 -1607
rect 9800 -1660 10070 -1607
rect 9800 -1667 9820 -1660
rect 7340 -1668 9820 -1667
rect 4755 -1726 4815 -1696
rect 4811 -2466 4815 -1726
rect 4755 -2496 4815 -2466
rect 4913 -1726 4973 -1696
rect 4969 -2466 4973 -1726
rect 4913 -2496 4973 -2466
rect 5071 -1726 5131 -1696
rect 5127 -2466 5131 -1726
rect 5071 -2496 5131 -2466
rect 5229 -1726 5289 -1696
rect 5285 -2466 5289 -1726
rect 5229 -2496 5289 -2466
rect 5387 -1726 5447 -1696
rect 5443 -2466 5447 -1726
rect 5387 -2496 5447 -2466
rect 5545 -1726 5605 -1696
rect 5601 -2466 5605 -1726
rect 5545 -2496 5605 -2466
rect 5703 -1726 5763 -1696
rect 5759 -2466 5763 -1726
rect 5703 -2496 5763 -2466
rect 5861 -1726 5921 -1696
rect 5917 -2466 5921 -1726
rect 5861 -2496 5921 -2466
rect 6019 -1726 6079 -1696
rect 6075 -2466 6079 -1726
rect 6019 -2496 6079 -2466
rect 6177 -1726 6237 -1696
rect 6233 -2466 6237 -1726
rect 6177 -2496 6237 -2466
rect 6335 -1726 6395 -1696
rect 6391 -2466 6395 -1726
rect 6335 -2496 6395 -2466
rect 6493 -1726 6553 -1696
rect 6549 -2466 6553 -1726
rect 6493 -2496 6553 -2466
rect 6651 -1726 6711 -1696
rect 6707 -2466 6711 -1726
rect 6651 -2496 6711 -2466
rect 6809 -1726 6869 -1696
rect 6865 -2466 6869 -1726
rect 6809 -2496 6869 -2466
rect 6967 -1726 7027 -1696
rect 7023 -2466 7027 -1726
rect 6967 -2496 7027 -2466
rect 7125 -1726 7185 -1696
rect 7181 -2466 7185 -1726
rect 7125 -2496 7185 -2466
rect 7283 -1726 7343 -1696
rect 7339 -2466 7343 -1726
rect 7283 -2496 7343 -2466
rect 7441 -1726 7501 -1696
rect 7497 -2466 7501 -1726
rect 7441 -2496 7501 -2466
rect 7599 -1726 7659 -1696
rect 7655 -2466 7659 -1726
rect 7599 -2496 7659 -2466
rect 7757 -1726 7817 -1696
rect 7813 -2466 7817 -1726
rect 7757 -2496 7817 -2466
rect 7915 -1726 7975 -1696
rect 7971 -2466 7975 -1726
rect 7915 -2496 7975 -2466
rect 8073 -1726 8133 -1696
rect 8129 -2466 8133 -1726
rect 8073 -2496 8133 -2466
rect 8231 -1726 8291 -1696
rect 8287 -2466 8291 -1726
rect 8231 -2496 8291 -2466
rect 8389 -1726 8449 -1696
rect 8445 -2466 8449 -1726
rect 8389 -2496 8449 -2466
rect 8547 -1726 8607 -1696
rect 8603 -2466 8607 -1726
rect 8547 -2496 8607 -2466
rect 8705 -1726 8765 -1696
rect 8761 -2466 8765 -1726
rect 8705 -2496 8765 -2466
rect 8863 -1726 8923 -1696
rect 8919 -2466 8923 -1726
rect 8863 -2496 8923 -2466
rect 9021 -1726 9081 -1696
rect 9077 -2466 9081 -1726
rect 9021 -2496 9081 -2466
rect 9179 -1726 9239 -1696
rect 9235 -2466 9239 -1726
rect 9179 -2496 9239 -2466
rect 9337 -1726 9397 -1696
rect 9393 -2466 9397 -1726
rect 9337 -2496 9397 -2466
rect 9495 -1726 9555 -1696
rect 9551 -2466 9555 -1726
rect 9495 -2496 9555 -2466
rect 9653 -1726 9713 -1696
rect 9709 -2466 9713 -1726
rect 9653 -2496 9713 -2466
rect 9811 -1726 9871 -1696
rect 9867 -2466 9871 -1726
rect 9811 -2496 9871 -2466
rect 10060 -2530 10070 -1660
rect 4560 -2590 4820 -2530
rect 5060 -2590 5140 -2530
rect 5380 -2590 5460 -2530
rect 5700 -2590 5770 -2530
rect 6010 -2590 6090 -2530
rect 6330 -2590 6400 -2530
rect 6640 -2590 6720 -2530
rect 6960 -2590 7040 -2530
rect 7280 -2590 7290 -2530
rect 4560 -2624 7290 -2590
rect 4560 -2680 4820 -2624
rect 4560 -3550 4570 -2680
rect 4810 -2684 4820 -2680
rect 5060 -2684 5140 -2624
rect 5380 -2684 5460 -2624
rect 5700 -2684 5770 -2624
rect 6010 -2684 6090 -2624
rect 6330 -2684 6400 -2624
rect 6640 -2684 6720 -2624
rect 6960 -2684 7040 -2624
rect 7280 -2684 7290 -2624
rect 7340 -2590 7350 -2530
rect 7590 -2590 7670 -2530
rect 7910 -2590 7980 -2530
rect 8220 -2590 8300 -2530
rect 8540 -2590 8620 -2530
rect 8860 -2590 8930 -2530
rect 9170 -2590 9250 -2530
rect 9490 -2590 9560 -2530
rect 9800 -2590 10070 -2530
rect 7340 -2624 10070 -2590
rect 7340 -2684 7350 -2624
rect 7590 -2684 7670 -2624
rect 7910 -2684 7980 -2624
rect 8220 -2684 8300 -2624
rect 8540 -2684 8620 -2624
rect 8860 -2684 8930 -2624
rect 9170 -2684 9250 -2624
rect 9490 -2684 9560 -2624
rect 9800 -2680 10070 -2624
rect 9800 -2684 9820 -2680
rect 4755 -2744 4815 -2714
rect 4811 -3484 4815 -2744
rect 4755 -3514 4815 -3484
rect 4913 -2744 4973 -2714
rect 4969 -3484 4973 -2744
rect 4913 -3514 4973 -3484
rect 5071 -2744 5131 -2714
rect 5127 -3484 5131 -2744
rect 5071 -3514 5131 -3484
rect 5229 -2744 5289 -2714
rect 5285 -3484 5289 -2744
rect 5229 -3514 5289 -3484
rect 5387 -2744 5447 -2714
rect 5443 -3484 5447 -2744
rect 5387 -3514 5447 -3484
rect 5545 -2744 5605 -2714
rect 5601 -3484 5605 -2744
rect 5545 -3514 5605 -3484
rect 5703 -2744 5763 -2714
rect 5759 -3484 5763 -2744
rect 5703 -3514 5763 -3484
rect 5861 -2744 5921 -2714
rect 5917 -3484 5921 -2744
rect 5861 -3514 5921 -3484
rect 6019 -2744 6079 -2714
rect 6075 -3484 6079 -2744
rect 6019 -3514 6079 -3484
rect 6177 -2744 6237 -2714
rect 6233 -3484 6237 -2744
rect 6177 -3514 6237 -3484
rect 6335 -2744 6395 -2714
rect 6391 -3484 6395 -2744
rect 6335 -3514 6395 -3484
rect 6493 -2744 6553 -2714
rect 6549 -3484 6553 -2744
rect 6493 -3514 6553 -3484
rect 6651 -2744 6711 -2714
rect 6707 -3484 6711 -2744
rect 6651 -3514 6711 -3484
rect 6809 -2744 6869 -2714
rect 6865 -3484 6869 -2744
rect 6809 -3514 6869 -3484
rect 6967 -2744 7027 -2714
rect 7023 -3484 7027 -2744
rect 6967 -3514 7027 -3484
rect 7125 -2744 7185 -2714
rect 7181 -3484 7185 -2744
rect 7125 -3514 7185 -3484
rect 7283 -2744 7343 -2714
rect 7339 -3484 7343 -2744
rect 7283 -3514 7343 -3484
rect 7441 -2744 7501 -2714
rect 7497 -3484 7501 -2744
rect 7441 -3514 7501 -3484
rect 7599 -2744 7659 -2714
rect 7655 -3484 7659 -2744
rect 7599 -3514 7659 -3484
rect 7757 -2744 7817 -2714
rect 7813 -3484 7817 -2744
rect 7757 -3514 7817 -3484
rect 7915 -2744 7975 -2714
rect 7971 -3484 7975 -2744
rect 7915 -3514 7975 -3484
rect 8073 -2744 8133 -2714
rect 8129 -3484 8133 -2744
rect 8073 -3514 8133 -3484
rect 8231 -2744 8291 -2714
rect 8287 -3484 8291 -2744
rect 8231 -3514 8291 -3484
rect 8389 -2744 8449 -2714
rect 8445 -3484 8449 -2744
rect 8389 -3514 8449 -3484
rect 8547 -2744 8607 -2714
rect 8603 -3484 8607 -2744
rect 8547 -3514 8607 -3484
rect 8705 -2744 8765 -2714
rect 8761 -3484 8765 -2744
rect 8705 -3514 8765 -3484
rect 8863 -2744 8923 -2714
rect 8919 -3484 8923 -2744
rect 8863 -3514 8923 -3484
rect 9021 -2744 9081 -2714
rect 9077 -3484 9081 -2744
rect 9021 -3514 9081 -3484
rect 9179 -2744 9239 -2714
rect 9235 -3484 9239 -2744
rect 9179 -3514 9239 -3484
rect 9337 -2744 9397 -2714
rect 9393 -3484 9397 -2744
rect 9337 -3514 9397 -3484
rect 9495 -2744 9555 -2714
rect 9551 -3484 9555 -2744
rect 9495 -3514 9555 -3484
rect 9653 -2744 9713 -2714
rect 9709 -3484 9713 -2744
rect 9653 -3514 9713 -3484
rect 9811 -2744 9871 -2714
rect 9867 -3484 9871 -2744
rect 9811 -3514 9871 -3484
rect 10060 -3550 10070 -2680
rect 4560 -3610 4820 -3550
rect 5060 -3610 5140 -3550
rect 5380 -3610 5460 -3550
rect 5700 -3610 5770 -3550
rect 6010 -3610 6090 -3550
rect 6330 -3610 6400 -3550
rect 6640 -3610 6720 -3550
rect 6960 -3610 7040 -3550
rect 7280 -3610 7290 -3550
rect 7340 -3610 7350 -3550
rect 7590 -3610 7670 -3550
rect 7910 -3610 7980 -3550
rect 8220 -3610 8300 -3550
rect 8540 -3610 8620 -3550
rect 8860 -3610 8930 -3550
rect 9170 -3610 9250 -3550
rect 9490 -3610 9560 -3550
rect 9800 -3610 10070 -3550
rect 10150 -3610 10160 430
rect 4470 -3630 4810 -3610
rect 9820 -3630 10160 -3610
rect 4200 -4140 4280 -4020
rect 10440 -4060 10520 -4020
rect 4360 -4140 4380 -4060
rect 10420 -4140 10520 -4060
<< via2 >>
rect 4660 580 9880 640
rect 4660 500 9880 580
rect 4480 -3610 4560 430
rect 4755 -430 4810 310
rect 4810 -430 4811 310
rect 4913 -430 4968 310
rect 4968 -430 4969 310
rect 5071 -430 5126 310
rect 5126 -430 5127 310
rect 5229 -430 5284 310
rect 5284 -430 5285 310
rect 5387 -430 5442 310
rect 5442 -430 5443 310
rect 5545 -430 5600 310
rect 5600 -430 5601 310
rect 5703 -430 5758 310
rect 5758 -430 5759 310
rect 5861 -430 5916 310
rect 5916 -430 5917 310
rect 6019 -430 6074 310
rect 6074 -430 6075 310
rect 6177 -430 6232 310
rect 6232 -430 6233 310
rect 6335 -430 6390 310
rect 6390 -430 6391 310
rect 6493 -430 6548 310
rect 6548 -430 6549 310
rect 6651 -430 6706 310
rect 6706 -430 6707 310
rect 6809 -430 6864 310
rect 6864 -430 6865 310
rect 6967 -430 7022 310
rect 7022 -430 7023 310
rect 7125 -430 7180 310
rect 7180 -430 7181 310
rect 7283 -430 7338 310
rect 7338 -430 7339 310
rect 7441 -430 7496 310
rect 7496 -430 7497 310
rect 7599 -430 7654 310
rect 7654 -430 7655 310
rect 7757 -430 7812 310
rect 7812 -430 7813 310
rect 7915 -430 7970 310
rect 7970 -430 7971 310
rect 8073 -430 8128 310
rect 8128 -430 8129 310
rect 8231 -430 8286 310
rect 8286 -430 8287 310
rect 8389 -430 8444 310
rect 8444 -430 8445 310
rect 8547 -430 8602 310
rect 8602 -430 8603 310
rect 8705 -430 8760 310
rect 8760 -430 8761 310
rect 8863 -430 8918 310
rect 8918 -430 8919 310
rect 9021 -430 9076 310
rect 9076 -430 9077 310
rect 9179 -430 9234 310
rect 9234 -430 9235 310
rect 9337 -430 9392 310
rect 9392 -430 9393 310
rect 9495 -430 9550 310
rect 9550 -430 9551 310
rect 9653 -430 9708 310
rect 9708 -430 9709 310
rect 9811 -430 9866 310
rect 9866 -430 9867 310
rect 4755 -1448 4810 -708
rect 4810 -1448 4811 -708
rect 4913 -1448 4968 -708
rect 4968 -1448 4969 -708
rect 5071 -1448 5126 -708
rect 5126 -1448 5127 -708
rect 5229 -1448 5284 -708
rect 5284 -1448 5285 -708
rect 5387 -1448 5442 -708
rect 5442 -1448 5443 -708
rect 5545 -1448 5600 -708
rect 5600 -1448 5601 -708
rect 5703 -1448 5758 -708
rect 5758 -1448 5759 -708
rect 5861 -1448 5916 -708
rect 5916 -1448 5917 -708
rect 6019 -1448 6074 -708
rect 6074 -1448 6075 -708
rect 6177 -1448 6232 -708
rect 6232 -1448 6233 -708
rect 6335 -1448 6390 -708
rect 6390 -1448 6391 -708
rect 6493 -1448 6548 -708
rect 6548 -1448 6549 -708
rect 6651 -1448 6706 -708
rect 6706 -1448 6707 -708
rect 6809 -1448 6864 -708
rect 6864 -1448 6865 -708
rect 6967 -1448 7022 -708
rect 7022 -1448 7023 -708
rect 7125 -1448 7180 -708
rect 7180 -1448 7181 -708
rect 7283 -1448 7338 -708
rect 7338 -1448 7339 -708
rect 7441 -1448 7496 -708
rect 7496 -1448 7497 -708
rect 7599 -1448 7654 -708
rect 7654 -1448 7655 -708
rect 7757 -1448 7812 -708
rect 7812 -1448 7813 -708
rect 7915 -1448 7970 -708
rect 7970 -1448 7971 -708
rect 8073 -1448 8128 -708
rect 8128 -1448 8129 -708
rect 8231 -1448 8286 -708
rect 8286 -1448 8287 -708
rect 8389 -1448 8444 -708
rect 8444 -1448 8445 -708
rect 8547 -1448 8602 -708
rect 8602 -1448 8603 -708
rect 8705 -1448 8760 -708
rect 8760 -1448 8761 -708
rect 8863 -1448 8918 -708
rect 8918 -1448 8919 -708
rect 9021 -1448 9076 -708
rect 9076 -1448 9077 -708
rect 9179 -1448 9234 -708
rect 9234 -1448 9235 -708
rect 9337 -1448 9392 -708
rect 9392 -1448 9393 -708
rect 9495 -1448 9550 -708
rect 9550 -1448 9551 -708
rect 9653 -1448 9708 -708
rect 9708 -1448 9709 -708
rect 9811 -1448 9866 -708
rect 9866 -1448 9867 -708
rect 4755 -2466 4810 -1726
rect 4810 -2466 4811 -1726
rect 4913 -2466 4968 -1726
rect 4968 -2466 4969 -1726
rect 5071 -2466 5126 -1726
rect 5126 -2466 5127 -1726
rect 5229 -2466 5284 -1726
rect 5284 -2466 5285 -1726
rect 5387 -2466 5442 -1726
rect 5442 -2466 5443 -1726
rect 5545 -2466 5600 -1726
rect 5600 -2466 5601 -1726
rect 5703 -2466 5758 -1726
rect 5758 -2466 5759 -1726
rect 5861 -2466 5916 -1726
rect 5916 -2466 5917 -1726
rect 6019 -2466 6074 -1726
rect 6074 -2466 6075 -1726
rect 6177 -2466 6232 -1726
rect 6232 -2466 6233 -1726
rect 6335 -2466 6390 -1726
rect 6390 -2466 6391 -1726
rect 6493 -2466 6548 -1726
rect 6548 -2466 6549 -1726
rect 6651 -2466 6706 -1726
rect 6706 -2466 6707 -1726
rect 6809 -2466 6864 -1726
rect 6864 -2466 6865 -1726
rect 6967 -2466 7022 -1726
rect 7022 -2466 7023 -1726
rect 7125 -2466 7180 -1726
rect 7180 -2466 7181 -1726
rect 7283 -2466 7338 -1726
rect 7338 -2466 7339 -1726
rect 7441 -2466 7496 -1726
rect 7496 -2466 7497 -1726
rect 7599 -2466 7654 -1726
rect 7654 -2466 7655 -1726
rect 7757 -2466 7812 -1726
rect 7812 -2466 7813 -1726
rect 7915 -2466 7970 -1726
rect 7970 -2466 7971 -1726
rect 8073 -2466 8128 -1726
rect 8128 -2466 8129 -1726
rect 8231 -2466 8286 -1726
rect 8286 -2466 8287 -1726
rect 8389 -2466 8444 -1726
rect 8444 -2466 8445 -1726
rect 8547 -2466 8602 -1726
rect 8602 -2466 8603 -1726
rect 8705 -2466 8760 -1726
rect 8760 -2466 8761 -1726
rect 8863 -2466 8918 -1726
rect 8918 -2466 8919 -1726
rect 9021 -2466 9076 -1726
rect 9076 -2466 9077 -1726
rect 9179 -2466 9234 -1726
rect 9234 -2466 9235 -1726
rect 9337 -2466 9392 -1726
rect 9392 -2466 9393 -1726
rect 9495 -2466 9550 -1726
rect 9550 -2466 9551 -1726
rect 9653 -2466 9708 -1726
rect 9708 -2466 9709 -1726
rect 9811 -2466 9866 -1726
rect 9866 -2466 9867 -1726
rect 4755 -3484 4810 -2744
rect 4810 -3484 4811 -2744
rect 4913 -3484 4968 -2744
rect 4968 -3484 4969 -2744
rect 5071 -3484 5126 -2744
rect 5126 -3484 5127 -2744
rect 5229 -3484 5284 -2744
rect 5284 -3484 5285 -2744
rect 5387 -3484 5442 -2744
rect 5442 -3484 5443 -2744
rect 5545 -3484 5600 -2744
rect 5600 -3484 5601 -2744
rect 5703 -3484 5758 -2744
rect 5758 -3484 5759 -2744
rect 5861 -3484 5916 -2744
rect 5916 -3484 5917 -2744
rect 6019 -3484 6074 -2744
rect 6074 -3484 6075 -2744
rect 6177 -3484 6232 -2744
rect 6232 -3484 6233 -2744
rect 6335 -3484 6390 -2744
rect 6390 -3484 6391 -2744
rect 6493 -3484 6548 -2744
rect 6548 -3484 6549 -2744
rect 6651 -3484 6706 -2744
rect 6706 -3484 6707 -2744
rect 6809 -3484 6864 -2744
rect 6864 -3484 6865 -2744
rect 6967 -3484 7022 -2744
rect 7022 -3484 7023 -2744
rect 7125 -3484 7180 -2744
rect 7180 -3484 7181 -2744
rect 7283 -3484 7338 -2744
rect 7338 -3484 7339 -2744
rect 7441 -3484 7496 -2744
rect 7496 -3484 7497 -2744
rect 7599 -3484 7654 -2744
rect 7654 -3484 7655 -2744
rect 7757 -3484 7812 -2744
rect 7812 -3484 7813 -2744
rect 7915 -3484 7970 -2744
rect 7970 -3484 7971 -2744
rect 8073 -3484 8128 -2744
rect 8128 -3484 8129 -2744
rect 8231 -3484 8286 -2744
rect 8286 -3484 8287 -2744
rect 8389 -3484 8444 -2744
rect 8444 -3484 8445 -2744
rect 8547 -3484 8602 -2744
rect 8602 -3484 8603 -2744
rect 8705 -3484 8760 -2744
rect 8760 -3484 8761 -2744
rect 8863 -3484 8918 -2744
rect 8918 -3484 8919 -2744
rect 9021 -3484 9076 -2744
rect 9076 -3484 9077 -2744
rect 9179 -3484 9234 -2744
rect 9234 -3484 9235 -2744
rect 9337 -3484 9392 -2744
rect 9392 -3484 9393 -2744
rect 9495 -3484 9550 -2744
rect 9550 -3484 9551 -2744
rect 9653 -3484 9708 -2744
rect 9708 -3484 9709 -2744
rect 9811 -3484 9866 -2744
rect 9866 -3484 9867 -2744
rect 10070 -3610 10150 430
<< metal3 >>
rect 4640 640 9920 660
rect 4640 500 4660 640
rect 9880 500 9920 640
rect 4640 480 9920 500
rect 4470 430 4570 450
rect 4470 -3610 4480 430
rect 4560 -3610 4570 430
rect 4750 310 4820 480
rect 4750 -430 4755 310
rect 4811 -430 4820 310
rect 4750 -708 4820 -430
rect 4750 -1448 4755 -708
rect 4811 -1448 4820 -708
rect 4750 -1726 4820 -1448
rect 4750 -2466 4755 -1726
rect 4811 -2466 4820 -1726
rect 4750 -2744 4820 -2466
rect 4750 -3484 4755 -2744
rect 4811 -3484 4820 -2744
rect 4750 -3520 4820 -3484
rect 4908 310 4978 340
rect 4908 -430 4913 310
rect 4969 -430 4978 310
rect 4908 -708 4978 -430
rect 4908 -1448 4913 -708
rect 4969 -1448 4978 -708
rect 4908 -1726 4978 -1448
rect 4908 -2466 4913 -1726
rect 4969 -2466 4978 -1726
rect 4908 -2744 4978 -2466
rect 4908 -3484 4913 -2744
rect 4969 -3484 4978 -2744
rect 4470 -3630 4570 -3610
rect 4908 -3680 4978 -3484
rect 5066 310 5136 480
rect 5066 -430 5071 310
rect 5127 -430 5136 310
rect 5066 -708 5136 -430
rect 5066 -1448 5071 -708
rect 5127 -1448 5136 -708
rect 5066 -1726 5136 -1448
rect 5066 -2466 5071 -1726
rect 5127 -2466 5136 -1726
rect 5066 -2744 5136 -2466
rect 5066 -3484 5071 -2744
rect 5127 -3484 5136 -2744
rect 5066 -3520 5136 -3484
rect 5224 310 5294 340
rect 5224 -430 5229 310
rect 5285 -430 5294 310
rect 5224 -708 5294 -430
rect 5224 -1448 5229 -708
rect 5285 -1448 5294 -708
rect 5224 -1726 5294 -1448
rect 5224 -2466 5229 -1726
rect 5285 -2466 5294 -1726
rect 5224 -2744 5294 -2466
rect 5224 -3484 5229 -2744
rect 5285 -3484 5294 -2744
rect 5224 -3680 5294 -3484
rect 5382 310 5452 480
rect 5382 -430 5387 310
rect 5443 -430 5452 310
rect 5382 -708 5452 -430
rect 5382 -1448 5387 -708
rect 5443 -1448 5452 -708
rect 5382 -1726 5452 -1448
rect 5382 -2466 5387 -1726
rect 5443 -2466 5452 -1726
rect 5382 -2744 5452 -2466
rect 5382 -3484 5387 -2744
rect 5443 -3484 5452 -2744
rect 5382 -3520 5452 -3484
rect 5540 310 5610 340
rect 5540 -430 5545 310
rect 5601 -430 5610 310
rect 5540 -708 5610 -430
rect 5540 -1448 5545 -708
rect 5601 -1448 5610 -708
rect 5540 -1726 5610 -1448
rect 5540 -2466 5545 -1726
rect 5601 -2466 5610 -1726
rect 5540 -2744 5610 -2466
rect 5540 -3484 5545 -2744
rect 5601 -3484 5610 -2744
rect 5540 -3680 5610 -3484
rect 5698 310 5768 480
rect 5698 -430 5703 310
rect 5759 -430 5768 310
rect 5698 -708 5768 -430
rect 5698 -1448 5703 -708
rect 5759 -1448 5768 -708
rect 5698 -1726 5768 -1448
rect 5698 -2466 5703 -1726
rect 5759 -2466 5768 -1726
rect 5698 -2744 5768 -2466
rect 5698 -3484 5703 -2744
rect 5759 -3484 5768 -2744
rect 5698 -3520 5768 -3484
rect 5856 310 5926 340
rect 5856 -430 5861 310
rect 5917 -430 5926 310
rect 5856 -708 5926 -430
rect 5856 -1448 5861 -708
rect 5917 -1448 5926 -708
rect 5856 -1726 5926 -1448
rect 5856 -2466 5861 -1726
rect 5917 -2466 5926 -1726
rect 5856 -2744 5926 -2466
rect 5856 -3484 5861 -2744
rect 5917 -3484 5926 -2744
rect 5856 -3680 5926 -3484
rect 6014 310 6084 480
rect 6014 -430 6019 310
rect 6075 -430 6084 310
rect 6014 -708 6084 -430
rect 6014 -1448 6019 -708
rect 6075 -1448 6084 -708
rect 6014 -1726 6084 -1448
rect 6014 -2466 6019 -1726
rect 6075 -2466 6084 -1726
rect 6014 -2744 6084 -2466
rect 6014 -3484 6019 -2744
rect 6075 -3484 6084 -2744
rect 6014 -3520 6084 -3484
rect 6172 310 6242 340
rect 6172 -430 6177 310
rect 6233 -430 6242 310
rect 6172 -708 6242 -430
rect 6172 -1448 6177 -708
rect 6233 -1448 6242 -708
rect 6172 -1726 6242 -1448
rect 6172 -2466 6177 -1726
rect 6233 -2466 6242 -1726
rect 6172 -2744 6242 -2466
rect 6172 -3484 6177 -2744
rect 6233 -3484 6242 -2744
rect 6172 -3680 6242 -3484
rect 6330 310 6400 480
rect 6330 -430 6335 310
rect 6391 -430 6400 310
rect 6330 -708 6400 -430
rect 6330 -1448 6335 -708
rect 6391 -1448 6400 -708
rect 6330 -1726 6400 -1448
rect 6330 -2466 6335 -1726
rect 6391 -2466 6400 -1726
rect 6330 -2744 6400 -2466
rect 6330 -3484 6335 -2744
rect 6391 -3484 6400 -2744
rect 6330 -3520 6400 -3484
rect 6488 310 6558 340
rect 6488 -430 6493 310
rect 6549 -430 6558 310
rect 6488 -708 6558 -430
rect 6488 -1448 6493 -708
rect 6549 -1448 6558 -708
rect 6488 -1726 6558 -1448
rect 6488 -2466 6493 -1726
rect 6549 -2466 6558 -1726
rect 6488 -2744 6558 -2466
rect 6488 -3484 6493 -2744
rect 6549 -3484 6558 -2744
rect 6488 -3680 6558 -3484
rect 6646 310 6716 480
rect 6646 -430 6651 310
rect 6707 -430 6716 310
rect 6646 -708 6716 -430
rect 6646 -1448 6651 -708
rect 6707 -1448 6716 -708
rect 6646 -1726 6716 -1448
rect 6646 -2466 6651 -1726
rect 6707 -2466 6716 -1726
rect 6646 -2744 6716 -2466
rect 6646 -3484 6651 -2744
rect 6707 -3484 6716 -2744
rect 6646 -3520 6716 -3484
rect 6804 310 6874 340
rect 6804 -430 6809 310
rect 6865 -430 6874 310
rect 6804 -708 6874 -430
rect 6804 -1448 6809 -708
rect 6865 -1448 6874 -708
rect 6804 -1726 6874 -1448
rect 6804 -2466 6809 -1726
rect 6865 -2466 6874 -1726
rect 6804 -2744 6874 -2466
rect 6804 -3484 6809 -2744
rect 6865 -3484 6874 -2744
rect 6804 -3680 6874 -3484
rect 6962 310 7032 480
rect 6962 -430 6967 310
rect 7023 -430 7032 310
rect 6962 -708 7032 -430
rect 6962 -1448 6967 -708
rect 7023 -1448 7032 -708
rect 6962 -1726 7032 -1448
rect 6962 -2466 6967 -1726
rect 7023 -2466 7032 -1726
rect 6962 -2744 7032 -2466
rect 6962 -3484 6967 -2744
rect 7023 -3484 7032 -2744
rect 6962 -3520 7032 -3484
rect 7120 310 7190 340
rect 7120 -430 7125 310
rect 7181 -430 7190 310
rect 7120 -708 7190 -430
rect 7120 -1448 7125 -708
rect 7181 -1448 7190 -708
rect 7120 -1726 7190 -1448
rect 7120 -2466 7125 -1726
rect 7181 -2466 7190 -1726
rect 7120 -2744 7190 -2466
rect 7120 -3484 7125 -2744
rect 7181 -3484 7190 -2744
rect 7120 -3680 7190 -3484
rect 7278 310 7348 480
rect 7278 -430 7283 310
rect 7339 -430 7348 310
rect 7278 -708 7348 -430
rect 7278 -1448 7283 -708
rect 7339 -1448 7348 -708
rect 7278 -1726 7348 -1448
rect 7278 -2466 7283 -1726
rect 7339 -2466 7348 -1726
rect 7278 -2744 7348 -2466
rect 7278 -3484 7283 -2744
rect 7339 -3484 7348 -2744
rect 7278 -3520 7348 -3484
rect 7436 310 7506 340
rect 7436 -430 7441 310
rect 7497 -430 7506 310
rect 7436 -708 7506 -430
rect 7436 -1448 7441 -708
rect 7497 -1448 7506 -708
rect 7436 -1726 7506 -1448
rect 7436 -2466 7441 -1726
rect 7497 -2466 7506 -1726
rect 7436 -2744 7506 -2466
rect 7436 -3484 7441 -2744
rect 7497 -3484 7506 -2744
rect 7436 -3680 7506 -3484
rect 7594 310 7664 480
rect 7594 -430 7599 310
rect 7655 -430 7664 310
rect 7594 -708 7664 -430
rect 7594 -1448 7599 -708
rect 7655 -1448 7664 -708
rect 7594 -1726 7664 -1448
rect 7594 -2466 7599 -1726
rect 7655 -2466 7664 -1726
rect 7594 -2744 7664 -2466
rect 7594 -3484 7599 -2744
rect 7655 -3484 7664 -2744
rect 7594 -3520 7664 -3484
rect 7752 310 7822 340
rect 7752 -430 7757 310
rect 7813 -430 7822 310
rect 7752 -708 7822 -430
rect 7752 -1448 7757 -708
rect 7813 -1448 7822 -708
rect 7752 -1726 7822 -1448
rect 7752 -2466 7757 -1726
rect 7813 -2466 7822 -1726
rect 7752 -2744 7822 -2466
rect 7752 -3484 7757 -2744
rect 7813 -3484 7822 -2744
rect 7752 -3680 7822 -3484
rect 7910 310 7980 480
rect 7910 -430 7915 310
rect 7971 -430 7980 310
rect 7910 -708 7980 -430
rect 7910 -1448 7915 -708
rect 7971 -1448 7980 -708
rect 7910 -1726 7980 -1448
rect 7910 -2466 7915 -1726
rect 7971 -2466 7980 -1726
rect 7910 -2744 7980 -2466
rect 7910 -3484 7915 -2744
rect 7971 -3484 7980 -2744
rect 7910 -3520 7980 -3484
rect 8068 310 8138 340
rect 8068 -430 8073 310
rect 8129 -430 8138 310
rect 8068 -708 8138 -430
rect 8068 -1448 8073 -708
rect 8129 -1448 8138 -708
rect 8068 -1726 8138 -1448
rect 8068 -2466 8073 -1726
rect 8129 -2466 8138 -1726
rect 8068 -2744 8138 -2466
rect 8068 -3484 8073 -2744
rect 8129 -3484 8138 -2744
rect 8068 -3680 8138 -3484
rect 8226 310 8296 480
rect 8226 -430 8231 310
rect 8287 -430 8296 310
rect 8226 -708 8296 -430
rect 8226 -1448 8231 -708
rect 8287 -1448 8296 -708
rect 8226 -1726 8296 -1448
rect 8226 -2466 8231 -1726
rect 8287 -2466 8296 -1726
rect 8226 -2744 8296 -2466
rect 8226 -3484 8231 -2744
rect 8287 -3484 8296 -2744
rect 8226 -3520 8296 -3484
rect 8384 310 8454 340
rect 8384 -430 8389 310
rect 8445 -430 8454 310
rect 8384 -708 8454 -430
rect 8384 -1448 8389 -708
rect 8445 -1448 8454 -708
rect 8384 -1726 8454 -1448
rect 8384 -2466 8389 -1726
rect 8445 -2466 8454 -1726
rect 8384 -2744 8454 -2466
rect 8384 -3484 8389 -2744
rect 8445 -3484 8454 -2744
rect 8384 -3680 8454 -3484
rect 8542 310 8612 480
rect 8542 -430 8547 310
rect 8603 -430 8612 310
rect 8542 -708 8612 -430
rect 8542 -1448 8547 -708
rect 8603 -1448 8612 -708
rect 8542 -1726 8612 -1448
rect 8542 -2466 8547 -1726
rect 8603 -2466 8612 -1726
rect 8542 -2744 8612 -2466
rect 8542 -3484 8547 -2744
rect 8603 -3484 8612 -2744
rect 8542 -3520 8612 -3484
rect 8700 310 8770 340
rect 8700 -430 8705 310
rect 8761 -430 8770 310
rect 8700 -708 8770 -430
rect 8700 -1448 8705 -708
rect 8761 -1448 8770 -708
rect 8700 -1726 8770 -1448
rect 8700 -2466 8705 -1726
rect 8761 -2466 8770 -1726
rect 8700 -2744 8770 -2466
rect 8700 -3484 8705 -2744
rect 8761 -3484 8770 -2744
rect 8700 -3680 8770 -3484
rect 8858 310 8928 480
rect 8858 -430 8863 310
rect 8919 -430 8928 310
rect 8858 -708 8928 -430
rect 8858 -1448 8863 -708
rect 8919 -1448 8928 -708
rect 8858 -1726 8928 -1448
rect 8858 -2466 8863 -1726
rect 8919 -2466 8928 -1726
rect 8858 -2744 8928 -2466
rect 8858 -3484 8863 -2744
rect 8919 -3484 8928 -2744
rect 8858 -3520 8928 -3484
rect 9016 310 9086 340
rect 9016 -430 9021 310
rect 9077 -430 9086 310
rect 9016 -708 9086 -430
rect 9016 -1448 9021 -708
rect 9077 -1448 9086 -708
rect 9016 -1726 9086 -1448
rect 9016 -2466 9021 -1726
rect 9077 -2466 9086 -1726
rect 9016 -2744 9086 -2466
rect 9016 -3484 9021 -2744
rect 9077 -3484 9086 -2744
rect 9016 -3680 9086 -3484
rect 9174 310 9244 480
rect 9174 -430 9179 310
rect 9235 -430 9244 310
rect 9174 -708 9244 -430
rect 9174 -1448 9179 -708
rect 9235 -1448 9244 -708
rect 9174 -1726 9244 -1448
rect 9174 -2466 9179 -1726
rect 9235 -2466 9244 -1726
rect 9174 -2744 9244 -2466
rect 9174 -3484 9179 -2744
rect 9235 -3484 9244 -2744
rect 9174 -3520 9244 -3484
rect 9332 310 9402 340
rect 9332 -430 9337 310
rect 9393 -430 9402 310
rect 9332 -708 9402 -430
rect 9332 -1448 9337 -708
rect 9393 -1448 9402 -708
rect 9332 -1726 9402 -1448
rect 9332 -2466 9337 -1726
rect 9393 -2466 9402 -1726
rect 9332 -2744 9402 -2466
rect 9332 -3484 9337 -2744
rect 9393 -3484 9402 -2744
rect 9332 -3680 9402 -3484
rect 9490 310 9560 480
rect 9490 -430 9495 310
rect 9551 -430 9560 310
rect 9490 -708 9560 -430
rect 9490 -1448 9495 -708
rect 9551 -1448 9560 -708
rect 9490 -1726 9560 -1448
rect 9490 -2466 9495 -1726
rect 9551 -2466 9560 -1726
rect 9490 -2744 9560 -2466
rect 9490 -3484 9495 -2744
rect 9551 -3484 9560 -2744
rect 9490 -3520 9560 -3484
rect 9648 310 9718 340
rect 9648 -430 9653 310
rect 9709 -430 9718 310
rect 9648 -708 9718 -430
rect 9648 -1448 9653 -708
rect 9709 -1448 9718 -708
rect 9648 -1726 9718 -1448
rect 9648 -2466 9653 -1726
rect 9709 -2466 9718 -1726
rect 9648 -2744 9718 -2466
rect 9648 -3484 9653 -2744
rect 9709 -3484 9718 -2744
rect 9648 -3680 9718 -3484
rect 9806 310 9876 480
rect 9806 -430 9811 310
rect 9867 -430 9876 310
rect 9806 -708 9876 -430
rect 9806 -1448 9811 -708
rect 9867 -1448 9876 -708
rect 9806 -1726 9876 -1448
rect 9806 -2466 9811 -1726
rect 9867 -2466 9876 -1726
rect 9806 -2744 9876 -2466
rect 9806 -3484 9811 -2744
rect 9867 -3484 9876 -2744
rect 9806 -3520 9876 -3484
rect 10060 430 10160 450
rect 10060 -3610 10070 430
rect 10150 -3610 10160 430
rect 10060 -3630 10160 -3610
rect 4908 -3780 9718 -3680
use sky130_fd_pr__nfet_03v3_nvt_EV757D  sky130_fd_pr__nfet_03v3_nvt_EV757D_0
timestamp 1660188747
transform 1 0 7312 0 1 -1590
box -2727 -2185 2727 2185
<< labels >>
rlabel metal3 4640 480 9920 660 1 SB
rlabel metal3 10060 -3630 10160 450 1 G1
rlabel metal3 4470 -3630 4570 450 1 G2
rlabel metal3 4900 -3780 9720 -3680 1 D
rlabel metal2 4160 860 10540 940 1 DNW
<< end >>
