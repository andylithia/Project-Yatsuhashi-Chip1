* SPICE3 file created from /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON/mimcap_1.ext - technology: sky130A

X0 top bot sky130_fd_pr__cap_mim_m3_1 l=1e+06u w=1e+07u
