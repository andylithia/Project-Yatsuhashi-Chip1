magic
tech sky130B
magscale 1 2
timestamp 1662258694
<< metal4 >>
rect -21700 -32300 -18700 -32100
rect -21700 -34500 -21500 -32300
rect -18900 -34500 -18700 -32300
rect -21700 -34700 -18700 -34500
rect -21700 -43900 -18900 -34700
<< via4 >>
rect -21500 -34500 -18900 -32300
<< metal5 >>
tri -29099 500 -27099 2500 se
rect -27099 500 -15501 2500
tri -15501 500 -13501 2500 sw
tri -30928 -1329 -29099 500 se
rect -29099 -100 -26871 500
tri -26871 -100 -26271 500 nw
tri -16329 -100 -15729 500 ne
rect -15729 -100 -13501 500
rect -29099 -949 -27720 -100
tri -27720 -949 -26871 -100 nw
tri -26871 -949 -26022 -100 se
rect -26022 -949 -16578 -100
tri -16578 -949 -15729 -100 sw
tri -15729 -949 -14880 -100 ne
rect -14880 -949 -13501 -100
rect -29099 -1329 -28100 -949
tri -28100 -1329 -27720 -949 nw
tri -27251 -1329 -26871 -949 se
rect -26871 -1251 -15729 -949
tri -15729 -1251 -15427 -949 sw
tri -14880 -1251 -14578 -949 ne
rect -14578 -1251 -13501 -949
rect -26871 -1329 -15427 -1251
tri -33528 -3929 -30928 -1329 se
rect -30928 -2178 -28949 -1329
tri -28949 -2178 -28100 -1329 nw
tri -28100 -2178 -27251 -1329 se
rect -27251 -2100 -15427 -1329
tri -15427 -2100 -14578 -1251 sw
tri -14578 -2100 -13729 -1251 ne
rect -13729 -2100 -13501 -1251
tri -13501 -2100 -10901 500 sw
rect -27251 -2178 -25794 -2100
rect -30928 -2406 -29177 -2178
tri -29177 -2406 -28949 -2178 nw
tri -28328 -2406 -28100 -2178 se
rect -28100 -2406 -25794 -2178
rect -30928 -3255 -30026 -2406
tri -30026 -3255 -29177 -2406 nw
tri -29177 -3255 -28328 -2406 se
rect -28328 -2700 -25794 -2406
tri -25794 -2700 -25194 -2100 nw
tri -17406 -2700 -16806 -2100 ne
rect -16806 -2700 -14578 -2100
rect -28328 -3255 -26349 -2700
tri -26349 -3255 -25794 -2700 nw
tri -25500 -3255 -24945 -2700 se
rect -24945 -3255 -17655 -2700
rect -30928 -3929 -30700 -3255
tri -30700 -3929 -30026 -3255 nw
tri -29851 -3929 -29177 -3255 se
rect -29177 -3929 -27198 -3255
tri -35300 -5701 -33528 -3929 se
rect -33528 -4778 -31549 -3929
tri -31549 -4778 -30700 -3929 nw
tri -30700 -4778 -29851 -3929 se
rect -29851 -4104 -27198 -3929
tri -27198 -4104 -26349 -3255 nw
tri -26349 -4104 -25500 -3255 se
rect -25500 -3549 -17655 -3255
tri -17655 -3549 -16806 -2700 sw
tri -16806 -3549 -15957 -2700 ne
rect -15957 -2949 -14578 -2700
tri -14578 -2949 -13729 -2100 sw
tri -13729 -2949 -12880 -2100 ne
rect -12880 -2949 -10901 -2100
rect -15957 -3002 -13729 -2949
tri -13729 -3002 -13676 -2949 sw
tri -12880 -3002 -12827 -2949 ne
rect -12827 -3002 -10901 -2949
rect -15957 -3549 -13676 -3002
rect -25500 -3851 -16806 -3549
tri -16806 -3851 -16504 -3549 sw
tri -15957 -3851 -15655 -3549 ne
rect -15655 -3851 -13676 -3549
tri -13676 -3851 -12827 -3002 sw
tri -12827 -3851 -11978 -3002 ne
rect -11978 -3851 -10901 -3002
rect -25500 -4104 -16504 -3851
rect -29851 -4700 -27794 -4104
tri -27794 -4700 -27198 -4104 nw
tri -26945 -4700 -26349 -4104 se
rect -26349 -4700 -16504 -4104
tri -16504 -4700 -15655 -3851 sw
tri -15655 -4700 -14806 -3851 ne
rect -14806 -4700 -12827 -3851
tri -12827 -4700 -11978 -3851 sw
tri -11978 -4700 -11129 -3851 ne
rect -11129 -4700 -10901 -3851
tri -10901 -4700 -8301 -2100 sw
rect -29851 -4778 -28100 -4700
rect -33528 -5006 -31777 -4778
tri -31777 -5006 -31549 -4778 nw
tri -30928 -5006 -30700 -4778 se
rect -30700 -5006 -28100 -4778
tri -28100 -5006 -27794 -4700 nw
tri -27251 -5006 -26945 -4700 se
rect -26945 -5006 -24717 -4700
rect -33528 -5701 -32626 -5006
rect -35300 -5855 -32626 -5701
tri -32626 -5855 -31777 -5006 nw
tri -31777 -5855 -30928 -5006 se
rect -30928 -5855 -28949 -5006
tri -28949 -5855 -28100 -5006 nw
tri -28100 -5855 -27251 -5006 se
rect -27251 -5300 -24717 -5006
tri -24717 -5300 -24117 -4700 nw
tri -18483 -5300 -17883 -4700 ne
rect -17883 -5300 -15655 -4700
rect -27251 -5855 -25500 -5300
rect -35300 -19000 -33300 -5855
tri -33300 -6529 -32626 -5855 nw
tri -31851 -5929 -31777 -5855 se
rect -31777 -5929 -29177 -5855
tri -32451 -6529 -31851 -5929 se
rect -31851 -6083 -29177 -5929
tri -29177 -6083 -28949 -5855 nw
tri -28328 -6083 -28100 -5855 se
rect -28100 -6083 -25500 -5855
tri -25500 -6083 -24717 -5300 nw
tri -24651 -6083 -23868 -5300 se
rect -23868 -6083 -18732 -5300
rect -31851 -6529 -30026 -6083
rect -37300 -21000 -33300 -19000
tri -32700 -6778 -32451 -6529 se
rect -32451 -6778 -30026 -6529
rect -32700 -6932 -30026 -6778
tri -30026 -6932 -29177 -6083 nw
tri -29177 -6932 -28328 -6083 se
rect -28328 -6932 -26349 -6083
tri -26349 -6932 -25500 -6083 nw
tri -25500 -6932 -24651 -6083 se
rect -24651 -6149 -18732 -6083
tri -18732 -6149 -17883 -5300 sw
tri -17883 -6149 -17034 -5300 ne
rect -17034 -5549 -15655 -5300
tri -15655 -5549 -14806 -4700 sw
tri -14806 -5549 -13957 -4700 ne
rect -13957 -5549 -11978 -4700
tri -11978 -5549 -11129 -4700 sw
tri -11129 -5549 -10280 -4700 ne
rect -10280 -5549 -8301 -4700
rect -17034 -5602 -14806 -5549
tri -14806 -5602 -14753 -5549 sw
tri -13957 -5602 -13904 -5549 ne
rect -13904 -5602 -11129 -5549
rect -17034 -6149 -14753 -5602
rect -24651 -6932 -17883 -6149
tri -17883 -6932 -17100 -6149 sw
tri -17034 -6932 -16251 -6149 ne
rect -16251 -6451 -14753 -6149
tri -14753 -6451 -13904 -5602 sw
tri -13904 -6451 -13055 -5602 ne
rect -13055 -5929 -11129 -5602
tri -11129 -5929 -10749 -5549 sw
tri -10280 -5929 -9900 -5549 ne
rect -9900 -5701 -8301 -5549
tri -8301 -5701 -7300 -4700 sw
rect -9900 -5929 -7300 -5701
rect -13055 -6451 -10749 -5929
rect -16251 -6932 -13904 -6451
rect -32700 -34832 -30700 -6932
tri -30700 -7606 -30026 -6932 nw
tri -29251 -7006 -29177 -6932 se
rect -29177 -7006 -26717 -6932
tri -29851 -7606 -29251 -7006 se
rect -29251 -7300 -26717 -7006
tri -26717 -7300 -26349 -6932 nw
tri -25868 -7300 -25500 -6932 se
rect -25500 -7300 -17100 -6932
tri -17100 -7300 -16732 -6932 sw
tri -16251 -7300 -15883 -6932 ne
rect -15883 -7300 -13904 -6932
tri -13904 -7300 -13055 -6451 sw
tri -13055 -7300 -12206 -6451 ne
rect -12206 -6778 -10749 -6451
tri -10749 -6778 -9900 -5929 sw
tri -9900 -6529 -9300 -5929 ne
rect -12206 -7300 -9900 -6778
rect -29251 -7606 -27500 -7300
tri -30100 -7855 -29851 -7606 se
rect -29851 -7855 -27500 -7606
rect -30100 -8083 -27500 -7855
tri -27500 -8083 -26717 -7300 nw
tri -26651 -8083 -25868 -7300 se
rect -25868 -8083 -25500 -7300
rect -30100 -33755 -28100 -8083
tri -28100 -8683 -27500 -8083 nw
tri -27500 -8932 -26651 -8083 se
rect -26651 -8932 -25500 -8083
rect -27500 -32907 -25500 -8932
tri -25500 -9760 -23040 -7300 nw
tri -19560 -9760 -17100 -7300 ne
rect -17100 -8083 -16732 -7300
tri -16732 -8083 -15949 -7300 sw
tri -15883 -8083 -15100 -7300 ne
rect -15100 -7855 -13055 -7300
tri -13055 -7855 -12500 -7300 sw
tri -12206 -7606 -11900 -7300 ne
rect -15100 -8083 -12500 -7855
rect -17100 -8932 -15949 -8083
tri -15949 -8932 -15100 -8083 sw
tri -15100 -8683 -14500 -8083 ne
tri -28100 -33755 -27500 -33155 sw
tri -27500 -33755 -26652 -32907 ne
rect -26652 -33755 -25500 -32907
rect -30100 -33984 -27500 -33755
tri -30700 -34832 -30100 -34232 sw
tri -30100 -34832 -29252 -33984 ne
rect -29252 -34588 -27500 -33984
tri -27500 -34588 -26667 -33755 sw
tri -26652 -34588 -25819 -33755 ne
rect -25819 -34588 -25500 -33755
rect -29252 -34832 -26667 -34588
rect -32700 -35061 -30100 -34832
tri -30100 -35061 -29871 -34832 sw
tri -29252 -35061 -29023 -34832 ne
rect -29023 -34907 -26667 -34832
tri -26667 -34907 -26348 -34588 sw
tri -25819 -34907 -25500 -34588 ne
tri -25500 -34907 -22671 -32078 sw
tri -18199 -32100 -17100 -31001 se
rect -17100 -31830 -15100 -8932
rect -17100 -32100 -15948 -31830
rect -21700 -32300 -15948 -32100
rect -21700 -34500 -21500 -32300
rect -18900 -32678 -15948 -32300
tri -15948 -32678 -15100 -31830 nw
tri -15100 -32678 -14500 -32078 se
rect -14500 -32678 -12500 -8083
rect -18900 -32982 -16252 -32678
tri -16252 -32982 -15948 -32678 nw
tri -15122 -32700 -15100 -32678 se
rect -15100 -32700 -12500 -32678
tri -15404 -32982 -15122 -32700 se
rect -15122 -32907 -12500 -32700
rect -15122 -32982 -13348 -32907
rect -18900 -33830 -17100 -32982
tri -17100 -33830 -16252 -32982 nw
tri -16252 -33830 -15404 -32982 se
rect -15404 -33755 -13348 -32982
tri -13348 -33755 -12500 -32907 nw
tri -12500 -33755 -11900 -33155 se
rect -11900 -33755 -9900 -7300
rect -15404 -33830 -13423 -33755
tri -13423 -33830 -13348 -33755 nw
tri -12575 -33830 -12500 -33755 se
rect -12500 -33830 -9900 -33755
rect -18900 -34500 -17948 -33830
rect -21700 -34678 -17948 -34500
tri -17948 -34678 -17100 -33830 nw
tri -17100 -34678 -16252 -33830 se
rect -16252 -34678 -14271 -33830
tri -14271 -34678 -13423 -33830 nw
tri -13423 -34678 -12575 -33830 se
rect -12575 -33984 -9900 -33830
rect -12575 -34678 -10748 -33984
rect -21700 -34700 -17970 -34678
tri -17970 -34700 -17948 -34678 nw
rect -29023 -35061 -26348 -34907
tri -32700 -37736 -30025 -35061 ne
rect -30025 -35909 -29871 -35061
tri -29871 -35909 -29023 -35061 sw
tri -29023 -35909 -28175 -35061 ne
rect -28175 -35755 -26348 -35061
tri -26348 -35755 -25500 -34907 sw
tri -25500 -35755 -24652 -34907 ne
rect -24652 -35300 -22671 -34907
tri -22671 -35300 -22278 -34907 sw
tri -17722 -35300 -17100 -34678 se
rect -17100 -35300 -14893 -34678
tri -14893 -35300 -14271 -34678 nw
tri -14045 -35300 -13423 -34678 se
rect -13423 -34832 -10748 -34678
tri -10748 -34832 -9900 -33984 nw
tri -9900 -34832 -9300 -34232 se
rect -9300 -34832 -7300 -5929
rect -13423 -34907 -10823 -34832
tri -10823 -34907 -10748 -34832 nw
tri -9975 -34907 -9900 -34832 se
rect -9900 -34907 -7300 -34832
rect -13423 -35300 -11671 -34907
rect -24652 -35755 -15348 -35300
tri -15348 -35755 -14893 -35300 nw
tri -14500 -35755 -14045 -35300 se
rect -14045 -35755 -11671 -35300
tri -11671 -35755 -10823 -34907 nw
tri -10823 -35755 -9975 -34907 se
rect -9975 -35061 -7300 -34907
rect -9975 -35755 -9300 -35061
rect -28175 -35909 -25500 -35755
rect -30025 -36757 -29023 -35909
tri -29023 -36757 -28175 -35909 sw
tri -28175 -36757 -27327 -35909 ne
rect -27327 -36452 -25500 -35909
tri -25500 -36452 -24803 -35755 sw
tri -24652 -36452 -23955 -35755 ne
rect -23955 -36452 -16045 -35755
tri -16045 -36452 -15348 -35755 nw
tri -15197 -36452 -14500 -35755 se
rect -14500 -35984 -11900 -35755
tri -11900 -35984 -11671 -35755 nw
tri -11052 -35984 -10823 -35755 se
rect -10823 -35984 -9300 -35755
rect -14500 -36452 -12748 -35984
rect -27327 -36757 -24803 -36452
rect -30025 -36888 -28175 -36757
tri -28175 -36888 -28044 -36757 sw
tri -27327 -36888 -27196 -36757 ne
rect -27196 -36888 -24803 -36757
rect -30025 -37736 -28044 -36888
tri -28044 -37736 -27196 -36888 sw
tri -27196 -37736 -26348 -36888 ne
rect -26348 -37300 -24803 -36888
tri -24803 -37300 -23955 -36452 sw
tri -23955 -37300 -23107 -36452 ne
rect -23107 -37300 -16893 -36452
tri -16893 -37300 -16045 -36452 nw
tri -16045 -37300 -15197 -36452 se
rect -15197 -36832 -12748 -36452
tri -12748 -36832 -11900 -35984 nw
tri -11900 -36832 -11052 -35984 se
rect -11052 -36832 -9300 -35984
rect -15197 -37052 -12968 -36832
tri -12968 -37052 -12748 -36832 nw
tri -12120 -37052 -11900 -36832 se
rect -11900 -37052 -9300 -36832
rect -15197 -37300 -13816 -37052
rect -26348 -37736 -23955 -37300
tri -30025 -40500 -27261 -37736 ne
rect -27261 -38584 -27196 -37736
tri -27196 -38584 -26348 -37736 sw
tri -26348 -38584 -25500 -37736 ne
rect -25500 -37900 -23955 -37736
tri -23955 -37900 -23355 -37300 sw
tri -16645 -37900 -16045 -37300 se
rect -16045 -37900 -13816 -37300
tri -13816 -37900 -12968 -37052 nw
tri -12968 -37900 -12120 -37052 se
rect -12120 -37061 -9300 -37052
tri -9300 -37061 -7300 -35061 nw
rect -12120 -37900 -11900 -37061
rect -25500 -38584 -14500 -37900
tri -14500 -38584 -13816 -37900 nw
tri -13652 -38584 -12968 -37900 se
rect -12968 -38584 -11900 -37900
rect -27261 -39052 -26348 -38584
tri -26348 -39052 -25880 -38584 sw
tri -25500 -39052 -25032 -38584 ne
rect -25032 -39052 -15348 -38584
rect -27261 -39900 -25880 -39052
tri -25880 -39900 -25032 -39052 sw
tri -25032 -39900 -24184 -39052 ne
rect -24184 -39432 -15348 -39052
tri -15348 -39432 -14500 -38584 nw
tri -14500 -39432 -13652 -38584 se
rect -13652 -39432 -11900 -38584
rect -24184 -39900 -15816 -39432
tri -15816 -39900 -15348 -39432 nw
tri -14968 -39900 -14500 -39432 se
rect -14500 -39661 -11900 -39432
tri -11900 -39661 -9300 -37061 nw
rect -27261 -40500 -25032 -39900
tri -25032 -40500 -24432 -39900 sw
tri -15568 -40500 -14968 -39900 se
rect -14968 -40500 -14500 -39900
tri -27261 -42500 -25261 -40500 ne
rect -25261 -42261 -14500 -40500
tri -14500 -42261 -11900 -39661 nw
rect -25261 -42500 -14739 -42261
tri -14739 -42500 -14500 -42261 nw
<< end >>
