magic
tech sky130B
timestamp 1662317335
<< metal4 >>
rect 17000 -6550 17300 -6100
rect 16500 -8650 16800 -6650
rect 17500 -6850 17800 -5950
rect 18000 -7300 18300 -6000
rect 17000 -9550 17300 -7300
rect 18500 -7700 18800 -6200
rect 0 -19550 300 -17400
rect 500 -19900 800 -17850
rect 0 -83850 300 -19950
rect 0 -94750 300 -84450
rect 500 -85250 800 -20300
rect 1000 -20350 1300 -18350
rect 500 -93200 800 -85700
rect 1000 -85950 1300 -20750
rect 1500 -20850 1800 -18850
rect 1000 -92000 1300 -86500
rect 1500 -86650 1800 -21300
rect 2000 -21400 2300 -19250
rect 2000 -25850 2300 -21850
rect 2500 -22050 2800 -19750
rect 2500 -24900 2800 -22500
rect 3000 -22600 3300 -20300
rect 3000 -24450 3300 -23150
rect 3500 -23300 3800 -20750
rect 3500 -23900 3800 -23600
rect 4000 -23700 4300 -20900
rect 4500 -23200 4800 -20900
rect 5000 -22650 5300 -20600
rect 5500 -22150 5800 -20150
rect 6000 -21700 6300 -19750
rect 6500 -21300 6800 -19350
rect 7000 -20900 7300 -18900
rect 7500 -20450 7800 -18500
rect 8000 -20000 8300 -18050
rect 8500 -19600 8800 -17600
rect 9000 -19200 9300 -17250
rect 9500 -18800 9800 -16850
rect 10000 -18400 10300 -16500
rect 10500 -17950 10800 -16150
rect 11000 -17600 11300 -15750
rect 11500 -17300 11800 -15250
rect 12000 -17050 12300 -14700
rect 12500 -16800 12800 -14150
rect 13000 -15550 13300 -13700
rect 13500 -15150 13800 -13200
rect 14000 -14750 14300 -12800
rect 14500 -14300 14800 -12350
rect 15000 -13950 15300 -12000
rect 15500 -13500 15800 -11650
rect 16000 -13100 16300 -11250
rect 16500 -12750 16800 -10850
rect 17000 -12350 17300 -10300
rect 17500 -12050 17800 -7950
rect 19000 -8000 19300 -6350
rect 18500 -8500 18800 -8150
rect 19500 -8200 19800 -6550
rect 20000 -8300 20300 -6650
rect 20500 -8350 20800 -6750
rect 18000 -11700 18300 -8550
rect 19000 -9000 19300 -8350
rect 21000 -8400 21300 -6800
rect 21500 -8450 21800 -6850
rect 22000 -8400 22300 -6850
rect 22500 -8300 22800 -6800
rect 23000 -8250 23300 -6750
rect 23500 -8200 23800 -6700
rect 24000 -8150 24300 -6700
rect 24500 -8050 24800 -6700
rect 25000 -8000 25300 -6650
rect 25500 -8000 25800 -6650
rect 26000 -8100 26300 -6700
rect 26500 -8150 26800 -6700
rect 27000 -8200 27300 -6700
rect 27500 -8250 27800 -6800
rect 28000 -8300 28300 -6850
rect 18500 -11400 18800 -9050
rect 19500 -9500 19800 -8500
rect 19000 -11200 19300 -9500
rect 20000 -9950 20300 -8650
rect 19500 -11000 19800 -10000
rect 20500 -10400 20800 -8750
rect 20000 -10850 20300 -10450
rect 21000 -10750 21300 -8800
rect 14000 -15700 14300 -15200
rect 14500 -15700 14800 -14800
rect 15000 -15700 15300 -14350
rect 15500 -15800 15800 -13950
rect 16000 -15950 16300 -13600
rect 13000 -16600 13300 -16250
rect 13500 -16600 13800 -16050
rect 2000 -76900 2300 -27700
rect 2500 -27950 2800 -26150
rect 2500 -71600 2800 -28500
rect 3000 -28750 3300 -25500
rect 3000 -68950 3300 -29200
rect 3500 -29300 3800 -24850
rect 4000 -29750 4300 -24300
rect 3500 -62850 3800 -29800
rect 4500 -30100 4800 -23700
rect 4000 -59800 4300 -30200
rect 5000 -30400 5300 -23200
rect 4500 -38750 4800 -30500
rect 5500 -30650 5800 -22700
rect 5000 -36250 5300 -30800
rect 6000 -31000 6300 -22200
rect 5500 -34350 5800 -31050
rect 6500 -31300 6800 -21750
rect 6000 -33300 6300 -31300
rect 6500 -32500 6800 -31600
rect 5500 -36250 5800 -35400
rect 6000 -35950 6300 -34100
rect 6500 -35350 6800 -33150
rect 7000 -34800 7300 -21350
rect 7500 -34300 7800 -20900
rect 8000 -33800 8300 -20500
rect 8500 -33400 8800 -20050
rect 9000 -33000 9300 -19650
rect 9500 -32650 9800 -19250
rect 10000 -32250 10300 -18800
rect 10500 -31900 10800 -18450
rect 11000 -31600 11300 -18050
rect 11500 -31350 11800 -17750
rect 12000 -31100 12300 -17450
rect 12500 -30900 12800 -17200
rect 13000 -30650 13300 -17000
rect 13500 -30450 13800 -16900
rect 14000 -30250 14300 -16000
rect 14500 -30100 14800 -16000
rect 15000 -30000 15300 -16000
rect 16500 -16200 16800 -13200
rect 15500 -30050 15800 -16200
rect 5000 -37550 5300 -37250
rect 4500 -42850 4800 -40450
rect 5000 -42750 5300 -38350
rect 5500 -42100 5800 -37400
rect 6000 -41600 6300 -36450
rect 6500 -41250 6800 -35950
rect 4500 -57500 4800 -43600
rect 5000 -55900 5300 -43300
rect 5500 -54250 5800 -42650
rect 6000 -53100 6300 -42050
rect 6500 -51900 6800 -44700
rect 7000 -45350 7300 -35300
rect 7000 -50800 7300 -46250
rect 7500 -46350 7800 -34850
rect 7500 -50100 7800 -47100
rect 8000 -47150 8300 -34350
rect 8500 -47800 8800 -33900
rect 8000 -49550 8300 -47800
rect 9000 -47950 9300 -33450
rect 9500 -48000 9800 -33000
rect 8500 -49000 8800 -48200
rect 9000 -48700 9300 -48250
rect 9500 -48600 9800 -48300
rect 10000 -48400 10300 -32700
rect 10500 -48050 10800 -32350
rect 11000 -47750 11300 -32000
rect 11500 -47550 11800 -31750
rect 12000 -47400 12300 -31450
rect 12500 -47500 12800 -31250
rect 13000 -47550 13300 -31000
rect 13500 -47650 13800 -30800
rect 14000 -47750 14300 -30600
rect 14500 -47850 14800 -30450
rect 15000 -47900 15300 -30350
rect 15500 -38650 15800 -30400
rect 16000 -38500 16300 -16300
rect 17000 -16450 17300 -12800
rect 16500 -38300 16800 -16500
rect 17000 -17600 17300 -16750
rect 17500 -17850 17800 -12400
rect 17000 -38050 17300 -17950
rect 18000 -18250 18300 -12100
rect 17500 -28650 17800 -18350
rect 18500 -18600 18800 -11800
rect 18000 -27800 18300 -18700
rect 19000 -18900 19300 -11600
rect 18500 -27000 18800 -19000
rect 19500 -19150 19800 -11400
rect 20000 -19300 20300 -11200
rect 20500 -19300 20800 -11100
rect 21000 -19250 21300 -11050
rect 21500 -19100 21800 -8800
rect 22000 -19000 22300 -8800
rect 22500 -18850 22800 -8700
rect 23000 -18750 23300 -8550
rect 23500 -18550 23800 -8500
rect 24000 -18400 24300 -8500
rect 24500 -18250 24800 -8400
rect 25000 -18000 25300 -8400
rect 25500 -17800 25800 -8400
rect 28500 -8450 28800 -6950
rect 26000 -17650 26300 -8500
rect 26500 -17550 26800 -8500
rect 27000 -17350 27300 -8500
rect 27500 -17350 27800 -8600
rect 29000 -8650 29300 -7100
rect 28000 -17650 28300 -8750
rect 29500 -8800 29800 -7200
rect 28500 -17000 28800 -8850
rect 30000 -8950 30300 -7350
rect 29000 -16300 29300 -9000
rect 30500 -9100 30800 -7500
rect 29500 -15700 29800 -9150
rect 31000 -9300 31300 -7700
rect 30000 -15150 30300 -9300
rect 31500 -9500 31800 -7850
rect 30500 -14650 30800 -9500
rect 31000 -14100 31300 -9650
rect 32000 -9800 32300 -8100
rect 31500 -13600 31800 -9900
rect 32500 -10050 32800 -8300
rect 32000 -13150 32300 -10150
rect 33000 -10350 33300 -8600
rect 32500 -12650 32800 -10450
rect 33500 -10800 33800 -8800
rect 33000 -12150 33300 -10800
rect 34000 -11200 34300 -9000
rect 34500 -10950 34800 -8950
rect 35000 -10600 35300 -8750
rect 35500 -10250 35800 -8450
rect 36000 -9950 36300 -8150
rect 36500 -9600 36800 -7800
rect 37000 -9300 37300 -7550
rect 37500 -9000 37800 -7250
rect 38000 -8700 38300 -7000
rect 38500 -8400 38800 -6700
rect 39000 -8150 39300 -6450
rect 39500 -7900 39800 -6200
rect 40000 -7650 40300 -6000
rect 40500 -7400 40800 -5750
rect 41000 -7200 41300 -5550
rect 41500 -6950 41800 -5300
rect 42000 -6750 42300 -5100
rect 42500 -6500 42800 -4850
rect 43000 -6250 43300 -4650
rect 43500 -6000 43800 -4500
rect 44000 -5800 44300 -4400
rect 44500 -5600 44800 -4300
rect 45000 -5400 45300 -4300
rect 45500 -5300 45800 -4450
rect 19000 -26400 19300 -19300
rect 19500 -25750 19800 -19500
rect 20000 -25200 20300 -19600
rect 20500 -24700 20800 -19600
rect 21000 -24250 21300 -19550
rect 21500 -23750 21800 -19450
rect 22000 -23350 22300 -19300
rect 22500 -22950 22800 -19200
rect 23000 -22500 23300 -19050
rect 23500 -22150 23800 -18850
rect 24000 -21750 24300 -18700
rect 24500 -21450 24800 -18550
rect 25000 -21150 25300 -18400
rect 25500 -20850 25800 -18200
rect 26000 -20450 26300 -18000
rect 26500 -19800 26800 -17850
rect 27000 -19150 27300 -17700
rect 27500 -18500 27800 -17650
rect 21500 -24650 21800 -24250
rect 22000 -24300 22300 -23800
rect 22500 -24050 22800 -23400
rect 23000 -23800 23300 -23000
rect 23500 -23550 23800 -22600
rect 24000 -23300 24300 -22200
rect 24500 -23150 24800 -21800
rect 25000 -22950 25300 -21500
rect 17500 -37700 17800 -29100
rect 18000 -37300 18300 -28400
rect 18500 -36750 18800 -27950
rect 19000 -36200 19300 -27150
rect 19500 -35700 19800 -26650
rect 20000 -35150 20300 -26100
rect 20500 -34550 20800 -25750
rect 21000 -34100 21300 -25300
rect 21500 -26700 21800 -25000
rect 22000 -26100 22300 -24700
rect 22500 -25500 22800 -24400
rect 23000 -25050 23300 -24150
rect 23500 -24650 23800 -23900
rect 24000 -24250 24300 -23650
rect 24500 -23950 24800 -23450
rect 25000 -23800 25300 -23250
rect 21500 -33600 21800 -27000
rect 22000 -33100 22300 -26500
rect 22500 -32600 22800 -25950
rect 23000 -32100 23300 -25450
rect 23500 -31550 23800 -25000
rect 24000 -31100 24300 -24600
rect 24500 -30700 24800 -24300
rect 25000 -30250 25300 -24100
rect 25500 -29900 25800 -21350
rect 26000 -29500 26300 -21250
rect 26500 -29150 26800 -20350
rect 27000 -28800 27300 -19700
rect 27500 -28500 27800 -19050
rect 28000 -28150 28300 -18300
rect 28500 -27850 28800 -17550
rect 29000 -27550 29300 -16850
rect 29500 -27150 29800 -16250
rect 30000 -26900 30300 -15700
rect 30500 -26650 30800 -15100
rect 31000 -26450 31300 -14600
rect 31500 -26250 31800 -14150
rect 32000 -26000 32300 -13650
rect 32500 -25800 32800 -13100
rect 33000 -25600 33300 -12650
rect 33500 -21200 33800 -12200
rect 34000 -20300 34300 -11800
rect 34500 -19350 34800 -11350
rect 35000 -18500 35300 -11000
rect 35500 -17700 35800 -10700
rect 36000 -16950 36300 -10350
rect 36500 -16200 36800 -10050
rect 37000 -15500 37300 -9700
rect 37500 -14800 37800 -9400
rect 38000 -14200 38300 -9100
rect 38500 -13600 38800 -8800
rect 39000 -12950 39300 -8500
rect 39500 -12400 39800 -8250
rect 40000 -11800 40300 -8000
rect 40500 -11250 40800 -7750
rect 41000 -10800 41300 -7600
rect 41500 -10350 41800 -7350
rect 42000 -10000 42300 -7150
rect 42500 -9600 42800 -6850
rect 43000 -9300 43300 -6600
rect 43500 -8950 43800 -6350
rect 34500 -21100 34800 -20050
rect 35000 -20200 35300 -19200
rect 35500 -19300 35800 -18400
rect 36000 -18650 36300 -17550
rect 36500 -18050 36800 -16800
rect 37000 -17600 37300 -16050
rect 37500 -17300 37800 -15350
rect 38000 -17300 38300 -14800
rect 35000 -20800 35300 -20500
rect 35500 -21450 35800 -19850
rect 34000 -23800 34300 -22200
rect 33500 -25450 33800 -24250
rect 34500 -24450 34800 -21550
rect 34000 -25250 34300 -24450
rect 35000 -24650 35300 -21600
rect 35500 -24700 35800 -21950
rect 36000 -24700 36300 -19100
rect 36500 -24700 36800 -18550
rect 37000 -24800 37300 -18000
rect 37500 -19750 37800 -17700
rect 38000 -19950 38300 -18700
rect 38500 -19750 38800 -14150
rect 39000 -19550 39300 -13550
rect 39500 -19350 39800 -12700
rect 40000 -19200 40300 -12300
rect 40500 -19150 40800 -11800
rect 41000 -19100 41300 -11300
rect 41500 -19100 41800 -10850
rect 15500 -47800 15800 -39050
rect 16500 -39250 16800 -38650
rect 16000 -47550 16300 -39400
rect 17000 -39450 17300 -38450
rect 17500 -39600 17800 -38150
rect 16500 -47300 16800 -39650
rect 18000 -39700 18300 -37750
rect 18500 -39800 18800 -37250
rect 17000 -47000 17300 -39800
rect 19000 -39850 19300 -36750
rect 19500 -39800 19800 -36200
rect 20000 -39800 20300 -35650
rect 17500 -46650 17800 -39950
rect 18000 -46250 18300 -40050
rect 18500 -44150 18800 -40150
rect 19000 -42100 19300 -40200
rect 19500 -40650 19800 -40350
rect 18500 -45950 18800 -45650
rect 11000 -48550 11300 -48250
rect 4000 -68450 4300 -63850
rect 4500 -68100 4800 -60550
rect 5000 -67950 5300 -57650
rect 5500 -67800 5800 -56100
rect 6000 -67750 6300 -54600
rect 6500 -67750 6800 -53650
rect 7000 -67750 7300 -52800
rect 7500 -67650 7800 -51850
rect 8000 -67650 8300 -51150
rect 8500 -67700 8800 -50550
rect 9000 -67700 9300 -50050
rect 9500 -67700 9800 -49400
rect 10000 -67700 10300 -49150
rect 10500 -67800 10800 -48900
rect 11000 -67800 11300 -48850
rect 11500 -67900 11800 -48250
rect 12000 -68000 12300 -48050
rect 16500 -48100 16800 -47750
rect 4500 -68750 4800 -68400
rect 5000 -68650 5300 -68250
rect 5500 -68550 5800 -68100
rect 6000 -68500 6300 -68050
rect 6500 -68400 6800 -68050
rect 7000 -68350 7300 -68050
rect 7500 -68350 7800 -68050
rect 8000 -68400 8300 -68100
rect 8500 -68400 8800 -68100
rect 9000 -68350 9300 -68050
rect 9500 -68350 9800 -68000
rect 10000 -68350 10300 -68000
rect 10500 -68400 10800 -68100
rect 11000 -68400 11300 -68100
rect 12500 -68150 12800 -48100
rect 13000 -68400 13300 -48150
rect 3000 -70950 3300 -70650
rect 3500 -70800 3800 -70300
rect 4000 -70550 4300 -69950
rect 4500 -70450 4800 -69650
rect 5000 -70350 5300 -69350
rect 5500 -70300 5800 -69150
rect 6000 -70200 6300 -69050
rect 6500 -70150 6800 -68950
rect 7000 -70150 7300 -68850
rect 7500 -70150 7800 -68850
rect 8000 -70200 8300 -68850
rect 8500 -70300 8800 -68850
rect 9000 -70450 9300 -68900
rect 4000 -71300 4300 -70900
rect 4500 -71150 4800 -70750
rect 5000 -71000 5300 -70650
rect 5500 -70900 5800 -70600
rect 6000 -70900 6300 -70600
rect 7000 -70750 7300 -70450
rect 7500 -70750 7800 -70450
rect 9500 -70650 9800 -68950
rect 10500 -69000 10800 -68700
rect 11000 -69000 11300 -68700
rect 11500 -69050 11800 -68550
rect 13500 -68600 13800 -48150
rect 10000 -70700 10300 -69050
rect 12000 -69100 12300 -68600
rect 14000 -68700 14300 -48250
rect 12500 -69100 12800 -68700
rect 13000 -69250 13300 -68800
rect 14500 -68900 14800 -48400
rect 13500 -69300 13800 -69000
rect 15000 -69150 15300 -48500
rect 17000 -48750 17300 -47400
rect 10500 -70800 10800 -69300
rect 11000 -70800 11300 -69300
rect 11500 -70900 11800 -69350
rect 15500 -69400 15800 -48800
rect 17500 -49150 17800 -47050
rect 16000 -67750 16300 -49150
rect 16500 -65500 16800 -49500
rect 18000 -49600 18300 -46850
rect 18500 -47200 18800 -46900
rect 17000 -64400 17300 -49650
rect 18500 -49750 18800 -48450
rect 19000 -49300 19300 -43400
rect 17500 -63450 17800 -49800
rect 18000 -62200 18300 -50100
rect 18500 -60100 18800 -50550
rect 19500 -51200 19800 -41550
rect 20000 -51300 20300 -40300
rect 20500 -51200 20800 -35100
rect 19000 -52750 19300 -51300
rect 19000 -53350 19300 -53050
rect 18500 -62850 18800 -61850
rect 19000 -62500 19300 -53650
rect 19500 -56500 19800 -52050
rect 19500 -60200 19800 -57200
rect 20000 -57850 20300 -52200
rect 20500 -52400 20800 -51500
rect 21000 -53400 21300 -34600
rect 21500 -53150 21800 -34100
rect 22000 -52750 22300 -33600
rect 22500 -52350 22800 -33000
rect 23000 -52000 23300 -32550
rect 23500 -51550 23800 -32150
rect 24000 -51100 24300 -31600
rect 24500 -50700 24800 -31150
rect 25000 -50400 25300 -30750
rect 25500 -49800 25800 -30350
rect 26000 -49550 26300 -29950
rect 26500 -49050 26800 -29600
rect 27000 -48600 27300 -29250
rect 27500 -48050 27800 -28900
rect 28000 -47600 28300 -28600
rect 28500 -42100 28800 -28250
rect 29000 -40100 29300 -27950
rect 29500 -40400 29800 -27650
rect 29000 -42100 29300 -40500
rect 30000 -40850 30300 -27300
rect 30500 -41200 30800 -27050
rect 29500 -42100 29800 -41200
rect 31000 -41450 31300 -26800
rect 31500 -41750 31800 -26600
rect 30000 -42100 30300 -41800
rect 32000 -42000 32300 -26350
rect 32500 -42050 32800 -26150
rect 33000 -41550 33300 -26000
rect 33500 -40900 33800 -25850
rect 34000 -40250 34300 -25800
rect 34500 -39600 34800 -25650
rect 35000 -34550 35300 -25500
rect 35500 -33850 35800 -25350
rect 36000 -33200 36300 -25250
rect 36500 -32700 36800 -25150
rect 37000 -32200 37300 -25100
rect 37500 -31700 37800 -20800
rect 38000 -24000 38300 -20450
rect 38500 -23750 38800 -20100
rect 39000 -23550 39300 -19850
rect 39500 -23250 39800 -19650
rect 40000 -22900 40300 -19500
rect 40500 -22150 40800 -19500
rect 41000 -20950 41300 -19400
rect 38000 -31350 38300 -24300
rect 38500 -30900 38800 -24050
rect 39000 -30500 39300 -23900
rect 39500 -30100 39800 -23700
rect 40000 -24350 40300 -24050
rect 40000 -24950 40300 -24650
rect 40000 -26950 40300 -25300
rect 40500 -25400 40800 -22900
rect 41000 -24450 41300 -21950
rect 41500 -23500 41800 -20300
rect 42000 -22550 42300 -10500
rect 42500 -21200 42800 -10100
rect 43000 -19750 43300 -9700
rect 43500 -9900 43800 -9600
rect 43500 -17550 43800 -10650
rect 44000 -14300 44300 -6150
rect 44500 -9500 44800 -6000
rect 44500 -10300 44800 -10000
rect 44500 -11100 44800 -10800
rect 42000 -24000 42300 -23300
rect 40000 -29700 40300 -27500
rect 40500 -29400 40800 -27000
rect 41000 -29100 41300 -26150
rect 41500 -28900 41800 -25150
rect 36000 -34550 36300 -33750
rect 36500 -34450 36800 -33200
rect 35000 -38850 35300 -35000
rect 35500 -38050 35800 -35050
rect 36000 -37200 36300 -34950
rect 37000 -37350 37300 -32700
rect 28500 -47100 28800 -42400
rect 33500 -42500 33800 -41550
rect 29000 -46550 29300 -42500
rect 29500 -45900 29800 -42600
rect 34000 -42700 34300 -40900
rect 30000 -45300 30300 -42750
rect 34500 -42850 34800 -40200
rect 35000 -42750 35300 -39500
rect 35500 -42550 35800 -38650
rect 36000 -42450 36300 -37800
rect 36500 -42300 36800 -37400
rect 37000 -42300 37300 -38400
rect 37500 -38700 37800 -32250
rect 37500 -42300 37800 -39400
rect 38000 -39550 38300 -31800
rect 38500 -40100 38800 -31400
rect 38000 -42350 38300 -40100
rect 39000 -40650 39300 -30950
rect 38500 -42500 38800 -40650
rect 39500 -41100 39800 -30550
rect 39000 -42700 39300 -41150
rect 30500 -44550 30800 -43200
rect 31000 -44100 31300 -43250
rect 36500 -43300 36800 -43000
rect 37000 -43350 37300 -42850
rect 31500 -43650 31800 -43350
rect 31500 -44850 31800 -44050
rect 32000 -44800 32300 -43500
rect 32500 -44450 32800 -43550
rect 33000 -44000 33300 -43700
rect 26000 -51350 26300 -50050
rect 20000 -58450 20300 -58150
rect 20500 -59400 20800 -53500
rect 21000 -60850 21300 -53900
rect 18000 -64950 18300 -63450
rect 18500 -64100 18800 -63150
rect 17500 -65400 17800 -65100
rect 12000 -70900 12300 -69400
rect 12500 -70950 12800 -69450
rect 2500 -73700 2800 -72100
rect 2000 -79450 2300 -78200
rect 2500 -83750 2800 -79550
rect 2500 -84400 2800 -84050
rect 1500 -91150 1800 -87100
rect 2000 -87250 2300 -85650
rect 2000 -90300 2300 -87750
rect 3000 -88300 3300 -74600
rect 3500 -88100 3800 -73150
rect 4000 -84500 4300 -72400
rect 4500 -84150 4800 -72000
rect 5000 -83800 5300 -71700
rect 5500 -83500 5800 -71500
rect 6000 -83250 6300 -71350
rect 6500 -83050 6800 -71200
rect 7000 -82850 7300 -71150
rect 7500 -82700 7800 -71100
rect 8000 -82550 8300 -71000
rect 8500 -82500 8800 -71000
rect 9000 -82400 9300 -71000
rect 9500 -82250 9800 -71050
rect 13000 -71100 13300 -69600
rect 10000 -82150 10300 -71100
rect 10500 -82000 10800 -71100
rect 13500 -71200 13800 -69650
rect 11000 -81900 11300 -71200
rect 11500 -81700 11800 -71300
rect 14000 -71400 14300 -69800
rect 12000 -81600 12300 -71450
rect 14500 -71550 14800 -69900
rect 12500 -81450 12800 -71600
rect 13000 -81250 13300 -71650
rect 15000 -71750 15300 -69950
rect 13500 -81050 13800 -71750
rect 14000 -80900 14300 -71900
rect 15500 -71950 15800 -70600
rect 14500 -80600 14800 -72100
rect 15000 -80200 15300 -72350
rect 15500 -79750 15800 -72850
rect 16500 -75700 16800 -73350
rect 16500 -78000 16800 -76500
rect 17000 -78800 17300 -72450
rect 17500 -78600 17800 -71800
rect 18000 -78400 18300 -70700
rect 18500 -78250 18800 -69400
rect 19000 -76550 19300 -68150
rect 19500 -76350 19800 -66900
rect 20000 -76100 20300 -64550
rect 20500 -75950 20800 -61500
rect 21000 -75500 21300 -61900
rect 21500 -62150 21800 -53600
rect 22000 -53950 22300 -53650
rect 22500 -54200 22800 -52800
rect 21500 -62750 21800 -62450
rect 21500 -75700 21800 -63050
rect 22000 -63150 22300 -54250
rect 23000 -54700 23300 -52400
rect 22000 -75450 22300 -63750
rect 22500 -64150 22800 -54750
rect 23500 -55150 23800 -52000
rect 26500 -52100 26800 -49550
rect 22500 -75100 22800 -64600
rect 23000 -65150 23300 -55150
rect 24000 -55650 24300 -52400
rect 27000 -52650 27300 -49000
rect 23000 -74750 23300 -65700
rect 23500 -65950 23800 -55700
rect 24500 -56050 24800 -53000
rect 27500 -53150 27800 -48550
rect 28000 -49500 28300 -48100
rect 28500 -50250 28800 -47600
rect 28000 -53500 28300 -50400
rect 29000 -50850 29300 -47000
rect 23500 -74450 23800 -66500
rect 24000 -66650 24300 -56100
rect 25000 -56500 25300 -53500
rect 28500 -53850 28800 -51050
rect 29500 -51450 29800 -46500
rect 24000 -74050 24300 -67050
rect 24500 -67300 24800 -56550
rect 25500 -56850 25800 -54000
rect 29000 -54300 29300 -51600
rect 30000 -52000 30300 -45800
rect 24500 -73800 24800 -67750
rect 25000 -67850 25300 -56900
rect 26000 -57200 26300 -54450
rect 29500 -54650 29800 -52150
rect 30500 -52500 30800 -45250
rect 30000 -54900 30300 -52700
rect 31000 -53000 31300 -45300
rect 31500 -46000 31800 -45700
rect 25000 -73550 25300 -68300
rect 25500 -68400 25800 -57300
rect 26500 -57550 26800 -54900
rect 30500 -55100 30800 -53200
rect 31500 -53550 31800 -48650
rect 32000 -48700 32300 -46550
rect 32500 -49200 32800 -45550
rect 31000 -55100 31300 -53700
rect 32000 -54050 32300 -49300
rect 33000 -49450 33300 -44900
rect 33500 -49600 33800 -44450
rect 34000 -49700 34300 -44050
rect 34500 -49700 34800 -44000
rect 35000 -49650 35300 -44250
rect 35500 -49550 35800 -44400
rect 36000 -49450 36300 -44550
rect 36500 -49200 36800 -44150
rect 37000 -49000 37300 -43800
rect 37500 -48700 37800 -42850
rect 38000 -48350 38300 -42900
rect 39500 -43000 39800 -41700
rect 40000 -41800 40300 -30150
rect 40500 -42000 40800 -29800
rect 41000 -41800 41300 -29450
rect 41500 -41550 41800 -29200
rect 42000 -41300 42300 -24300
rect 42500 -40450 42800 -22200
rect 43000 -39650 43300 -20650
rect 43500 -38700 43800 -18950
rect 44000 -37700 44300 -16600
rect 44500 -36600 44800 -11550
rect 45000 -35950 45300 -8300
rect 45500 -15550 45800 -6200
rect 46000 -11800 46300 -4700
rect 46500 -8450 46800 -5300
rect 46000 -15950 46300 -13050
rect 45500 -34000 45800 -16000
rect 46500 -16400 46800 -14300
rect 56500 -14700 56800 -11450
rect 57000 -11650 57300 -11300
rect 57500 -11600 57800 -11300
rect 58000 -11600 58300 -11300
rect 58500 -11650 58800 -11350
rect 59000 -11850 59300 -11450
rect 62000 -11600 62300 -11300
rect 62500 -11600 62800 -11300
rect 59500 -12350 59800 -11750
rect 63000 -11800 63300 -11300
rect 63500 -11700 63800 -11300
rect 64000 -11600 64300 -11300
rect 64500 -11600 64800 -11300
rect 60000 -14200 60300 -12500
rect 47000 -16450 47300 -14750
rect 38500 -47950 38800 -43050
rect 39000 -47400 39300 -43200
rect 40000 -43550 40300 -42100
rect 39500 -46700 39800 -43550
rect 40500 -44400 40800 -42300
rect 40000 -44950 40300 -44650
rect 40000 -47550 40300 -47250
rect 40500 -47950 40800 -45900
rect 41000 -47750 41300 -42100
rect 41500 -47450 41800 -41950
rect 42000 -47200 42300 -41700
rect 42500 -42800 42800 -40950
rect 43000 -41750 43300 -40000
rect 43500 -40300 43800 -40000
rect 43000 -43600 43300 -42600
rect 43500 -43700 43800 -41200
rect 42500 -47100 42800 -43800
rect 44000 -43850 44300 -39800
rect 44500 -43850 44800 -37750
rect 45000 -43800 45300 -36250
rect 45500 -43800 45800 -34550
rect 46000 -43750 46300 -16450
rect 47500 -16800 47800 -15050
rect 46500 -43600 46800 -16850
rect 48000 -17200 48300 -15400
rect 47000 -43500 47300 -17400
rect 48500 -17650 48800 -15700
rect 49000 -17800 49300 -16050
rect 47500 -43350 47800 -17900
rect 48000 -19100 48300 -18000
rect 48500 -19350 48800 -18100
rect 49500 -18150 49800 -16400
rect 48000 -43150 48300 -19400
rect 49000 -19650 49300 -18300
rect 50000 -18450 50300 -16700
rect 48500 -43000 48800 -19850
rect 49500 -20200 49800 -18550
rect 50500 -18750 50800 -16950
rect 49000 -42850 49300 -20350
rect 49500 -42350 49800 -20850
rect 50000 -20950 50300 -18850
rect 51000 -19100 51300 -17300
rect 50000 -41700 50300 -21550
rect 50500 -21650 50800 -19150
rect 51500 -19400 51800 -17550
rect 50500 -40650 50800 -22300
rect 51000 -22500 51300 -19500
rect 52000 -19800 52300 -17900
rect 56500 -18350 56800 -15000
rect 57000 -15450 57300 -15000
rect 57500 -15400 57800 -15050
rect 58000 -15450 58300 -15050
rect 58500 -16150 58800 -15000
rect 59000 -15300 59300 -14900
rect 59500 -14950 59800 -14400
rect 59000 -17050 59300 -16400
rect 59500 -18050 59800 -17350
rect 63300 -18000 63600 -12000
rect 67000 -12350 67300 -11700
rect 67500 -11800 67800 -11400
rect 68000 -11600 68300 -11300
rect 68500 -11600 68800 -11300
rect 69000 -11700 69300 -11350
rect 69500 -12100 69800 -11600
rect 66500 -13700 66800 -12400
rect 70000 -12850 70300 -12150
rect 67000 -14300 67300 -13650
rect 67500 -14750 67800 -14300
rect 68000 -15050 68300 -14650
rect 68500 -15300 68800 -14900
rect 69000 -15600 69300 -15150
rect 69500 -16100 69800 -15500
rect 66500 -17750 66800 -17300
rect 51000 -39150 51300 -23150
rect 51500 -38850 51800 -19800
rect 52500 -20250 52800 -18400
rect 60000 -18500 60300 -18200
rect 62000 -18750 62300 -18350
rect 62500 -18750 62800 -18350
rect 63000 -18750 63300 -18200
rect 63500 -18750 63800 -18250
rect 64000 -18750 64300 -18350
rect 64500 -18750 64800 -18350
rect 67000 -18400 67300 -17850
rect 70000 -17900 70300 -16150
rect 67500 -18700 67800 -18300
rect 68000 -18800 68300 -18400
rect 68500 -18800 68800 -18400
rect 69000 -18700 69300 -18300
rect 69500 -18400 69800 -17950
rect 72000 -18200 72300 -11550
rect 75000 -17850 75300 -11450
rect 82500 -11950 82800 -11500
rect 83000 -11600 83300 -11300
rect 83500 -11550 83800 -11250
rect 84000 -11600 84300 -11300
rect 84500 -11950 84800 -11500
rect 77000 -15450 77300 -15150
rect 77500 -15450 77800 -15150
rect 78000 -15450 78300 -15150
rect 78500 -15450 78800 -15150
rect 79000 -15450 79300 -15150
rect 79500 -15450 79800 -15150
rect 80000 -15450 80300 -15150
rect 72500 -18600 72800 -18150
rect 73000 -18750 73300 -18400
rect 73500 -18800 73800 -18400
rect 74000 -18700 74300 -18300
rect 74500 -18450 74800 -17950
rect 82000 -18100 82300 -11950
rect 84500 -14400 84800 -14000
rect 82500 -16050 82800 -15550
rect 83000 -15600 83300 -15200
rect 83500 -15250 83800 -14800
rect 84000 -14850 84300 -14400
rect 82500 -18500 82800 -18100
rect 83000 -18750 83300 -18350
rect 83500 -18800 83800 -18400
rect 84000 -18750 84300 -18350
rect 84500 -18550 84800 -18100
rect 85000 -18150 85300 -11900
rect 88500 -12500 88800 -11650
rect 94500 -11750 94800 -11450
rect 88000 -13500 88300 -12650
rect 94000 -12700 94300 -11900
rect 93500 -13650 93800 -12900
rect 87000 -17950 87300 -14800
rect 87500 -15150 87800 -13650
rect 88000 -14800 88300 -14450
rect 88500 -14700 88800 -14400
rect 89000 -14800 89300 -14450
rect 93000 -14650 93300 -13850
rect 89500 -15050 89800 -14650
rect 87500 -18500 87800 -18050
rect 88000 -18750 88300 -18350
rect 88500 -18800 88800 -18400
rect 89000 -18750 89300 -18350
rect 89500 -18550 89800 -18100
rect 90000 -18150 90300 -15000
rect 92500 -15550 92800 -14800
rect 92000 -16600 92300 -15700
rect 92500 -16600 92800 -16300
rect 93000 -16600 93300 -16300
rect 93500 -16600 93800 -16300
rect 94000 -16650 94300 -16300
rect 94500 -18450 94800 -14350
rect 95000 -16600 95300 -16300
rect 43000 -47200 43300 -43950
rect 48000 -44000 48300 -43550
rect 32500 -54550 32800 -49750
rect 33000 -54900 33300 -50000
rect 33500 -55150 33800 -50200
rect 25500 -71950 25800 -68800
rect 26000 -68900 26300 -57650
rect 27000 -57850 27300 -55200
rect 34000 -55300 34300 -50300
rect 34500 -55400 34800 -50300
rect 35000 -55300 35300 -50300
rect 35500 -55250 35800 -50200
rect 36000 -52050 36300 -50100
rect 36500 -52300 36800 -49950
rect 37000 -52350 37300 -49750
rect 36000 -55200 36300 -52350
rect 37500 -52400 37800 -49500
rect 36500 -55100 36800 -52600
rect 37000 -55000 37300 -52650
rect 37500 -54900 37800 -52800
rect 38000 -54850 38300 -49200
rect 38500 -54750 38800 -48850
rect 39000 -54700 39300 -48450
rect 39500 -54650 39800 -48100
rect 40000 -54600 40300 -48250
rect 40500 -54400 40800 -48500
rect 41000 -54350 41300 -48400
rect 41500 -50500 41800 -47900
rect 42000 -49000 42300 -47600
rect 42500 -49800 42800 -47450
rect 42000 -50800 42300 -50500
rect 42500 -50650 42800 -50350
rect 41500 -54200 41800 -51250
rect 42000 -54100 42300 -51150
rect 42500 -53900 42800 -50950
rect 43000 -53650 43300 -48000
rect 43500 -48250 43800 -44050
rect 48500 -44100 48800 -43350
rect 49000 -44050 49300 -43150
rect 49500 -44000 49800 -42850
rect 50000 -43100 50300 -42350
rect 50500 -43250 50800 -42400
rect 51000 -43000 51300 -40950
rect 51500 -42600 51800 -39150
rect 52000 -41900 52300 -20250
rect 52500 -40950 52800 -20650
rect 53000 -20750 53300 -18800
rect 53000 -39600 53300 -21250
rect 53500 -21300 53800 -19200
rect 53500 -38000 53800 -21800
rect 54000 -21900 54300 -19650
rect 54000 -36100 54300 -22450
rect 54500 -22550 54800 -20200
rect 55000 -23100 55300 -20750
rect 54500 -30800 54800 -23150
rect 55500 -23450 55800 -21350
rect 55000 -24350 55300 -23500
rect 56000 -23700 56300 -21850
rect 55500 -24800 55800 -24500
rect 56000 -24800 56300 -24200
rect 56500 -24800 56800 -22350
rect 57000 -24750 57300 -22750
rect 57500 -24800 57800 -23100
rect 54500 -32800 54800 -32300
rect 44000 -47450 44300 -44150
rect 44500 -46400 44800 -44300
rect 50500 -44400 50800 -43750
rect 51000 -44250 51300 -43400
rect 51500 -43550 51800 -43100
rect 45000 -45150 45300 -44850
rect 46000 -47800 46300 -47300
rect 44500 -49000 44800 -48650
rect 45000 -48850 45300 -48400
rect 45500 -48450 45800 -47850
rect 43500 -53350 43800 -49450
rect 44000 -49650 44300 -49200
rect 44500 -50600 44800 -49300
rect 44000 -52950 44300 -50600
rect 45000 -50850 45300 -49200
rect 45500 -51000 45800 -49000
rect 46000 -50200 46300 -48300
rect 46500 -49450 46800 -47650
rect 47000 -48800 47300 -46850
rect 47500 -47050 47800 -46050
rect 48500 -47300 48800 -46650
rect 49000 -46900 49300 -45200
rect 49500 -46400 49800 -44650
rect 50000 -45650 50300 -44650
rect 50500 -45200 50800 -44900
rect 48000 -47750 48300 -47450
rect 47500 -48200 47800 -47800
rect 48500 -48350 48800 -48050
rect 49000 -48600 49300 -47550
rect 46000 -51000 46300 -50550
rect 46500 -50900 46800 -50150
rect 47000 -50700 47300 -49650
rect 47500 -50550 47800 -49050
rect 48000 -50250 48300 -48750
rect 49500 -49000 49800 -47050
rect 50000 -48650 50300 -46450
rect 50500 -47950 50800 -45800
rect 51000 -46550 51300 -45700
rect 51500 -45800 51800 -44400
rect 48500 -50000 48800 -49050
rect 44500 -52300 44800 -51150
rect 26000 -71900 26300 -69350
rect 26500 -69400 26800 -58050
rect 27500 -58200 27800 -55700
rect 27000 -69850 27300 -58400
rect 28000 -58500 28300 -56050
rect 34000 -56200 34300 -55900
rect 34500 -56250 34800 -55800
rect 26500 -71750 26800 -69850
rect 27500 -70200 27800 -58750
rect 28500 -58800 28800 -56350
rect 35000 -56400 35300 -55750
rect 27000 -71700 27300 -70200
rect 28000 -70600 28300 -59100
rect 29000 -59200 29300 -56600
rect 29500 -59450 29800 -56750
rect 28500 -68500 28800 -59450
rect 29000 -68550 29300 -59750
rect 30000 -59800 30300 -57750
rect 34500 -58100 34800 -56750
rect 30500 -60050 30800 -58650
rect 35000 -59200 35300 -56700
rect 29500 -68900 29800 -60050
rect 31000 -60400 31300 -59200
rect 28500 -69500 28800 -68950
rect 29000 -69500 29300 -68900
rect 27500 -71600 27800 -70600
rect 28500 -70900 28800 -69900
rect 28000 -71500 28300 -70900
rect 29000 -71100 29300 -69900
rect 29500 -70900 29800 -69450
rect 30000 -70100 30300 -60450
rect 31500 -60650 31800 -59750
rect 30500 -68850 30800 -60750
rect 31000 -68100 31300 -61000
rect 31500 -66600 31800 -61300
rect 32000 -65150 32300 -61550
rect 32500 -62850 32800 -61700
rect 33000 -61900 33300 -61600
rect 33500 -62350 33800 -59950
rect 34000 -63050 34300 -60500
rect 35500 -60650 35800 -55700
rect 36000 -56500 36300 -55550
rect 36500 -56550 36800 -55400
rect 37000 -56700 37300 -55300
rect 37500 -56750 37800 -55200
rect 33500 -63750 33800 -63200
rect 30500 -69450 30800 -69150
rect 28500 -71500 28800 -71200
rect 30000 -71400 30300 -70950
rect 30500 -71400 30800 -69750
rect 31000 -71400 31300 -68400
rect 31500 -71150 31800 -67700
rect 32000 -67750 32300 -65600
rect 32500 -68000 32800 -64250
rect 33000 -67700 33300 -63900
rect 34000 -64000 34300 -63700
rect 34500 -63900 34800 -61250
rect 36000 -61950 36300 -56800
rect 33500 -67200 33800 -64100
rect 34000 -66100 34300 -64300
rect 35000 -64500 35300 -62100
rect 36500 -62900 36800 -56850
rect 38000 -56950 38300 -55150
rect 35500 -65700 35800 -63000
rect 37000 -63650 37300 -57000
rect 34000 -67650 34300 -66400
rect 34500 -67400 34800 -65700
rect 35000 -66500 35300 -65950
rect 36000 -66550 36300 -64000
rect 36500 -64500 36800 -64200
rect 37500 -64400 37800 -57050
rect 38500 -57100 38800 -55100
rect 39000 -55700 39300 -55400
rect 39000 -56750 39300 -56450
rect 39500 -56650 39800 -54950
rect 38000 -65100 38300 -57250
rect 40000 -57500 40300 -54900
rect 39000 -58050 39300 -57750
rect 38500 -65200 38800 -58150
rect 39000 -65200 39300 -58350
rect 39500 -58400 39800 -58100
rect 40500 -58250 40800 -54700
rect 39500 -65200 39800 -58700
rect 40000 -65100 40300 -58900
rect 41000 -58950 41300 -54650
rect 40500 -65050 40800 -59350
rect 41500 -59650 41800 -54500
rect 41000 -65050 41300 -60100
rect 42000 -60350 42300 -54400
rect 42500 -60750 42800 -54200
rect 43000 -60400 43300 -54000
rect 43500 -59950 43800 -53750
rect 44000 -59400 44300 -53400
rect 44500 -58850 44800 -52800
rect 45000 -58200 45300 -52150
rect 45500 -57500 45800 -51600
rect 46000 -56850 46300 -51500
rect 46500 -56150 46800 -51450
rect 47000 -55200 47300 -51350
rect 47500 -54400 47800 -51200
rect 48000 -53250 48300 -50950
rect 42000 -61750 42300 -61200
rect 42500 -63500 42800 -61250
rect 41500 -65000 41800 -64150
rect 43000 -65000 43300 -60900
rect 43500 -64950 43800 -60500
rect 44000 -64950 44300 -60000
rect 44500 -64950 44800 -59450
rect 45000 -65100 45300 -58800
rect 45500 -65350 45800 -58100
rect 46000 -62300 46300 -57450
rect 46500 -62000 46800 -56750
rect 47000 -58800 47300 -55950
rect 47500 -58050 47800 -55000
rect 48000 -55400 48300 -54950
rect 48500 -55050 48800 -50650
rect 49000 -54450 49300 -50350
rect 49500 -53600 49800 -49950
rect 50000 -52750 50300 -49500
rect 50500 -51900 50800 -48950
rect 51000 -51000 51300 -48200
rect 51500 -50050 51800 -46950
rect 52000 -49100 52300 -43600
rect 52500 -48100 52800 -42700
rect 53000 -47050 53300 -40700
rect 53500 -45750 53800 -39300
rect 54000 -44350 54300 -39350
rect 53500 -48650 53800 -47400
rect 54000 -48200 54300 -45900
rect 54500 -47850 54800 -35300
rect 55000 -47400 55300 -24800
rect 58000 -24850 58300 -23250
rect 58500 -24950 58800 -23450
rect 59000 -25000 59300 -23500
rect 59500 -25050 59800 -23600
rect 55500 -47000 55800 -25100
rect 56000 -33250 56300 -25100
rect 56000 -34100 56300 -33800
rect 56000 -46550 56300 -34400
rect 56500 -34600 56800 -25100
rect 56500 -46050 56800 -35400
rect 57000 -36000 57300 -25100
rect 57000 -36900 57300 -36600
rect 57000 -45500 57300 -37200
rect 57500 -37750 57800 -25150
rect 57500 -38350 57800 -38050
rect 58000 -38200 58300 -25200
rect 58500 -37550 58800 -25250
rect 60000 -25300 60300 -23700
rect 60500 -25250 60800 -23750
rect 59000 -36600 59300 -25300
rect 61000 -25350 61300 -23900
rect 59500 -36200 59800 -25350
rect 61500 -25500 61800 -24000
rect 60000 -35900 60300 -25600
rect 60500 -35450 60800 -25600
rect 62000 -25650 62300 -24150
rect 61000 -35050 61300 -25700
rect 62500 -25800 62800 -24300
rect 61500 -34600 61800 -25800
rect 63000 -26000 63300 -24450
rect 62000 -34250 62300 -26000
rect 62500 -34000 62800 -26150
rect 63500 -26250 63800 -24650
rect 63000 -33650 63300 -26400
rect 64000 -26500 64300 -24850
rect 63500 -33300 63800 -26600
rect 64500 -26700 64800 -25050
rect 64000 -33000 64300 -26850
rect 65000 -26900 65300 -25300
rect 64500 -32750 64800 -27100
rect 65500 -27150 65800 -25500
rect 65000 -32500 65300 -27350
rect 66000 -27500 66300 -25750
rect 65500 -32250 65800 -27650
rect 66500 -27700 66800 -25950
rect 66000 -31900 66300 -27850
rect 67000 -27950 67300 -26200
rect 67500 -28100 67800 -26400
rect 66500 -31700 66800 -28100
rect 68000 -28300 68300 -26600
rect 67000 -31500 67300 -28300
rect 68500 -28450 68800 -26750
rect 67500 -31300 67800 -28500
rect 69000 -28600 69300 -26900
rect 68000 -31150 68300 -28650
rect 69500 -28750 69800 -27050
rect 70000 -28850 70300 -27150
rect 68500 -30900 68800 -28850
rect 70500 -28900 70800 -27250
rect 71000 -28950 71300 -27350
rect 69000 -30600 69300 -28950
rect 71500 -29000 71800 -27450
rect 72000 -29050 72300 -27550
rect 72500 -28950 72800 -27600
rect 73000 -28850 73300 -27750
rect 73500 -28900 73800 -27900
rect 69500 -30400 69800 -29100
rect 70000 -30100 70300 -29200
rect 70500 -29850 70800 -29350
rect 71000 -29700 71300 -29400
rect 61000 -35850 61300 -35550
rect 61500 -35900 61800 -35100
rect 62000 -36100 62300 -34700
rect 57500 -40200 57800 -39900
rect 57500 -44650 57800 -40550
rect 58000 -40950 58300 -38900
rect 58500 -39900 58800 -38150
rect 59000 -40050 59300 -37500
rect 59500 -40200 59800 -36850
rect 60000 -38050 60300 -36400
rect 60500 -37700 60800 -36300
rect 61000 -37300 61300 -36200
rect 61500 -36850 61800 -36250
rect 60000 -40100 60300 -38400
rect 61000 -38750 61300 -37700
rect 60500 -39900 60800 -38750
rect 61000 -39650 61300 -39200
rect 61500 -39300 61800 -37350
rect 58500 -41150 58800 -40300
rect 58500 -42200 58800 -41650
rect 59000 -42000 59300 -40550
rect 59500 -41850 59800 -40500
rect 60000 -41700 60300 -40450
rect 60500 -41150 60800 -40250
rect 61000 -41000 61300 -40000
rect 61500 -40800 61800 -39750
rect 62000 -40450 62300 -36900
rect 62500 -40100 62800 -34350
rect 63000 -39700 63300 -34000
rect 63500 -39250 63800 -33700
rect 64000 -38850 64300 -33450
rect 64500 -38400 64800 -33100
rect 65000 -37900 65300 -32850
rect 65500 -37400 65800 -32600
rect 66000 -36900 66300 -32350
rect 66500 -36400 66800 -32050
rect 67000 -35850 67300 -31850
rect 67500 -35350 67800 -31650
rect 68000 -34750 68300 -31450
rect 68500 -34150 68800 -31200
rect 69000 -33600 69300 -31000
rect 69500 -33050 69800 -30800
rect 70000 -32450 70300 -30550
rect 70500 -31600 70800 -30350
rect 71000 -31050 71300 -30150
rect 71500 -30550 71800 -29400
rect 72000 -30050 72300 -29400
rect 53000 -49000 53300 -48650
rect 52000 -50800 52300 -50500
rect 48000 -57550 48300 -55700
rect 48500 -57150 48800 -55950
rect 49000 -56850 49300 -55150
rect 49500 -56550 49800 -54250
rect 50000 -56100 50300 -53500
rect 50500 -55500 50800 -52600
rect 51000 -54700 51300 -51650
rect 51500 -53850 51800 -50800
rect 52000 -53050 52300 -51150
rect 52500 -52400 52800 -50150
rect 53000 -51800 53300 -49600
rect 53500 -51300 53800 -49100
rect 54000 -50750 54300 -48700
rect 54500 -50250 54800 -48250
rect 55000 -49800 55300 -47850
rect 55500 -49400 55800 -47450
rect 56000 -48950 56300 -47050
rect 56500 -48500 56800 -46600
rect 57000 -48100 57300 -45950
rect 57500 -47600 57800 -45500
rect 58000 -47050 58300 -43750
rect 58500 -46450 58800 -42550
rect 59000 -45500 59300 -42400
rect 59500 -44500 59800 -42200
rect 60000 -43850 60300 -42050
rect 60500 -43450 60800 -41800
rect 61000 -43200 61300 -41550
rect 61500 -42900 61800 -41250
rect 62000 -42650 62300 -40950
rect 62500 -42350 62800 -40550
rect 63000 -42000 63300 -40150
rect 63500 -41700 63800 -39750
rect 64000 -41200 64300 -39300
rect 64500 -40850 64800 -38850
rect 65000 -40400 65300 -38400
rect 65500 -39950 65800 -37950
rect 66000 -39500 66300 -37450
rect 66500 -39050 66800 -36900
rect 67000 -38550 67300 -36350
rect 67500 -38050 67800 -35850
rect 68000 -37500 68300 -35300
rect 68500 -37000 68800 -34700
rect 69000 -36350 69300 -34050
rect 69500 -35850 69800 -33600
rect 70000 -35250 70300 -33200
rect 70500 -34750 70800 -32550
rect 71000 -34200 71300 -31800
rect 71500 -33650 71800 -31200
rect 72000 -33000 72300 -30700
rect 72500 -32450 72800 -30200
rect 73000 -31800 73300 -29800
rect 73500 -31250 73800 -29450
rect 74000 -30600 74300 -28300
rect 47000 -61700 47300 -59700
rect 47500 -61400 47800 -59550
rect 48000 -61150 48300 -59300
rect 48500 -60850 48800 -59050
rect 49000 -60600 49300 -58800
rect 49500 -60300 49800 -58500
rect 50000 -60000 50300 -58250
rect 50500 -59700 50800 -58000
rect 51000 -59400 51300 -57800
rect 51500 -59150 51800 -57600
rect 52000 -58850 52300 -57500
rect 52500 -58600 52800 -57500
rect 53000 -58600 53300 -57550
rect 35000 -67100 35300 -66800
rect 35000 -67750 35300 -67400
rect 32000 -68800 32300 -68150
rect 32000 -71400 32300 -69100
rect 32500 -71450 32800 -68500
rect 33000 -71450 33300 -68200
rect 33500 -71500 33800 -67850
rect 34000 -71300 34300 -67950
rect 34500 -70950 34800 -67950
rect 35000 -70550 35300 -68250
rect 35500 -68950 35800 -66600
rect 36500 -67000 36800 -66150
rect 37000 -67600 37300 -65550
rect 38500 -65800 38800 -65500
rect 39000 -65800 39300 -65500
rect 39500 -65800 39800 -65500
rect 40000 -65800 40300 -65400
rect 40500 -65800 40800 -65500
rect 37500 -67400 37800 -66200
rect 38000 -66650 38300 -66350
rect 38500 -66550 38800 -66100
rect 36000 -68850 36300 -68100
rect 25500 -73300 25800 -72450
rect 26500 -72550 26800 -72050
rect 27000 -72700 27300 -72000
rect 26000 -73050 26300 -72700
rect 27500 -72800 27800 -71900
rect 23000 -75500 23300 -75150
rect 23500 -75450 23800 -75150
rect 24500 -75800 24800 -74950
rect 19000 -77250 19300 -76950
rect 19000 -78100 19300 -77650
rect 19500 -77800 19800 -76650
rect 4500 -85500 4800 -84500
rect 4000 -87400 4300 -85500
rect 5000 -85700 5300 -84200
rect 4500 -86750 4800 -85800
rect 5500 -86000 5800 -83900
rect 5000 -86300 5300 -86000
rect 2500 -89450 2800 -89150
rect 0 -99050 300 -96450
rect 500 -99200 800 -93700
rect 1000 -99400 1300 -92300
rect 1500 -99500 1800 -91700
rect 2000 -99600 2300 -90900
rect 2500 -98750 2800 -89900
rect 3000 -98750 3300 -89200
rect 3500 -98900 3800 -88600
rect 4000 -99000 4300 -87950
rect 4500 -99050 4800 -87500
rect 2500 -99700 2800 -99050
rect 3000 -99700 3300 -99050
rect 5000 -99200 5300 -87050
rect 5500 -99200 5800 -86600
rect 3500 -99800 3800 -99200
rect 6000 -99300 6300 -83650
rect 4000 -99850 4300 -99300
rect 6500 -99450 6800 -83400
rect 7000 -99450 7300 -83200
rect 7500 -99400 7800 -83000
rect 8000 -99450 8300 -82850
rect 8500 -99400 8800 -82800
rect 9000 -99400 9300 -82700
rect 9500 -99300 9800 -82550
rect 10000 -99200 10300 -82450
rect 10500 -99200 10800 -82300
rect 11000 -99250 11300 -82200
rect 11500 -99550 11800 -82050
rect 15500 -87450 15800 -80250
rect 16000 -85900 16300 -79900
rect 16500 -84750 16800 -79550
rect 17000 -83900 17300 -79200
rect 17500 -82900 17800 -78900
rect 15500 -89900 15800 -88100
rect 16000 -89900 16300 -86250
rect 16500 -89700 16800 -85100
rect 17000 -89550 17300 -84250
rect 17500 -89400 17800 -83400
rect 18000 -89550 18300 -78700
rect 17500 -99650 17800 -89700
rect 18000 -98350 18300 -90050
rect 18500 -91550 18800 -78550
rect 18500 -92150 18800 -91850
rect 18000 -99200 18300 -98650
rect 18500 -98950 18800 -92450
rect 19000 -92850 19300 -78500
rect 19000 -98550 19300 -93450
rect 19500 -93750 19800 -78300
rect 19500 -98150 19800 -94250
rect 20000 -94450 20300 -76500
rect 20000 -97700 20300 -94950
rect 20500 -95100 20800 -76300
rect 21000 -77000 21300 -76500
rect 21500 -77200 21800 -76250
rect 20500 -97150 20800 -95550
rect 21000 -95600 21300 -77300
rect 21500 -96100 21800 -77500
rect 21000 -96850 21300 -96100
rect 22000 -96350 22300 -75950
rect 22500 -76500 22800 -75850
rect 25000 -75900 25300 -74600
rect 25500 -75800 25800 -74250
rect 26000 -75800 26300 -73950
rect 22500 -86250 22800 -77050
rect 23000 -84050 23300 -76550
rect 23500 -82100 23800 -75950
rect 24000 -79550 24300 -75950
rect 24500 -78500 24800 -76100
rect 25000 -77250 25300 -76200
rect 24000 -80350 24300 -80050
rect 23000 -84700 23300 -84350
rect 23000 -86550 23300 -85300
rect 22500 -96150 22800 -86550
rect 23500 -86800 23800 -82850
rect 23000 -95900 23300 -86900
rect 24000 -87050 24300 -80700
rect 23500 -95600 23800 -87100
rect 24500 -87250 24800 -79300
rect 24000 -95300 24300 -87350
rect 25000 -87500 25300 -78350
rect 24500 -94950 24800 -87600
rect 25500 -87700 25800 -77600
rect 25000 -93650 25300 -87850
rect 26000 -87900 26300 -76500
rect 25500 -93250 25800 -88050
rect 26500 -88100 26800 -73700
rect 26000 -92850 26300 -88200
rect 27000 -88250 27300 -73500
rect 27500 -88400 27800 -73250
rect 26500 -92400 26800 -88400
rect 28000 -88550 28300 -71900
rect 27000 -92150 27300 -88600
rect 28500 -88700 28800 -71900
rect 29000 -88700 29300 -71800
rect 29500 -88600 29800 -71800
rect 30000 -88450 30300 -71900
rect 30500 -88400 30800 -71800
rect 31000 -88250 31300 -71850
rect 31500 -88150 31800 -71900
rect 32000 -88050 32300 -72000
rect 32500 -87900 32800 -72150
rect 33000 -87700 33300 -72100
rect 33500 -87450 33800 -72050
rect 34000 -87500 34300 -71800
rect 34500 -87550 34800 -71400
rect 35000 -87700 35300 -71000
rect 35500 -87800 35800 -70550
rect 36000 -87800 36300 -69900
rect 36500 -87700 36800 -68900
rect 37000 -87500 37300 -68650
rect 37500 -87550 37800 -67800
rect 38000 -87500 38300 -67700
rect 38500 -87300 38800 -67600
rect 39000 -87150 39300 -66950
rect 39500 -86950 39800 -67000
rect 40000 -86800 40300 -66600
rect 40500 -86550 40800 -66250
rect 41000 -86350 41300 -65900
rect 41500 -86100 41800 -65700
rect 42000 -85850 42300 -65550
rect 42500 -85600 42800 -65500
rect 43000 -85350 43300 -65500
rect 46000 -65650 46300 -62800
rect 46500 -63300 46800 -62350
rect 43500 -69950 43800 -65650
rect 44000 -69900 44300 -65700
rect 44500 -69850 44800 -65900
rect 46500 -65950 46800 -63700
rect 47000 -64500 47300 -62050
rect 45000 -69800 45300 -66000
rect 47000 -66200 47300 -65350
rect 47500 -65700 47800 -61800
rect 45500 -69400 45800 -66400
rect 46000 -66550 46300 -66250
rect 46000 -67150 46300 -66850
rect 46000 -69750 46300 -67450
rect 46500 -69050 46800 -66500
rect 48000 -66900 48300 -61500
rect 47000 -68800 47300 -67250
rect 47500 -67500 47800 -67050
rect 48000 -67600 48300 -67250
rect 46500 -70450 46800 -70150
rect 47000 -70400 47300 -69800
rect 43500 -85000 43800 -70750
rect 44000 -77650 44300 -70500
rect 44500 -77350 44800 -70450
rect 45000 -77150 45300 -70450
rect 45500 -76900 45800 -70450
rect 46000 -76550 46300 -70500
rect 47500 -70550 47800 -68000
rect 48000 -68200 48300 -67900
rect 48500 -68200 48800 -61200
rect 49000 -63100 49300 -60950
rect 49500 -62850 49800 -60650
rect 50000 -62600 50300 -60350
rect 50500 -62350 50800 -60050
rect 51000 -62050 51300 -59750
rect 51500 -62050 51800 -59500
rect 50000 -63400 50300 -62900
rect 50500 -63150 50800 -62650
rect 51000 -62950 51300 -62650
rect 52000 -62900 52300 -59200
rect 48000 -69500 48300 -68900
rect 48000 -70700 48300 -70150
rect 46500 -76250 46800 -70750
rect 47000 -75550 47300 -70700
rect 47500 -74550 47800 -70900
rect 48500 -70950 48800 -68900
rect 49000 -69400 49300 -63900
rect 50000 -64550 50300 -64250
rect 49500 -69600 49800 -64600
rect 50000 -65150 50300 -64850
rect 50500 -65050 50800 -63450
rect 51000 -65850 51300 -63350
rect 51500 -64950 51800 -63300
rect 52000 -64800 52300 -64000
rect 52500 -64150 52800 -59000
rect 53500 -59550 53800 -57750
rect 51500 -65550 51800 -65250
rect 50000 -69350 50300 -66150
rect 50500 -69100 50800 -66550
rect 51000 -68800 51300 -66400
rect 51500 -68550 51800 -66150
rect 52000 -68300 52300 -65900
rect 52500 -68050 52800 -65700
rect 53000 -67800 53300 -59700
rect 54000 -60800 54300 -58000
rect 53500 -67550 53800 -60950
rect 54500 -62000 54800 -58450
rect 54000 -67300 54300 -62150
rect 55000 -62900 55300 -58700
rect 55500 -61400 55800 -58700
rect 56000 -60450 56300 -58500
rect 56500 -59850 56800 -58300
rect 57000 -59500 57300 -58100
rect 57500 -59300 57800 -58000
rect 58000 -59250 58300 -57950
rect 58500 -59250 58800 -58000
rect 59000 -59400 59300 -58050
rect 55500 -62050 55800 -61750
rect 54500 -67050 54800 -63300
rect 55500 -64400 55800 -62600
rect 55000 -66800 55300 -64600
rect 56000 -65700 56300 -61000
rect 55500 -66500 55800 -65950
rect 48000 -73400 48300 -71050
rect 48500 -71900 48800 -71350
rect 48000 -75400 48300 -74000
rect 47000 -76700 47300 -76150
rect 46500 -77700 46800 -76850
rect 47000 -77700 47300 -77400
rect 44000 -84650 44300 -77950
rect 44500 -84200 44800 -77800
rect 47500 -77900 47800 -75650
rect 45000 -83800 45300 -77900
rect 45500 -83300 45800 -77900
rect 46000 -82900 46300 -77900
rect 46500 -82500 46800 -78150
rect 48000 -78300 48300 -77350
rect 47000 -82150 47300 -78350
rect 48500 -78550 48800 -72550
rect 47500 -81600 47800 -78550
rect 48000 -81000 48300 -78700
rect 49000 -78900 49300 -70000
rect 48500 -80500 48800 -78900
rect 49500 -79550 49800 -70100
rect 49000 -80000 49300 -79600
rect 47000 -82850 47300 -82550
rect 46000 -84450 46300 -83300
rect 47000 -83850 47300 -83200
rect 47500 -84050 47800 -82050
rect 48000 -83800 48300 -81450
rect 48500 -83450 48800 -80950
rect 49000 -83150 49300 -80450
rect 49500 -82750 49800 -79950
rect 50000 -82400 50300 -70000
rect 50500 -82000 50800 -69700
rect 51000 -81450 51300 -69400
rect 51500 -80700 51800 -69150
rect 52000 -69200 52300 -68900
rect 52500 -69300 52800 -68650
rect 52000 -80050 52300 -69500
rect 53000 -69700 53300 -68450
rect 52500 -79100 52800 -69850
rect 53500 -70000 53800 -68200
rect 53000 -77900 53300 -70200
rect 54000 -70300 54300 -67950
rect 53500 -76700 53800 -70650
rect 54500 -71100 54800 -67700
rect 55000 -70850 55300 -67400
rect 55500 -69850 55800 -67200
rect 56000 -67550 56300 -66900
rect 56000 -69850 56300 -68150
rect 56500 -68300 56800 -60350
rect 57000 -68400 57300 -59900
rect 57500 -64750 57800 -59600
rect 58000 -64200 58300 -59550
rect 58500 -64150 58800 -59550
rect 59500 -59750 59800 -58200
rect 59000 -64350 59300 -59800
rect 60000 -60200 60300 -58450
rect 54000 -75200 54300 -71150
rect 55000 -71450 55300 -71150
rect 55000 -76100 55300 -72700
rect 49500 -84750 49800 -83850
rect 50000 -84600 50300 -83350
rect 50500 -83500 50800 -83200
rect 27500 -92300 27800 -88750
rect 28000 -91700 28300 -88850
rect 28500 -91150 28800 -89000
rect 29000 -90750 29300 -89000
rect 27000 -92750 27300 -92450
rect 25000 -94700 25300 -93950
rect 25500 -94350 25800 -93650
rect 26000 -93900 26300 -93250
rect 26500 -93450 26800 -92900
rect 27500 -93300 27800 -92850
rect 28000 -93800 28300 -92350
rect 28500 -93950 28800 -91800
rect 29000 -92850 29300 -91050
rect 29500 -92300 29800 -88900
rect 30000 -91900 30300 -88800
rect 30500 -91500 30800 -88700
rect 31000 -91100 31300 -88600
rect 31500 -90700 31800 -88500
rect 32000 -90300 32300 -88400
rect 32500 -89900 32800 -88200
rect 33000 -89500 33300 -88100
rect 33500 -89100 33800 -87900
rect 34000 -88550 34300 -87850
rect 29500 -94400 29800 -92700
rect 30000 -94100 30300 -92300
rect 30500 -93800 30800 -91900
rect 31000 -93400 31300 -91500
rect 31500 -93050 31800 -91100
rect 32000 -92650 32300 -90700
rect 32500 -92300 32800 -90350
rect 33000 -92000 33300 -89950
rect 33500 -91650 33800 -89500
rect 34000 -91250 34300 -89050
rect 34500 -89200 34800 -88500
rect 35500 -89700 35800 -88850
rect 37000 -89550 37300 -89150
rect 37500 -89400 37800 -88750
rect 38500 -89050 38800 -88150
rect 39000 -88950 39300 -88000
rect 39500 -88900 39800 -87750
rect 40000 -88700 40300 -87600
rect 40500 -88700 40800 -87450
rect 41000 -88700 41300 -87000
rect 34500 -90850 34800 -89900
rect 35000 -91950 35300 -91450
rect 35500 -91700 35800 -91200
rect 36000 -91450 36300 -90700
rect 36500 -91200 36800 -90150
rect 37000 -91000 37300 -89950
rect 37500 -90800 37800 -89700
rect 38000 -90600 38300 -89500
rect 38500 -90450 38800 -89350
rect 39000 -89550 39300 -89250
rect 39500 -89550 39800 -89250
rect 39000 -90250 39300 -89850
rect 39500 -90150 39800 -89850
rect 40000 -89950 40300 -89000
rect 40500 -89750 40800 -89000
rect 41000 -89550 41300 -89000
rect 41500 -89250 41800 -86700
rect 42000 -89100 42300 -86500
rect 42500 -88850 42800 -86250
rect 43000 -88700 43300 -85950
rect 43500 -88600 43800 -85550
rect 44000 -88450 44300 -85750
rect 44500 -86150 44800 -84900
rect 44500 -87050 44800 -86750
rect 45000 -87050 45300 -84800
rect 44500 -88350 44800 -87350
rect 45500 -88150 45800 -85100
rect 49000 -85200 49300 -84900
rect 46000 -88200 46300 -85500
rect 46500 -88100 46800 -85900
rect 48500 -86000 48800 -85650
rect 47000 -88100 47300 -86400
rect 47500 -88000 47800 -86200
rect 48000 -87850 48300 -86450
rect 48500 -86900 48800 -86600
rect 48500 -88000 48800 -87700
rect 49000 -87900 49300 -86200
rect 49500 -87600 49800 -85600
rect 50000 -87700 50300 -85000
rect 50500 -86550 50800 -84550
rect 51500 -85250 51800 -81700
rect 52000 -81800 52300 -80950
rect 52500 -81000 52800 -80150
rect 53000 -80350 53300 -79300
rect 53500 -79750 53800 -78100
rect 54000 -79150 54300 -76500
rect 54500 -78650 54800 -76100
rect 55000 -78200 55300 -76800
rect 55500 -77000 55800 -70200
rect 55500 -77800 55800 -77500
rect 56000 -77650 56300 -70200
rect 52000 -82400 52300 -82100
rect 52500 -82200 52800 -81500
rect 53000 -81900 53300 -80800
rect 53500 -81800 53800 -80200
rect 52000 -83950 52300 -82850
rect 52500 -83050 52800 -82550
rect 51000 -86100 51300 -85800
rect 51000 -87500 51300 -87200
rect 51500 -87850 51800 -85550
rect 52000 -88200 52300 -84500
rect 52500 -88250 52800 -83700
rect 53000 -88100 53300 -82800
rect 53500 -87900 53800 -82200
rect 54000 -87700 54300 -79700
rect 54500 -82700 54800 -79150
rect 55000 -81850 55300 -78650
rect 55500 -81200 55800 -78200
rect 56000 -80700 56300 -77950
rect 55000 -82750 55300 -82450
rect 55500 -82700 55800 -81700
rect 56000 -82600 56300 -81050
rect 54500 -87600 54800 -83200
rect 55000 -87500 55300 -83100
rect 55500 -87400 55800 -83000
rect 56000 -83400 56300 -83100
rect 56000 -84500 56300 -83700
rect 56000 -85150 56300 -84850
rect 56000 -87300 56300 -85450
rect 56500 -86250 56800 -68650
rect 57000 -73050 57300 -69100
rect 57500 -70100 57800 -65300
rect 58000 -70750 58300 -64600
rect 57500 -71500 57800 -70750
rect 58000 -71400 58300 -71100
rect 57000 -75800 57300 -73500
rect 57000 -76400 57300 -76100
rect 57000 -86600 57300 -76700
rect 57500 -77800 57800 -71950
rect 57500 -86600 57800 -78300
rect 58000 -78850 58300 -71700
rect 58000 -86550 58300 -79450
rect 58500 -79700 58800 -64450
rect 59000 -72250 59300 -64900
rect 59500 -65000 59800 -60250
rect 59500 -72650 59800 -65550
rect 60000 -65700 60300 -60700
rect 60500 -60750 60800 -58800
rect 60000 -71700 60300 -66250
rect 60500 -66450 60800 -61200
rect 61000 -61250 61300 -59200
rect 60500 -71750 60800 -67000
rect 61000 -67150 61300 -61700
rect 61500 -61800 61800 -59650
rect 61000 -72100 61300 -67700
rect 61500 -67950 61800 -62250
rect 62000 -62450 62300 -60200
rect 61500 -71700 61800 -68500
rect 62000 -68850 62300 -63100
rect 62500 -63400 62800 -60650
rect 63000 -63500 63300 -61000
rect 63500 -62850 63800 -61250
rect 64000 -62600 64300 -61350
rect 64500 -62600 64800 -61450
rect 62000 -70900 62300 -69750
rect 62500 -70350 62800 -64300
rect 63000 -70750 63300 -64400
rect 61500 -72300 61800 -72000
rect 62000 -72150 62300 -71450
rect 62500 -71750 62800 -71450
rect 58500 -86400 58800 -80100
rect 59000 -80200 59300 -72650
rect 60000 -73000 60300 -72350
rect 59000 -86500 59300 -80550
rect 59500 -86550 59800 -73000
rect 60500 -73450 60800 -72650
rect 60000 -86500 60300 -73450
rect 61000 -73800 61300 -72700
rect 61500 -73450 61800 -73150
rect 60500 -82200 60800 -73850
rect 61000 -82200 61300 -74250
rect 61500 -74300 61800 -73750
rect 62000 -74750 62300 -72550
rect 61500 -82200 61800 -74750
rect 62000 -81900 62300 -75200
rect 62500 -75250 62800 -72050
rect 63000 -75750 63300 -71150
rect 63500 -71350 63800 -63250
rect 63500 -76450 63800 -71950
rect 64000 -72350 64300 -62900
rect 62500 -81200 62800 -76750
rect 63000 -80150 63300 -76800
rect 63500 -78450 63800 -77000
rect 64000 -78350 64300 -73050
rect 64500 -73650 64800 -63100
rect 65000 -63300 65300 -61700
rect 64500 -77550 64800 -74050
rect 65000 -75300 65300 -63950
rect 65500 -64500 65800 -61950
rect 65000 -76600 65300 -76200
rect 65000 -77200 65300 -76900
rect 65500 -77450 65800 -65000
rect 66000 -65900 66300 -62400
rect 64500 -78600 64800 -78000
rect 63000 -80750 63300 -80450
rect 60500 -82900 60800 -82600
rect 61000 -82800 61300 -82500
rect 60500 -86400 60800 -83200
rect 61000 -86300 61300 -83200
rect 61500 -86200 61800 -82500
rect 62000 -86100 62300 -82200
rect 62500 -86100 62800 -81700
rect 63000 -86100 63300 -81050
rect 63500 -86050 63800 -78750
rect 64000 -82000 64300 -78650
rect 64000 -86000 64300 -82600
rect 64500 -82650 64800 -79500
rect 65000 -82900 65300 -78500
rect 65500 -82900 65800 -77900
rect 66000 -82650 66300 -66600
rect 66500 -67700 66800 -63050
rect 66500 -71400 66800 -68700
rect 67000 -70900 67300 -64050
rect 66500 -82200 66800 -71700
rect 67500 -71800 67800 -65400
rect 68000 -71450 68300 -67300
rect 68500 -71200 68800 -69100
rect 69000 -71000 69300 -69600
rect 69500 -71000 69800 -69850
rect 67000 -77350 67300 -72950
rect 67000 -81650 67300 -77700
rect 67500 -77750 67800 -72800
rect 67500 -79450 67800 -78550
rect 67500 -80200 67800 -79900
rect 64500 -86000 64800 -83000
rect 65000 -86000 65300 -83200
rect 65500 -85700 65800 -83200
rect 66000 -85150 66300 -83000
rect 66500 -85050 66800 -82650
rect 67000 -84600 67300 -82000
rect 67500 -83850 67800 -80700
rect 68000 -83250 68300 -71800
rect 68500 -82100 68800 -71500
rect 69000 -82550 69300 -71350
rect 69500 -81250 69800 -71400
rect 70000 -71850 70300 -70100
rect 70000 -72750 70300 -72350
rect 70000 -77700 70300 -73550
rect 70000 -79150 70300 -78500
rect 70000 -79750 70300 -79450
rect 67000 -85950 67300 -85150
rect 67500 -86050 67800 -84700
rect 68000 -86100 68300 -84800
rect 68500 -86100 68800 -84150
rect 69000 -86000 69300 -83250
rect 69500 -85850 69800 -81550
rect 70000 -85600 70300 -80050
rect 70500 -85250 70800 -70400
rect 71000 -84850 71300 -71000
rect 71500 -80150 71800 -72050
rect 71500 -84500 71800 -81750
rect 72000 -84050 72300 -81750
rect 72500 -83650 72800 -81500
rect 73000 -83200 73300 -81150
rect 73500 -82600 73800 -80850
rect 74000 -82250 74300 -80450
rect 74500 -82000 74800 -80100
rect 75000 -81600 75300 -79700
rect 75500 -81200 75800 -79350
rect 76000 -80850 76300 -78900
rect 76500 -80450 76800 -78500
rect 77000 -80050 77300 -78100
rect 77500 -79600 77800 -77700
rect 78000 -79250 78300 -77300
rect 78500 -78800 78800 -76900
rect 79000 -78400 79300 -76600
rect 79500 -78000 79800 -76400
rect 80000 -77550 80300 -76250
rect 80500 -77050 80800 -76250
rect 56500 -87200 56800 -86750
rect 31500 -95000 31800 -93450
rect 22500 -96800 22800 -96500
rect 23000 -96550 23300 -96250
rect 21000 -99800 21300 -97400
rect 21500 -99550 21800 -97000
rect 22000 -99300 22300 -97100
rect 32000 -97350 32300 -93100
rect 32000 -98200 32300 -97650
rect 47000 -99850 47300 -88600
rect 49500 -88700 49800 -88400
rect 47500 -99150 47800 -88850
rect 48000 -98400 48300 -88800
rect 48500 -97650 48800 -89350
rect 49000 -95050 49300 -89100
rect 49500 -94850 49800 -89750
rect 50500 -90100 50800 -89800
rect 50000 -94550 50300 -90100
rect 50500 -93800 50800 -91800
rect 51000 -91900 51300 -89500
rect 51000 -94600 51300 -92400
rect 49000 -97000 49300 -95350
rect 49500 -96350 49800 -95150
rect 48500 -99200 48800 -98200
rect 49000 -98550 49300 -97450
rect 50000 -98450 50300 -97750
rect 50500 -98300 50800 -96000
rect 51000 -98100 51300 -95600
rect 51500 -97900 51800 -89400
rect 52000 -97600 52300 -88850
rect 52500 -97350 52800 -88650
rect 53000 -97050 53300 -88450
rect 53500 -96800 53800 -88250
rect 54000 -96450 54300 -88100
rect 54500 -96100 54800 -87900
rect 55000 -95750 55300 -87800
rect 55500 -95300 55800 -87700
rect 56000 -94850 56300 -87600
rect 56500 -94400 56800 -87500
rect 57000 -93950 57300 -87400
rect 57500 -93550 57800 -87400
rect 58000 -93150 58300 -87300
rect 58500 -92750 58800 -87150
rect 59000 -92400 59300 -87100
rect 59500 -91950 59800 -86950
rect 60000 -91550 60300 -86850
rect 60500 -91200 60800 -86700
rect 61000 -90800 61300 -86600
rect 61500 -90400 61800 -86600
rect 62000 -90050 62300 -86500
rect 62500 -89600 62800 -86450
rect 63000 -89250 63300 -86400
rect 63500 -88850 63800 -86350
rect 64000 -88300 64300 -86300
rect 64500 -87800 64800 -86300
rect 65000 -87450 65300 -86300
rect 65500 -87100 65800 -86300
rect 66000 -86700 66300 -86300
rect 68000 -87200 68300 -86650
rect 68500 -86900 68800 -86600
rect 72000 -97150 72300 -84700
rect 72500 -97900 72800 -84350
rect 73000 -96950 73300 -83900
rect 73500 -96900 73800 -83350
rect 74000 -96900 74300 -82850
rect 74500 -96900 74800 -82400
rect 75000 -96900 75300 -82200
rect 75500 -96900 75800 -81850
rect 76000 -96950 76300 -81200
rect 76500 -91800 76800 -80850
rect 77000 -91650 77300 -80450
rect 76500 -97150 76800 -92450
rect 77500 -94700 77800 -80100
rect 77000 -96300 77300 -94800
rect 77000 -97000 77300 -96600
rect 77500 -97100 77800 -95000
rect 73000 -98400 73300 -97250
rect 73500 -98700 73800 -97200
rect 74000 -99050 74300 -97200
rect 74500 -99400 74800 -97200
rect 75000 -99600 75300 -97200
rect 75500 -99800 75800 -97200
rect 78000 -97450 78300 -79650
rect 78500 -98000 78800 -79200
rect 79000 -94250 79300 -78800
rect 79500 -91400 79800 -78400
rect 79000 -94850 79300 -94550
rect 79000 -95700 79300 -95300
rect 79000 -96500 79300 -96100
rect 79500 -97400 79800 -92850
rect 80000 -92900 80300 -77950
rect 81000 -79250 81300 -76350
rect 81000 -80400 81300 -79550
rect 81500 -80250 81800 -76600
rect 82000 -80350 82300 -77100
rect 82500 -80300 82800 -77750
rect 83000 -80250 83300 -78250
rect 83500 -80100 83800 -78450
rect 84000 -80050 84300 -78500
rect 84500 -80000 84800 -78500
rect 85000 -79950 85300 -78400
rect 85500 -79900 85800 -78400
rect 86000 -79900 86300 -78350
rect 86500 -79850 86800 -78300
rect 87000 -79750 87300 -78250
rect 87500 -79700 87800 -78200
rect 88000 -79650 88300 -78150
rect 88500 -79600 88800 -78100
rect 89000 -79600 89300 -78050
rect 89500 -79550 89800 -78000
rect 90000 -79550 90300 -78000
rect 90500 -79550 90800 -78000
rect 91000 -79550 91300 -78000
rect 91500 -79550 91800 -78000
rect 92000 -79550 92300 -77950
rect 92500 -79500 92800 -77900
rect 93000 -79500 93300 -77900
rect 93500 -79500 93800 -77900
rect 94000 -79500 94300 -77900
rect 94500 -79500 94800 -77900
rect 95000 -79500 95300 -77900
rect 95500 -79450 95800 -77850
rect 96000 -79400 96300 -77800
rect 96500 -79300 96800 -77700
rect 97000 -79200 97300 -77600
rect 97500 -79100 97800 -77550
rect 98500 -78850 98800 -77250
rect 99000 -78700 99300 -77100
rect 99500 -78600 99800 -76950
rect 81500 -81050 81800 -80700
rect 82000 -81050 82300 -80750
rect 80000 -93950 80300 -93450
rect 80000 -97300 80300 -94500
rect 78000 -98400 78300 -98100
rect 78500 -99300 78800 -98500
<< end >>
