magic
tech sky130B
magscale 1 2
timestamp 1663444684
<< locali >>
rect -30 12410 4250 12420
rect -30 12370 40 12410
rect 4180 12370 4250 12410
rect -30 12360 4250 12370
rect -30 12170 30 12190
rect -30 230 -20 12170
rect 20 230 30 12170
rect -30 210 30 230
rect 4190 12170 4250 12190
rect 4190 230 4200 12170
rect 4240 230 4250 12170
rect 4190 210 4250 230
rect -30 20 4250 30
rect -30 -20 40 20
rect 4180 -20 4250 20
rect -30 -30 4250 -20
<< viali >>
rect 40 12370 4180 12410
rect -20 230 20 12170
rect 4200 230 4240 12170
rect 40 -20 4180 20
<< metal1 >>
rect -30 12410 4250 12420
rect -30 12370 40 12410
rect 4180 12370 4250 12410
rect -30 12360 4250 12370
rect -30 12170 30 12360
rect 150 12240 170 12310
rect 4050 12240 4070 12310
rect 164 12222 4058 12240
rect -30 30 30 230
rect 101 12173 167 12193
rect 101 193 167 213
rect 259 12173 325 12193
rect 259 193 325 213
rect 417 12173 483 12193
rect 417 193 483 213
rect 575 12173 641 12193
rect 575 193 641 213
rect 733 12173 799 12193
rect 733 193 799 213
rect 891 12173 957 12193
rect 891 193 957 213
rect 1049 12173 1115 12193
rect 1049 193 1115 213
rect 1207 12173 1273 12193
rect 1207 193 1273 213
rect 1365 12173 1431 12193
rect 1365 193 1431 213
rect 1523 12173 1589 12193
rect 1523 193 1589 213
rect 1681 12173 1747 12193
rect 1681 193 1747 213
rect 1839 12173 1905 12193
rect 1839 193 1905 213
rect 1997 12173 2063 12193
rect 1997 193 2063 213
rect 2155 12173 2221 12193
rect 2155 193 2221 213
rect 2313 12173 2379 12193
rect 2313 193 2379 213
rect 2471 12173 2537 12193
rect 2471 193 2537 213
rect 2629 12173 2695 12193
rect 2629 193 2695 213
rect 2787 12173 2853 12193
rect 2787 193 2853 213
rect 2945 12173 3011 12193
rect 2945 193 3011 213
rect 3103 12173 3169 12193
rect 3103 193 3169 213
rect 3261 12173 3327 12193
rect 3261 193 3327 213
rect 3419 12173 3485 12193
rect 3419 193 3485 213
rect 3577 12173 3643 12193
rect 3577 193 3643 213
rect 3735 12173 3801 12193
rect 3735 193 3801 213
rect 3893 12173 3959 12193
rect 3893 193 3959 213
rect 4051 12173 4117 12193
rect 4051 193 4117 213
rect 4190 12170 4250 12360
rect 162 150 4056 162
rect 150 80 170 150
rect 4050 80 4070 150
rect 4190 30 4250 230
rect -30 20 4250 30
rect -30 -20 40 20
rect 4180 -20 4250 20
rect -30 -30 4250 -20
<< via1 >>
rect 170 12240 4050 12310
rect -30 230 -20 12170
rect -20 230 20 12170
rect 20 230 30 12170
rect 101 213 167 12173
rect 259 213 325 12173
rect 417 213 483 12173
rect 575 213 641 12173
rect 733 213 799 12173
rect 891 213 957 12173
rect 1049 213 1115 12173
rect 1207 213 1273 12173
rect 1365 213 1431 12173
rect 1523 213 1589 12173
rect 1681 213 1747 12173
rect 1839 213 1905 12173
rect 1997 213 2063 12173
rect 2155 213 2221 12173
rect 2313 213 2379 12173
rect 2471 213 2537 12173
rect 2629 213 2695 12173
rect 2787 213 2853 12173
rect 2945 213 3011 12173
rect 3103 213 3169 12173
rect 3261 213 3327 12173
rect 3419 213 3485 12173
rect 3577 213 3643 12173
rect 3735 213 3801 12173
rect 3893 213 3959 12173
rect 4051 213 4117 12173
rect 4190 230 4200 12170
rect 4200 230 4240 12170
rect 4240 230 4250 12170
rect 170 80 4050 150
<< metal2 >>
rect 10 12240 170 12310
rect 4050 12240 4070 12310
rect -30 12170 30 12190
rect -30 210 30 230
rect 101 12173 167 12193
rect 101 193 167 213
rect 259 12173 325 12193
rect 259 193 325 213
rect 417 12173 483 12193
rect 417 193 483 213
rect 575 12173 641 12193
rect 575 193 641 213
rect 733 12173 799 12193
rect 733 193 799 213
rect 891 12173 957 12193
rect 891 193 957 213
rect 1049 12173 1115 12193
rect 1049 193 1115 213
rect 1207 12173 1273 12193
rect 1207 193 1273 213
rect 1365 12173 1431 12193
rect 1365 193 1431 213
rect 1523 12173 1589 12193
rect 1523 193 1589 213
rect 1681 12173 1747 12193
rect 1681 193 1747 213
rect 1839 12173 1905 12193
rect 1839 193 1905 213
rect 1997 12173 2063 12193
rect 1997 193 2063 213
rect 2155 12173 2221 12193
rect 2155 193 2221 213
rect 2313 12173 2379 12193
rect 2313 193 2379 213
rect 2471 12173 2537 12193
rect 2471 193 2537 213
rect 2629 12173 2695 12193
rect 2629 193 2695 213
rect 2787 12173 2853 12193
rect 2787 193 2853 213
rect 2945 12173 3011 12193
rect 2945 193 3011 213
rect 3103 12173 3169 12193
rect 3103 193 3169 213
rect 3261 12173 3327 12193
rect 3261 193 3327 213
rect 3419 12173 3485 12193
rect 3419 193 3485 213
rect 3577 12173 3643 12193
rect 3577 193 3643 213
rect 3735 12173 3801 12193
rect 3735 193 3801 213
rect 3893 12173 3959 12193
rect 3893 193 3959 213
rect 4051 12173 4117 12193
rect 4051 193 4117 213
rect 4190 12170 4250 12190
rect 4190 210 4250 230
rect 10 80 170 150
rect 4050 80 4070 150
<< via2 >>
rect 101 6420 167 12173
rect 259 213 325 5966
rect 417 6420 483 12173
rect 575 213 641 5966
rect 733 6420 799 12173
rect 891 213 957 5966
rect 1049 6420 1115 12173
rect 1207 213 1273 5966
rect 1365 6420 1431 12173
rect 1523 213 1589 5966
rect 1681 6420 1747 12173
rect 1839 213 1905 5966
rect 1997 6420 2063 12173
rect 2155 213 2221 5966
rect 2313 6420 2379 12173
rect 2471 213 2537 5966
rect 2629 6420 2695 12173
rect 2787 213 2853 5966
rect 2945 6420 3011 12173
rect 3103 213 3169 5966
rect 3261 6420 3327 12173
rect 3419 213 3485 5966
rect 3577 6420 3643 12173
rect 3735 213 3801 5966
rect 3893 6420 3959 12173
rect 4051 213 4117 5966
<< metal3 >>
rect 0 12173 4200 12200
rect 0 6420 101 12173
rect 167 6420 417 12173
rect 483 6420 733 12173
rect 799 6420 1049 12173
rect 1115 6420 1365 12173
rect 1431 6420 1681 12173
rect 1747 6420 1997 12173
rect 2063 6420 2313 12173
rect 2379 6420 2629 12173
rect 2695 6420 2945 12173
rect 3011 6420 3261 12173
rect 3327 6420 3577 12173
rect 3643 6420 3893 12173
rect 3959 6420 4200 12173
rect 0 6400 4200 6420
rect 0 5966 4200 6000
rect 0 213 259 5966
rect 325 213 575 5966
rect 641 213 891 5966
rect 957 213 1207 5966
rect 1273 213 1523 5966
rect 1589 213 1839 5966
rect 1905 213 2155 5966
rect 2221 213 2471 5966
rect 2537 213 2787 5966
rect 2853 213 3103 5966
rect 3169 213 3419 5966
rect 3485 213 3735 5966
rect 3801 213 4051 5966
rect 4117 213 4200 5966
rect 0 200 4200 213
use sky130_fd_pr__nfet_g5v0d10v5_NJL6SH  sky130_fd_pr__nfet_g5v0d10v5_NJL6SH_0
timestamp 1663433502
transform 1 0 2109 0 1 6193
box -2174 -6258 2174 6258
<< labels >>
rlabel metal2 50 12240 80 12310 1 G
rlabel metal1 -30 -30 20 30 1 SUB
rlabel metal3 40 6400 90 12200 1 SD1
rlabel metal3 40 200 90 6000 1 SD2
<< end >>
