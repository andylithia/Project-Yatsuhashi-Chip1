magic
tech sky130B
magscale 1 2
timestamp 1659923628
<< error_p >>
rect -401 407 -355 419
rect -293 407 -247 419
rect -185 407 -139 419
rect -77 407 -31 419
rect 31 407 77 419
rect 139 407 185 419
rect 247 407 293 419
rect 355 407 401 419
rect -401 367 -395 407
rect -293 367 -287 407
rect -185 367 -179 407
rect -77 367 -71 407
rect 31 367 37 407
rect 139 367 145 407
rect 247 367 253 407
rect 355 367 361 407
rect -401 355 -355 367
rect -293 355 -247 367
rect -185 355 -139 367
rect -77 355 -31 367
rect 31 355 77 367
rect 139 355 185 367
rect 247 355 293 367
rect 355 355 401 367
rect -401 -367 -355 -355
rect -293 -367 -247 -355
rect -185 -367 -139 -355
rect -77 -367 -31 -355
rect 31 -367 77 -355
rect 139 -367 185 -355
rect 247 -367 293 -355
rect 355 -367 401 -355
rect -401 -407 -395 -367
rect -293 -407 -287 -367
rect -185 -407 -179 -367
rect -77 -407 -71 -367
rect 31 -407 37 -367
rect 139 -407 145 -367
rect 247 -407 253 -367
rect 355 -407 361 -367
rect -401 -419 -355 -407
rect -293 -419 -247 -407
rect -185 -419 -139 -407
rect -77 -419 -31 -407
rect 31 -419 77 -407
rect 139 -419 185 -407
rect 247 -419 293 -407
rect 355 -419 401 -407
<< pwell >>
rect -577 -589 577 589
<< psubdiff >>
rect -541 519 -445 553
rect 445 519 541 553
rect -541 457 -507 519
rect 507 457 541 519
rect -541 -519 -507 -457
rect 507 -519 541 -457
rect -541 -553 -445 -519
rect 445 -553 541 -519
<< psubdiffcont >>
rect -445 519 445 553
rect -541 -457 -507 457
rect 507 -457 541 457
rect -445 -553 445 -519
<< poly >>
rect -411 407 -345 423
rect -411 373 -395 407
rect -361 373 -345 407
rect -411 350 -345 373
rect -411 -373 -345 -350
rect -411 -407 -395 -373
rect -361 -407 -345 -373
rect -411 -423 -345 -407
rect -303 407 -237 423
rect -303 373 -287 407
rect -253 373 -237 407
rect -303 350 -237 373
rect -303 -373 -237 -350
rect -303 -407 -287 -373
rect -253 -407 -237 -373
rect -303 -423 -237 -407
rect -195 407 -129 423
rect -195 373 -179 407
rect -145 373 -129 407
rect -195 350 -129 373
rect -195 -373 -129 -350
rect -195 -407 -179 -373
rect -145 -407 -129 -373
rect -195 -423 -129 -407
rect -87 407 -21 423
rect -87 373 -71 407
rect -37 373 -21 407
rect -87 350 -21 373
rect -87 -373 -21 -350
rect -87 -407 -71 -373
rect -37 -407 -21 -373
rect -87 -423 -21 -407
rect 21 407 87 423
rect 21 373 37 407
rect 71 373 87 407
rect 21 350 87 373
rect 21 -373 87 -350
rect 21 -407 37 -373
rect 71 -407 87 -373
rect 21 -423 87 -407
rect 129 407 195 423
rect 129 373 145 407
rect 179 373 195 407
rect 129 350 195 373
rect 129 -373 195 -350
rect 129 -407 145 -373
rect 179 -407 195 -373
rect 129 -423 195 -407
rect 237 407 303 423
rect 237 373 253 407
rect 287 373 303 407
rect 237 350 303 373
rect 237 -373 303 -350
rect 237 -407 253 -373
rect 287 -407 303 -373
rect 237 -423 303 -407
rect 345 407 411 423
rect 345 373 361 407
rect 395 373 411 407
rect 345 350 411 373
rect 345 -373 411 -350
rect 345 -407 361 -373
rect 395 -407 411 -373
rect 345 -423 411 -407
<< polycont >>
rect -395 373 -361 407
rect -395 -407 -361 -373
rect -287 373 -253 407
rect -287 -407 -253 -373
rect -179 373 -145 407
rect -179 -407 -145 -373
rect -71 373 -37 407
rect -71 -407 -37 -373
rect 37 373 71 407
rect 37 -407 71 -373
rect 145 373 179 407
rect 145 -407 179 -373
rect 253 373 287 407
rect 253 -407 287 -373
rect 361 373 395 407
rect 361 -407 395 -373
<< npolyres >>
rect -411 -350 -345 350
rect -303 -350 -237 350
rect -195 -350 -129 350
rect -87 -350 -21 350
rect 21 -350 87 350
rect 129 -350 195 350
rect 237 -350 303 350
rect 345 -350 411 350
<< locali >>
rect -541 519 -445 553
rect 445 519 541 553
rect -541 457 -507 519
rect 507 457 541 519
rect -411 373 -395 407
rect -361 373 -345 407
rect -303 373 -287 407
rect -253 373 -237 407
rect -195 373 -179 407
rect -145 373 -129 407
rect -87 373 -71 407
rect -37 373 -21 407
rect 21 373 37 407
rect 71 373 87 407
rect 129 373 145 407
rect 179 373 195 407
rect 237 373 253 407
rect 287 373 303 407
rect 345 373 361 407
rect 395 373 411 407
rect -411 -407 -395 -373
rect -361 -407 -345 -373
rect -303 -407 -287 -373
rect -253 -407 -237 -373
rect -195 -407 -179 -373
rect -145 -407 -129 -373
rect -87 -407 -71 -373
rect -37 -407 -21 -373
rect 21 -407 37 -373
rect 71 -407 87 -373
rect 129 -407 145 -373
rect 179 -407 195 -373
rect 237 -407 253 -373
rect 287 -407 303 -373
rect 345 -407 361 -373
rect 395 -407 411 -373
rect -541 -519 -507 -457
rect 507 -519 541 -457
rect -541 -553 -445 -519
rect 445 -553 541 -519
<< viali >>
rect -395 373 -361 407
rect -287 373 -253 407
rect -179 373 -145 407
rect -71 373 -37 407
rect 37 373 71 407
rect 145 373 179 407
rect 253 373 287 407
rect 361 373 395 407
rect -395 367 -361 373
rect -287 367 -253 373
rect -179 367 -145 373
rect -71 367 -37 373
rect 37 367 71 373
rect 145 367 179 373
rect 253 367 287 373
rect 361 367 395 373
rect -395 -373 -361 -367
rect -287 -373 -253 -367
rect -179 -373 -145 -367
rect -71 -373 -37 -367
rect 37 -373 71 -367
rect 145 -373 179 -367
rect 253 -373 287 -367
rect 361 -373 395 -367
rect -395 -407 -361 -373
rect -287 -407 -253 -373
rect -179 -407 -145 -373
rect -71 -407 -37 -373
rect 37 -407 71 -373
rect 145 -407 179 -373
rect 253 -407 287 -373
rect 361 -407 395 -373
<< metal1 >>
rect -401 407 -355 419
rect -401 367 -395 407
rect -361 367 -355 407
rect -401 355 -355 367
rect -293 407 -247 419
rect -293 367 -287 407
rect -253 367 -247 407
rect -293 355 -247 367
rect -185 407 -139 419
rect -185 367 -179 407
rect -145 367 -139 407
rect -185 355 -139 367
rect -77 407 -31 419
rect -77 367 -71 407
rect -37 367 -31 407
rect -77 355 -31 367
rect 31 407 77 419
rect 31 367 37 407
rect 71 367 77 407
rect 31 355 77 367
rect 139 407 185 419
rect 139 367 145 407
rect 179 367 185 407
rect 139 355 185 367
rect 247 407 293 419
rect 247 367 253 407
rect 287 367 293 407
rect 247 355 293 367
rect 355 407 401 419
rect 355 367 361 407
rect 395 367 401 407
rect 355 355 401 367
rect -401 -367 -355 -355
rect -401 -407 -395 -367
rect -361 -407 -355 -367
rect -401 -419 -355 -407
rect -293 -367 -247 -355
rect -293 -407 -287 -367
rect -253 -407 -247 -367
rect -293 -419 -247 -407
rect -185 -367 -139 -355
rect -185 -407 -179 -367
rect -145 -407 -139 -367
rect -185 -419 -139 -407
rect -77 -367 -31 -355
rect -77 -407 -71 -367
rect -37 -407 -31 -367
rect -77 -419 -31 -407
rect 31 -367 77 -355
rect 31 -407 37 -367
rect 71 -407 77 -367
rect 31 -419 77 -407
rect 139 -367 185 -355
rect 139 -407 145 -367
rect 179 -407 185 -367
rect 139 -419 185 -407
rect 247 -367 293 -355
rect 247 -407 253 -367
rect 287 -407 293 -367
rect 247 -419 293 -407
rect 355 -367 401 -355
rect 355 -407 361 -367
rect 395 -407 401 -367
rect 355 -419 401 -407
<< properties >>
string FIXED_BBOX -524 -536 524 536
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 3.5 m 1 nx 8 wmin 0.330 lmin 1.650 rho 48.2 val 511.212 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
