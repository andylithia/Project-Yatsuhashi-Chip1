magic
tech sky130B
magscale 1 2
timestamp 1663443203
<< locali >>
rect -30 12410 4250 12420
rect -30 12370 40 12410
rect 4180 12370 4250 12410
rect -30 12360 4250 12370
rect -30 12170 30 12190
rect -30 230 -20 12170
rect 20 230 30 12170
rect -30 210 30 230
rect 4190 12170 4250 12190
rect 4190 230 4200 12170
rect 4240 230 4250 12170
rect 4190 210 4250 230
rect -30 20 4250 30
rect -30 -20 40 20
rect 4180 -20 4250 20
rect -30 -30 4250 -20
<< viali >>
rect 40 12370 4180 12410
rect -20 230 20 12170
rect 4200 230 4240 12170
rect 40 -20 4180 20
<< metal1 >>
rect -30 12410 4250 12420
rect -30 12370 40 12410
rect 4180 12370 4250 12410
rect -30 12360 4250 12370
rect -30 12170 30 12360
rect 150 12240 170 12310
rect 4050 12240 4070 12310
rect 164 12222 4058 12240
rect -30 30 30 230
rect 101 12173 167 12193
rect 101 193 167 213
rect 259 12173 325 12193
rect 259 193 325 213
rect 417 12173 483 12193
rect 417 193 483 213
rect 575 12173 641 12193
rect 575 193 641 213
rect 733 12173 799 12193
rect 733 193 799 213
rect 891 12173 957 12193
rect 891 193 957 213
rect 1049 12173 1115 12193
rect 1049 193 1115 213
rect 1207 12173 1273 12193
rect 1207 193 1273 213
rect 1365 12173 1431 12193
rect 1365 193 1431 213
rect 1523 12173 1589 12193
rect 1523 193 1589 213
rect 1681 12173 1747 12193
rect 1681 193 1747 213
rect 1839 12173 1905 12193
rect 1839 193 1905 213
rect 1997 12173 2063 12193
rect 1997 193 2063 213
rect 2155 12173 2221 12193
rect 2155 193 2221 213
rect 2313 12173 2379 12193
rect 2313 193 2379 213
rect 2471 12173 2537 12193
rect 2471 193 2537 213
rect 2629 12173 2695 12193
rect 2629 193 2695 213
rect 2787 12173 2853 12193
rect 2787 193 2853 213
rect 2945 12173 3011 12193
rect 2945 193 3011 213
rect 3103 12173 3169 12193
rect 3103 193 3169 213
rect 3261 12173 3327 12193
rect 3261 193 3327 213
rect 3419 12173 3485 12193
rect 3419 193 3485 213
rect 3577 12173 3643 12193
rect 3577 193 3643 213
rect 3735 12173 3801 12193
rect 3735 193 3801 213
rect 3893 12173 3959 12193
rect 3893 193 3959 213
rect 4051 12173 4117 12193
rect 4051 193 4117 213
rect 4190 12170 4250 12360
rect 162 150 4056 162
rect 150 80 170 150
rect 4050 80 4070 150
rect 4190 30 4250 230
rect -30 20 4250 30
rect -30 -20 40 20
rect 4180 -20 4250 20
rect -30 -30 4250 -20
<< via1 >>
rect 170 12240 4050 12310
rect -30 230 -20 12170
rect -20 230 20 12170
rect 20 230 30 12170
rect 101 213 167 12173
rect 259 213 325 12173
rect 417 213 483 12173
rect 575 213 641 12173
rect 733 213 799 12173
rect 891 213 957 12173
rect 1049 213 1115 12173
rect 1207 213 1273 12173
rect 1365 213 1431 12173
rect 1523 213 1589 12173
rect 1681 213 1747 12173
rect 1839 213 1905 12173
rect 1997 213 2063 12173
rect 2155 213 2221 12173
rect 2313 213 2379 12173
rect 2471 213 2537 12173
rect 2629 213 2695 12173
rect 2787 213 2853 12173
rect 2945 213 3011 12173
rect 3103 213 3169 12173
rect 3261 213 3327 12173
rect 3419 213 3485 12173
rect 3577 213 3643 12173
rect 3735 213 3801 12173
rect 3893 213 3959 12173
rect 4051 213 4117 12173
rect 4190 230 4200 12170
rect 4200 230 4240 12170
rect 4240 230 4250 12170
rect 170 80 4050 150
<< metal2 >>
rect 10 12240 170 12310
rect 4050 12240 4070 12310
rect -30 12170 30 12190
rect -30 210 30 230
rect 101 12173 167 12193
rect 101 193 167 213
rect 259 12173 325 12193
rect 259 193 325 213
rect 417 12173 483 12193
rect 417 193 483 213
rect 575 12173 641 12193
rect 575 193 641 213
rect 733 12173 799 12193
rect 733 193 799 213
rect 891 12173 957 12193
rect 891 193 957 213
rect 1049 12173 1115 12193
rect 1049 193 1115 213
rect 1207 12173 1273 12193
rect 1207 193 1273 213
rect 1365 12173 1431 12193
rect 1365 193 1431 213
rect 1523 12173 1589 12193
rect 1523 193 1589 213
rect 1681 12173 1747 12193
rect 1681 193 1747 213
rect 1839 12173 1905 12193
rect 1839 193 1905 213
rect 1997 12173 2063 12193
rect 1997 193 2063 213
rect 2155 12173 2221 12193
rect 2155 193 2221 213
rect 2313 12173 2379 12193
rect 2313 193 2379 213
rect 2471 12173 2537 12193
rect 2471 193 2537 213
rect 2629 12173 2695 12193
rect 2629 193 2695 213
rect 2787 12173 2853 12193
rect 2787 193 2853 213
rect 2945 12173 3011 12193
rect 2945 193 3011 213
rect 3103 12173 3169 12193
rect 3103 193 3169 213
rect 3261 12173 3327 12193
rect 3261 193 3327 213
rect 3419 12173 3485 12193
rect 3419 193 3485 213
rect 3577 12173 3643 12193
rect 3577 193 3643 213
rect 3735 12173 3801 12193
rect 3735 193 3801 213
rect 3893 12173 3959 12193
rect 3893 193 3959 213
rect 4051 12173 4117 12193
rect 4051 193 4117 213
rect 4190 12170 4250 12190
rect 4190 210 4250 230
rect 10 80 170 150
rect 4050 80 4070 150
<< via2 >>
rect 101 233 167 12153
rect 259 233 325 12153
rect 417 233 483 12153
rect 575 233 641 12153
rect 733 233 799 12153
rect 891 233 957 12153
rect 1049 233 1115 12153
rect 1207 233 1273 12153
rect 1365 233 1431 12153
rect 1523 233 1589 12153
rect 1681 233 1747 12153
rect 1839 233 1905 12153
rect 1997 233 2063 12153
rect 2155 233 2221 12153
rect 2313 233 2379 12153
rect 2471 233 2537 12153
rect 2629 233 2695 12153
rect 2787 233 2853 12153
rect 2945 233 3011 12153
rect 3103 233 3169 12153
rect 3261 233 3327 12153
rect 3419 233 3485 12153
rect 3577 233 3643 12153
rect 3735 233 3801 12153
rect 3893 233 3959 12153
rect 4051 233 4117 12153
<< metal3 >>
rect 88 12340 4130 12430
rect 88 12153 180 12340
rect 88 233 101 12153
rect 167 233 180 12153
rect 88 213 180 233
rect 246 12153 338 12173
rect 246 233 259 12153
rect 325 233 338 12153
rect 246 46 338 233
rect 404 12153 496 12340
rect 404 233 417 12153
rect 483 233 496 12153
rect 404 213 496 233
rect 562 12153 654 12173
rect 562 233 575 12153
rect 641 233 654 12153
rect 562 46 654 233
rect 720 12153 812 12340
rect 720 233 733 12153
rect 799 233 812 12153
rect 720 213 812 233
rect 878 12153 970 12173
rect 878 233 891 12153
rect 957 233 970 12153
rect 878 46 970 233
rect 1036 12153 1128 12340
rect 1036 233 1049 12153
rect 1115 233 1128 12153
rect 1036 213 1128 233
rect 1194 12153 1286 12173
rect 1194 233 1207 12153
rect 1273 233 1286 12153
rect 1194 46 1286 233
rect 1352 12153 1444 12340
rect 1352 233 1365 12153
rect 1431 233 1444 12153
rect 1352 213 1444 233
rect 1510 12153 1602 12173
rect 1510 233 1523 12153
rect 1589 233 1602 12153
rect 1510 46 1602 233
rect 1668 12153 1760 12340
rect 1668 233 1681 12153
rect 1747 233 1760 12153
rect 1668 213 1760 233
rect 1826 12153 1918 12173
rect 1826 233 1839 12153
rect 1905 233 1918 12153
rect 1826 46 1918 233
rect 1984 12153 2076 12340
rect 1984 233 1997 12153
rect 2063 233 2076 12153
rect 1984 213 2076 233
rect 2142 12153 2234 12173
rect 2142 233 2155 12153
rect 2221 233 2234 12153
rect 2142 46 2234 233
rect 2300 12153 2392 12340
rect 2300 233 2313 12153
rect 2379 233 2392 12153
rect 2300 213 2392 233
rect 2458 12153 2550 12173
rect 2458 233 2471 12153
rect 2537 233 2550 12153
rect 2458 46 2550 233
rect 2616 12153 2708 12340
rect 2616 233 2629 12153
rect 2695 233 2708 12153
rect 2616 213 2708 233
rect 2774 12153 2866 12173
rect 2774 233 2787 12153
rect 2853 233 2866 12153
rect 2774 46 2866 233
rect 2932 12153 3024 12340
rect 2932 233 2945 12153
rect 3011 233 3024 12153
rect 2932 213 3024 233
rect 3090 12153 3182 12173
rect 3090 233 3103 12153
rect 3169 233 3182 12153
rect 3090 46 3182 233
rect 3248 12153 3340 12340
rect 3248 233 3261 12153
rect 3327 233 3340 12153
rect 3248 213 3340 233
rect 3406 12153 3498 12173
rect 3406 233 3419 12153
rect 3485 233 3498 12153
rect 3406 46 3498 233
rect 3564 12153 3656 12340
rect 3564 233 3577 12153
rect 3643 233 3656 12153
rect 3564 213 3656 233
rect 3722 12153 3814 12173
rect 3722 233 3735 12153
rect 3801 233 3814 12153
rect 3722 46 3814 233
rect 3880 12153 3972 12340
rect 3880 233 3893 12153
rect 3959 233 3972 12153
rect 3880 213 3972 233
rect 4038 12153 4130 12173
rect 4038 233 4051 12153
rect 4117 233 4130 12153
rect 4038 46 4130 233
rect 88 -44 4130 46
use sky130_fd_pr__nfet_g5v0d10v5_NJL6SH  sky130_fd_pr__nfet_g5v0d10v5_NJL6SH_0
timestamp 1663433502
transform 1 0 2109 0 1 6193
box -2174 -6258 2174 6258
<< labels >>
rlabel metal2 50 12240 80 12310 1 G
rlabel metal3 90 12420 170 12430 1 SD1
rlabel metal3 240 -40 320 -30 1 SD2
rlabel metal1 -30 -30 20 30 1 SUB
<< end >>
