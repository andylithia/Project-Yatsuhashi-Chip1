magic
tech sky130B
timestamp 1659290390
<< metal4 >>
rect 2400 4050 3100 6900
rect 2400 3350 2450 4050
rect 3050 3350 3100 4050
rect 2400 3300 3100 3350
rect -200 750 500 800
rect -200 50 -150 750
rect 450 50 500 750
rect -200 -200 500 50
<< via4 >>
rect 2450 3350 3050 4050
rect -150 50 450 750
<< metal5 >>
rect 0 6000 6500 6500
rect 0 950 500 6000
rect -50 900 500 950
rect -100 850 500 900
rect -150 800 500 850
rect -200 750 500 800
rect -200 50 -150 750
rect 450 50 500 750
rect -200 0 500 50
rect 800 5200 5700 5700
rect 800 500 1300 5200
rect 1600 4400 4900 4900
rect 1600 1300 2100 4400
rect 2400 4050 3100 4100
rect 2400 3350 2450 4050
rect 3050 3350 3100 4050
rect 2400 3300 3100 3350
rect 2400 3250 3050 3300
rect 2400 3200 3000 3250
rect 2400 3150 2950 3200
rect 2400 2100 2900 3150
rect 4400 2100 4900 4400
rect 2400 1600 4900 2100
rect 5200 1300 5700 5200
rect 1600 800 5700 1300
rect 6000 500 6500 6000
rect 800 0 6500 500
<< end >>
