magic
tech sky130B
magscale 1 2
timestamp 1660708745
<< metal5 >>
rect -23000 47000 17000 48000
rect -23000 16000 -22000 47000
rect 16000 33000 17000 47000
rect 16000 32000 71000 33000
rect 70000 5000 71000 32000
rect 66000 -9000 71000 5000
rect 64000 -11000 71000 -9000
rect 70000 -26000 71000 -11000
rect 26231 -27000 71000 -26000
use PA_complete_without_ind  PA_complete_without_ind_0
timestamp 1660708695
transform 1 0 1 0 1 0
box -23000 -42000 71000 48000
use octa_ind_3t_140_160_flat  octa_ind_3t_140_160_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1660524083
transform 0 -1 -23000 1 0 47900
box -39300 -34000 -5300 -6000
use octa_ind_thick_1p8n_flat  octa_ind_thick_1p8n_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1659752630
transform -1 0 20600 0 -1 -16800
box -51300 -45000 3200 5000
<< end >>
