magic
tech sky130A
timestamp 1660275339
<< metal1 >>
rect 50 -310 300 -300
rect 50 -345 125 -310
rect 225 -345 300 -310
rect 50 -350 300 -345
rect 50 -360 110 -350
rect 240 -360 300 -350
rect 50 -375 100 -360
rect 50 -475 60 -375
rect 95 -475 100 -375
rect 50 -490 100 -475
rect 250 -375 300 -360
rect 250 -475 255 -375
rect 290 -475 300 -375
rect 250 -490 300 -475
rect 50 -500 110 -490
rect 240 -500 300 -490
rect 50 -505 300 -500
rect 50 -540 125 -505
rect 225 -540 300 -505
rect 50 -550 300 -540
<< via1 >>
rect 125 -345 225 -310
rect 60 -475 95 -375
rect 255 -475 290 -375
rect 125 -540 225 -505
<< metal2 >>
rect 120 -310 230 -300
rect 120 -345 125 -310
rect 225 -345 230 -310
rect 120 -370 230 -345
rect 50 -375 300 -370
rect 50 -475 60 -375
rect 95 -475 255 -375
rect 290 -475 300 -375
rect 50 -480 300 -475
rect 120 -505 230 -480
rect 120 -540 125 -505
rect 225 -540 230 -505
rect 120 -550 230 -540
<< end >>
