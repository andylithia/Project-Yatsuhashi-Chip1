magic
tech sky130B
timestamp 1662577679
<< metal2 >>
rect -1100 4300 -800 4400
<< metal4 >>
rect 1700 -1700 2900 -600
rect 1400 -6700 2900 -1700
<< via4 >>
rect -350 -2300 550 -1200
<< metal5 >>
rect -4550 -2000 -3050 1500
rect -4650 -2100 -3050 -2000
rect -750 -1200 650 -1100
rect -4750 -2200 -3150 -2100
rect -4850 -2300 -3250 -2200
rect -750 -2300 -350 -1200
rect 550 -2300 650 -1200
rect -4850 -6200 -3350 -2300
rect -750 -2500 650 -2300
rect -1250 -2600 350 -2500
rect -1350 -2700 250 -2600
rect -1450 -2800 150 -2700
rect -1450 -6200 50 -2800
rect -4850 -7200 50 -6200
use lna_complete_2_wo_ind  lna_complete_2_wo_ind_0
timestamp 1662577679
transform 1 0 0 0 1 0
box -10500 -7100 5450 11950
use octa_2t_190_170_flat  octa_2t_190_170_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1661314321
transform 1 0 21550 0 1 11400
box -19700 -19500 -2700 -500
use octa_thick_3t_250_250_flat  octa_thick_3t_250_250_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1661315583
transform 0 -1 -13400 1 0 33650
box -23550 -22500 1450 2500
<< end >>
