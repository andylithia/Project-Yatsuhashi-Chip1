magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< poly >>
rect 2166 387 2196 648
rect 2790 511 2820 648
rect 3414 387 3444 648
rect 4038 511 4068 648
rect 4662 387 4692 648
rect 5286 511 5316 648
rect 5910 387 5940 648
rect 6534 511 6564 648
rect 7158 387 7188 648
rect 7782 511 7812 648
rect 8406 387 8436 648
rect 9030 511 9060 648
rect 9654 387 9684 648
rect 10278 511 10308 648
rect 10902 387 10932 648
rect 11526 511 11556 648
rect 12150 387 12180 648
rect 12774 511 12804 648
rect 13398 387 13428 648
rect 14022 511 14052 648
rect 14646 387 14676 648
rect 15270 511 15300 648
rect 15894 387 15924 648
rect 16518 511 16548 648
rect 17142 387 17172 648
rect 17766 511 17796 648
rect 18390 387 18420 648
rect 19014 511 19044 648
rect 19638 387 19668 648
rect 20262 511 20292 648
rect 20886 387 20916 648
rect 21510 511 21540 648
rect 22134 387 22164 648
rect 22758 511 22788 648
rect 23382 387 23412 648
rect 24006 511 24036 648
rect 24630 387 24660 648
rect 25254 511 25284 648
rect 25878 387 25908 648
rect 26502 511 26532 648
rect 27126 387 27156 648
rect 27750 511 27780 648
rect 28374 387 28404 648
rect 28998 511 29028 648
rect 29622 387 29652 648
rect 30246 511 30276 648
rect 30870 387 30900 648
rect 31494 511 31524 648
<< metal1 >>
rect 1949 1880 1977 1936
rect 2413 1880 2441 1936
rect 2545 1880 2573 1936
rect 3009 1880 3037 1936
rect 3197 1880 3225 1936
rect 3661 1880 3689 1936
rect 3793 1880 3821 1936
rect 4257 1880 4285 1936
rect 4445 1880 4473 1936
rect 4909 1880 4937 1936
rect 5041 1880 5069 1936
rect 5505 1880 5533 1936
rect 5693 1880 5721 1936
rect 6157 1880 6185 1936
rect 6289 1880 6317 1936
rect 6753 1880 6781 1936
rect 6941 1880 6969 1936
rect 7405 1880 7433 1936
rect 7537 1880 7565 1936
rect 8001 1880 8029 1936
rect 8189 1880 8217 1936
rect 8653 1880 8681 1936
rect 8785 1880 8813 1936
rect 9249 1880 9277 1936
rect 9437 1880 9465 1936
rect 9901 1880 9929 1936
rect 10033 1880 10061 1936
rect 10497 1880 10525 1936
rect 10685 1880 10713 1936
rect 11149 1880 11177 1936
rect 11281 1880 11309 1936
rect 11745 1880 11773 1936
rect 11933 1880 11961 1936
rect 12397 1880 12425 1936
rect 12529 1880 12557 1936
rect 12993 1880 13021 1936
rect 13181 1880 13209 1936
rect 13645 1880 13673 1936
rect 13777 1880 13805 1936
rect 14241 1880 14269 1936
rect 14429 1880 14457 1936
rect 14893 1880 14921 1936
rect 15025 1880 15053 1936
rect 15489 1880 15517 1936
rect 15677 1880 15705 1936
rect 16141 1880 16169 1936
rect 16273 1880 16301 1936
rect 16737 1880 16765 1936
rect 16925 1880 16953 1936
rect 17389 1880 17417 1936
rect 17521 1880 17549 1936
rect 17985 1880 18013 1936
rect 18173 1880 18201 1936
rect 18637 1880 18665 1936
rect 18769 1880 18797 1936
rect 19233 1880 19261 1936
rect 19421 1880 19449 1936
rect 19885 1880 19913 1936
rect 20017 1880 20045 1936
rect 20481 1880 20509 1936
rect 20669 1880 20697 1936
rect 21133 1880 21161 1936
rect 21265 1880 21293 1936
rect 21729 1880 21757 1936
rect 21917 1880 21945 1936
rect 22381 1880 22409 1936
rect 22513 1880 22541 1936
rect 22977 1880 23005 1936
rect 23165 1880 23193 1936
rect 23629 1880 23657 1936
rect 23761 1880 23789 1936
rect 24225 1880 24253 1936
rect 24413 1880 24441 1936
rect 24877 1880 24905 1936
rect 25009 1880 25037 1936
rect 25473 1880 25501 1936
rect 25661 1880 25689 1936
rect 26125 1880 26153 1936
rect 26257 1880 26285 1936
rect 26721 1880 26749 1936
rect 26909 1880 26937 1936
rect 27373 1880 27401 1936
rect 27505 1880 27533 1936
rect 27969 1880 27997 1936
rect 28157 1880 28185 1936
rect 28621 1880 28649 1936
rect 28753 1880 28781 1936
rect 29217 1880 29245 1936
rect 29405 1880 29433 1936
rect 29869 1880 29897 1936
rect 30001 1880 30029 1936
rect 30465 1880 30493 1936
rect 30653 1880 30681 1936
rect 31117 1880 31145 1936
rect 31249 1880 31277 1936
rect 31713 1880 31741 1936
rect 2461 1257 2525 1309
rect 3709 1257 3773 1309
rect 4957 1257 5021 1309
rect 6205 1257 6269 1309
rect 7453 1257 7517 1309
rect 8701 1257 8765 1309
rect 9949 1257 10013 1309
rect 11197 1257 11261 1309
rect 12445 1257 12509 1309
rect 13693 1257 13757 1309
rect 14941 1257 15005 1309
rect 16189 1257 16253 1309
rect 17437 1257 17501 1309
rect 18685 1257 18749 1309
rect 19933 1257 19997 1309
rect 21181 1257 21245 1309
rect 22429 1257 22493 1309
rect 23677 1257 23741 1309
rect 24925 1257 24989 1309
rect 26173 1257 26237 1309
rect 27421 1257 27485 1309
rect 28669 1257 28733 1309
rect 29917 1257 29981 1309
rect 31165 1257 31229 1309
rect 1949 274 1977 620
rect 2163 376 2227 428
rect 1931 222 1995 274
rect 2413 150 2441 620
rect 2545 150 2573 620
rect 2759 500 2823 552
rect 3009 274 3037 620
rect 3197 274 3225 620
rect 3411 376 3475 428
rect 2991 222 3055 274
rect 3179 222 3243 274
rect 3661 150 3689 620
rect 3793 150 3821 620
rect 4007 500 4071 552
rect 4257 274 4285 620
rect 4445 274 4473 620
rect 4659 376 4723 428
rect 4239 222 4303 274
rect 4427 222 4491 274
rect 4909 150 4937 620
rect 5041 150 5069 620
rect 5255 500 5319 552
rect 5505 274 5533 620
rect 5693 274 5721 620
rect 5907 376 5971 428
rect 5487 222 5551 274
rect 5675 222 5739 274
rect 6157 150 6185 620
rect 6289 150 6317 620
rect 6503 500 6567 552
rect 6753 274 6781 620
rect 6941 274 6969 620
rect 7155 376 7219 428
rect 6735 222 6799 274
rect 6923 222 6987 274
rect 7405 150 7433 620
rect 7537 150 7565 620
rect 7751 500 7815 552
rect 8001 274 8029 620
rect 8189 274 8217 620
rect 8403 376 8467 428
rect 7983 222 8047 274
rect 8171 222 8235 274
rect 8653 150 8681 620
rect 8785 150 8813 620
rect 8999 500 9063 552
rect 9249 274 9277 620
rect 9437 274 9465 620
rect 9651 376 9715 428
rect 9231 222 9295 274
rect 9419 222 9483 274
rect 9901 150 9929 620
rect 10033 150 10061 620
rect 10247 500 10311 552
rect 10497 274 10525 620
rect 10685 274 10713 620
rect 10899 376 10963 428
rect 10479 222 10543 274
rect 10667 222 10731 274
rect 11149 150 11177 620
rect 11281 150 11309 620
rect 11495 500 11559 552
rect 11745 274 11773 620
rect 11933 274 11961 620
rect 12147 376 12211 428
rect 11727 222 11791 274
rect 11915 222 11979 274
rect 12397 150 12425 620
rect 12529 150 12557 620
rect 12743 500 12807 552
rect 12993 274 13021 620
rect 13181 274 13209 620
rect 13395 376 13459 428
rect 12975 222 13039 274
rect 13163 222 13227 274
rect 13645 150 13673 620
rect 13777 150 13805 620
rect 13991 500 14055 552
rect 14241 274 14269 620
rect 14429 274 14457 620
rect 14643 376 14707 428
rect 14223 222 14287 274
rect 14411 222 14475 274
rect 14893 150 14921 620
rect 15025 150 15053 620
rect 15239 500 15303 552
rect 15489 274 15517 620
rect 15677 274 15705 620
rect 15891 376 15955 428
rect 15471 222 15535 274
rect 15659 222 15723 274
rect 16141 150 16169 620
rect 16273 150 16301 620
rect 16487 500 16551 552
rect 16737 274 16765 620
rect 16925 274 16953 620
rect 17139 376 17203 428
rect 16719 222 16783 274
rect 16907 222 16971 274
rect 17389 150 17417 620
rect 17521 150 17549 620
rect 17735 500 17799 552
rect 17985 274 18013 620
rect 18173 274 18201 620
rect 18387 376 18451 428
rect 17967 222 18031 274
rect 18155 222 18219 274
rect 18637 150 18665 620
rect 18769 150 18797 620
rect 18983 500 19047 552
rect 19233 274 19261 620
rect 19421 274 19449 620
rect 19635 376 19699 428
rect 19215 222 19279 274
rect 19403 222 19467 274
rect 19885 150 19913 620
rect 20017 150 20045 620
rect 20231 500 20295 552
rect 20481 274 20509 620
rect 20669 274 20697 620
rect 20883 376 20947 428
rect 20463 222 20527 274
rect 20651 222 20715 274
rect 21133 150 21161 620
rect 21265 150 21293 620
rect 21479 500 21543 552
rect 21729 274 21757 620
rect 21917 274 21945 620
rect 22131 376 22195 428
rect 21711 222 21775 274
rect 21899 222 21963 274
rect 22381 150 22409 620
rect 22513 150 22541 620
rect 22727 500 22791 552
rect 22977 274 23005 620
rect 23165 274 23193 620
rect 23379 376 23443 428
rect 22959 222 23023 274
rect 23147 222 23211 274
rect 23629 150 23657 620
rect 23761 150 23789 620
rect 23975 500 24039 552
rect 24225 274 24253 620
rect 24413 274 24441 620
rect 24627 376 24691 428
rect 24207 222 24271 274
rect 24395 222 24459 274
rect 24877 150 24905 620
rect 25009 150 25037 620
rect 25223 500 25287 552
rect 25473 274 25501 620
rect 25661 274 25689 620
rect 25875 376 25939 428
rect 25455 222 25519 274
rect 25643 222 25707 274
rect 26125 150 26153 620
rect 26257 150 26285 620
rect 26471 500 26535 552
rect 26721 274 26749 620
rect 26909 274 26937 620
rect 27123 376 27187 428
rect 26703 222 26767 274
rect 26891 222 26955 274
rect 27373 150 27401 620
rect 27505 150 27533 620
rect 27719 500 27783 552
rect 27969 274 27997 620
rect 28157 274 28185 620
rect 28371 376 28435 428
rect 27951 222 28015 274
rect 28139 222 28203 274
rect 28621 150 28649 620
rect 28753 150 28781 620
rect 28967 500 29031 552
rect 29217 274 29245 620
rect 29405 274 29433 620
rect 29619 376 29683 428
rect 29199 222 29263 274
rect 29387 222 29451 274
rect 29869 150 29897 620
rect 30001 150 30029 620
rect 30215 500 30279 552
rect 30465 274 30493 620
rect 30653 274 30681 620
rect 30867 376 30931 428
rect 30447 222 30511 274
rect 30635 222 30699 274
rect 31117 150 31145 620
rect 31249 150 31277 620
rect 31463 500 31527 552
rect 31713 274 31741 620
rect 31695 222 31759 274
rect 2395 98 2459 150
rect 2527 98 2591 150
rect 3643 98 3707 150
rect 3775 98 3839 150
rect 4891 98 4955 150
rect 5023 98 5087 150
rect 6139 98 6203 150
rect 6271 98 6335 150
rect 7387 98 7451 150
rect 7519 98 7583 150
rect 8635 98 8699 150
rect 8767 98 8831 150
rect 9883 98 9947 150
rect 10015 98 10079 150
rect 11131 98 11195 150
rect 11263 98 11327 150
rect 12379 98 12443 150
rect 12511 98 12575 150
rect 13627 98 13691 150
rect 13759 98 13823 150
rect 14875 98 14939 150
rect 15007 98 15071 150
rect 16123 98 16187 150
rect 16255 98 16319 150
rect 17371 98 17435 150
rect 17503 98 17567 150
rect 18619 98 18683 150
rect 18751 98 18815 150
rect 19867 98 19931 150
rect 19999 98 20063 150
rect 21115 98 21179 150
rect 21247 98 21311 150
rect 22363 98 22427 150
rect 22495 98 22559 150
rect 23611 98 23675 150
rect 23743 98 23807 150
rect 24859 98 24923 150
rect 24991 98 25055 150
rect 26107 98 26171 150
rect 26239 98 26303 150
rect 27355 98 27419 150
rect 27487 98 27551 150
rect 28603 98 28667 150
rect 28735 98 28799 150
rect 29851 98 29915 150
rect 29983 98 30047 150
rect 31099 98 31163 150
rect 31231 98 31295 150
<< metal2 >>
rect 2465 1259 2521 1307
rect 3713 1259 3769 1307
rect 4961 1259 5017 1307
rect 6209 1259 6265 1307
rect 7457 1259 7513 1307
rect 8705 1259 8761 1307
rect 9953 1259 10009 1307
rect 11201 1259 11257 1307
rect 12449 1259 12505 1307
rect 13697 1259 13753 1307
rect 14945 1259 15001 1307
rect 16193 1259 16249 1307
rect 17441 1259 17497 1307
rect 18689 1259 18745 1307
rect 19937 1259 19993 1307
rect 21185 1259 21241 1307
rect 22433 1259 22489 1307
rect 23681 1259 23737 1307
rect 24929 1259 24985 1307
rect 26177 1259 26233 1307
rect 27425 1259 27481 1307
rect 28673 1259 28729 1307
rect 29921 1259 29977 1307
rect 31169 1259 31225 1307
rect 2763 502 2819 550
rect 4011 502 4067 550
rect 5259 502 5315 550
rect 6507 502 6563 550
rect 7755 502 7811 550
rect 9003 502 9059 550
rect 10251 502 10307 550
rect 11499 502 11555 550
rect 12747 502 12803 550
rect 13995 502 14051 550
rect 15243 502 15299 550
rect 16491 502 16547 550
rect 17739 502 17795 550
rect 18987 502 19043 550
rect 20235 502 20291 550
rect 21483 502 21539 550
rect 22731 502 22787 550
rect 23979 502 24035 550
rect 25227 502 25283 550
rect 26475 502 26531 550
rect 27723 502 27779 550
rect 28971 502 29027 550
rect 30219 502 30275 550
rect 31467 502 31523 550
rect 2167 378 2223 426
rect 3415 378 3471 426
rect 4663 378 4719 426
rect 5911 378 5967 426
rect 7159 378 7215 426
rect 8407 378 8463 426
rect 9655 378 9711 426
rect 10903 378 10959 426
rect 12151 378 12207 426
rect 13399 378 13455 426
rect 14647 378 14703 426
rect 15895 378 15951 426
rect 17143 378 17199 426
rect 18391 378 18447 426
rect 19639 378 19695 426
rect 20887 378 20943 426
rect 22135 378 22191 426
rect 23383 378 23439 426
rect 24631 378 24687 426
rect 25879 378 25935 426
rect 27127 378 27183 426
rect 28375 378 28431 426
rect 29623 378 29679 426
rect 30871 378 30927 426
rect 1935 224 1991 272
rect 2995 224 3051 272
rect 3183 224 3239 272
rect 4243 224 4299 272
rect 4431 224 4487 272
rect 5491 224 5547 272
rect 5679 224 5735 272
rect 6739 224 6795 272
rect 6927 224 6983 272
rect 7987 224 8043 272
rect 8175 224 8231 272
rect 9235 224 9291 272
rect 9423 224 9479 272
rect 10483 224 10539 272
rect 10671 224 10727 272
rect 11731 224 11787 272
rect 11919 224 11975 272
rect 12979 224 13035 272
rect 13167 224 13223 272
rect 14227 224 14283 272
rect 14415 224 14471 272
rect 15475 224 15531 272
rect 15663 224 15719 272
rect 16723 224 16779 272
rect 16911 224 16967 272
rect 17971 224 18027 272
rect 18159 224 18215 272
rect 19219 224 19275 272
rect 19407 224 19463 272
rect 20467 224 20523 272
rect 20655 224 20711 272
rect 21715 224 21771 272
rect 21903 224 21959 272
rect 22963 224 23019 272
rect 23151 224 23207 272
rect 24211 224 24267 272
rect 24399 224 24455 272
rect 25459 224 25515 272
rect 25647 224 25703 272
rect 26707 224 26763 272
rect 26895 224 26951 272
rect 27955 224 28011 272
rect 28143 224 28199 272
rect 29203 224 29259 272
rect 29391 224 29447 272
rect 30451 224 30507 272
rect 30639 224 30695 272
rect 31699 224 31755 272
rect 2399 100 2455 148
rect 2531 100 2587 148
rect 3647 100 3703 148
rect 3779 100 3835 148
rect 4895 100 4951 148
rect 5027 100 5083 148
rect 6143 100 6199 148
rect 6275 100 6331 148
rect 7391 100 7447 148
rect 7523 100 7579 148
rect 8639 100 8695 148
rect 8771 100 8827 148
rect 9887 100 9943 148
rect 10019 100 10075 148
rect 11135 100 11191 148
rect 11267 100 11323 148
rect 12383 100 12439 148
rect 12515 100 12571 148
rect 13631 100 13687 148
rect 13763 100 13819 148
rect 14879 100 14935 148
rect 15011 100 15067 148
rect 16127 100 16183 148
rect 16259 100 16315 148
rect 17375 100 17431 148
rect 17507 100 17563 148
rect 18623 100 18679 148
rect 18755 100 18811 148
rect 19871 100 19927 148
rect 20003 100 20059 148
rect 21119 100 21175 148
rect 21251 100 21307 148
rect 22367 100 22423 148
rect 22499 100 22555 148
rect 23615 100 23671 148
rect 23747 100 23803 148
rect 24863 100 24919 148
rect 24995 100 25051 148
rect 26111 100 26167 148
rect 26243 100 26299 148
rect 27359 100 27415 148
rect 27491 100 27547 148
rect 28607 100 28663 148
rect 28739 100 28795 148
rect 29855 100 29911 148
rect 29987 100 30043 148
rect 31103 100 31159 148
rect 31235 100 31291 148
<< metal3 >>
rect 33 1250 31244 1316
rect 0 496 31821 556
rect 0 372 31821 432
rect 1963 218 3023 278
rect 3211 218 4271 278
rect 4459 218 5519 278
rect 5707 218 6767 278
rect 6955 218 8015 278
rect 8203 218 9263 278
rect 9451 218 10511 278
rect 10699 218 11759 278
rect 11947 218 13007 278
rect 13195 218 14255 278
rect 14443 218 15503 278
rect 15691 218 16751 278
rect 16939 218 17999 278
rect 18187 218 19247 278
rect 19435 218 20495 278
rect 20683 218 21743 278
rect 21931 218 22991 278
rect 23179 218 24239 278
rect 24427 218 25487 278
rect 25675 218 26735 278
rect 26923 218 27983 278
rect 28171 218 29231 278
rect 29419 218 30479 278
rect 30667 218 31727 278
rect 2427 94 2559 154
rect 3675 94 3807 154
rect 4923 94 5055 154
rect 6171 94 6303 154
rect 7419 94 7551 154
rect 8667 94 8799 154
rect 9915 94 10047 154
rect 11163 94 11295 154
rect 12411 94 12543 154
rect 13659 94 13791 154
rect 14907 94 15039 154
rect 16155 94 16287 154
rect 17403 94 17535 154
rect 18651 94 18783 154
rect 19899 94 20031 154
rect 21147 94 21279 154
rect 22395 94 22527 154
rect 23643 94 23775 154
rect 24891 94 25023 154
rect 26139 94 26271 154
rect 27387 94 27519 154
rect 28635 94 28767 154
rect 29883 94 30015 154
rect 31131 94 31263 154
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_0
timestamp 1661296025
transform -1 0 31821 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_1
timestamp 1661296025
transform 1 0 30573 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_2
timestamp 1661296025
transform -1 0 30573 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_3
timestamp 1661296025
transform 1 0 29325 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_4
timestamp 1661296025
transform -1 0 29325 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_5
timestamp 1661296025
transform 1 0 28077 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_6
timestamp 1661296025
transform -1 0 28077 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_7
timestamp 1661296025
transform 1 0 26829 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_8
timestamp 1661296025
transform -1 0 26829 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_9
timestamp 1661296025
transform 1 0 25581 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_10
timestamp 1661296025
transform -1 0 25581 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_11
timestamp 1661296025
transform 1 0 24333 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_12
timestamp 1661296025
transform -1 0 24333 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_13
timestamp 1661296025
transform 1 0 23085 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_14
timestamp 1661296025
transform -1 0 23085 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_15
timestamp 1661296025
transform 1 0 21837 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_16
timestamp 1661296025
transform -1 0 21837 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_17
timestamp 1661296025
transform 1 0 20589 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_18
timestamp 1661296025
transform -1 0 20589 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_19
timestamp 1661296025
transform 1 0 19341 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_20
timestamp 1661296025
transform -1 0 19341 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_21
timestamp 1661296025
transform 1 0 18093 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_22
timestamp 1661296025
transform -1 0 18093 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_23
timestamp 1661296025
transform 1 0 16845 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_24
timestamp 1661296025
transform -1 0 16845 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_25
timestamp 1661296025
transform 1 0 15597 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_26
timestamp 1661296025
transform -1 0 15597 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_27
timestamp 1661296025
transform 1 0 14349 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_28
timestamp 1661296025
transform -1 0 14349 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_29
timestamp 1661296025
transform 1 0 13101 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_30
timestamp 1661296025
transform -1 0 13101 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_31
timestamp 1661296025
transform 1 0 11853 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_32
timestamp 1661296025
transform -1 0 11853 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_33
timestamp 1661296025
transform 1 0 10605 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_34
timestamp 1661296025
transform -1 0 10605 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_35
timestamp 1661296025
transform 1 0 9357 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_36
timestamp 1661296025
transform -1 0 9357 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_37
timestamp 1661296025
transform 1 0 8109 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_38
timestamp 1661296025
transform -1 0 8109 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_39
timestamp 1661296025
transform 1 0 6861 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_40
timestamp 1661296025
transform -1 0 6861 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_41
timestamp 1661296025
transform 1 0 5613 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_42
timestamp 1661296025
transform -1 0 5613 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_43
timestamp 1661296025
transform 1 0 4365 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_44
timestamp 1661296025
transform -1 0 4365 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_45
timestamp 1661296025
transform 1 0 3117 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_46
timestamp 1661296025
transform -1 0 3117 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_column_mux  sky130_sram_1r1w_24x128_8_column_mux_47
timestamp 1661296025
transform 1 0 1869 0 1 620
box 65 0 675 1316
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_0
timestamp 1661296025
transform 1 0 31165 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_1
timestamp 1661296025
transform 1 0 31165 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_2
timestamp 1661296025
transform 1 0 29917 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_3
timestamp 1661296025
transform 1 0 29917 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_4
timestamp 1661296025
transform 1 0 28669 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_5
timestamp 1661296025
transform 1 0 28669 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_6
timestamp 1661296025
transform 1 0 27421 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_7
timestamp 1661296025
transform 1 0 27421 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_8
timestamp 1661296025
transform 1 0 26173 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_9
timestamp 1661296025
transform 1 0 26173 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_10
timestamp 1661296025
transform 1 0 24925 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_11
timestamp 1661296025
transform 1 0 24925 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_12
timestamp 1661296025
transform 1 0 23677 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_13
timestamp 1661296025
transform 1 0 23677 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_14
timestamp 1661296025
transform 1 0 22429 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_15
timestamp 1661296025
transform 1 0 22429 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_16
timestamp 1661296025
transform 1 0 21181 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_17
timestamp 1661296025
transform 1 0 21181 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_18
timestamp 1661296025
transform 1 0 19933 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_19
timestamp 1661296025
transform 1 0 19933 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_20
timestamp 1661296025
transform 1 0 18685 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_21
timestamp 1661296025
transform 1 0 18685 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_22
timestamp 1661296025
transform 1 0 17437 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_23
timestamp 1661296025
transform 1 0 17437 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_24
timestamp 1661296025
transform 1 0 16189 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_25
timestamp 1661296025
transform 1 0 16189 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_26
timestamp 1661296025
transform 1 0 14941 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_27
timestamp 1661296025
transform 1 0 14941 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_28
timestamp 1661296025
transform 1 0 13693 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_29
timestamp 1661296025
transform 1 0 13693 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_30
timestamp 1661296025
transform 1 0 12445 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_31
timestamp 1661296025
transform 1 0 12445 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_32
timestamp 1661296025
transform 1 0 11197 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_33
timestamp 1661296025
transform 1 0 11197 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_34
timestamp 1661296025
transform 1 0 9949 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_35
timestamp 1661296025
transform 1 0 9949 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_36
timestamp 1661296025
transform 1 0 8701 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_37
timestamp 1661296025
transform 1 0 8701 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_38
timestamp 1661296025
transform 1 0 7453 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_39
timestamp 1661296025
transform 1 0 7453 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_40
timestamp 1661296025
transform 1 0 6205 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_41
timestamp 1661296025
transform 1 0 6205 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_42
timestamp 1661296025
transform 1 0 4957 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_43
timestamp 1661296025
transform 1 0 4957 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_44
timestamp 1661296025
transform 1 0 3709 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_45
timestamp 1661296025
transform 1 0 3709 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_46
timestamp 1661296025
transform 1 0 2461 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_47
timestamp 1661296025
transform 1 0 2461 0 1 1251
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_0
timestamp 1661296025
transform 1 0 31164 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_1
timestamp 1661296025
transform 1 0 31164 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_2
timestamp 1661296025
transform 1 0 29916 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_3
timestamp 1661296025
transform 1 0 29916 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_4
timestamp 1661296025
transform 1 0 28668 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_5
timestamp 1661296025
transform 1 0 28668 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_6
timestamp 1661296025
transform 1 0 27420 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_7
timestamp 1661296025
transform 1 0 27420 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_8
timestamp 1661296025
transform 1 0 26172 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_9
timestamp 1661296025
transform 1 0 26172 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_10
timestamp 1661296025
transform 1 0 24924 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_11
timestamp 1661296025
transform 1 0 24924 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_12
timestamp 1661296025
transform 1 0 23676 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_13
timestamp 1661296025
transform 1 0 23676 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_14
timestamp 1661296025
transform 1 0 22428 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_15
timestamp 1661296025
transform 1 0 22428 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_16
timestamp 1661296025
transform 1 0 21180 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_17
timestamp 1661296025
transform 1 0 21180 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_18
timestamp 1661296025
transform 1 0 19932 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_19
timestamp 1661296025
transform 1 0 19932 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_20
timestamp 1661296025
transform 1 0 18684 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_21
timestamp 1661296025
transform 1 0 18684 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_22
timestamp 1661296025
transform 1 0 17436 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_23
timestamp 1661296025
transform 1 0 17436 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_24
timestamp 1661296025
transform 1 0 16188 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_25
timestamp 1661296025
transform 1 0 16188 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_26
timestamp 1661296025
transform 1 0 14940 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_27
timestamp 1661296025
transform 1 0 14940 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_28
timestamp 1661296025
transform 1 0 13692 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_29
timestamp 1661296025
transform 1 0 13692 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_30
timestamp 1661296025
transform 1 0 12444 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_31
timestamp 1661296025
transform 1 0 12444 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_32
timestamp 1661296025
transform 1 0 11196 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_33
timestamp 1661296025
transform 1 0 11196 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_34
timestamp 1661296025
transform 1 0 9948 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_35
timestamp 1661296025
transform 1 0 9948 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_36
timestamp 1661296025
transform 1 0 8700 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_37
timestamp 1661296025
transform 1 0 8700 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_38
timestamp 1661296025
transform 1 0 7452 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_39
timestamp 1661296025
transform 1 0 7452 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_40
timestamp 1661296025
transform 1 0 6204 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_41
timestamp 1661296025
transform 1 0 6204 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_42
timestamp 1661296025
transform 1 0 4956 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_43
timestamp 1661296025
transform 1 0 4956 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_44
timestamp 1661296025
transform 1 0 3708 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_45
timestamp 1661296025
transform 1 0 3708 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_46
timestamp 1661296025
transform 1 0 2460 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_47
timestamp 1661296025
transform 1 0 2460 0 1 1246
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_0
timestamp 1661296025
transform 1 0 31462 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_1
timestamp 1661296025
transform 1 0 30866 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_2
timestamp 1661296025
transform 1 0 30214 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_3
timestamp 1661296025
transform 1 0 29618 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_4
timestamp 1661296025
transform 1 0 28966 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_5
timestamp 1661296025
transform 1 0 28370 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_6
timestamp 1661296025
transform 1 0 27718 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_7
timestamp 1661296025
transform 1 0 27122 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_8
timestamp 1661296025
transform 1 0 26470 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_9
timestamp 1661296025
transform 1 0 25874 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_10
timestamp 1661296025
transform 1 0 25222 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_11
timestamp 1661296025
transform 1 0 24626 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_12
timestamp 1661296025
transform 1 0 23974 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_13
timestamp 1661296025
transform 1 0 23378 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_14
timestamp 1661296025
transform 1 0 22726 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_15
timestamp 1661296025
transform 1 0 22130 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_16
timestamp 1661296025
transform 1 0 21478 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_17
timestamp 1661296025
transform 1 0 20882 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_18
timestamp 1661296025
transform 1 0 20230 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_19
timestamp 1661296025
transform 1 0 19634 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_20
timestamp 1661296025
transform 1 0 18982 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_21
timestamp 1661296025
transform 1 0 18386 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_22
timestamp 1661296025
transform 1 0 17734 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_23
timestamp 1661296025
transform 1 0 17138 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_24
timestamp 1661296025
transform 1 0 16486 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_25
timestamp 1661296025
transform 1 0 15890 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_26
timestamp 1661296025
transform 1 0 15238 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_27
timestamp 1661296025
transform 1 0 14642 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_28
timestamp 1661296025
transform 1 0 13990 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_29
timestamp 1661296025
transform 1 0 13394 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_30
timestamp 1661296025
transform 1 0 12742 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_31
timestamp 1661296025
transform 1 0 12146 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_32
timestamp 1661296025
transform 1 0 11494 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_33
timestamp 1661296025
transform 1 0 10898 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_34
timestamp 1661296025
transform 1 0 10246 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_35
timestamp 1661296025
transform 1 0 9650 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_36
timestamp 1661296025
transform 1 0 8998 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_37
timestamp 1661296025
transform 1 0 8402 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_38
timestamp 1661296025
transform 1 0 7750 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_39
timestamp 1661296025
transform 1 0 7154 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_40
timestamp 1661296025
transform 1 0 6502 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_41
timestamp 1661296025
transform 1 0 5906 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_42
timestamp 1661296025
transform 1 0 5254 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_43
timestamp 1661296025
transform 1 0 4658 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_44
timestamp 1661296025
transform 1 0 4006 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_45
timestamp 1661296025
transform 1 0 3410 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_46
timestamp 1661296025
transform 1 0 2758 0 1 493
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_24  sky130_sram_1r1w_24x128_8_contact_24_47
timestamp 1661296025
transform 1 0 2162 0 1 369
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_0
timestamp 1661296025
transform 1 0 31466 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_1
timestamp 1661296025
transform 1 0 30870 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_2
timestamp 1661296025
transform 1 0 30218 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_3
timestamp 1661296025
transform 1 0 29622 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_4
timestamp 1661296025
transform 1 0 28970 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_5
timestamp 1661296025
transform 1 0 28374 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_6
timestamp 1661296025
transform 1 0 27722 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_7
timestamp 1661296025
transform 1 0 27126 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_8
timestamp 1661296025
transform 1 0 26474 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_9
timestamp 1661296025
transform 1 0 25878 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_10
timestamp 1661296025
transform 1 0 25226 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_11
timestamp 1661296025
transform 1 0 24630 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_12
timestamp 1661296025
transform 1 0 23978 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_13
timestamp 1661296025
transform 1 0 23382 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_14
timestamp 1661296025
transform 1 0 22730 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_15
timestamp 1661296025
transform 1 0 22134 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_16
timestamp 1661296025
transform 1 0 21482 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_17
timestamp 1661296025
transform 1 0 20886 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_18
timestamp 1661296025
transform 1 0 20234 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_19
timestamp 1661296025
transform 1 0 19638 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_20
timestamp 1661296025
transform 1 0 18986 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_21
timestamp 1661296025
transform 1 0 18390 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_22
timestamp 1661296025
transform 1 0 17738 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_23
timestamp 1661296025
transform 1 0 17142 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_24
timestamp 1661296025
transform 1 0 16490 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_25
timestamp 1661296025
transform 1 0 15894 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_26
timestamp 1661296025
transform 1 0 15242 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_27
timestamp 1661296025
transform 1 0 14646 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_28
timestamp 1661296025
transform 1 0 13994 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_29
timestamp 1661296025
transform 1 0 13398 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_30
timestamp 1661296025
transform 1 0 12746 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_31
timestamp 1661296025
transform 1 0 12150 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_32
timestamp 1661296025
transform 1 0 11498 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_33
timestamp 1661296025
transform 1 0 10902 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_34
timestamp 1661296025
transform 1 0 10250 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_35
timestamp 1661296025
transform 1 0 9654 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_36
timestamp 1661296025
transform 1 0 9002 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_37
timestamp 1661296025
transform 1 0 8406 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_38
timestamp 1661296025
transform 1 0 7754 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_39
timestamp 1661296025
transform 1 0 7158 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_40
timestamp 1661296025
transform 1 0 6506 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_41
timestamp 1661296025
transform 1 0 5910 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_42
timestamp 1661296025
transform 1 0 5258 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_43
timestamp 1661296025
transform 1 0 4662 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_44
timestamp 1661296025
transform 1 0 4010 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_45
timestamp 1661296025
transform 1 0 3414 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_46
timestamp 1661296025
transform 1 0 2762 0 1 493
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_25  sky130_sram_1r1w_24x128_8_contact_25_47
timestamp 1661296025
transform 1 0 2166 0 1 369
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_0
timestamp 1661296025
transform 1 0 31231 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_1
timestamp 1661296025
transform 1 0 31695 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_2
timestamp 1661296025
transform 1 0 31099 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_3
timestamp 1661296025
transform 1 0 30635 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_4
timestamp 1661296025
transform 1 0 29983 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_5
timestamp 1661296025
transform 1 0 30447 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_6
timestamp 1661296025
transform 1 0 29851 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_7
timestamp 1661296025
transform 1 0 29387 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_8
timestamp 1661296025
transform 1 0 28735 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_9
timestamp 1661296025
transform 1 0 29199 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_10
timestamp 1661296025
transform 1 0 28603 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_11
timestamp 1661296025
transform 1 0 28139 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_12
timestamp 1661296025
transform 1 0 27487 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_13
timestamp 1661296025
transform 1 0 27951 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_14
timestamp 1661296025
transform 1 0 27355 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_15
timestamp 1661296025
transform 1 0 26891 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_16
timestamp 1661296025
transform 1 0 26239 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_17
timestamp 1661296025
transform 1 0 26703 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_18
timestamp 1661296025
transform 1 0 26107 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_19
timestamp 1661296025
transform 1 0 25643 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_20
timestamp 1661296025
transform 1 0 24991 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_21
timestamp 1661296025
transform 1 0 25455 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_22
timestamp 1661296025
transform 1 0 24859 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_23
timestamp 1661296025
transform 1 0 24395 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_24
timestamp 1661296025
transform 1 0 23743 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_25
timestamp 1661296025
transform 1 0 24207 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_26
timestamp 1661296025
transform 1 0 23611 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_27
timestamp 1661296025
transform 1 0 23147 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_28
timestamp 1661296025
transform 1 0 22495 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_29
timestamp 1661296025
transform 1 0 22959 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_30
timestamp 1661296025
transform 1 0 22363 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_31
timestamp 1661296025
transform 1 0 21899 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_32
timestamp 1661296025
transform 1 0 21247 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_33
timestamp 1661296025
transform 1 0 21711 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_34
timestamp 1661296025
transform 1 0 21115 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_35
timestamp 1661296025
transform 1 0 20651 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_36
timestamp 1661296025
transform 1 0 19999 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_37
timestamp 1661296025
transform 1 0 20463 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_38
timestamp 1661296025
transform 1 0 19867 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_39
timestamp 1661296025
transform 1 0 19403 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_40
timestamp 1661296025
transform 1 0 18751 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_41
timestamp 1661296025
transform 1 0 19215 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_42
timestamp 1661296025
transform 1 0 18619 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_43
timestamp 1661296025
transform 1 0 18155 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_44
timestamp 1661296025
transform 1 0 17503 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_45
timestamp 1661296025
transform 1 0 17967 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_46
timestamp 1661296025
transform 1 0 17371 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_47
timestamp 1661296025
transform 1 0 16907 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_48
timestamp 1661296025
transform 1 0 16255 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_49
timestamp 1661296025
transform 1 0 16719 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_50
timestamp 1661296025
transform 1 0 16123 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_51
timestamp 1661296025
transform 1 0 15659 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_52
timestamp 1661296025
transform 1 0 15007 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_53
timestamp 1661296025
transform 1 0 15471 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_54
timestamp 1661296025
transform 1 0 14875 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_55
timestamp 1661296025
transform 1 0 14411 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_56
timestamp 1661296025
transform 1 0 13759 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_57
timestamp 1661296025
transform 1 0 14223 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_58
timestamp 1661296025
transform 1 0 13627 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_59
timestamp 1661296025
transform 1 0 13163 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_60
timestamp 1661296025
transform 1 0 12511 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_61
timestamp 1661296025
transform 1 0 12975 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_62
timestamp 1661296025
transform 1 0 12379 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_63
timestamp 1661296025
transform 1 0 11915 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_64
timestamp 1661296025
transform 1 0 11263 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_65
timestamp 1661296025
transform 1 0 11727 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_66
timestamp 1661296025
transform 1 0 11131 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_67
timestamp 1661296025
transform 1 0 10667 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_68
timestamp 1661296025
transform 1 0 10015 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_69
timestamp 1661296025
transform 1 0 10479 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_70
timestamp 1661296025
transform 1 0 9883 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_71
timestamp 1661296025
transform 1 0 9419 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_72
timestamp 1661296025
transform 1 0 8767 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_73
timestamp 1661296025
transform 1 0 9231 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_74
timestamp 1661296025
transform 1 0 8635 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_75
timestamp 1661296025
transform 1 0 8171 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_76
timestamp 1661296025
transform 1 0 7519 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_77
timestamp 1661296025
transform 1 0 7983 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_78
timestamp 1661296025
transform 1 0 7387 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_79
timestamp 1661296025
transform 1 0 6923 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_80
timestamp 1661296025
transform 1 0 6271 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_81
timestamp 1661296025
transform 1 0 6735 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_82
timestamp 1661296025
transform 1 0 6139 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_83
timestamp 1661296025
transform 1 0 5675 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_84
timestamp 1661296025
transform 1 0 5023 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_85
timestamp 1661296025
transform 1 0 5487 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_86
timestamp 1661296025
transform 1 0 4891 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_87
timestamp 1661296025
transform 1 0 4427 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_88
timestamp 1661296025
transform 1 0 3775 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_89
timestamp 1661296025
transform 1 0 4239 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_90
timestamp 1661296025
transform 1 0 3643 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_91
timestamp 1661296025
transform 1 0 3179 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_92
timestamp 1661296025
transform 1 0 2527 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_93
timestamp 1661296025
transform 1 0 2991 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_94
timestamp 1661296025
transform 1 0 2395 0 1 92
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_95
timestamp 1661296025
transform 1 0 1931 0 1 216
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_96
timestamp 1661296025
transform 1 0 31463 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_97
timestamp 1661296025
transform 1 0 30867 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_98
timestamp 1661296025
transform 1 0 30215 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_99
timestamp 1661296025
transform 1 0 29619 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_100
timestamp 1661296025
transform 1 0 28967 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_101
timestamp 1661296025
transform 1 0 28371 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_102
timestamp 1661296025
transform 1 0 27719 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_103
timestamp 1661296025
transform 1 0 27123 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_104
timestamp 1661296025
transform 1 0 26471 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_105
timestamp 1661296025
transform 1 0 25875 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_106
timestamp 1661296025
transform 1 0 25223 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_107
timestamp 1661296025
transform 1 0 24627 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_108
timestamp 1661296025
transform 1 0 23975 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_109
timestamp 1661296025
transform 1 0 23379 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_110
timestamp 1661296025
transform 1 0 22727 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_111
timestamp 1661296025
transform 1 0 22131 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_112
timestamp 1661296025
transform 1 0 21479 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_113
timestamp 1661296025
transform 1 0 20883 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_114
timestamp 1661296025
transform 1 0 20231 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_115
timestamp 1661296025
transform 1 0 19635 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_116
timestamp 1661296025
transform 1 0 18983 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_117
timestamp 1661296025
transform 1 0 18387 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_118
timestamp 1661296025
transform 1 0 17735 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_119
timestamp 1661296025
transform 1 0 17139 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_120
timestamp 1661296025
transform 1 0 16487 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_121
timestamp 1661296025
transform 1 0 15891 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_122
timestamp 1661296025
transform 1 0 15239 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_123
timestamp 1661296025
transform 1 0 14643 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_124
timestamp 1661296025
transform 1 0 13991 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_125
timestamp 1661296025
transform 1 0 13395 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_126
timestamp 1661296025
transform 1 0 12743 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_127
timestamp 1661296025
transform 1 0 12147 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_128
timestamp 1661296025
transform 1 0 11495 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_129
timestamp 1661296025
transform 1 0 10899 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_130
timestamp 1661296025
transform 1 0 10247 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_131
timestamp 1661296025
transform 1 0 9651 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_132
timestamp 1661296025
transform 1 0 8999 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_133
timestamp 1661296025
transform 1 0 8403 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_134
timestamp 1661296025
transform 1 0 7751 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_135
timestamp 1661296025
transform 1 0 7155 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_136
timestamp 1661296025
transform 1 0 6503 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_137
timestamp 1661296025
transform 1 0 5907 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_138
timestamp 1661296025
transform 1 0 5255 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_139
timestamp 1661296025
transform 1 0 4659 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_140
timestamp 1661296025
transform 1 0 4007 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_141
timestamp 1661296025
transform 1 0 3411 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_142
timestamp 1661296025
transform 1 0 2759 0 1 494
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_26  sky130_sram_1r1w_24x128_8_contact_26_143
timestamp 1661296025
transform 1 0 2163 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_0
timestamp 1661296025
transform 1 0 31230 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_1
timestamp 1661296025
transform 1 0 31694 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_2
timestamp 1661296025
transform 1 0 31098 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_3
timestamp 1661296025
transform 1 0 30634 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_4
timestamp 1661296025
transform 1 0 29982 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_5
timestamp 1661296025
transform 1 0 30446 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_6
timestamp 1661296025
transform 1 0 29850 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_7
timestamp 1661296025
transform 1 0 29386 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_8
timestamp 1661296025
transform 1 0 28734 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_9
timestamp 1661296025
transform 1 0 29198 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_10
timestamp 1661296025
transform 1 0 28602 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_11
timestamp 1661296025
transform 1 0 28138 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_12
timestamp 1661296025
transform 1 0 27486 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_13
timestamp 1661296025
transform 1 0 27950 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_14
timestamp 1661296025
transform 1 0 27354 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_15
timestamp 1661296025
transform 1 0 26890 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_16
timestamp 1661296025
transform 1 0 26238 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_17
timestamp 1661296025
transform 1 0 26702 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_18
timestamp 1661296025
transform 1 0 26106 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_19
timestamp 1661296025
transform 1 0 25642 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_20
timestamp 1661296025
transform 1 0 24990 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_21
timestamp 1661296025
transform 1 0 25454 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_22
timestamp 1661296025
transform 1 0 24858 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_23
timestamp 1661296025
transform 1 0 24394 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_24
timestamp 1661296025
transform 1 0 23742 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_25
timestamp 1661296025
transform 1 0 24206 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_26
timestamp 1661296025
transform 1 0 23610 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_27
timestamp 1661296025
transform 1 0 23146 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_28
timestamp 1661296025
transform 1 0 22494 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_29
timestamp 1661296025
transform 1 0 22958 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_30
timestamp 1661296025
transform 1 0 22362 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_31
timestamp 1661296025
transform 1 0 21898 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_32
timestamp 1661296025
transform 1 0 21246 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_33
timestamp 1661296025
transform 1 0 21710 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_34
timestamp 1661296025
transform 1 0 21114 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_35
timestamp 1661296025
transform 1 0 20650 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_36
timestamp 1661296025
transform 1 0 19998 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_37
timestamp 1661296025
transform 1 0 20462 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_38
timestamp 1661296025
transform 1 0 19866 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_39
timestamp 1661296025
transform 1 0 19402 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_40
timestamp 1661296025
transform 1 0 18750 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_41
timestamp 1661296025
transform 1 0 19214 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_42
timestamp 1661296025
transform 1 0 18618 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_43
timestamp 1661296025
transform 1 0 18154 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_44
timestamp 1661296025
transform 1 0 17502 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_45
timestamp 1661296025
transform 1 0 17966 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_46
timestamp 1661296025
transform 1 0 17370 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_47
timestamp 1661296025
transform 1 0 16906 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_48
timestamp 1661296025
transform 1 0 16254 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_49
timestamp 1661296025
transform 1 0 16718 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_50
timestamp 1661296025
transform 1 0 16122 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_51
timestamp 1661296025
transform 1 0 15658 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_52
timestamp 1661296025
transform 1 0 15006 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_53
timestamp 1661296025
transform 1 0 15470 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_54
timestamp 1661296025
transform 1 0 14874 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_55
timestamp 1661296025
transform 1 0 14410 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_56
timestamp 1661296025
transform 1 0 13758 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_57
timestamp 1661296025
transform 1 0 14222 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_58
timestamp 1661296025
transform 1 0 13626 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_59
timestamp 1661296025
transform 1 0 13162 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_60
timestamp 1661296025
transform 1 0 12510 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_61
timestamp 1661296025
transform 1 0 12974 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_62
timestamp 1661296025
transform 1 0 12378 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_63
timestamp 1661296025
transform 1 0 11914 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_64
timestamp 1661296025
transform 1 0 11262 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_65
timestamp 1661296025
transform 1 0 11726 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_66
timestamp 1661296025
transform 1 0 11130 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_67
timestamp 1661296025
transform 1 0 10666 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_68
timestamp 1661296025
transform 1 0 10014 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_69
timestamp 1661296025
transform 1 0 10478 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_70
timestamp 1661296025
transform 1 0 9882 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_71
timestamp 1661296025
transform 1 0 9418 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_72
timestamp 1661296025
transform 1 0 8766 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_73
timestamp 1661296025
transform 1 0 9230 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_74
timestamp 1661296025
transform 1 0 8634 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_75
timestamp 1661296025
transform 1 0 8170 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_76
timestamp 1661296025
transform 1 0 7518 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_77
timestamp 1661296025
transform 1 0 7982 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_78
timestamp 1661296025
transform 1 0 7386 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_79
timestamp 1661296025
transform 1 0 6922 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_80
timestamp 1661296025
transform 1 0 6270 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_81
timestamp 1661296025
transform 1 0 6734 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_82
timestamp 1661296025
transform 1 0 6138 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_83
timestamp 1661296025
transform 1 0 5674 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_84
timestamp 1661296025
transform 1 0 5022 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_85
timestamp 1661296025
transform 1 0 5486 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_86
timestamp 1661296025
transform 1 0 4890 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_87
timestamp 1661296025
transform 1 0 4426 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_88
timestamp 1661296025
transform 1 0 3774 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_89
timestamp 1661296025
transform 1 0 4238 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_90
timestamp 1661296025
transform 1 0 3642 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_91
timestamp 1661296025
transform 1 0 3178 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_92
timestamp 1661296025
transform 1 0 2526 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_93
timestamp 1661296025
transform 1 0 2990 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_94
timestamp 1661296025
transform 1 0 2394 0 1 87
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_95
timestamp 1661296025
transform 1 0 1930 0 1 211
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_96
timestamp 1661296025
transform 1 0 31462 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_97
timestamp 1661296025
transform 1 0 30866 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_98
timestamp 1661296025
transform 1 0 30214 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_99
timestamp 1661296025
transform 1 0 29618 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_100
timestamp 1661296025
transform 1 0 28966 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_101
timestamp 1661296025
transform 1 0 28370 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_102
timestamp 1661296025
transform 1 0 27718 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_103
timestamp 1661296025
transform 1 0 27122 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_104
timestamp 1661296025
transform 1 0 26470 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_105
timestamp 1661296025
transform 1 0 25874 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_106
timestamp 1661296025
transform 1 0 25222 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_107
timestamp 1661296025
transform 1 0 24626 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_108
timestamp 1661296025
transform 1 0 23974 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_109
timestamp 1661296025
transform 1 0 23378 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_110
timestamp 1661296025
transform 1 0 22726 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_111
timestamp 1661296025
transform 1 0 22130 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_112
timestamp 1661296025
transform 1 0 21478 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_113
timestamp 1661296025
transform 1 0 20882 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_114
timestamp 1661296025
transform 1 0 20230 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_115
timestamp 1661296025
transform 1 0 19634 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_116
timestamp 1661296025
transform 1 0 18982 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_117
timestamp 1661296025
transform 1 0 18386 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_118
timestamp 1661296025
transform 1 0 17734 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_119
timestamp 1661296025
transform 1 0 17138 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_120
timestamp 1661296025
transform 1 0 16486 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_121
timestamp 1661296025
transform 1 0 15890 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_122
timestamp 1661296025
transform 1 0 15238 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_123
timestamp 1661296025
transform 1 0 14642 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_124
timestamp 1661296025
transform 1 0 13990 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_125
timestamp 1661296025
transform 1 0 13394 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_126
timestamp 1661296025
transform 1 0 12742 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_127
timestamp 1661296025
transform 1 0 12146 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_128
timestamp 1661296025
transform 1 0 11494 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_129
timestamp 1661296025
transform 1 0 10898 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_130
timestamp 1661296025
transform 1 0 10246 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_131
timestamp 1661296025
transform 1 0 9650 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_132
timestamp 1661296025
transform 1 0 8998 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_133
timestamp 1661296025
transform 1 0 8402 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_134
timestamp 1661296025
transform 1 0 7750 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_135
timestamp 1661296025
transform 1 0 7154 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_136
timestamp 1661296025
transform 1 0 6502 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_137
timestamp 1661296025
transform 1 0 5906 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_138
timestamp 1661296025
transform 1 0 5254 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_139
timestamp 1661296025
transform 1 0 4658 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_140
timestamp 1661296025
transform 1 0 4006 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_141
timestamp 1661296025
transform 1 0 3410 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_142
timestamp 1661296025
transform 1 0 2758 0 1 489
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_27  sky130_sram_1r1w_24x128_8_contact_27_143
timestamp 1661296025
transform 1 0 2162 0 1 365
box 0 0 66 74
<< labels >>
rlabel metal3 s 0 372 31821 432 4 sel_0
port 1 nsew
rlabel metal3 s 0 496 31821 556 4 sel_1
port 2 nsew
rlabel metal1 s 1949 248 1977 620 4 bl_out_0
port 3 nsew
rlabel metal1 s 2413 124 2441 620 4 br_out_0
port 4 nsew
rlabel metal1 s 3197 248 3225 620 4 bl_out_1
port 5 nsew
rlabel metal1 s 3661 124 3689 620 4 br_out_1
port 6 nsew
rlabel metal1 s 4445 248 4473 620 4 bl_out_2
port 7 nsew
rlabel metal1 s 4909 124 4937 620 4 br_out_2
port 8 nsew
rlabel metal1 s 5693 248 5721 620 4 bl_out_3
port 9 nsew
rlabel metal1 s 6157 124 6185 620 4 br_out_3
port 10 nsew
rlabel metal1 s 6941 248 6969 620 4 bl_out_4
port 11 nsew
rlabel metal1 s 7405 124 7433 620 4 br_out_4
port 12 nsew
rlabel metal1 s 8189 248 8217 620 4 bl_out_5
port 13 nsew
rlabel metal1 s 8653 124 8681 620 4 br_out_5
port 14 nsew
rlabel metal1 s 9437 248 9465 620 4 bl_out_6
port 15 nsew
rlabel metal1 s 9901 124 9929 620 4 br_out_6
port 16 nsew
rlabel metal1 s 10685 248 10713 620 4 bl_out_7
port 17 nsew
rlabel metal1 s 11149 124 11177 620 4 br_out_7
port 18 nsew
rlabel metal1 s 11933 248 11961 620 4 bl_out_8
port 19 nsew
rlabel metal1 s 12397 124 12425 620 4 br_out_8
port 20 nsew
rlabel metal1 s 13181 248 13209 620 4 bl_out_9
port 21 nsew
rlabel metal1 s 13645 124 13673 620 4 br_out_9
port 22 nsew
rlabel metal1 s 14429 248 14457 620 4 bl_out_10
port 23 nsew
rlabel metal1 s 14893 124 14921 620 4 br_out_10
port 24 nsew
rlabel metal1 s 15677 248 15705 620 4 bl_out_11
port 25 nsew
rlabel metal1 s 16141 124 16169 620 4 br_out_11
port 26 nsew
rlabel metal1 s 16925 248 16953 620 4 bl_out_12
port 27 nsew
rlabel metal1 s 17389 124 17417 620 4 br_out_12
port 28 nsew
rlabel metal1 s 18173 248 18201 620 4 bl_out_13
port 29 nsew
rlabel metal1 s 18637 124 18665 620 4 br_out_13
port 30 nsew
rlabel metal1 s 19421 248 19449 620 4 bl_out_14
port 31 nsew
rlabel metal1 s 19885 124 19913 620 4 br_out_14
port 32 nsew
rlabel metal1 s 20669 248 20697 620 4 bl_out_15
port 33 nsew
rlabel metal1 s 21133 124 21161 620 4 br_out_15
port 34 nsew
rlabel metal1 s 21917 248 21945 620 4 bl_out_16
port 35 nsew
rlabel metal1 s 22381 124 22409 620 4 br_out_16
port 36 nsew
rlabel metal1 s 23165 248 23193 620 4 bl_out_17
port 37 nsew
rlabel metal1 s 23629 124 23657 620 4 br_out_17
port 38 nsew
rlabel metal1 s 24413 248 24441 620 4 bl_out_18
port 39 nsew
rlabel metal1 s 24877 124 24905 620 4 br_out_18
port 40 nsew
rlabel metal1 s 25661 248 25689 620 4 bl_out_19
port 41 nsew
rlabel metal1 s 26125 124 26153 620 4 br_out_19
port 42 nsew
rlabel metal1 s 26909 248 26937 620 4 bl_out_20
port 43 nsew
rlabel metal1 s 27373 124 27401 620 4 br_out_20
port 44 nsew
rlabel metal1 s 28157 248 28185 620 4 bl_out_21
port 45 nsew
rlabel metal1 s 28621 124 28649 620 4 br_out_21
port 46 nsew
rlabel metal1 s 29405 248 29433 620 4 bl_out_22
port 47 nsew
rlabel metal1 s 29869 124 29897 620 4 br_out_22
port 48 nsew
rlabel metal1 s 30653 248 30681 620 4 bl_out_23
port 49 nsew
rlabel metal1 s 31117 124 31145 620 4 br_out_23
port 50 nsew
rlabel metal3 s 33 1250 31244 1316 4 gnd
port 51 nsew
rlabel metal1 s 1949 1880 1977 1936 4 bl_0
port 52 nsew
rlabel metal1 s 2413 1880 2441 1936 4 br_0
port 53 nsew
rlabel metal1 s 3009 1880 3037 1936 4 bl_1
port 54 nsew
rlabel metal1 s 2545 1880 2573 1936 4 br_1
port 55 nsew
rlabel metal1 s 3197 1880 3225 1936 4 bl_2
port 56 nsew
rlabel metal1 s 3661 1880 3689 1936 4 br_2
port 57 nsew
rlabel metal1 s 4257 1880 4285 1936 4 bl_3
port 58 nsew
rlabel metal1 s 3793 1880 3821 1936 4 br_3
port 59 nsew
rlabel metal1 s 4445 1880 4473 1936 4 bl_4
port 60 nsew
rlabel metal1 s 4909 1880 4937 1936 4 br_4
port 61 nsew
rlabel metal1 s 5505 1880 5533 1936 4 bl_5
port 62 nsew
rlabel metal1 s 5041 1880 5069 1936 4 br_5
port 63 nsew
rlabel metal1 s 5693 1880 5721 1936 4 bl_6
port 64 nsew
rlabel metal1 s 6157 1880 6185 1936 4 br_6
port 65 nsew
rlabel metal1 s 6753 1880 6781 1936 4 bl_7
port 66 nsew
rlabel metal1 s 6289 1880 6317 1936 4 br_7
port 67 nsew
rlabel metal1 s 6941 1880 6969 1936 4 bl_8
port 68 nsew
rlabel metal1 s 7405 1880 7433 1936 4 br_8
port 69 nsew
rlabel metal1 s 8001 1880 8029 1936 4 bl_9
port 70 nsew
rlabel metal1 s 7537 1880 7565 1936 4 br_9
port 71 nsew
rlabel metal1 s 8189 1880 8217 1936 4 bl_10
port 72 nsew
rlabel metal1 s 8653 1880 8681 1936 4 br_10
port 73 nsew
rlabel metal1 s 9249 1880 9277 1936 4 bl_11
port 74 nsew
rlabel metal1 s 8785 1880 8813 1936 4 br_11
port 75 nsew
rlabel metal1 s 9437 1880 9465 1936 4 bl_12
port 76 nsew
rlabel metal1 s 9901 1880 9929 1936 4 br_12
port 77 nsew
rlabel metal1 s 10497 1880 10525 1936 4 bl_13
port 78 nsew
rlabel metal1 s 10033 1880 10061 1936 4 br_13
port 79 nsew
rlabel metal1 s 10685 1880 10713 1936 4 bl_14
port 80 nsew
rlabel metal1 s 11149 1880 11177 1936 4 br_14
port 81 nsew
rlabel metal1 s 11745 1880 11773 1936 4 bl_15
port 82 nsew
rlabel metal1 s 11281 1880 11309 1936 4 br_15
port 83 nsew
rlabel metal1 s 11933 1880 11961 1936 4 bl_16
port 84 nsew
rlabel metal1 s 12397 1880 12425 1936 4 br_16
port 85 nsew
rlabel metal1 s 12993 1880 13021 1936 4 bl_17
port 86 nsew
rlabel metal1 s 12529 1880 12557 1936 4 br_17
port 87 nsew
rlabel metal1 s 13181 1880 13209 1936 4 bl_18
port 88 nsew
rlabel metal1 s 13645 1880 13673 1936 4 br_18
port 89 nsew
rlabel metal1 s 14241 1880 14269 1936 4 bl_19
port 90 nsew
rlabel metal1 s 13777 1880 13805 1936 4 br_19
port 91 nsew
rlabel metal1 s 14429 1880 14457 1936 4 bl_20
port 92 nsew
rlabel metal1 s 14893 1880 14921 1936 4 br_20
port 93 nsew
rlabel metal1 s 15489 1880 15517 1936 4 bl_21
port 94 nsew
rlabel metal1 s 15025 1880 15053 1936 4 br_21
port 95 nsew
rlabel metal1 s 15677 1880 15705 1936 4 bl_22
port 96 nsew
rlabel metal1 s 16141 1880 16169 1936 4 br_22
port 97 nsew
rlabel metal1 s 16737 1880 16765 1936 4 bl_23
port 98 nsew
rlabel metal1 s 16273 1880 16301 1936 4 br_23
port 99 nsew
rlabel metal1 s 16925 1880 16953 1936 4 bl_24
port 100 nsew
rlabel metal1 s 17389 1880 17417 1936 4 br_24
port 101 nsew
rlabel metal1 s 17985 1880 18013 1936 4 bl_25
port 102 nsew
rlabel metal1 s 17521 1880 17549 1936 4 br_25
port 103 nsew
rlabel metal1 s 18173 1880 18201 1936 4 bl_26
port 104 nsew
rlabel metal1 s 18637 1880 18665 1936 4 br_26
port 105 nsew
rlabel metal1 s 19233 1880 19261 1936 4 bl_27
port 106 nsew
rlabel metal1 s 18769 1880 18797 1936 4 br_27
port 107 nsew
rlabel metal1 s 19421 1880 19449 1936 4 bl_28
port 108 nsew
rlabel metal1 s 19885 1880 19913 1936 4 br_28
port 109 nsew
rlabel metal1 s 20481 1880 20509 1936 4 bl_29
port 110 nsew
rlabel metal1 s 20017 1880 20045 1936 4 br_29
port 111 nsew
rlabel metal1 s 20669 1880 20697 1936 4 bl_30
port 112 nsew
rlabel metal1 s 21133 1880 21161 1936 4 br_30
port 113 nsew
rlabel metal1 s 21729 1880 21757 1936 4 bl_31
port 114 nsew
rlabel metal1 s 21265 1880 21293 1936 4 br_31
port 115 nsew
rlabel metal1 s 21917 1880 21945 1936 4 bl_32
port 116 nsew
rlabel metal1 s 22381 1880 22409 1936 4 br_32
port 117 nsew
rlabel metal1 s 22977 1880 23005 1936 4 bl_33
port 118 nsew
rlabel metal1 s 22513 1880 22541 1936 4 br_33
port 119 nsew
rlabel metal1 s 23165 1880 23193 1936 4 bl_34
port 120 nsew
rlabel metal1 s 23629 1880 23657 1936 4 br_34
port 121 nsew
rlabel metal1 s 24225 1880 24253 1936 4 bl_35
port 122 nsew
rlabel metal1 s 23761 1880 23789 1936 4 br_35
port 123 nsew
rlabel metal1 s 24413 1880 24441 1936 4 bl_36
port 124 nsew
rlabel metal1 s 24877 1880 24905 1936 4 br_36
port 125 nsew
rlabel metal1 s 25473 1880 25501 1936 4 bl_37
port 126 nsew
rlabel metal1 s 25009 1880 25037 1936 4 br_37
port 127 nsew
rlabel metal1 s 25661 1880 25689 1936 4 bl_38
port 128 nsew
rlabel metal1 s 26125 1880 26153 1936 4 br_38
port 129 nsew
rlabel metal1 s 26721 1880 26749 1936 4 bl_39
port 130 nsew
rlabel metal1 s 26257 1880 26285 1936 4 br_39
port 131 nsew
rlabel metal1 s 26909 1880 26937 1936 4 bl_40
port 132 nsew
rlabel metal1 s 27373 1880 27401 1936 4 br_40
port 133 nsew
rlabel metal1 s 27969 1880 27997 1936 4 bl_41
port 134 nsew
rlabel metal1 s 27505 1880 27533 1936 4 br_41
port 135 nsew
rlabel metal1 s 28157 1880 28185 1936 4 bl_42
port 136 nsew
rlabel metal1 s 28621 1880 28649 1936 4 br_42
port 137 nsew
rlabel metal1 s 29217 1880 29245 1936 4 bl_43
port 138 nsew
rlabel metal1 s 28753 1880 28781 1936 4 br_43
port 139 nsew
rlabel metal1 s 29405 1880 29433 1936 4 bl_44
port 140 nsew
rlabel metal1 s 29869 1880 29897 1936 4 br_44
port 141 nsew
rlabel metal1 s 30465 1880 30493 1936 4 bl_45
port 142 nsew
rlabel metal1 s 30001 1880 30029 1936 4 br_45
port 143 nsew
rlabel metal1 s 30653 1880 30681 1936 4 bl_46
port 144 nsew
rlabel metal1 s 31117 1880 31145 1936 4 br_46
port 145 nsew
rlabel metal1 s 31713 1880 31741 1936 4 bl_47
port 146 nsew
rlabel metal1 s 31249 1880 31277 1936 4 br_47
port 147 nsew
<< properties >>
string FIXED_BBOX 0 0 29952 1936
<< end >>
