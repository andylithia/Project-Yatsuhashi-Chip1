magic
tech sky130B
timestamp 1659145761
<< metal4 >>
rect -200 2350 3400 2400
rect -200 1650 -150 2350
rect 450 2300 3400 2350
rect 450 2200 3500 2300
rect 6400 2250 7200 2300
rect 450 1650 3600 2200
rect -200 1600 3600 1650
rect 2800 -400 3600 1600
rect 6400 1650 6450 2250
rect 7150 1650 7200 2250
rect 6400 -400 7200 1650
<< via4 >>
rect -150 1650 450 2350
rect 6450 1650 7150 2250
<< metal5 >>
rect 0 9500 10000 10000
rect 0 2550 500 9500
rect -50 2500 500 2550
rect -100 2450 500 2500
rect -150 2400 500 2450
rect -200 2350 500 2400
rect -200 1650 -150 2350
rect 450 1650 500 2350
rect -200 1600 500 1650
rect 800 8700 9200 9200
rect 800 500 1300 8700
rect 1600 7900 8400 8400
rect 1600 1300 2100 7900
rect 6400 2250 7200 2300
rect 6400 1650 6450 2250
rect 7150 2200 7250 2250
rect 7150 2150 7300 2200
rect 7150 2100 7350 2150
rect 7900 2100 8400 7900
rect 7150 1650 8400 2100
rect 6400 1600 8400 1650
rect 8700 1300 9200 8700
rect 1600 800 9200 1300
rect 9500 500 10000 9500
rect 800 0 10000 500
<< labels >>
rlabel metal4 6400 -400 7200 -100 1 B
rlabel metal4 2800 -400 3600 -100 1 A
<< end >>
