magic
tech sky130B
timestamp 1660959839
<< metal1 >>
rect -1000 3500 0 3700
rect -1000 -100 -900 3500
rect -100 2200 0 3500
rect 2400 3500 3400 3700
rect 2400 2200 2500 3500
rect -100 -100 2500 2200
rect 3300 -100 3400 3500
rect -1000 -300 3400 -100
<< via1 >>
rect -900 -100 -100 3500
rect 2500 -100 3300 3500
<< metal2 >>
rect -1000 3500 0 3700
rect -1000 -100 -900 3500
rect -100 2200 0 3500
rect 2400 3500 3400 3700
rect 2400 2200 2500 3500
rect -100 -100 2500 2200
rect 3300 -100 3400 3500
rect -1000 -300 3400 -100
<< via2 >>
rect -900 -100 -100 3500
rect 2500 -100 3300 3500
<< metal3 >>
rect -1000 3500 0 3700
rect -1000 -100 -900 3500
rect -100 2200 0 3500
rect 2400 3500 3400 3700
rect 2400 2200 2500 3500
rect -100 -100 2500 2200
rect 3300 -100 3400 3500
rect -1000 -300 3400 -100
<< via3 >>
rect -900 -100 -100 3500
rect 2500 -100 3300 3500
<< metal4 >>
rect -1000 3500 0 3700
rect -1000 -100 -900 3500
rect -100 -100 0 3500
rect -1000 -300 0 -100
rect 2400 3500 3400 3700
rect 2400 -100 2500 3500
rect 3300 -100 3400 3500
rect 2400 -300 3400 -100
<< via4 >>
rect -900 -100 -100 3500
rect 2500 -100 3300 3500
<< metal5 >>
rect -1000 3500 0 3700
rect -1000 -100 -900 3500
rect -100 -100 0 3500
rect -1000 -300 0 -100
rect 300 -300 2100 3700
rect 2400 3500 3400 3700
rect 2400 -100 2500 3500
rect 3300 -100 3400 3500
rect 2400 -300 3400 -100
<< end >>
