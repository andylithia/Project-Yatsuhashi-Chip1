magic
tech sky130A
timestamp 1659498593
<< metal4 >>
rect 260 -110 740 150
rect 0 -590 1000 -110
rect 260 -850 740 -590
<< end >>
