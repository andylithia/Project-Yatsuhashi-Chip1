magic
tech sky130A
magscale 1 2
timestamp 1665275356
<< metal4 >>
rect 14000 1863 41000 1975
rect 14000 -3913 14112 1863
rect 19888 -3913 35112 1863
rect 40888 -3913 41000 1863
rect 14000 -4025 41000 -3913
<< via4 >>
rect 14112 -3913 19888 1863
rect 35112 -3913 40888 1863
<< metal5 >>
tri -28000 20477 -25477 23000 se
rect -25477 20477 18477 23000
tri 18477 20477 21000 23000 sw
tri -31477 17000 -28000 20477 se
rect -28000 17000 21000 20477
tri 21000 17000 24477 20477 sw
tri -35000 13477 -31477 17000 se
rect -31477 16000 -23991 17000
tri -23991 16000 -22991 17000 nw
tri 15991 16000 16991 17000 ne
rect 16991 16000 24477 17000
rect -31477 14586 -25405 16000
tri -25405 14586 -23991 16000 nw
tri -23991 14586 -22577 16000 se
rect -22577 14586 15577 16000
tri 15577 14586 16991 16000 sw
tri 16991 14586 18405 16000 ne
rect 18405 14586 24477 16000
rect -31477 13477 -26586 14586
tri -36486 11991 -35000 13477 se
rect -35000 13405 -26586 13477
tri -26586 13405 -25405 14586 nw
tri -25172 13405 -23991 14586 se
rect -23991 13405 16991 14586
rect -35000 11991 -28000 13405
tri -28000 11991 -26586 13405 nw
tri -26586 11991 -25172 13405 se
rect -25172 13172 16991 13405
tri 16991 13172 18405 14586 sw
tri 18405 13172 19819 14586 ne
rect 19819 13172 24477 14586
rect -25172 12828 18405 13172
tri 18405 12828 18749 13172 sw
tri 19819 12828 20163 13172 ne
rect 20163 12828 24477 13172
rect -25172 11991 18749 12828
tri -41000 7477 -36486 11991 se
rect -36486 10577 -29414 11991
tri -29414 10577 -28000 11991 nw
tri -28000 10577 -26586 11991 se
rect -26586 11414 18749 11991
tri 18749 11414 20163 12828 sw
tri 20163 11414 21577 12828 ne
rect 21577 11414 24477 12828
rect -26586 10577 20163 11414
tri 20163 10577 21000 11414 sw
tri 21577 10577 22414 11414 ne
rect 22414 10577 24477 11414
rect -36486 10000 -29991 10577
tri -29991 10000 -29414 10577 nw
tri -28577 10000 -28000 10577 se
rect -28000 10000 21000 10577
tri 21000 10000 21577 10577 sw
tri 22414 10000 22991 10577 ne
rect 22991 10000 24477 10577
tri 24477 10000 31477 17000 sw
rect -36486 9092 -30899 10000
tri -30899 9092 -29991 10000 nw
tri -29485 9092 -28577 10000 se
rect -28577 9092 -21000 10000
tri -21000 9092 -20092 10000 nw
tri 13092 9092 14000 10000 ne
rect 14000 9092 21577 10000
rect -36486 7678 -32313 9092
tri -32313 7678 -30899 9092 nw
tri -30899 7678 -29485 9092 se
rect -29485 7678 -22414 9092
tri -22414 7678 -21000 9092 nw
tri 14000 9000 14092 9092 ne
rect 14092 9000 21577 9092
tri -21000 7678 -19678 9000 se
rect -19678 7678 12678 9000
tri 12678 7678 14000 9000 sw
tri 14092 7678 15414 9000 ne
rect 15414 8586 21577 9000
tri 21577 8586 22991 10000 sw
tri 22991 8586 24405 10000 ne
rect 24405 8586 31477 10000
rect 15414 7678 22991 8586
rect -36486 7477 -32586 7678
rect -41000 7405 -32586 7477
tri -32586 7405 -32313 7678 nw
tri -31172 7405 -30899 7678 se
rect -30899 7405 -23828 7678
rect -41000 5991 -34000 7405
tri -34000 5991 -32586 7405 nw
tri -32586 5991 -31172 7405 se
rect -31172 6264 -23828 7405
tri -23828 6264 -22414 7678 nw
tri -22414 6264 -21000 7678 se
rect -21000 7586 14000 7678
tri 14000 7586 14092 7678 sw
tri 15414 7586 15506 7678 ne
rect 15506 7586 22991 7678
rect -21000 6264 14092 7586
rect -31172 5991 -25242 6264
rect -41000 3000 -35000 5991
tri -35000 4991 -34000 5991 nw
tri -33586 4991 -32586 5991 se
rect -32586 4991 -25242 5991
rect -47000 -3000 -35000 3000
tri -34000 4577 -33586 4991 se
rect -33586 4850 -25242 4991
tri -25242 4850 -23828 6264 nw
tri -23828 4850 -22414 6264 se
rect -22414 6172 14092 6264
tri 14092 6172 15506 7586 sw
tri 15506 6172 16920 7586 ne
rect 16920 7405 22991 7586
tri 22991 7405 24172 8586 sw
tri 24405 7405 25586 8586 ne
rect 25586 7477 31477 8586
tri 31477 7477 34000 10000 sw
rect 25586 7405 34000 7477
rect 16920 6172 24172 7405
rect -22414 5828 15506 6172
tri 15506 5828 15850 6172 sw
tri 16920 5828 17264 6172 ne
rect 17264 5991 24172 6172
tri 24172 5991 25586 7405 sw
tri 25586 5991 27000 7405 ne
rect 27000 5991 34000 7405
rect 17264 5828 25586 5991
rect -22414 4850 15850 5828
rect -33586 4577 -25586 4850
rect -34000 4506 -25586 4577
tri -25586 4506 -25242 4850 nw
tri -24172 4506 -23828 4850 se
rect -23828 4506 15850 4850
rect -34000 3092 -27000 4506
tri -27000 3092 -25586 4506 nw
tri -25586 3092 -24172 4506 se
rect -24172 4414 15850 4506
tri 15850 4414 17264 5828 sw
tri 17264 4414 18678 5828 ne
rect 18678 4991 25586 5828
tri 25586 4991 26586 5991 sw
tri 27000 4991 28000 5991 ne
rect 18678 4577 26586 4991
tri 26586 4577 27000 4991 sw
rect 18678 4414 27000 4577
rect -24172 3092 17264 4414
rect -34000 3000 -27092 3092
tri -27092 3000 -27000 3092 nw
tri -25678 3000 -25586 3092 se
rect -25586 3000 17264 3092
tri 17264 3000 18678 4414 sw
tri 18678 3000 20092 4414 ne
rect 20092 3000 27000 4414
rect -34000 -8042 -28000 3000
tri -28000 2092 -27092 3000 nw
tri -26586 2092 -25678 3000 se
rect -25678 2092 -21000 3000
tri -27000 1678 -26586 2092 se
rect -26586 1678 -21000 2092
rect -27000 -6627 -21000 1678
tri -21000 -808 -17192 3000 nw
tri 10192 -808 14000 3000 ne
rect 14000 2092 18678 3000
tri 18678 2092 19586 3000 sw
tri 20092 2092 21000 3000 ne
rect 14000 1975 19586 2092
tri 19586 1975 19703 2092 sw
rect 14000 1863 20000 1975
rect 14000 -3913 14112 1863
rect 19888 -3913 20000 1863
rect 14000 -4025 20000 -3913
tri -27000 -7042 -26585 -6627 ne
rect -26585 -7042 -21000 -6627
tri -28000 -8042 -27000 -7042 sw
tri -26585 -8042 -25585 -7042 ne
rect -25585 -8042 -21000 -7042
rect -34000 -8585 -27000 -8042
tri -27000 -8585 -26457 -8042 sw
tri -25585 -8585 -25042 -8042 ne
rect -25042 -8585 -21000 -8042
rect -34000 -9527 -26457 -8585
tri -34000 -10000 -33527 -9527 ne
rect -33527 -10000 -26457 -9527
tri -26457 -10000 -25042 -8585 sw
tri -25042 -10000 -23627 -8585 ne
rect -23627 -10000 -21000 -8585
tri -21000 -10000 -15142 -4142 sw
tri 15142 -10000 21000 -4142 se
rect 21000 -6627 27000 3000
rect 21000 -7042 26585 -6627
tri 26585 -7042 27000 -6627 nw
rect 21000 -8042 25585 -7042
tri 25585 -8042 26585 -7042 nw
tri 27000 -8042 28000 -7042 se
rect 28000 -8042 34000 5991
rect 35000 1863 41000 1975
rect 35000 -3913 35112 1863
rect 40888 -3913 41000 1863
rect 35000 -4025 41000 -3913
rect 21000 -8585 25042 -8042
tri 25042 -8585 25585 -8042 nw
tri 26457 -8585 27000 -8042 se
rect 27000 -8585 34000 -8042
rect 21000 -10000 23627 -8585
tri 23627 -10000 25042 -8585 nw
tri 25042 -10000 26457 -8585 se
rect 26457 -9527 34000 -8585
rect 26457 -10000 29485 -9527
tri -33527 -17000 -26527 -10000 ne
rect -26527 -11415 -25042 -10000
tri -25042 -11415 -23627 -10000 sw
tri -23627 -11415 -22212 -10000 ne
rect -22212 -11212 22415 -10000
tri 22415 -11212 23627 -10000 nw
tri 23830 -11212 25042 -10000 se
rect 25042 -11212 29485 -10000
rect -22212 -11415 21000 -11212
rect -26527 -12830 -23627 -11415
tri -23627 -12830 -22212 -11415 sw
tri -22212 -12830 -20797 -11415 ne
rect -20797 -12627 21000 -11415
tri 21000 -12627 22415 -11212 nw
tri 22415 -12627 23830 -11212 se
rect 23830 -12627 29485 -11212
rect -20797 -12830 19585 -12627
rect -26527 -13170 -22212 -12830
tri -22212 -13170 -21872 -12830 sw
tri -20797 -13170 -20457 -12830 ne
rect -20457 -13170 19585 -12830
rect -26527 -14585 -21872 -13170
tri -21872 -14585 -20457 -13170 sw
tri -20457 -14585 -19042 -13170 ne
rect -19042 -14042 19585 -13170
tri 19585 -14042 21000 -12627 nw
tri 21000 -14042 22415 -12627 se
rect 22415 -14042 29485 -12627
tri 29485 -14042 34000 -9527 nw
rect -19042 -14585 19042 -14042
tri 19042 -14585 19585 -14042 nw
tri 20457 -14585 21000 -14042 se
rect 21000 -14585 28000 -14042
rect -26527 -16000 -20457 -14585
tri -20457 -16000 -19042 -14585 sw
tri -19042 -16000 -17627 -14585 ne
rect -17627 -16000 17627 -14585
tri 17627 -16000 19042 -14585 nw
tri 19042 -16000 20457 -14585 se
rect 20457 -15527 28000 -14585
tri 28000 -15527 29485 -14042 nw
rect 20457 -16000 26527 -15527
rect -26527 -17000 -19042 -16000
tri -19042 -17000 -18042 -16000 sw
tri 18042 -17000 19042 -16000 se
rect 19042 -17000 26527 -16000
tri 26527 -17000 28000 -15527 nw
tri -26527 -22527 -21000 -17000 ne
rect -21000 -22527 21000 -17000
tri 21000 -22527 26527 -17000 nw
tri -21000 -23000 -20527 -22527 ne
rect -20527 -23000 20527 -22527
tri 20527 -23000 21000 -22527 nw
<< end >>
