magic
tech sky130B
timestamp 1666844558
<< end >>
