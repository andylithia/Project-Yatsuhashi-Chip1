** sch_path:
*+ /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA5_with_output_buf_4_SP_PEX.sch
**.subckt LNA5_with_output_buf_4_SP_PEX
V1 VDD GND 1.8
V2 net3 GND dc 0.9 ac 1 portnum 1 z0 50
I0 VDDI Vref 2m
XM1 Vref Vref GNDI GNDI sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=2
XC7 Vref GNDI sky130_fd_pr__cap_mim_m3_1 W=20 L=30 MF=1 m=1
Ldeg5 net1 VDDI 2n m=1
R3 net1 VDD 3 m=1
Ldeg6 net2 GND 2n m=1
R4 net2 GNDI 3 m=1
C17 net7 net4 0.3p m=1
L2 VDDI net4 2.5n m=1
XC3 net12 GNDI sky130_fd_pr__cap_mim_m3_1 W=40 L=60 MF=8 m=8
C8 GNDI GND 200f m=1
C19 VDD VDDI 200f m=1
R2 net12 VDDI 5 m=1
C1 net5 net3 1n m=1
Ldeg1 net6 net5 2n m=1
L1 net10 vmid 0.7n m=1
Ldeg2 net11 net6 0.5n m=1
XC4 net13 GNDI sky130_fd_pr__cap_mim_m3_1 W=40 L=60 MF=8 m=8
R8 net13 VDDI 5 m=1
L4 net9 GNDI 0.15n m=1
V3 net7 GNDI dc 0.9 ac 1 portnum 2 z0 50
R7 net8 VDDI 5k m=1
C5 GNDI net8 50f m=1
x1 VDDI net4 GNDI VDDI GNDI GNDI __UNCONNECTED_PIN__0 VDDI __UNCONNECTED_PIN__1 net10 vmid net9 Vref
+ net11 GNDI LNA_complete_2_wo_ind_PEX
**** begin user architecture code


.subckt sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=4.242e+12p
+ ps=3.198e+07u w=5.05e+06u l=150000u
X1 SOURCE SUBSTRATE SUBSTRATE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.03e+12p
+ ps=2.14e+07u w=5.05e+06u l=150000u
X2 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X5 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends
.sp dec 1000 0.1e9 100e9 1
* .ac dec 1000 0.01e9 100e9
.control
run
display
let z11=50*(1+s_1_1)/(1-s_1_1)
let z22=50*(1+s_2_2)/(1-s_2_2)
let S11 = S_1_1
let S21 = S_2_1
let S12 = S_1_2
let S22 = S_2_2

* Stability
let delta=S11*S22-S12*S21
let K    = (1-mag(S11)^2-mag(S22)^2+mag(delta)^2)/(2*mag(S12*S21))
let mu   = (1-mag(S11)^2)/(mag(S22-conj(S11)*delta)+mag(S21*S12))
* plot real(z11) real(z22)
* plot imag(z11) imag(z22)
plot db(S_1_1) db(S_2_2) db(S_2_1)

plot db(K)
plot mag(delta)
plot db(mu)
plot NF NFmin
.endc


.lib /home/andylithia/openmpw/pdk_1/sky130B/libs.tech/ngspice/sky130.lib.spice tt
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130B/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

**** end user architecture code
**.ends

* expanding   symbol:  LNA_complete_2_wo_ind_PEX.sym # of pins=15
** sym_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA_complete_2_wo_ind_PEX.sym
** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/LNA_complete_2_wo_ind_PEX.sch
.subckt LNA_complete_2_wo_ind_PEX  VHI VOUT G4 G8 G2 G1 RFB_MID G_TOP BIAS_TOP S1 D1 SS BIAS_BOT VIN
+ VLO
*.iopin VHI
*.iopin VLO
*.iopin VOUT
*.iopin VIN
*.iopin SS
*.iopin D1
*.iopin S1
*.iopin BIAS_BOT
*.iopin BIAS_TOP
*.iopin G_TOP
*.iopin G2
*.iopin G8
*.iopin G4
*.iopin G1
*.iopin RFB_MID
**** begin user architecture code

X0 S1.t11 G_TOP VOUT.t2 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X1 SS.t7 VIN D1.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X2 VHI VLO sky130_fd_pr__cap_mim_m3_2 l=4.4e+07u w=5e+07u
X3 VOUT.t5 G_TOP S1.t10 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SS.t6 VIN D1.t3 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X5 D1.t0 VIN SS.t5 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X6 VHI a_n6328_16092.t2 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2.5e+06u
X7 D1.t2 VIN SS.t4 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X8 S1.t9 G_TOP VOUT.t4 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X9 SS.t3 VIN D1.t5 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X10 D1.t4 VIN SS.t2 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X11 VLO VHI sky130_fd_pr__cap_mim_m3_1 l=4.4e+07u w=5e+07u
X12 S1.t8 G_TOP VOUT.t7 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X13 VOUT.t8 G_TOP S1.t7 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X14 D1.t6 VIN SS.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X15 VOUT.t3 G_TOP S1.t6 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X16 a_n6328_16092.t1 G1 VOUT.t12 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X17 a_n5540_16092.t1 G4 VOUT.t16 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X18 S1.t5 G_TOP VOUT.t11 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X19 VOUT.t15 G2 a_n6722_16092.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X20 VOUT.t18 G8 a_n5934_16092.t2 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X21 VOUT.t0 G_TOP S1.t4 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X22 S1.t3 G_TOP VOUT.t9 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X23 VOUT.t10 G_TOP S1.t2 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X24 VOUT.t6 G_TOP S1.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X25 S1.t0 G_TOP VOUT.t1 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X26 VHI a_n5934_16092.t0 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=8e+06u
X27 VOUT.t13 G1 a_n6328_16092.t0 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X28 VOUT.t17 G4 a_n5540_16092.t0 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X29 a_n5934_16092.t1 G8 VOUT.t19 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X30 VHI a_n5540_16092.t2 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=4e+06u
X31 VHI a_n6722_16092.t2 sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=2.5e+06u
X32 a_n6722_16092.t0 G2 VOUT.t14 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X33 SS.t0 VIN D1.t7 VLO sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R0 VOUT.n135 VOUT.n722 9.305
R1 VOUT.n136 VOUT.n603 9.305
R2 VOUT.n137 VOUT.n663 9.305
R3 VOUT.n724 VOUT.n725 9.3
R4 VOUT.n85 VOUT.n737 9.3
R5 VOUT.n15 VOUT.n748 9.3
R6 VOUT.n75 VOUT.n728 9.3
R7 VOUT.n731 VOUT.n730 9.3
R8 VOUT.n84 VOUT.n734 9.3
R9 VOUT.n85 VOUT.n736 9.3
R10 VOUT.n119 VOUT.n740 9.3
R11 VOUT.n120 VOUT.n743 9.3
R12 VOUT.n120 VOUT.n742 9.3
R13 VOUT.n138 VOUT.n746 9.3
R14 VOUT.n86 VOUT.n721 9.3
R15 VOUT.n15 VOUT.n749 9.3
R16 VOUT.n88 VOUT.n618 9.3
R17 VOUT.n87 VOUT.n615 9.3
R18 VOUT.n121 VOUT.n621 9.3
R19 VOUT.n612 VOUT.n611 9.3
R20 VOUT.n72 VOUT.n609 9.3
R21 VOUT.n605 VOUT.n606 9.3
R22 VOUT.n122 VOUT.n624 9.3
R23 VOUT.n14 VOUT.n630 9.3
R24 VOUT.n14 VOUT.n629 9.3
R25 VOUT.n89 VOUT.n602 9.3
R26 VOUT.n139 VOUT.n627 9.3
R27 VOUT.n122 VOUT.n623 9.3
R28 VOUT.n88 VOUT.n617 9.3
R29 VOUT.n92 VOUT.n682 9.3
R30 VOUT.n125 VOUT.n704 9.3
R31 VOUT.n124 VOUT.n701 9.3
R32 VOUT.n13 VOUT.n710 9.3
R33 VOUT.n13 VOUT.n709 9.3
R34 VOUT.n140 VOUT.n707 9.3
R35 VOUT.n91 VOUT.n698 9.3
R36 VOUT.n91 VOUT.n697 9.3
R37 VOUT.n90 VOUT.n695 9.3
R38 VOUT.n692 VOUT.n691 9.3
R39 VOUT.n74 VOUT.n689 9.3
R40 VOUT.n685 VOUT.n686 9.3
R41 VOUT.n123 VOUT.n683 9.3
R42 VOUT.n125 VOUT.n703 9.3
R43 VOUT.n665 VOUT.n666 9.3
R44 VOUT.n672 VOUT.n671 9.3
R45 VOUT.n93 VOUT.n659 9.3
R46 VOUT.n12 VOUT.n647 9.3
R47 VOUT.n94 VOUT.n662 9.3
R48 VOUT.n93 VOUT.n660 9.3
R49 VOUT.n126 VOUT.n657 9.3
R50 VOUT.n642 VOUT.n641 9.3
R51 VOUT.n655 VOUT.n654 9.3
R52 VOUT.n141 VOUT.n645 9.3
R53 VOUT.n95 VOUT.n635 9.3
R54 VOUT.n12 VOUT.n648 9.3
R55 VOUT.n73 VOUT.n669 9.3
R56 VOUT.n108 VOUT.n513 9.3
R57 VOUT.n63 VOUT.n501 9.3
R58 VOUT.n109 VOUT.n490 9.3
R59 VOUT.n127 VOUT.n494 9.3
R60 VOUT.n127 VOUT.n495 9.3
R61 VOUT.n498 VOUT.n497 9.3
R62 VOUT.n62 VOUT.n500 9.3
R63 VOUT.n63 VOUT.n503 9.3
R64 VOUT.n145 VOUT.n504 9.3
R65 VOUT.n144 VOUT.n505 9.3
R66 VOUT.n144 VOUT.n507 9.3
R67 VOUT.n10 VOUT.n509 9.3
R68 VOUT.n108 VOUT.n511 9.3
R69 VOUT.n38 VOUT.n515 9.3
R70 VOUT.n1 VOUT.n517 9.3
R71 VOUT.n29 VOUT.n518 9.3
R72 VOUT.n80 VOUT.n450 9.3
R73 VOUT.n24 VOUT.n472 9.3
R74 VOUT.n97 VOUT.n485 9.3
R75 VOUT.n96 VOUT.n484 9.3
R76 VOUT.n96 VOUT.n483 9.3
R77 VOUT.n40 VOUT.n464 9.3
R78 VOUT.n41 VOUT.n465 9.3
R79 VOUT.n39 VOUT.n468 9.3
R80 VOUT.n459 VOUT.n469 9.3
R81 VOUT.n24 VOUT.n473 9.3
R82 VOUT.n25 VOUT.n474 9.3
R83 VOUT.n489 VOUT.n488 9.3
R84 VOUT.n109 VOUT.n491 9.3
R85 VOUT.n110 VOUT.n440 9.3
R86 VOUT.n65 VOUT.n428 9.3
R87 VOUT.n111 VOUT.n417 9.3
R88 VOUT.n128 VOUT.n421 9.3
R89 VOUT.n128 VOUT.n422 9.3
R90 VOUT.n425 VOUT.n424 9.3
R91 VOUT.n64 VOUT.n427 9.3
R92 VOUT.n65 VOUT.n430 9.3
R93 VOUT.n147 VOUT.n431 9.3
R94 VOUT.n146 VOUT.n432 9.3
R95 VOUT.n146 VOUT.n434 9.3
R96 VOUT.n9 VOUT.n436 9.3
R97 VOUT.n110 VOUT.n438 9.3
R98 VOUT.n42 VOUT.n442 9.3
R99 VOUT.n2 VOUT.n444 9.3
R100 VOUT.n30 VOUT.n445 9.3
R101 VOUT.n79 VOUT.n377 9.3
R102 VOUT.n22 VOUT.n399 9.3
R103 VOUT.n99 VOUT.n412 9.3
R104 VOUT.n98 VOUT.n411 9.3
R105 VOUT.n98 VOUT.n410 9.3
R106 VOUT.n44 VOUT.n391 9.3
R107 VOUT.n45 VOUT.n392 9.3
R108 VOUT.n43 VOUT.n395 9.3
R109 VOUT.n386 VOUT.n396 9.3
R110 VOUT.n22 VOUT.n400 9.3
R111 VOUT.n23 VOUT.n401 9.3
R112 VOUT.n416 VOUT.n415 9.3
R113 VOUT.n111 VOUT.n418 9.3
R114 VOUT.n112 VOUT.n220 9.3
R115 VOUT.n67 VOUT.n208 9.3
R116 VOUT.n113 VOUT.n197 9.3
R117 VOUT.n129 VOUT.n201 9.3
R118 VOUT.n129 VOUT.n202 9.3
R119 VOUT.n205 VOUT.n204 9.3
R120 VOUT.n66 VOUT.n207 9.3
R121 VOUT.n67 VOUT.n210 9.3
R122 VOUT.n149 VOUT.n211 9.3
R123 VOUT.n148 VOUT.n212 9.3
R124 VOUT.n148 VOUT.n214 9.3
R125 VOUT.n8 VOUT.n216 9.3
R126 VOUT.n112 VOUT.n218 9.3
R127 VOUT.n46 VOUT.n222 9.3
R128 VOUT.n3 VOUT.n224 9.3
R129 VOUT.n31 VOUT.n225 9.3
R130 VOUT.n76 VOUT.n157 9.3
R131 VOUT.n20 VOUT.n179 9.3
R132 VOUT.n101 VOUT.n192 9.3
R133 VOUT.n100 VOUT.n191 9.3
R134 VOUT.n100 VOUT.n190 9.3
R135 VOUT.n48 VOUT.n171 9.3
R136 VOUT.n49 VOUT.n172 9.3
R137 VOUT.n47 VOUT.n175 9.3
R138 VOUT.n166 VOUT.n176 9.3
R139 VOUT.n20 VOUT.n180 9.3
R140 VOUT.n21 VOUT.n181 9.3
R141 VOUT.n196 VOUT.n195 9.3
R142 VOUT.n113 VOUT.n198 9.3
R143 VOUT.n114 VOUT.n293 9.3
R144 VOUT.n69 VOUT.n281 9.3
R145 VOUT.n115 VOUT.n270 9.3
R146 VOUT.n130 VOUT.n274 9.3
R147 VOUT.n130 VOUT.n275 9.3
R148 VOUT.n278 VOUT.n277 9.3
R149 VOUT.n68 VOUT.n280 9.3
R150 VOUT.n69 VOUT.n283 9.3
R151 VOUT.n151 VOUT.n284 9.3
R152 VOUT.n150 VOUT.n285 9.3
R153 VOUT.n150 VOUT.n287 9.3
R154 VOUT.n7 VOUT.n289 9.3
R155 VOUT.n114 VOUT.n291 9.3
R156 VOUT.n50 VOUT.n295 9.3
R157 VOUT.n4 VOUT.n297 9.3
R158 VOUT.n32 VOUT.n298 9.3
R159 VOUT.n77 VOUT.n230 9.3
R160 VOUT.n18 VOUT.n252 9.3
R161 VOUT.n103 VOUT.n265 9.3
R162 VOUT.n102 VOUT.n264 9.3
R163 VOUT.n102 VOUT.n263 9.3
R164 VOUT.n52 VOUT.n244 9.3
R165 VOUT.n53 VOUT.n245 9.3
R166 VOUT.n51 VOUT.n248 9.3
R167 VOUT.n239 VOUT.n249 9.3
R168 VOUT.n18 VOUT.n253 9.3
R169 VOUT.n19 VOUT.n254 9.3
R170 VOUT.n269 VOUT.n268 9.3
R171 VOUT.n115 VOUT.n271 9.3
R172 VOUT.n116 VOUT.n366 9.3
R173 VOUT.n71 VOUT.n354 9.3
R174 VOUT.n117 VOUT.n343 9.3
R175 VOUT.n131 VOUT.n347 9.3
R176 VOUT.n131 VOUT.n348 9.3
R177 VOUT.n351 VOUT.n350 9.3
R178 VOUT.n70 VOUT.n353 9.3
R179 VOUT.n71 VOUT.n356 9.3
R180 VOUT.n153 VOUT.n357 9.3
R181 VOUT.n152 VOUT.n358 9.3
R182 VOUT.n152 VOUT.n360 9.3
R183 VOUT.n6 VOUT.n362 9.3
R184 VOUT.n116 VOUT.n364 9.3
R185 VOUT.n54 VOUT.n368 9.3
R186 VOUT.n5 VOUT.n370 9.3
R187 VOUT.n33 VOUT.n371 9.3
R188 VOUT.n78 VOUT.n303 9.3
R189 VOUT.n16 VOUT.n325 9.3
R190 VOUT.n105 VOUT.n338 9.3
R191 VOUT.n104 VOUT.n337 9.3
R192 VOUT.n104 VOUT.n336 9.3
R193 VOUT.n56 VOUT.n317 9.3
R194 VOUT.n57 VOUT.n318 9.3
R195 VOUT.n55 VOUT.n321 9.3
R196 VOUT.n312 VOUT.n322 9.3
R197 VOUT.n16 VOUT.n326 9.3
R198 VOUT.n17 VOUT.n327 9.3
R199 VOUT.n342 VOUT.n341 9.3
R200 VOUT.n117 VOUT.n344 9.3
R201 VOUT.n106 VOUT.n586 9.3
R202 VOUT.n61 VOUT.n573 9.3
R203 VOUT.n107 VOUT.n559 9.3
R204 VOUT.n118 VOUT.n566 9.3
R205 VOUT.n118 VOUT.n567 9.3
R206 VOUT.n60 VOUT.n572 9.3
R207 VOUT.n143 VOUT.n577 9.3
R208 VOUT.n142 VOUT.n578 9.3
R209 VOUT.n11 VOUT.n582 9.3
R210 VOUT.n34 VOUT.n588 9.3
R211 VOUT.n28 VOUT.n592 9.3
R212 VOUT.n26 VOUT.n539 9.3
R213 VOUT.n83 VOUT.n554 9.3
R214 VOUT.n82 VOUT.n553 9.3
R215 VOUT.n37 VOUT.n531 9.3
R216 VOUT.n526 VOUT.n536 9.3
R217 VOUT.n27 VOUT.n542 9.3
R218 VOUT.n107 VOUT.n560 9.3
R219 VOUT.n570 VOUT.n569 9.3
R220 VOUT.n61 VOUT.n575 9.3
R221 VOUT.n142 VOUT.n580 9.3
R222 VOUT.n106 VOUT.n584 9.3
R223 VOUT.n0 VOUT.n591 9.3
R224 VOUT.n81 VOUT.n524 9.3
R225 VOUT.n82 VOUT.n552 9.3
R226 VOUT.n36 VOUT.n529 9.3
R227 VOUT.n35 VOUT.n534 9.3
R228 VOUT.n26 VOUT.n540 9.3
R229 VOUT.n558 VOUT.n557 9.3
R230 VOUT.n123 VOUT.n684 9
R231 VOUT.n74 VOUT.n690 9
R232 VOUT.n90 VOUT.n696 9
R233 VOUT.n89 VOUT.n598 9
R234 VOUT.n86 VOUT.n717 9
R235 VOUT.n72 VOUT.n610 9
R236 VOUT.n136 VOUT.n604 9
R237 VOUT.n75 VOUT.n729 9
R238 VOUT.n84 VOUT.n735 9
R239 VOUT.n119 VOUT.n741 9
R240 VOUT.n92 VOUT.n678 9
R241 VOUT.n95 VOUT.n636 9
R242 VOUT.n94 VOUT.n652 9
R243 VOUT.n126 VOUT.n653 9
R244 VOUT.n13 VOUT.n711 9
R245 VOUT.n12 VOUT.n649 9
R246 VOUT.n141 VOUT.n646 9
R247 VOUT.n140 VOUT.n708 9
R248 VOUT.n124 VOUT.n702 9
R249 VOUT.n73 VOUT.n670 9
R250 VOUT.n14 VOUT.n631 9
R251 VOUT.n15 VOUT.n750 9
R252 VOUT.n138 VOUT.n747 9
R253 VOUT.n139 VOUT.n628 9
R254 VOUT.n121 VOUT.n622 9
R255 VOUT.n135 VOUT.n723 9
R256 VOUT.n87 VOUT.n616 9
R257 VOUT.n137 VOUT.n664 9
R258 VOUT.n80 VOUT.n451 9
R259 VOUT.n1 VOUT.n452 9
R260 VOUT.n10 VOUT.n510 9
R261 VOUT.n145 VOUT.n453 9
R262 VOUT.n62 VOUT.n499 9
R263 VOUT.n493 VOUT.n455 9
R264 VOUT.n40 VOUT.n461 9
R265 VOUT.n39 VOUT.n460 9
R266 VOUT.n25 VOUT.n458 9
R267 VOUT.n97 VOUT.n486 9
R268 VOUT.n492 VOUT.n456 9
R269 VOUT.n79 VOUT.n378 9
R270 VOUT.n2 VOUT.n379 9
R271 VOUT.n9 VOUT.n437 9
R272 VOUT.n147 VOUT.n380 9
R273 VOUT.n64 VOUT.n426 9
R274 VOUT.n420 VOUT.n382 9
R275 VOUT.n44 VOUT.n388 9
R276 VOUT.n43 VOUT.n387 9
R277 VOUT.n23 VOUT.n385 9
R278 VOUT.n99 VOUT.n413 9
R279 VOUT.n419 VOUT.n383 9
R280 VOUT.n76 VOUT.n158 9
R281 VOUT.n3 VOUT.n159 9
R282 VOUT.n8 VOUT.n217 9
R283 VOUT.n149 VOUT.n160 9
R284 VOUT.n66 VOUT.n206 9
R285 VOUT.n200 VOUT.n162 9
R286 VOUT.n48 VOUT.n168 9
R287 VOUT.n47 VOUT.n167 9
R288 VOUT.n21 VOUT.n165 9
R289 VOUT.n101 VOUT.n193 9
R290 VOUT.n199 VOUT.n163 9
R291 VOUT.n77 VOUT.n231 9
R292 VOUT.n4 VOUT.n232 9
R293 VOUT.n7 VOUT.n290 9
R294 VOUT.n151 VOUT.n233 9
R295 VOUT.n68 VOUT.n279 9
R296 VOUT.n273 VOUT.n235 9
R297 VOUT.n52 VOUT.n241 9
R298 VOUT.n51 VOUT.n240 9
R299 VOUT.n19 VOUT.n238 9
R300 VOUT.n103 VOUT.n266 9
R301 VOUT.n272 VOUT.n236 9
R302 VOUT.n78 VOUT.n304 9
R303 VOUT.n5 VOUT.n305 9
R304 VOUT.n6 VOUT.n363 9
R305 VOUT.n153 VOUT.n306 9
R306 VOUT.n70 VOUT.n352 9
R307 VOUT.n346 VOUT.n308 9
R308 VOUT.n56 VOUT.n314 9
R309 VOUT.n55 VOUT.n313 9
R310 VOUT.n17 VOUT.n311 9
R311 VOUT.n105 VOUT.n339 9
R312 VOUT.n345 VOUT.n309 9
R313 VOUT.n81 VOUT.n525 9
R314 VOUT.n0 VOUT.n589 9
R315 VOUT.n11 VOUT.n583 9
R316 VOUT.n143 VOUT.n576 9
R317 VOUT.n60 VOUT.n571 9
R318 VOUT.n565 VOUT.n564 9
R319 VOUT.n36 VOUT.n530 9
R320 VOUT.n35 VOUT.n535 9
R321 VOUT.n27 VOUT.n541 9
R322 VOUT.n83 VOUT.n555 9
R323 VOUT.n562 VOUT.n561 9
R324 VOUT.n455 VOUT.n454 8.282
R325 VOUT.n382 VOUT.n381 8.282
R326 VOUT.n162 VOUT.n161 8.282
R327 VOUT.n235 VOUT.n234 8.282
R328 VOUT.n308 VOUT.n307 8.282
R329 VOUT.n564 VOUT.n563 8.282
R330 VOUT.n523 VOUT.n522 7.854
R331 VOUT.n449 VOUT.n448 7.853
R332 VOUT.n376 VOUT.n375 7.853
R333 VOUT.n156 VOUT.n155 7.853
R334 VOUT.n229 VOUT.n228 7.853
R335 VOUT.n302 VOUT.n301 7.853
R336 VOUT.n463 VOUT.n462 7.851
R337 VOUT.n390 VOUT.n389 7.851
R338 VOUT.n170 VOUT.n169 7.851
R339 VOUT.n243 VOUT.n242 7.851
R340 VOUT.n316 VOUT.n315 7.851
R341 VOUT.n528 VOUT.n527 7.851
R342 VOUT.n478 VOUT.n477 4.65
R343 VOUT.n405 VOUT.n404 4.65
R344 VOUT.n185 VOUT.n184 4.65
R345 VOUT.n258 VOUT.n257 4.65
R346 VOUT.n331 VOUT.n330 4.65
R347 VOUT.n546 VOUT.n545 4.65
R348 VOUT.n650 VOUT.n640 4.61
R349 VOUT.n677 VOUT.n676 4.574
R350 VOUT.n597 VOUT.n596 4.574
R351 VOUT.n716 VOUT.n715 4.574
R352 VOUT.n479 VOUT.n457 4.574
R353 VOUT.n406 VOUT.n384 4.574
R354 VOUT.n186 VOUT.n164 4.574
R355 VOUT.n259 VOUT.n237 4.574
R356 VOUT.n332 VOUT.n310 4.574
R357 VOUT.n548 VOUT.n547 4.574
R358 VOUT.n715 VOUT.n714 3.388
R359 VOUT.n596 VOUT.n595 3.388
R360 VOUT.n676 VOUT.n675 3.388
R361 VOUT.n640 VOUT.n639 3.388
R362 VOUT.n718 VOUT.t16 3.326
R363 VOUT.n718 VOUT.t17 3.326
R364 VOUT.n599 VOUT.t19 3.326
R365 VOUT.n599 VOUT.t18 3.326
R366 VOUT.n679 VOUT.t12 3.326
R367 VOUT.n679 VOUT.t13 3.326
R368 VOUT.n633 VOUT.t14 3.326
R369 VOUT.n633 VOUT.t15 3.326
R370 VOUT.n447 VOUT.t2 3.326
R371 VOUT.n447 VOUT.t5 3.326
R372 VOUT.n374 VOUT.t7 3.326
R373 VOUT.n374 VOUT.t6 3.326
R374 VOUT.n154 VOUT.t11 3.326
R375 VOUT.n154 VOUT.t8 3.326
R376 VOUT.n227 VOUT.t1 3.326
R377 VOUT.n227 VOUT.t10 3.326
R378 VOUT.n300 VOUT.t9 3.326
R379 VOUT.n300 VOUT.t3 3.326
R380 VOUT.n521 VOUT.t4 3.326
R381 VOUT.n521 VOUT.t0 3.326
R382 VOUT.n513 VOUT.n512 3.191
R383 VOUT.n440 VOUT.n439 3.191
R384 VOUT.n220 VOUT.n219 3.191
R385 VOUT.n293 VOUT.n292 3.191
R386 VOUT.n366 VOUT.n365 3.191
R387 VOUT.n586 VOUT.n585 3.191
R388 VOUT.n519 VOUT.n80 3.055
R389 VOUT.n446 VOUT.n79 3.055
R390 VOUT.n226 VOUT.n76 3.055
R391 VOUT.n299 VOUT.n77 3.055
R392 VOUT.n372 VOUT.n78 3.055
R393 VOUT.n593 VOUT.n81 3.055
R394 VOUT.n651 VOUT.n650 2.989
R395 VOUT.n651 VOUT.n637 2.987
R396 VOUT.n651 VOUT.n673 2.979
R397 VOUT.n472 VOUT.n471 2.814
R398 VOUT.n399 VOUT.n398 2.814
R399 VOUT.n179 VOUT.n178 2.814
R400 VOUT.n252 VOUT.n251 2.814
R401 VOUT.n325 VOUT.n324 2.814
R402 VOUT.n539 VOUT.n538 2.814
R403 VOUT.n132 VOUT.n712 2.231
R404 VOUT.n134 VOUT.n751 2.231
R405 VOUT.n133 VOUT.n632 2.231
R406 VOUT.n448 VOUT.n447 2.082
R407 VOUT.n375 VOUT.n374 2.082
R408 VOUT.n155 VOUT.n154 2.082
R409 VOUT.n228 VOUT.n227 2.082
R410 VOUT.n301 VOUT.n300 2.082
R411 VOUT.n522 VOUT.n521 2.082
R412 VOUT.n634 VOUT.n633 1.155
R413 VOUT.n719 VOUT.n718 1.155
R414 VOUT.n600 VOUT.n599 1.155
R415 VOUT.n680 VOUT.n679 1.155
R416 VOUT.n637 VOUT.n634 0.921
R417 VOUT.n601 VOUT.n600 0.921
R418 VOUT.n681 VOUT.n680 0.921
R419 VOUT.n720 VOUT.n719 0.903
R420 VOUT.n497 VOUT.n496 0.536
R421 VOUT.n488 VOUT.n487 0.536
R422 VOUT.n424 VOUT.n423 0.536
R423 VOUT.n415 VOUT.n414 0.536
R424 VOUT.n204 VOUT.n203 0.536
R425 VOUT.n195 VOUT.n194 0.536
R426 VOUT.n277 VOUT.n276 0.536
R427 VOUT.n268 VOUT.n267 0.536
R428 VOUT.n350 VOUT.n349 0.536
R429 VOUT.n341 VOUT.n340 0.536
R430 VOUT.n569 VOUT.n568 0.536
R431 VOUT.n557 VOUT.n556 0.536
R432 VOUT.n715 VOUT.n713 0.506
R433 VOUT.n596 VOUT.n594 0.506
R434 VOUT.n676 VOUT.n674 0.506
R435 VOUT.n640 VOUT.n638 0.506
R436 VOUT.n503 VOUT.n502 0.506
R437 VOUT.n483 VOUT.n482 0.506
R438 VOUT.n430 VOUT.n429 0.506
R439 VOUT.n410 VOUT.n409 0.506
R440 VOUT.n210 VOUT.n209 0.506
R441 VOUT.n190 VOUT.n189 0.506
R442 VOUT.n283 VOUT.n282 0.506
R443 VOUT.n263 VOUT.n262 0.506
R444 VOUT.n356 VOUT.n355 0.506
R445 VOUT.n336 VOUT.n335 0.506
R446 VOUT.n552 VOUT.n551 0.506
R447 VOUT.n575 VOUT.n574 0.506
R448 VOUT.n746 VOUT.n745 0.476
R449 VOUT.n627 VOUT.n626 0.476
R450 VOUT.n707 VOUT.n706 0.476
R451 VOUT.n645 VOUT.n644 0.476
R452 VOUT.n507 VOUT.n506 0.476
R453 VOUT.n477 VOUT.n476 0.476
R454 VOUT.n434 VOUT.n433 0.476
R455 VOUT.n404 VOUT.n403 0.476
R456 VOUT.n214 VOUT.n213 0.476
R457 VOUT.n184 VOUT.n183 0.476
R458 VOUT.n287 VOUT.n286 0.476
R459 VOUT.n257 VOUT.n256 0.476
R460 VOUT.n360 VOUT.n359 0.476
R461 VOUT.n330 VOUT.n329 0.476
R462 VOUT.n545 VOUT.n544 0.476
R463 VOUT.n580 VOUT.n579 0.475
R464 VOUT.n740 VOUT.n739 0.445
R465 VOUT.n621 VOUT.n620 0.445
R466 VOUT.n701 VOUT.n700 0.445
R467 VOUT.n657 VOUT.n656 0.445
R468 VOUT.n734 VOUT.n733 0.414
R469 VOUT.n615 VOUT.n614 0.414
R470 VOUT.n695 VOUT.n694 0.414
R471 VOUT.n662 VOUT.n661 0.414
R472 VOUT.n517 VOUT.n516 0.414
R473 VOUT.n468 VOUT.n467 0.414
R474 VOUT.n444 VOUT.n443 0.414
R475 VOUT.n395 VOUT.n394 0.414
R476 VOUT.n224 VOUT.n223 0.414
R477 VOUT.n175 VOUT.n174 0.414
R478 VOUT.n297 VOUT.n296 0.414
R479 VOUT.n248 VOUT.n247 0.414
R480 VOUT.n370 VOUT.n369 0.414
R481 VOUT.n321 VOUT.n320 0.414
R482 VOUT.n534 VOUT.n533 0.414
R483 VOUT.n591 VOUT.n590 0.413
R484 VOUT.n728 VOUT.n727 0.382
R485 VOUT.n609 VOUT.n608 0.382
R486 VOUT.n689 VOUT.n688 0.382
R487 VOUT.n669 VOUT.n668 0.382
R488 VOUT.n520 VOUT.n519 0.271
R489 VOUT.n373 VOUT.n372 0.271
R490 VOUT.n752 VOUT.n134 0.246
R491 VOUT.n520 VOUT.n446 0.228
R492 VOUT.n58 VOUT.n226 0.228
R493 VOUT.n373 VOUT.n299 0.228
R494 VOUT.n59 VOUT.n593 0.228
R495 VOUT.n752 VOUT.n59 0.19
R496 VOUT.n132 VOUT.n651 0.103
R497 VOUT.n28 VOUT.n0 0.079
R498 VOUT.n587 VOUT.n106 0.079
R499 VOUT.n546 VOUT.n543 0.079
R500 VOUT.n26 VOUT.n537 0.079
R501 VOUT.n532 VOUT.n37 0.079
R502 VOUT.n29 VOUT.n1 0.079
R503 VOUT.n514 VOUT.n108 0.079
R504 VOUT.n478 VOUT.n475 0.079
R505 VOUT.n24 VOUT.n470 0.079
R506 VOUT.n466 VOUT.n41 0.079
R507 VOUT.n30 VOUT.n2 0.079
R508 VOUT.n441 VOUT.n110 0.079
R509 VOUT.n405 VOUT.n402 0.079
R510 VOUT.n22 VOUT.n397 0.079
R511 VOUT.n393 VOUT.n45 0.079
R512 VOUT.n31 VOUT.n3 0.079
R513 VOUT.n221 VOUT.n112 0.079
R514 VOUT.n185 VOUT.n182 0.079
R515 VOUT.n20 VOUT.n177 0.079
R516 VOUT.n173 VOUT.n49 0.079
R517 VOUT.n32 VOUT.n4 0.079
R518 VOUT.n294 VOUT.n114 0.079
R519 VOUT.n258 VOUT.n255 0.079
R520 VOUT.n18 VOUT.n250 0.079
R521 VOUT.n246 VOUT.n53 0.079
R522 VOUT.n33 VOUT.n5 0.079
R523 VOUT.n367 VOUT.n116 0.079
R524 VOUT.n331 VOUT.n328 0.079
R525 VOUT.n16 VOUT.n323 0.079
R526 VOUT.n319 VOUT.n57 0.079
R527 VOUT.n581 VOUT.n142 0.076
R528 VOUT.n508 VOUT.n144 0.076
R529 VOUT.n435 VOUT.n146 0.076
R530 VOUT.n215 VOUT.n148 0.076
R531 VOUT.n288 VOUT.n150 0.076
R532 VOUT.n361 VOUT.n152 0.076
R533 VOUT.n738 VOUT.n85 0.073
R534 VOUT.n619 VOUT.n88 0.073
R535 VOUT.n699 VOUT.n91 0.073
R536 VOUT.n93 VOUT.n658 0.073
R537 VOUT.n75 VOUT.n726 0.073
R538 VOUT.n72 VOUT.n607 0.073
R539 VOUT.n74 VOUT.n687 0.073
R540 VOUT.n73 VOUT.n667 0.073
R541 VOUT.n613 VOUT.n612 0.072
R542 VOUT.n650 VOUT.n12 0.072
R543 VOUT.n732 VOUT.n731 0.072
R544 VOUT.n693 VOUT.n692 0.072
R545 VOUT.n673 VOUT.n672 0.072
R546 VOUT.n744 VOUT.n120 0.068
R547 VOUT.n625 VOUT.n122 0.068
R548 VOUT.n705 VOUT.n125 0.068
R549 VOUT.n643 VOUT.n642 0.068
R550 VOUT.n82 VOUT.n550 0.064
R551 VOUT.n96 VOUT.n481 0.064
R552 VOUT.n98 VOUT.n408 0.064
R553 VOUT.n100 VOUT.n188 0.064
R554 VOUT.n102 VOUT.n261 0.064
R555 VOUT.n104 VOUT.n334 0.064
R556 VOUT.n143 VOUT.n61 0.126
R557 VOUT.n145 VOUT.n63 0.126
R558 VOUT.n147 VOUT.n65 0.126
R559 VOUT.n149 VOUT.n67 0.126
R560 VOUT.n151 VOUT.n69 0.126
R561 VOUT.n153 VOUT.n71 0.126
R562 VOUT.n673 VOUT.n94 0.057
R563 VOUT.n84 VOUT.n732 0.057
R564 VOUT.n90 VOUT.n693 0.057
R565 VOUT.n87 VOUT.n613 0.057
R566 VOUT.n726 VOUT.n724 0.054
R567 VOUT.n607 VOUT.n605 0.054
R568 VOUT.n687 VOUT.n685 0.054
R569 VOUT.n667 VOUT.n665 0.054
R570 VOUT.n712 VOUT.n677 0.054
R571 VOUT.n751 VOUT.n716 0.054
R572 VOUT.n632 VOUT.n597 0.054
R573 VOUT.n632 VOUT.n14 0.054
R574 VOUT.n751 VOUT.n15 0.054
R575 VOUT.n712 VOUT.n13 0.054
R576 VOUT.n86 VOUT.n720 0.053
R577 VOUT VOUT.n752 0.053
R578 VOUT.n565 VOUT.n562 0.106
R579 VOUT.n493 VOUT.n492 0.106
R580 VOUT.n420 VOUT.n419 0.106
R581 VOUT.n200 VOUT.n199 0.106
R582 VOUT.n273 VOUT.n272 0.106
R583 VOUT.n346 VOUT.n345 0.106
R584 VOUT.n558 VOUT.n83 0.112
R585 VOUT.n489 VOUT.n97 0.112
R586 VOUT.n416 VOUT.n99 0.112
R587 VOUT.n196 VOUT.n101 0.112
R588 VOUT.n269 VOUT.n103 0.112
R589 VOUT.n342 VOUT.n105 0.112
R590 VOUT.n138 VOUT.n744 0.048
R591 VOUT.n139 VOUT.n625 0.048
R592 VOUT.n140 VOUT.n705 0.048
R593 VOUT.n141 VOUT.n643 0.048
R594 VOUT.n60 VOUT.n570 0.109
R595 VOUT.n62 VOUT.n498 0.109
R596 VOUT.n64 VOUT.n425 0.109
R597 VOUT.n66 VOUT.n205 0.109
R598 VOUT.n68 VOUT.n278 0.109
R599 VOUT.n70 VOUT.n351 0.109
R600 VOUT.n133 VOUT.n132 0.109
R601 VOUT.n134 VOUT.n133 0.103
R602 VOUT.n5 VOUT.n54 0.066
R603 VOUT.n4 VOUT.n50 0.066
R604 VOUT.n3 VOUT.n46 0.066
R605 VOUT.n2 VOUT.n42 0.066
R606 VOUT.n1 VOUT.n38 0.066
R607 VOUT.n0 VOUT.n34 0.066
R608 VOUT.n11 VOUT.n581 0.062
R609 VOUT.n10 VOUT.n508 0.062
R610 VOUT.n9 VOUT.n435 0.062
R611 VOUT.n8 VOUT.n215 0.062
R612 VOUT.n7 VOUT.n288 0.062
R613 VOUT.n6 VOUT.n361 0.062
R614 VOUT.n78 VOUT.n33 0.061
R615 VOUT.n77 VOUT.n32 0.061
R616 VOUT.n76 VOUT.n31 0.061
R617 VOUT.n79 VOUT.n30 0.061
R618 VOUT.n80 VOUT.n29 0.061
R619 VOUT.n81 VOUT.n28 0.061
R620 VOUT.n543 VOUT.n27 0.061
R621 VOUT.n475 VOUT.n25 0.061
R622 VOUT.n402 VOUT.n23 0.061
R623 VOUT.n182 VOUT.n21 0.061
R624 VOUT.n255 VOUT.n19 0.061
R625 VOUT.n328 VOUT.n17 0.061
R626 VOUT.n57 VOUT.n56 0.059
R627 VOUT.n53 VOUT.n52 0.059
R628 VOUT.n49 VOUT.n48 0.059
R629 VOUT.n45 VOUT.n44 0.059
R630 VOUT.n41 VOUT.n40 0.059
R631 VOUT.n37 VOUT.n36 0.059
R632 VOUT.n15 VOUT.n138 0.058
R633 VOUT.n14 VOUT.n139 0.058
R634 VOUT.n13 VOUT.n140 0.058
R635 VOUT.n12 VOUT.n141 0.058
R636 VOUT.n71 VOUT.n70 0.056
R637 VOUT.n69 VOUT.n68 0.056
R638 VOUT.n67 VOUT.n66 0.056
R639 VOUT.n65 VOUT.n64 0.056
R640 VOUT.n63 VOUT.n62 0.056
R641 VOUT.n61 VOUT.n60 0.056
R642 VOUT.n105 VOUT.n104 0.054
R643 VOUT.n103 VOUT.n102 0.054
R644 VOUT.n101 VOUT.n100 0.054
R645 VOUT.n99 VOUT.n98 0.054
R646 VOUT.n97 VOUT.n96 0.054
R647 VOUT.n94 VOUT.n93 0.054
R648 VOUT.n91 VOUT.n90 0.054
R649 VOUT.n88 VOUT.n87 0.054
R650 VOUT.n716 VOUT.n86 0.054
R651 VOUT.n85 VOUT.n84 0.054
R652 VOUT.n83 VOUT.n82 0.054
R653 VOUT.n637 VOUT.n95 0.05
R654 VOUT.n92 VOUT.n681 0.05
R655 VOUT.n89 VOUT.n601 0.05
R656 VOUT.n124 VOUT.n699 0.048
R657 VOUT.n121 VOUT.n619 0.048
R658 VOUT.n119 VOUT.n738 0.048
R659 VOUT.n36 VOUT.n528 0.043
R660 VOUT.n40 VOUT.n463 0.043
R661 VOUT.n44 VOUT.n390 0.043
R662 VOUT.n48 VOUT.n170 0.043
R663 VOUT.n52 VOUT.n243 0.043
R664 VOUT.n56 VOUT.n316 0.043
R665 VOUT.n58 VOUT.n373 0.043
R666 VOUT.n59 VOUT.n520 0.043
R667 VOUT.n59 VOUT.n58 0.042
R668 VOUT.n731 VOUT.n75 0.041
R669 VOUT.n692 VOUT.n74 0.041
R670 VOUT.n672 VOUT.n73 0.041
R671 VOUT.n612 VOUT.n72 0.041
R672 VOUT.n597 VOUT.n89 0.04
R673 VOUT.n677 VOUT.n92 0.04
R674 VOUT.n81 VOUT.n523 0.04
R675 VOUT.n548 VOUT.n546 0.04
R676 VOUT.n80 VOUT.n449 0.04
R677 VOUT.n479 VOUT.n478 0.04
R678 VOUT.n79 VOUT.n376 0.04
R679 VOUT.n406 VOUT.n405 0.04
R680 VOUT.n76 VOUT.n156 0.04
R681 VOUT.n186 VOUT.n185 0.04
R682 VOUT.n77 VOUT.n229 0.04
R683 VOUT.n259 VOUT.n258 0.04
R684 VOUT.n78 VOUT.n302 0.04
R685 VOUT.n332 VOUT.n331 0.04
R686 VOUT.n152 VOUT.n153 0.04
R687 VOUT.n150 VOUT.n151 0.04
R688 VOUT.n148 VOUT.n149 0.04
R689 VOUT.n146 VOUT.n147 0.04
R690 VOUT.n144 VOUT.n145 0.04
R691 VOUT.n142 VOUT.n143 0.04
R692 VOUT.n351 VOUT.n131 0.04
R693 VOUT.n278 VOUT.n130 0.04
R694 VOUT.n205 VOUT.n129 0.04
R695 VOUT.n425 VOUT.n128 0.04
R696 VOUT.n498 VOUT.n127 0.04
R697 VOUT.n126 VOUT.n655 0.04
R698 VOUT.n125 VOUT.n124 0.04
R699 VOUT.n685 VOUT.n123 0.04
R700 VOUT.n122 VOUT.n121 0.04
R701 VOUT.n120 VOUT.n119 0.04
R702 VOUT.n570 VOUT.n118 0.04
R703 VOUT.n345 VOUT.n117 0.04
R704 VOUT.n116 VOUT.n6 0.04
R705 VOUT.n272 VOUT.n115 0.04
R706 VOUT.n114 VOUT.n7 0.04
R707 VOUT.n199 VOUT.n113 0.04
R708 VOUT.n112 VOUT.n8 0.04
R709 VOUT.n419 VOUT.n111 0.04
R710 VOUT.n110 VOUT.n9 0.04
R711 VOUT.n492 VOUT.n109 0.04
R712 VOUT.n108 VOUT.n10 0.04
R713 VOUT.n562 VOUT.n107 0.04
R714 VOUT.n106 VOUT.n11 0.04
R715 VOUT.n17 VOUT.n16 0.04
R716 VOUT.n19 VOUT.n18 0.04
R717 VOUT.n21 VOUT.n20 0.04
R718 VOUT.n23 VOUT.n22 0.04
R719 VOUT.n25 VOUT.n24 0.04
R720 VOUT.n27 VOUT.n26 0.04
R721 VOUT.n312 VOUT.n55 0.04
R722 VOUT.n239 VOUT.n51 0.04
R723 VOUT.n166 VOUT.n47 0.04
R724 VOUT.n386 VOUT.n43 0.04
R725 VOUT.n459 VOUT.n39 0.04
R726 VOUT.n526 VOUT.n35 0.04
R727 VOUT.n658 VOUT.n126 0.039
R728 VOUT.n34 VOUT.n587 0.036
R729 VOUT.n38 VOUT.n514 0.036
R730 VOUT.n42 VOUT.n441 0.036
R731 VOUT.n46 VOUT.n221 0.036
R732 VOUT.n50 VOUT.n294 0.036
R733 VOUT.n54 VOUT.n367 0.036
R734 VOUT.n665 VOUT.n137 0.036
R735 VOUT.n605 VOUT.n136 0.036
R736 VOUT.n724 VOUT.n135 0.036
R737 VOUT.n549 VOUT.n548 0.033
R738 VOUT.n537 VOUT.n526 0.033
R739 VOUT.n480 VOUT.n479 0.033
R740 VOUT.n470 VOUT.n459 0.033
R741 VOUT.n407 VOUT.n406 0.033
R742 VOUT.n397 VOUT.n386 0.033
R743 VOUT.n187 VOUT.n186 0.033
R744 VOUT.n177 VOUT.n166 0.033
R745 VOUT.n260 VOUT.n259 0.033
R746 VOUT.n250 VOUT.n239 0.033
R747 VOUT.n333 VOUT.n332 0.033
R748 VOUT.n323 VOUT.n312 0.033
R749 VOUT.n118 VOUT.n565 0.031
R750 VOUT.n127 VOUT.n493 0.031
R751 VOUT.n128 VOUT.n420 0.031
R752 VOUT.n129 VOUT.n200 0.031
R753 VOUT.n130 VOUT.n273 0.031
R754 VOUT.n131 VOUT.n346 0.031
R755 VOUT.n107 VOUT.n558 0.028
R756 VOUT.n550 VOUT.n549 0.028
R757 VOUT.n35 VOUT.n532 0.028
R758 VOUT.n109 VOUT.n489 0.028
R759 VOUT.n481 VOUT.n480 0.028
R760 VOUT.n39 VOUT.n466 0.028
R761 VOUT.n111 VOUT.n416 0.028
R762 VOUT.n408 VOUT.n407 0.028
R763 VOUT.n43 VOUT.n393 0.028
R764 VOUT.n113 VOUT.n196 0.028
R765 VOUT.n188 VOUT.n187 0.028
R766 VOUT.n47 VOUT.n173 0.028
R767 VOUT.n115 VOUT.n269 0.028
R768 VOUT.n261 VOUT.n260 0.028
R769 VOUT.n51 VOUT.n246 0.028
R770 VOUT.n117 VOUT.n342 0.028
R771 VOUT.n334 VOUT.n333 0.028
R772 VOUT.n55 VOUT.n319 0.028
R773 S1.n3 S1.t10 5.393
R774 S1.n8 S1.t3 5.393
R775 S1.n7 S1.t6 3.326
R776 S1.n7 S1.t0 3.326
R777 S1.n6 S1.t2 3.326
R778 S1.n6 S1.t5 3.326
R779 S1.n0 S1.t7 3.326
R780 S1.n0 S1.t9 3.326
R781 S1.n1 S1.t4 3.326
R782 S1.n1 S1.t8 3.326
R783 S1.n2 S1.t1 3.326
R784 S1.n2 S1.t11 3.326
R785 S1.n8 S1.n7 1.79
R786 S1.n9 S1.n6 1.79
R787 S1.n5 S1.n0 1.79
R788 S1.n4 S1.n1 1.79
R789 S1.n3 S1.n2 1.79
R790 S1.n9 S1.n8 0.307
R791 S1.n5 S1.n4 0.307
R792 S1.n4 S1.n3 0.307
R793 S1.n10 S1.n9 0.296
R794 S1 S1.n10 0.085
R795 S1.n10 S1.n5 0.011
R796 D1.n2 D1.t0 5.416
R797 D1.n5 D1.t1 5.414
R798 D1.n4 D1.t5 3.326
R799 D1.n4 D1.t2 3.326
R800 D1.n3 D1.t3 3.326
R801 D1.n3 D1.t6 3.326
R802 D1.n1 D1.t7 3.326
R803 D1.n1 D1.t4 3.326
R804 D1.n5 D1.n4 1.766
R805 D1.n0 D1.n3 1.766
R806 D1.n2 D1.n1 1.766
R807 D1.n0 D1.n5 0.352
R808 D1.n0 D1.n2 0.35
R809 D1 D1.n0 0.261
R810 SS.n32 SS.n31 9.3
R811 SS.n52 SS.n51 9.3
R812 SS.n74 SS.n73 9.3
R813 SS.n3 SS.n14 9.3
R814 SS.n18 SS.n17 9.3
R815 SS.n23 SS.n22 9.3
R816 SS.n28 SS.n27 9.3
R817 SS.n34 SS.n33 9.3
R818 SS.n38 SS.n37 9.3
R819 SS.n50 SS.n49 9.3
R820 SS.n54 SS.n53 9.3
R821 SS.n61 SS.n60 9.3
R822 SS.n63 SS.n62 9.3
R823 SS.n65 SS.n64 9.3
R824 SS.n88 SS.n87 9.3
R825 SS.n5 SS.n93 9.3
R826 SS.n103 SS.n102 9.3
R827 SS.n106 SS.n105 9.3
R828 SS.n109 SS.n108 9.3
R829 SS.n125 SS.n124 9.3
R830 SS.n119 SS.n118 9.3
R831 SS.n115 SS.n114 9.3
R832 SS.n99 SS.n98 9.3
R833 SS.n5 SS.n95 9.3
R834 SS.n4 SS.n92 9.3
R835 SS.n85 SS.n84 9.3
R836 SS.n83 SS.n82 9.3
R837 SS.n77 SS.n76 9.3
R838 SS.n72 SS.n71 9.3
R839 SS.n385 SS.n384 9.3
R840 SS.n405 SS.n404 9.3
R841 SS.n427 SS.n426 9.3
R842 SS.n6 SS.n367 9.3
R843 SS.n371 SS.n370 9.3
R844 SS.n376 SS.n375 9.3
R845 SS.n381 SS.n380 9.3
R846 SS.n387 SS.n386 9.3
R847 SS.n391 SS.n390 9.3
R848 SS.n403 SS.n402 9.3
R849 SS.n407 SS.n406 9.3
R850 SS.n414 SS.n413 9.3
R851 SS.n416 SS.n415 9.3
R852 SS.n418 SS.n417 9.3
R853 SS.n441 SS.n440 9.3
R854 SS.n8 SS.n446 9.3
R855 SS.n456 SS.n455 9.3
R856 SS.n459 SS.n458 9.3
R857 SS.n462 SS.n461 9.3
R858 SS.n478 SS.n477 9.3
R859 SS.n472 SS.n471 9.3
R860 SS.n468 SS.n467 9.3
R861 SS.n452 SS.n451 9.3
R862 SS.n8 SS.n448 9.3
R863 SS.n7 SS.n445 9.3
R864 SS.n438 SS.n437 9.3
R865 SS.n436 SS.n435 9.3
R866 SS.n430 SS.n429 9.3
R867 SS.n425 SS.n424 9.3
R868 SS.n268 SS.n267 9.3
R869 SS.n288 SS.n287 9.3
R870 SS.n310 SS.n309 9.3
R871 SS.n301 SS.n300 9.3
R872 SS.n299 SS.n298 9.3
R873 SS.n297 SS.n296 9.3
R874 SS.n290 SS.n289 9.3
R875 SS.n286 SS.n285 9.3
R876 SS.n274 SS.n273 9.3
R877 SS.n270 SS.n269 9.3
R878 SS.n264 SS.n263 9.3
R879 SS.n259 SS.n258 9.3
R880 SS.n254 SS.n253 9.3
R881 SS.n9 SS.n250 9.3
R882 SS.n342 SS.n341 9.3
R883 SS.n11 SS.n329 9.3
R884 SS.n319 SS.n318 9.3
R885 SS.n321 SS.n320 9.3
R886 SS.n324 SS.n323 9.3
R887 SS.n361 SS.n360 9.3
R888 SS.n355 SS.n354 9.3
R889 SS.n351 SS.n350 9.3
R890 SS.n345 SS.n344 9.3
R891 SS.n339 SS.n338 9.3
R892 SS.n335 SS.n334 9.3
R893 SS.n11 SS.n331 9.3
R894 SS.n10 SS.n328 9.3
R895 SS.n313 SS.n312 9.3
R896 SS.n308 SS.n307 9.3
R897 SS.n149 SS.n148 9.3
R898 SS.n169 SS.n168 9.3
R899 SS.n191 SS.n190 9.3
R900 SS.n135 SS.n134 9.3
R901 SS.n145 SS.n144 9.3
R902 SS.n155 SS.n154 9.3
R903 SS.n171 SS.n170 9.3
R904 SS.n180 SS.n179 9.3
R905 SS.n182 SS.n181 9.3
R906 SS.n2 SS.n210 9.3
R907 SS.n223 SS.n222 9.3
R908 SS.n226 SS.n225 9.3
R909 SS.n236 SS.n235 9.3
R910 SS.n216 SS.n215 9.3
R911 SS.n1 SS.n209 9.3
R912 SS.n202 SS.n201 9.3
R913 SS.n200 SS.n199 9.3
R914 SS.n189 SS.n188 9.3
R915 SS.n0 SS.n131 9.3
R916 SS.n140 SS.n139 9.3
R917 SS.n151 SS.n150 9.3
R918 SS.n167 SS.n166 9.3
R919 SS.n178 SS.n177 9.3
R920 SS.n205 SS.n204 9.3
R921 SS.n220 SS.n219 9.3
R922 SS.n242 SS.n241 9.3
R923 SS.n232 SS.n231 9.3
R924 SS.n2 SS.n212 9.3
R925 SS.n194 SS.n193 9.3
R926 SS.n127 SS.n120 9
R927 SS.n16 SS.n15 9
R928 SS.n25 SS.n24 9
R929 SS.n36 SS.n35 9
R930 SS.n56 SS.n55 9
R931 SS.n67 SS.n66 9
R932 SS.n81 SS.n80 9
R933 SS.n112 SS.n111 9
R934 SS.n101 SS.n100 9
R935 SS.n4 SS.n91 9
R936 SS.n70 SS.n69 9
R937 SS.n480 SS.n473 9
R938 SS.n369 SS.n368 9
R939 SS.n378 SS.n377 9
R940 SS.n389 SS.n388 9
R941 SS.n409 SS.n408 9
R942 SS.n420 SS.n419 9
R943 SS.n434 SS.n433 9
R944 SS.n465 SS.n464 9
R945 SS.n454 SS.n453 9
R946 SS.n7 SS.n444 9
R947 SS.n423 SS.n422 9
R948 SS.n252 SS.n251 9
R949 SS.n261 SS.n260 9
R950 SS.n272 SS.n271 9
R951 SS.n292 SS.n291 9
R952 SS.n303 SS.n302 9
R953 SS.n363 SS.n356 9
R954 SS.n348 SS.n347 9
R955 SS.n337 SS.n336 9
R956 SS.n317 SS.n316 9
R957 SS.n10 SS.n327 9
R958 SS.n306 SS.n305 9
R959 SS.n244 SS.n237 9
R960 SS.n133 SS.n132 9
R961 SS.n142 SS.n141 9
R962 SS.n153 SS.n152 9
R963 SS.n173 SS.n172 9
R964 SS.n184 SS.n183 9
R965 SS.n198 SS.n197 9
R966 SS.n229 SS.n228 9
R967 SS.n218 SS.n217 9
R968 SS.n1 SS.n208 9
R969 SS.n187 SS.n186 9
R970 SS.n69 SS.n68 8.282
R971 SS.n422 SS.n421 8.282
R972 SS.n305 SS.n304 8.282
R973 SS.n186 SS.n185 8.282
R974 SS.n123 SS.n122 7.853
R975 SS.n476 SS.n475 7.853
R976 SS.n359 SS.n358 7.853
R977 SS.n240 SS.n239 7.853
R978 SS.n130 SS.n129 7.852
R979 SS.n13 SS.n12 7.851
R980 SS.n366 SS.n365 7.851
R981 SS.n249 SS.n248 7.851
R982 SS.n43 SS.n42 4.65
R983 SS.n396 SS.n395 4.65
R984 SS.n279 SS.n278 4.65
R985 SS.n160 SS.n159 4.65
R986 SS.n45 SS.n44 4.574
R987 SS.n398 SS.n397 4.574
R988 SS.n281 SS.n280 4.574
R989 SS.n162 SS.n161 4.574
R990 SS.n121 SS.t5 3.326
R991 SS.n121 SS.t0 3.326
R992 SS.n474 SS.t1 3.326
R993 SS.n474 SS.t3 3.326
R994 SS.n357 SS.t4 3.326
R995 SS.n357 SS.t7 3.326
R996 SS.n238 SS.t2 3.326
R997 SS.n238 SS.t6 3.326
R998 SS.n105 SS.n104 3.191
R999 SS.n458 SS.n457 3.191
R1000 SS.n341 SS.n340 3.191
R1001 SS.n222 SS.n221 3.191
R1002 SS.n31 SS.n30 2.814
R1003 SS.n384 SS.n383 2.814
R1004 SS.n267 SS.n266 2.814
R1005 SS.n148 SS.n147 2.814
R1006 SS.n122 SS.n121 2.082
R1007 SS.n475 SS.n474 2.082
R1008 SS.n358 SS.n357 2.082
R1009 SS.n239 SS.n238 2.082
R1010 SS.n484 SS.n247 0.777
R1011 SS.n484 SS.n483 0.751
R1012 SS.n60 SS.n59 0.536
R1013 SS.n76 SS.n75 0.536
R1014 SS.n413 SS.n412 0.536
R1015 SS.n429 SS.n428 0.536
R1016 SS.n296 SS.n295 0.536
R1017 SS.n312 SS.n311 0.536
R1018 SS.n193 SS.n192 0.536
R1019 SS.n177 SS.n176 0.536
R1020 SS.n49 SS.n48 0.506
R1021 SS.n87 SS.n86 0.506
R1022 SS.n402 SS.n401 0.506
R1023 SS.n440 SS.n439 0.506
R1024 SS.n285 SS.n284 0.506
R1025 SS.n323 SS.n322 0.506
R1026 SS.n204 SS.n203 0.506
R1027 SS.n166 SS.n165 0.506
R1028 SS.n42 SS.n41 0.476
R1029 SS.n95 SS.n94 0.476
R1030 SS.n395 SS.n394 0.476
R1031 SS.n448 SS.n447 0.476
R1032 SS.n278 SS.n277 0.476
R1033 SS.n331 SS.n330 0.476
R1034 SS.n212 SS.n211 0.476
R1035 SS.n159 SS.n158 0.475
R1036 SS.n22 SS.n21 0.414
R1037 SS.n114 SS.n113 0.414
R1038 SS.n375 SS.n374 0.414
R1039 SS.n467 SS.n466 0.414
R1040 SS.n258 SS.n257 0.414
R1041 SS.n350 SS.n349 0.414
R1042 SS.n231 SS.n230 0.414
R1043 SS.n139 SS.n138 0.413
R1044 SS.n247 SS.n128 0.18
R1045 SS.n482 SS.n481 0.18
R1046 SS.n483 SS.n364 0.18
R1047 SS.n246 SS.n245 0.18
R1048 SS.n137 SS.n136 0.079
R1049 SS.n149 SS.n146 0.079
R1050 SS.n160 SS.n157 0.079
R1051 SS.n224 SS.n223 0.079
R1052 SS.n234 SS.n233 0.079
R1053 SS.n20 SS.n19 0.079
R1054 SS.n32 SS.n29 0.079
R1055 SS.n43 SS.n40 0.079
R1056 SS.n107 SS.n106 0.079
R1057 SS.n117 SS.n116 0.079
R1058 SS.n373 SS.n372 0.079
R1059 SS.n385 SS.n382 0.079
R1060 SS.n396 SS.n393 0.079
R1061 SS.n460 SS.n459 0.079
R1062 SS.n470 SS.n469 0.079
R1063 SS.n256 SS.n255 0.079
R1064 SS.n268 SS.n265 0.079
R1065 SS.n279 SS.n276 0.079
R1066 SS.n343 SS.n342 0.079
R1067 SS.n353 SS.n352 0.079
R1068 SS.n213 SS.n2 0.076
R1069 SS.n96 SS.n5 0.076
R1070 SS.n449 SS.n8 0.076
R1071 SS.n332 SS.n11 0.076
R1072 SS.n247 SS.n246 0.071
R1073 SS.n483 SS.n482 0.071
R1074 SS.n167 SS.n164 0.064
R1075 SS.n50 SS.n47 0.064
R1076 SS.n403 SS.n400 0.064
R1077 SS.n286 SS.n283 0.064
R1078 SS.n206 SS.n205 0.062
R1079 SS.n89 SS.n88 0.062
R1080 SS.n442 SS.n441 0.062
R1081 SS.n325 SS.n324 0.062
R1082 SS.n187 SS.n184 0.106
R1083 SS.n70 SS.n67 0.106
R1084 SS.n423 SS.n420 0.106
R1085 SS.n306 SS.n303 0.106
R1086 SS.n178 SS.n175 0.05
R1087 SS.n61 SS.n58 0.05
R1088 SS.n414 SS.n411 0.05
R1089 SS.n297 SS.n294 0.05
R1090 SS.n195 SS.n194 0.048
R1091 SS.n78 SS.n77 0.048
R1092 SS.n431 SS.n430 0.048
R1093 SS.n314 SS.n313 0.048
R1094 SS.n198 SS.n196 0.045
R1095 SS.n81 SS.n79 0.045
R1096 SS.n434 SS.n432 0.045
R1097 SS.n317 SS.n315 0.045
R1098 SS.n0 SS.n130 0.043
R1099 SS.n174 SS.n173 0.043
R1100 SS.n3 SS.n13 0.043
R1101 SS.n57 SS.n56 0.043
R1102 SS.n6 SS.n366 0.043
R1103 SS.n410 SS.n409 0.043
R1104 SS.n9 SS.n249 0.043
R1105 SS.n293 SS.n292 0.043
R1106 SS.n162 SS.n160 0.04
R1107 SS.n242 SS.n240 0.04
R1108 SS.n45 SS.n43 0.04
R1109 SS.n125 SS.n123 0.04
R1110 SS.n398 SS.n396 0.04
R1111 SS.n478 SS.n476 0.04
R1112 SS.n281 SS.n279 0.04
R1113 SS.n361 SS.n359 0.04
R1114 SS.n157 SS.n156 0.038
R1115 SS.n40 SS.n39 0.038
R1116 SS.n393 SS.n392 0.038
R1117 SS.n276 SS.n275 0.038
R1118 SS.n214 SS.n213 0.036
R1119 SS.n226 SS.n224 0.036
R1120 SS.n97 SS.n96 0.036
R1121 SS.n109 SS.n107 0.036
R1122 SS.n450 SS.n449 0.036
R1123 SS.n462 SS.n460 0.036
R1124 SS.n333 SS.n332 0.036
R1125 SS.n345 SS.n343 0.036
R1126 SS.n146 SS.n145 0.033
R1127 SS.n163 SS.n162 0.033
R1128 SS.n29 SS.n28 0.033
R1129 SS.n46 SS.n45 0.033
R1130 SS.n382 SS.n381 0.033
R1131 SS.n399 SS.n398 0.033
R1132 SS.n265 SS.n264 0.033
R1133 SS.n282 SS.n281 0.033
R1134 SS.n189 SS.n187 0.031
R1135 SS.n194 SS.n191 0.031
R1136 SS.n72 SS.n70 0.031
R1137 SS.n77 SS.n74 0.031
R1138 SS.n425 SS.n423 0.031
R1139 SS.n430 SS.n427 0.031
R1140 SS.n308 SS.n306 0.031
R1141 SS.n313 SS.n310 0.031
R1142 SS.n140 SS.n137 0.028
R1143 SS.n164 SS.n163 0.028
R1144 SS.n180 SS.n178 0.028
R1145 SS.n184 SS.n182 0.028
R1146 SS.n220 SS.n218 0.028
R1147 SS.n23 SS.n20 0.028
R1148 SS.n47 SS.n46 0.028
R1149 SS.n63 SS.n61 0.028
R1150 SS.n67 SS.n65 0.028
R1151 SS.n103 SS.n101 0.028
R1152 SS.n376 SS.n373 0.028
R1153 SS.n400 SS.n399 0.028
R1154 SS.n416 SS.n414 0.028
R1155 SS.n420 SS.n418 0.028
R1156 SS.n456 SS.n454 0.028
R1157 SS.n259 SS.n256 0.028
R1158 SS.n283 SS.n282 0.028
R1159 SS.n299 SS.n297 0.028
R1160 SS.n303 SS.n301 0.028
R1161 SS.n339 SS.n337 0.028
R1162 SS.n135 SS.n133 0.026
R1163 SS.n153 SS.n151 0.026
R1164 SS.n171 SS.n169 0.026
R1165 SS.n207 SS.n206 0.026
R1166 SS.n233 SS.n232 0.026
R1167 SS.n244 SS.n236 0.026
R1168 SS SS.n484 0.026
R1169 SS.n18 SS.n16 0.026
R1170 SS.n36 SS.n34 0.026
R1171 SS.n54 SS.n52 0.026
R1172 SS.n90 SS.n89 0.026
R1173 SS.n116 SS.n115 0.026
R1174 SS.n127 SS.n119 0.026
R1175 SS.n371 SS.n369 0.026
R1176 SS.n389 SS.n387 0.026
R1177 SS.n407 SS.n405 0.026
R1178 SS.n443 SS.n442 0.026
R1179 SS.n469 SS.n468 0.026
R1180 SS.n480 SS.n472 0.026
R1181 SS.n254 SS.n252 0.026
R1182 SS.n272 SS.n270 0.026
R1183 SS.n290 SS.n288 0.026
R1184 SS.n326 SS.n325 0.026
R1185 SS.n352 SS.n351 0.026
R1186 SS.n363 SS.n355 0.026
R1187 SS.n202 SS.n200 0.024
R1188 SS.n85 SS.n83 0.024
R1189 SS.n438 SS.n436 0.024
R1190 SS.n321 SS.n319 0.024
R1191 SS.n236 SS.n234 0.021
R1192 SS.n119 SS.n117 0.021
R1193 SS.n472 SS.n470 0.021
R1194 SS.n355 SS.n353 0.021
R1195 SS.n136 SS.n135 0.019
R1196 SS.n142 SS.n140 0.019
R1197 SS.n175 SS.n174 0.019
R1198 SS.n232 SS.n229 0.019
R1199 SS.n19 SS.n18 0.019
R1200 SS.n25 SS.n23 0.019
R1201 SS.n58 SS.n57 0.019
R1202 SS.n115 SS.n112 0.019
R1203 SS.n372 SS.n371 0.019
R1204 SS.n378 SS.n376 0.019
R1205 SS.n411 SS.n410 0.019
R1206 SS.n468 SS.n465 0.019
R1207 SS.n255 SS.n254 0.019
R1208 SS.n261 SS.n259 0.019
R1209 SS.n294 SS.n293 0.019
R1210 SS.n351 SS.n348 0.019
R1211 SS.n196 SS.n195 0.016
R1212 SS.n200 SS.n198 0.016
R1213 SS.n205 SS.n202 0.016
R1214 SS.n79 SS.n78 0.016
R1215 SS.n83 SS.n81 0.016
R1216 SS.n88 SS.n85 0.016
R1217 SS.n432 SS.n431 0.016
R1218 SS.n436 SS.n434 0.016
R1219 SS.n441 SS.n438 0.016
R1220 SS.n315 SS.n314 0.016
R1221 SS.n319 SS.n317 0.016
R1222 SS.n324 SS.n321 0.016
R1223 SS.n145 SS.n143 0.014
R1224 SS.n151 SS.n149 0.014
R1225 SS.n155 SS.n153 0.014
R1226 SS.n169 SS.n167 0.014
R1227 SS.n173 SS.n171 0.014
R1228 SS.n216 SS.n214 0.014
R1229 SS.n28 SS.n26 0.014
R1230 SS.n34 SS.n32 0.014
R1231 SS.n38 SS.n36 0.014
R1232 SS.n52 SS.n50 0.014
R1233 SS.n56 SS.n54 0.014
R1234 SS.n99 SS.n97 0.014
R1235 SS.n381 SS.n379 0.014
R1236 SS.n387 SS.n385 0.014
R1237 SS.n391 SS.n389 0.014
R1238 SS.n405 SS.n403 0.014
R1239 SS.n409 SS.n407 0.014
R1240 SS.n452 SS.n450 0.014
R1241 SS.n264 SS.n262 0.014
R1242 SS.n270 SS.n268 0.014
R1243 SS.n274 SS.n272 0.014
R1244 SS.n288 SS.n286 0.014
R1245 SS.n292 SS.n290 0.014
R1246 SS.n335 SS.n333 0.014
R1247 SS.n182 SS.n180 0.012
R1248 SS.n218 SS.n216 0.012
R1249 SS.n223 SS.n220 0.012
R1250 SS.n229 SS.n227 0.012
R1251 SS.n65 SS.n63 0.012
R1252 SS.n101 SS.n99 0.012
R1253 SS.n106 SS.n103 0.012
R1254 SS.n112 SS.n110 0.012
R1255 SS.n418 SS.n416 0.012
R1256 SS.n454 SS.n452 0.012
R1257 SS.n459 SS.n456 0.012
R1258 SS.n465 SS.n463 0.012
R1259 SS.n301 SS.n299 0.012
R1260 SS.n337 SS.n335 0.012
R1261 SS.n342 SS.n339 0.012
R1262 SS.n348 SS.n346 0.012
R1263 SS.n156 SS.n155 0.009
R1264 SS.n191 SS.n189 0.009
R1265 SS.n227 SS.n226 0.009
R1266 SS.n39 SS.n38 0.009
R1267 SS.n74 SS.n72 0.009
R1268 SS.n110 SS.n109 0.009
R1269 SS.n392 SS.n391 0.009
R1270 SS.n427 SS.n425 0.009
R1271 SS.n463 SS.n462 0.009
R1272 SS.n275 SS.n274 0.009
R1273 SS.n310 SS.n308 0.009
R1274 SS.n346 SS.n345 0.009
R1275 SS.n143 SS.n142 0.007
R1276 SS.n244 SS.n243 0.007
R1277 SS.n243 SS.n242 0.007
R1278 SS.n26 SS.n25 0.007
R1279 SS.n127 SS.n126 0.007
R1280 SS.n126 SS.n125 0.007
R1281 SS.n128 SS.n127 3.055
R1282 SS.n379 SS.n378 0.007
R1283 SS.n480 SS.n479 0.007
R1284 SS.n479 SS.n478 0.007
R1285 SS.n481 SS.n480 3.055
R1286 SS.n262 SS.n261 0.007
R1287 SS.n363 SS.n362 0.007
R1288 SS.n362 SS.n361 0.007
R1289 SS.n364 SS.n363 3.055
R1290 SS.n245 SS.n244 3.055
R1291 SS.n11 SS.n10 0.04
R1292 SS.n8 SS.n7 0.04
R1293 SS.n5 SS.n4 0.04
R1294 SS.n2 SS.n1 0.04
R1295 SS.n10 SS.n326 0.038
R1296 SS.n7 SS.n443 0.038
R1297 SS.n4 SS.n90 0.038
R1298 SS.n1 SS.n207 0.038
R1299 SS.n252 SS.n9 0.014
R1300 SS.n369 SS.n6 0.014
R1301 SS.n16 SS.n3 0.014
R1302 SS.n133 SS.n0 0.014
R1303 a_n6328_16092.n12 a_n6328_16092.n74 9.3
R1304 a_n6328_16092.n13 a_n6328_16092.n80 9.3
R1305 a_n6328_16092.n5 a_n6328_16092.n82 9.3
R1306 a_n6328_16092.n5 a_n6328_16092.n83 9.3
R1307 a_n6328_16092.n6 a_n6328_16092.n87 9.3
R1308 a_n6328_16092.n12 a_n6328_16092.n75 9.3
R1309 a_n6328_16092.n65 a_n6328_16092.n64 9.3
R1310 a_n6328_16092.n101 a_n6328_16092.n100 9.3
R1311 a_n6328_16092.n103 a_n6328_16092.n107 9.3
R1312 a_n6328_16092.n110 a_n6328_16092.n109 9.3
R1313 a_n6328_16092.n10 a_n6328_16092.n112 9.3
R1314 a_n6328_16092.n1 a_n6328_16092.n96 9.3
R1315 a_n6328_16092.n92 a_n6328_16092.n91 9.3
R1316 a_n6328_16092.n90 a_n6328_16092.n89 9.3
R1317 a_n6328_16092.n14 a_n6328_16092.n47 9.3
R1318 a_n6328_16092.n9 a_n6328_16092.n45 9.3
R1319 a_n6328_16092.n9 a_n6328_16092.n44 9.3
R1320 a_n6328_16092.n36 a_n6328_16092.n35 9.3
R1321 a_n6328_16092.n31 a_n6328_16092.n30 9.3
R1322 a_n6328_16092.n39 a_n6328_16092.n38 9.3
R1323 a_n6328_16092.n41 a_n6328_16092.n40 9.3
R1324 a_n6328_16092.n14 a_n6328_16092.n48 9.3
R1325 a_n6328_16092.n58 a_n6328_16092.n57 9.3
R1326 a_n6328_16092.n66 a_n6328_16092.n63 9
R1327 a_n6328_16092.n11 a_n6328_16092.n111 9
R1328 a_n6328_16092.n104 a_n6328_16092.n102 9
R1329 a_n6328_16092.n97 a_n6328_16092.n93 9
R1330 a_n6328_16092.n6 a_n6328_16092.n88 9
R1331 a_n6328_16092.n13 a_n6328_16092.n81 9
R1332 a_n6328_16092.n76 a_n6328_16092.n73 9
R1333 a_n6328_16092.n50 a_n6328_16092.n49 9
R1334 a_n6328_16092.n114 a_n6328_16092.n113 9
R1335 a_n6328_16092.n118 a_n6328_16092.n22 8.473
R1336 a_n6328_16092.n118 a_n6328_16092.n25 8.096
R1337 a_n6328_16092.n118 a_n6328_16092.n20 8.069
R1338 a_n6328_16092.n118 a_n6328_16092.n28 8.043
R1339 a_n6328_16092.n118 a_n6328_16092.n17 8.016
R1340 a_n6328_16092.n72 a_n6328_16092.n71 4.574
R1341 a_n6328_16092.n55 a_n6328_16092.n54 4.574
R1342 a_n6328_16092.n71 a_n6328_16092.n69 3.388
R1343 a_n6328_16092.n54 a_n6328_16092.n52 3.388
R1344 a_n6328_16092.n59 a_n6328_16092.t0 3.326
R1345 a_n6328_16092.t1 a_n6328_16092.n118 3.326
R1346 a_n6328_16092.n2 a_n6328_16092.n66 3
R1347 a_n6328_16092.n0 a_n6328_16092.n6 3
R1348 a_n6328_16092.n4 a_n6328_16092.n13 3
R1349 a_n6328_16092.n4 a_n6328_16092.n76 3
R1350 a_n6328_16092.n2 a_n6328_16092.n72 3
R1351 a_n6328_16092.n98 a_n6328_16092.n97 3
R1352 a_n6328_16092.n7 a_n6328_16092.n104 3
R1353 a_n6328_16092.n8 a_n6328_16092.n11 3
R1354 a_n6328_16092.n114 a_n6328_16092.n2 3
R1355 a_n6328_16092.n19 a_n6328_16092.n18 2.258
R1356 a_n6328_16092.n24 a_n6328_16092.n23 2.258
R1357 a_n6328_16092.n27 a_n6328_16092.n26 1.505
R1358 a_n6328_16092.n22 a_n6328_16092.n21 1.505
R1359 a_n6328_16092.n60 a_n6328_16092.n59 1.155
R1360 a_n6328_16092.n118 a_n6328_16092.n117 1.155
R1361 a_n6328_16092.n61 a_n6328_16092.n60 0.893
R1362 a_n6328_16092.n117 a_n6328_16092.n116 0.893
R1363 a_n6328_16092.n16 a_n6328_16092.n15 0.752
R1364 a_n6328_16092.n71 a_n6328_16092.n70 0.506
R1365 a_n6328_16092.n54 a_n6328_16092.n53 0.506
R1366 a_n6328_16092.n80 a_n6328_16092.n79 0.476
R1367 a_n6328_16092.n17 a_n6328_16092.n16 0.476
R1368 a_n6328_16092.n28 a_n6328_16092.n27 0.445
R1369 a_n6328_16092.n87 a_n6328_16092.n86 0.445
R1370 a_n6328_16092.n96 a_n6328_16092.n95 0.414
R1371 a_n6328_16092.n20 a_n6328_16092.n19 0.413
R1372 a_n6328_16092.n107 a_n6328_16092.n106 0.382
R1373 a_n6328_16092.n25 a_n6328_16092.n24 0.382
R1374 a_n6328_16092.n8 a_n6328_16092.t2 0.224
R1375 a_n6328_16092.n42 a_n6328_16092.n41 0.06
R1376 a_n6328_16092.n33 a_n6328_16092.n32 0.06
R1377 a_n6328_16092.n72 a_n6328_16092.n68 0.053
R1378 a_n6328_16092.n55 a_n6328_16092.n51 0.053
R1379 a_n6328_16092.n51 a_n6328_16092.n50 0.053
R1380 a_n6328_16092.n66 a_n6328_16092.n62 0.043
R1381 a_n6328_16092.n103 a_n6328_16092.n105 0.043
R1382 a_n6328_16092.n115 a_n6328_16092.n114 0.043
R1383 a_n6328_16092.n34 a_n6328_16092.n33 0.043
R1384 a_n6328_16092.n14 a_n6328_16092.n46 0.091
R1385 a_n6328_16092.n46 a_n6328_16092.n9 0.069
R1386 a_n6328_16092.n13 a_n6328_16092.n78 0.044
R1387 a_n6328_16092.n36 a_n6328_16092.n34 0.04
R1388 a_n6328_16092.n31 a_n6328_16092.n29 0.04
R1389 a_n6328_16092.n1 a_n6328_16092.n94 0.036
R1390 a_n6328_16092.n9 a_n6328_16092.n43 0.066
R1391 a_n6328_16092.n7 a_n6328_16092.n8 0.042
R1392 a_n6328_16092.n6 a_n6328_16092.n5 0.04
R1393 a_n6328_16092.n6 a_n6328_16092.n85 0.035
R1394 a_n6328_16092.n98 a_n6328_16092.n7 0.033
R1395 a_n6328_16092.n2 a_n6328_16092.n4 0.031
R1396 a_n6328_16092.n85 a_n6328_16092.n84 0.026
R1397 a_n6328_16092.n97 a_n6328_16092.n92 0.026
R1398 a_n6328_16092.n104 a_n6328_16092.n101 0.026
R1399 a_n6328_16092.n43 a_n6328_16092.n42 0.026
R1400 a_n6328_16092.n39 a_n6328_16092.n37 0.148
R1401 a_n6328_16092.n3 a_n6328_16092.n0 0.032
R1402 a_n6328_16092.n97 a_n6328_16092.n1 0.026
R1403 a_n6328_16092.n110 a_n6328_16092.n108 0.024
R1404 a_n6328_16092.n11 a_n6328_16092.n110 0.024
R1405 a_n6328_16092.n32 a_n6328_16092.n31 0.024
R1406 a_n6328_16092.n50 a_n6328_16092.n14 0.023
R1407 a_n6328_16092.n76 a_n6328_16092.n12 0.023
R1408 a_n6328_16092.n4 a_n6328_16092.n3 0.023
R1409 a_n6328_16092.n72 a_n6328_16092.n67 0.021
R1410 a_n6328_16092.n56 a_n6328_16092.n55 0.021
R1411 a_n6328_16092.n0 a_n6328_16092.n98 0.02
R1412 a_n6328_16092.n62 a_n6328_16092.n61 0.019
R1413 a_n6328_16092.n101 a_n6328_16092.n99 0.019
R1414 a_n6328_16092.n116 a_n6328_16092.n115 0.019
R1415 a_n6328_16092.n58 a_n6328_16092.n56 0.019
R1416 a_n6328_16092.n37 a_n6328_16092.n36 0.019
R1417 a_n6328_16092.n78 a_n6328_16092.n77 0.016
R1418 a_n6328_16092.n11 a_n6328_16092.n10 0.016
R1419 a_n6328_16092.n104 a_n6328_16092.n103 0.014
R1420 a_n6328_16092.n66 a_n6328_16092.n65 0.014
R1421 a_n6328_16092.n92 a_n6328_16092.n90 0.014
R1422 a_n6328_16092.n114 a_n6328_16092.n58 0.014
R1423 a_n6328_16092.n41 a_n6328_16092.n39 0.014
R1424 a_n5540_16092.n23 a_n5540_16092.n21 9.469
R1425 a_n5540_16092.n43 a_n5540_16092.n42 9.3
R1426 a_n5540_16092.n4 a_n5540_16092.n79 9.3
R1427 a_n5540_16092.n5 a_n5540_16092.n77 9.3
R1428 a_n5540_16092.n1 a_n5540_16092.n49 9.3
R1429 a_n5540_16092.n1 a_n5540_16092.n50 9.3
R1430 a_n5540_16092.n2 a_n5540_16092.n53 9.3
R1431 a_n5540_16092.n38 a_n5540_16092.n46 9.3
R1432 a_n5540_16092.n48 a_n5540_16092.n47 9.3
R1433 a_n5540_16092.n63 a_n5540_16092.n62 9.3
R1434 a_n5540_16092.n58 a_n5540_16092.n57 9.3
R1435 a_n5540_16092.n56 a_n5540_16092.n55 9.3
R1436 a_n5540_16092.n4 a_n5540_16092.n80 9.3
R1437 a_n5540_16092.n69 a_n5540_16092.n68 9.3
R1438 a_n5540_16092.n0 a_n5540_16092.n41 9.3
R1439 a_n5540_16092.n6 a_n5540_16092.n33 9.3
R1440 a_n5540_16092.n3 a_n5540_16092.n32 9.3
R1441 a_n5540_16092.n23 a_n5540_16092.n22 9.3
R1442 a_n5540_16092.n28 a_n5540_16092.n27 9.3
R1443 a_n5540_16092.n30 a_n5540_16092.n29 9.3
R1444 a_n5540_16092.n3 a_n5540_16092.n31 9.3
R1445 a_n5540_16092.n6 a_n5540_16092.n34 9.3
R1446 a_n5540_16092.n96 a_n5540_16092.n95 9.3
R1447 a_n5540_16092.n60 a_n5540_16092.n59 9
R1448 a_n5540_16092.n39 a_n5540_16092.n37 9
R1449 a_n5540_16092.n2 a_n5540_16092.n51 9
R1450 a_n5540_16092.n0 a_n5540_16092.n40 9
R1451 a_n5540_16092.n70 a_n5540_16092.n67 9
R1452 a_n5540_16092.n5 a_n5540_16092.n78 9
R1453 a_n5540_16092.n81 a_n5540_16092.n74 9
R1454 a_n5540_16092.n36 a_n5540_16092.n35 9
R1455 a_n5540_16092.n98 a_n5540_16092.n97 9
R1456 a_n5540_16092.n101 a_n5540_16092.n14 8.473
R1457 a_n5540_16092.n101 a_n5540_16092.n17 8.097
R1458 a_n5540_16092.n101 a_n5540_16092.n12 8.069
R1459 a_n5540_16092.n101 a_n5540_16092.n20 8.043
R1460 a_n5540_16092.n101 a_n5540_16092.n9 8.016
R1461 a_n5540_16092.n86 a_n5540_16092.n85 4.574
R1462 a_n5540_16092.n93 a_n5540_16092.n92 4.574
R1463 a_n5540_16092.n85 a_n5540_16092.n83 3.388
R1464 a_n5540_16092.n92 a_n5540_16092.n90 3.388
R1465 a_n5540_16092.n71 a_n5540_16092.t0 3.326
R1466 a_n5540_16092.t1 a_n5540_16092.n101 3.326
R1467 a_n5540_16092.n88 a_n5540_16092.n64 3.008
R1468 a_n5540_16092.n66 a_n5540_16092.n87 2.989
R1469 a_n5540_16092.n66 a_n5540_16092.n73 2.987
R1470 a_n5540_16092.n89 a_n5540_16092.n88 2.287
R1471 a_n5540_16092.n11 a_n5540_16092.n10 2.258
R1472 a_n5540_16092.n16 a_n5540_16092.n15 2.258
R1473 a_n5540_16092.n19 a_n5540_16092.n18 1.505
R1474 a_n5540_16092.n14 a_n5540_16092.n13 1.505
R1475 a_n5540_16092.n72 a_n5540_16092.n71 1.155
R1476 a_n5540_16092.n101 a_n5540_16092.n100 1.155
R1477 a_n5540_16092.n73 a_n5540_16092.n72 0.921
R1478 a_n5540_16092.n100 a_n5540_16092.n99 0.903
R1479 a_n5540_16092.n8 a_n5540_16092.n7 0.752
R1480 a_n5540_16092.n85 a_n5540_16092.n84 0.506
R1481 a_n5540_16092.n92 a_n5540_16092.n91 0.506
R1482 a_n5540_16092.n77 a_n5540_16092.n76 0.476
R1483 a_n5540_16092.n9 a_n5540_16092.n8 0.476
R1484 a_n5540_16092.n20 a_n5540_16092.n19 0.445
R1485 a_n5540_16092.n53 a_n5540_16092.n52 0.445
R1486 a_n5540_16092.n62 a_n5540_16092.n61 0.414
R1487 a_n5540_16092.n12 a_n5540_16092.n11 0.414
R1488 a_n5540_16092.n17 a_n5540_16092.n16 0.382
R1489 a_n5540_16092.n46 a_n5540_16092.n45 0.382
R1490 a_n5540_16092.n6 a_n5540_16092.n3 0.161
R1491 a_n5540_16092.n88 a_n5540_16092.t2 0.158
R1492 a_n5540_16092.n56 a_n5540_16092.n54 0.073
R1493 a_n5540_16092.n3 a_n5540_16092.n30 0.153
R1494 a_n5540_16092.n38 a_n5540_16092.n44 0.073
R1495 a_n5540_16092.n64 a_n5540_16092.n48 0.072
R1496 a_n5540_16092.n24 a_n5540_16092.n23 0.072
R1497 a_n5540_16092.n87 a_n5540_16092.n81 0.071
R1498 a_n5540_16092.n64 a_n5540_16092.n63 0.057
R1499 a_n5540_16092.n25 a_n5540_16092.n24 0.057
R1500 a_n5540_16092.n44 a_n5540_16092.n43 0.054
R1501 a_n5540_16092.n93 a_n5540_16092.n89 0.054
R1502 a_n5540_16092.n89 a_n5540_16092.n36 0.054
R1503 a_n5540_16092.n99 a_n5540_16092.n98 0.053
R1504 a_n5540_16092.n88 a_n5540_16092.n66 0.052
R1505 a_n5540_16092.n2 a_n5540_16092.n1 0.049
R1506 a_n5540_16092.n5 a_n5540_16092.n75 0.048
R1507 a_n5540_16092.n43 a_n5540_16092.n0 0.041
R1508 a_n5540_16092.n54 a_n5540_16092.n2 0.039
R1509 a_n5540_16092.n87 a_n5540_16092.n86 0.036
R1510 a_n5540_16092.n73 a_n5540_16092.n70 0.036
R1511 a_n5540_16092.n4 a_n5540_16092.n5 0.035
R1512 a_n5540_16092.n60 a_n5540_16092.n58 0.026
R1513 a_n5540_16092.n48 a_n5540_16092.n39 0.026
R1514 a_n5540_16092.n28 a_n5540_16092.n26 0.026
R1515 a_n5540_16092.n36 a_n5540_16092.n6 0.023
R1516 a_n5540_16092.n81 a_n5540_16092.n4 0.023
R1517 a_n5540_16092.n86 a_n5540_16092.n82 0.021
R1518 a_n5540_16092.n94 a_n5540_16092.n93 0.021
R1519 a_n5540_16092.n96 a_n5540_16092.n94 0.019
R1520 a_n5540_16092.n39 a_n5540_16092.n38 0.015
R1521 a_n5540_16092.n70 a_n5540_16092.n69 0.014
R1522 a_n5540_16092.n58 a_n5540_16092.n56 0.014
R1523 a_n5540_16092.n63 a_n5540_16092.n60 0.014
R1524 a_n5540_16092.n98 a_n5540_16092.n96 0.014
R1525 a_n5540_16092.n30 a_n5540_16092.n28 0.014
R1526 a_n5540_16092.n26 a_n5540_16092.n25 0.014
R1527 a_n5540_16092.n66 a_n5540_16092.n65 0.014
R1528 a_n6722_16092.n78 a_n6722_16092.n76 9.468
R1529 a_n6722_16092.n4 a_n6722_16092.n65 9.3
R1530 a_n6722_16092.n5 a_n6722_16092.n63 9.3
R1531 a_n6722_16092.n2 a_n6722_16092.n27 9.3
R1532 a_n6722_16092.n1 a_n6722_16092.n23 9.3
R1533 a_n6722_16092.n1 a_n6722_16092.n24 9.3
R1534 a_n6722_16092.n49 a_n6722_16092.n48 9.3
R1535 a_n6722_16092.n39 a_n6722_16092.n47 9.3
R1536 a_n6722_16092.n44 a_n6722_16092.n43 9.3
R1537 a_n6722_16092.n0 a_n6722_16092.n42 9.3
R1538 a_n6722_16092.n37 a_n6722_16092.n36 9.3
R1539 a_n6722_16092.n32 a_n6722_16092.n31 9.3
R1540 a_n6722_16092.n30 a_n6722_16092.n29 9.3
R1541 a_n6722_16092.n4 a_n6722_16092.n66 9.3
R1542 a_n6722_16092.n57 a_n6722_16092.n56 9.3
R1543 a_n6722_16092.n6 a_n6722_16092.n83 9.3
R1544 a_n6722_16092.n3 a_n6722_16092.n82 9.3
R1545 a_n6722_16092.n3 a_n6722_16092.n81 9.3
R1546 a_n6722_16092.n6 a_n6722_16092.n84 9.3
R1547 a_n6722_16092.n94 a_n6722_16092.n93 9.3
R1548 a_n6722_16092.n78 a_n6722_16092.n77 9.3
R1549 a_n6722_16092.n80 a_n6722_16092.n79 9.3
R1550 a_n6722_16092.n0 a_n6722_16092.n41 9
R1551 a_n6722_16092.n40 a_n6722_16092.n38 9
R1552 a_n6722_16092.n34 a_n6722_16092.n33 9
R1553 a_n6722_16092.n2 a_n6722_16092.n25 9
R1554 a_n6722_16092.n5 a_n6722_16092.n64 9
R1555 a_n6722_16092.n67 a_n6722_16092.n60 9
R1556 a_n6722_16092.n58 a_n6722_16092.n55 9
R1557 a_n6722_16092.n96 a_n6722_16092.n95 9
R1558 a_n6722_16092.n86 a_n6722_16092.n85 9
R1559 a_n6722_16092.n99 a_n6722_16092.n17 8.473
R1560 a_n6722_16092.n99 a_n6722_16092.n20 8.096
R1561 a_n6722_16092.n99 a_n6722_16092.n15 8.069
R1562 a_n6722_16092.n99 a_n6722_16092.n12 8.042
R1563 a_n6722_16092.n99 a_n6722_16092.n9 8.016
R1564 a_n6722_16092.n72 a_n6722_16092.n71 4.574
R1565 a_n6722_16092.n91 a_n6722_16092.n90 4.574
R1566 a_n6722_16092.n71 a_n6722_16092.n69 3.388
R1567 a_n6722_16092.n90 a_n6722_16092.n88 3.388
R1568 a_n6722_16092.n53 a_n6722_16092.t0 3.326
R1569 a_n6722_16092.t1 a_n6722_16092.n99 3.326
R1570 a_n6722_16092.n74 a_n6722_16092.n50 3.009
R1571 a_n6722_16092.n52 a_n6722_16092.n73 2.989
R1572 a_n6722_16092.n52 a_n6722_16092.n59 2.987
R1573 a_n6722_16092.n97 a_n6722_16092.n22 2.987
R1574 a_n6722_16092.n14 a_n6722_16092.n13 2.258
R1575 a_n6722_16092.n19 a_n6722_16092.n18 2.258
R1576 a_n6722_16092.n11 a_n6722_16092.n10 1.505
R1577 a_n6722_16092.n17 a_n6722_16092.n16 1.505
R1578 a_n6722_16092.n99 a_n6722_16092.n98 1.155
R1579 a_n6722_16092.n54 a_n6722_16092.n53 1.155
R1580 a_n6722_16092.n98 a_n6722_16092.n97 0.921
R1581 a_n6722_16092.n59 a_n6722_16092.n54 0.921
R1582 a_n6722_16092.n8 a_n6722_16092.n7 0.752
R1583 a_n6722_16092.n71 a_n6722_16092.n70 0.506
R1584 a_n6722_16092.n90 a_n6722_16092.n89 0.506
R1585 a_n6722_16092.n63 a_n6722_16092.n62 0.476
R1586 a_n6722_16092.n9 a_n6722_16092.n8 0.476
R1587 a_n6722_16092.n27 a_n6722_16092.n26 0.445
R1588 a_n6722_16092.n12 a_n6722_16092.n11 0.445
R1589 a_n6722_16092.n36 a_n6722_16092.n35 0.414
R1590 a_n6722_16092.n15 a_n6722_16092.n14 0.414
R1591 a_n6722_16092.n47 a_n6722_16092.n46 0.382
R1592 a_n6722_16092.n20 a_n6722_16092.n19 0.382
R1593 a_n6722_16092.n6 a_n6722_16092.n3 0.161
R1594 a_n6722_16092.n100 a_n6722_16092.t2 0.127
R1595 a_n6722_16092.n30 a_n6722_16092.n28 0.073
R1596 a_n6722_16092.n3 a_n6722_16092.n80 0.153
R1597 a_n6722_16092.n39 a_n6722_16092.n45 0.073
R1598 a_n6722_16092.n50 a_n6722_16092.n49 0.072
R1599 a_n6722_16092.n73 a_n6722_16092.n67 0.071
R1600 a_n6722_16092.n87 a_n6722_16092.n86 0.071
R1601 a_n6722_16092.n50 a_n6722_16092.n37 0.057
R1602 a_n6722_16092.n74 a_n6722_16092.n52 0.055
R1603 a_n6722_16092.n45 a_n6722_16092.n44 0.054
R1604 a_n6722_16092.n2 a_n6722_16092.n1 0.049
R1605 a_n6722_16092.n5 a_n6722_16092.n61 0.048
R1606 a_n6722_16092.n44 a_n6722_16092.n0 0.041
R1607 a_n6722_16092.n28 a_n6722_16092.n2 0.039
R1608 a_n6722_16092.n21 a_n6722_16092.n74 0.039
R1609 a_n6722_16092.n74 a_n6722_16092.n100 0.037
R1610 a_n6722_16092.n73 a_n6722_16092.n72 0.036
R1611 a_n6722_16092.n91 a_n6722_16092.n87 0.036
R1612 a_n6722_16092.n59 a_n6722_16092.n58 0.036
R1613 a_n6722_16092.n97 a_n6722_16092.n96 0.036
R1614 a_n6722_16092.n4 a_n6722_16092.n5 0.035
R1615 a_n6722_16092.n34 a_n6722_16092.n32 0.026
R1616 a_n6722_16092.n49 a_n6722_16092.n40 0.026
R1617 a_n6722_16092.n86 a_n6722_16092.n6 0.023
R1618 a_n6722_16092.n67 a_n6722_16092.n4 0.023
R1619 a_n6722_16092.n72 a_n6722_16092.n68 0.021
R1620 a_n6722_16092.n92 a_n6722_16092.n91 0.021
R1621 a_n6722_16092.n94 a_n6722_16092.n92 0.019
R1622 a_n6722_16092.n40 a_n6722_16092.n39 0.015
R1623 a_n6722_16092.n58 a_n6722_16092.n57 0.014
R1624 a_n6722_16092.n32 a_n6722_16092.n30 0.014
R1625 a_n6722_16092.n37 a_n6722_16092.n34 0.014
R1626 a_n6722_16092.n96 a_n6722_16092.n94 0.014
R1627 a_n6722_16092.n80 a_n6722_16092.n78 0.014
R1628 a_n6722_16092.n52 a_n6722_16092.n51 0.014
R1629 a_n6722_16092.n22 a_n6722_16092.n21 0.014
R1630 a_n6722_16092.n22 a_n6722_16092.n75 0.014
R1631 a_n5934_16092.n5 a_n5934_16092.n93 9.3
R1632 a_n5934_16092.n7 a_n5934_16092.n85 9.3
R1633 a_n5934_16092.n8 a_n5934_16092.n83 9.3
R1634 a_n5934_16092.n2 a_n5934_16092.n79 9.3
R1635 a_n5934_16092.n73 a_n5934_16092.n72 9.3
R1636 a_n5934_16092.n2 a_n5934_16092.n78 9.3
R1637 a_n5934_16092.n3 a_n5934_16092.n77 9.3
R1638 a_n5934_16092.n71 a_n5934_16092.n70 9.3
R1639 a_n5934_16092.n0 a_n5934_16092.n67 9.3
R1640 a_n5934_16092.n63 a_n5934_16092.n62 9.3
R1641 a_n5934_16092.n57 a_n5934_16092.n61 9.3
R1642 a_n5934_16092.n7 a_n5934_16092.n86 9.3
R1643 a_n5934_16092.n49 a_n5934_16092.n48 9.3
R1644 a_n5934_16092.n4 a_n5934_16092.n94 9.3
R1645 a_n5934_16092.n1 a_n5934_16092.n35 9.3
R1646 a_n5934_16092.n31 a_n5934_16092.n30 9.3
R1647 a_n5934_16092.n6 a_n5934_16092.n37 9.3
R1648 a_n5934_16092.n103 a_n5934_16092.n102 9.3
R1649 a_n5934_16092.n26 a_n5934_16092.n25 9.3
R1650 a_n5934_16092.n29 a_n5934_16092.n28 9.3
R1651 a_n5934_16092.n1 a_n5934_16092.n34 9.3
R1652 a_n5934_16092.n6 a_n5934_16092.n38 9.3
R1653 a_n5934_16092.n47 a_n5934_16092.n46 9
R1654 a_n5934_16092.n3 a_n5934_16092.n55 9
R1655 a_n5934_16092.n69 a_n5934_16092.n68 9
R1656 a_n5934_16092.n58 a_n5934_16092.n56 9
R1657 a_n5934_16092.n8 a_n5934_16092.n84 9
R1658 a_n5934_16092.n88 a_n5934_16092.n87 9
R1659 a_n5934_16092.n4 a_n5934_16092.n95 9
R1660 a_n5934_16092.n105 a_n5934_16092.n104 9
R1661 a_n5934_16092.n40 a_n5934_16092.n39 9
R1662 a_n5934_16092.n110 a_n5934_16092.n17 8.473
R1663 a_n5934_16092.n110 a_n5934_16092.n20 8.097
R1664 a_n5934_16092.n110 a_n5934_16092.n15 8.069
R1665 a_n5934_16092.n110 a_n5934_16092.n23 8.043
R1666 a_n5934_16092.n110 a_n5934_16092.n12 8.016
R1667 a_n5934_16092.n54 a_n5934_16092.n53 4.574
R1668 a_n5934_16092.n100 a_n5934_16092.n99 4.574
R1669 a_n5934_16092.n53 a_n5934_16092.n51 3.388
R1670 a_n5934_16092.n99 a_n5934_16092.n97 3.388
R1671 a_n5934_16092.n41 a_n5934_16092.t2 3.326
R1672 a_n5934_16092.t1 a_n5934_16092.n110 3.326
R1673 a_n5934_16092.n9 a_n5934_16092.n5 2.561
R1674 a_n5934_16092.n96 a_n5934_16092.n90 2.473
R1675 a_n5934_16092.n14 a_n5934_16092.n13 2.258
R1676 a_n5934_16092.n19 a_n5934_16092.n18 2.258
R1677 a_n5934_16092.n90 a_n5934_16092.n89 1.94
R1678 a_n5934_16092.n22 a_n5934_16092.n21 1.505
R1679 a_n5934_16092.n17 a_n5934_16092.n16 1.505
R1680 a_n5934_16092.n42 a_n5934_16092.n41 1.155
R1681 a_n5934_16092.n110 a_n5934_16092.n109 1.155
R1682 a_n5934_16092.n43 a_n5934_16092.n42 0.852
R1683 a_n5934_16092.n109 a_n5934_16092.n108 0.852
R1684 a_n5934_16092.n11 a_n5934_16092.n10 0.752
R1685 a_n5934_16092.n99 a_n5934_16092.n98 0.506
R1686 a_n5934_16092.n53 a_n5934_16092.n52 0.506
R1687 a_n5934_16092.n83 a_n5934_16092.n82 0.476
R1688 a_n5934_16092.n12 a_n5934_16092.n11 0.476
R1689 a_n5934_16092.n23 a_n5934_16092.n22 0.445
R1690 a_n5934_16092.n77 a_n5934_16092.n76 0.445
R1691 a_n5934_16092.n67 a_n5934_16092.n66 0.414
R1692 a_n5934_16092.n15 a_n5934_16092.n14 0.414
R1693 a_n5934_16092.n20 a_n5934_16092.n19 0.382
R1694 a_n5934_16092.n61 a_n5934_16092.n60 0.382
R1695 a_n5934_16092.n9 a_n5934_16092.t0 0.179
R1696 a_n5934_16092.n32 a_n5934_16092.n31 0.06
R1697 a_n5934_16092.n80 a_n5934_16092.n2 0.06
R1698 a_n5934_16092.n74 a_n5934_16092.n73 0.06
R1699 a_n5934_16092.n65 a_n5934_16092.n64 0.06
R1700 a_n5934_16092.n90 a_n5934_16092.n9 0.056
R1701 a_n5934_16092.n89 a_n5934_16092.n54 0.054
R1702 a_n5934_16092.n100 a_n5934_16092.n96 0.054
R1703 a_n5934_16092.n96 a_n5934_16092.n40 0.053
R1704 a_n5934_16092.n89 a_n5934_16092.n88 0.053
R1705 a_n5934_16092.n57 a_n5934_16092.n59 0.043
R1706 a_n5934_16092.n108 a_n5934_16092.n107 0.04
R1707 a_n5934_16092.n106 a_n5934_16092.n105 0.04
R1708 a_n5934_16092.n6 a_n5934_16092.n36 0.091
R1709 a_n5934_16092.n26 a_n5934_16092.n24 9.474
R1710 a_n5934_16092.n36 a_n5934_16092.n1 0.069
R1711 a_n5934_16092.n44 a_n5934_16092.n43 0.04
R1712 a_n5934_16092.n47 a_n5934_16092.n45 0.04
R1713 a_n5934_16092.n8 a_n5934_16092.n81 0.04
R1714 a_n5934_16092.n5 a_n5934_16092.n4 0.04
R1715 a_n5934_16092.n2 a_n5934_16092.n3 0.04
R1716 a_n5934_16092.n0 a_n5934_16092.n65 0.036
R1717 a_n5934_16092.n7 a_n5934_16092.n8 0.035
R1718 a_n5934_16092.n3 a_n5934_16092.n75 0.035
R1719 a_n5934_16092.n1 a_n5934_16092.n33 0.066
R1720 a_n5934_16092.n9 a_n5934_16092.n91 0.027
R1721 a_n5934_16092.n33 a_n5934_16092.n32 0.026
R1722 a_n5934_16092.n29 a_n5934_16092.n27 0.148
R1723 a_n5934_16092.n75 a_n5934_16092.n74 0.026
R1724 a_n5934_16092.n71 a_n5934_16092.n69 0.026
R1725 a_n5934_16092.n63 a_n5934_16092.n58 0.026
R1726 a_n5934_16092.n69 a_n5934_16092.n0 0.026
R1727 a_n5934_16092.n5 a_n5934_16092.n92 0.024
R1728 a_n5934_16092.n88 a_n5934_16092.n7 0.023
R1729 a_n5934_16092.n40 a_n5934_16092.n6 0.023
R1730 a_n5934_16092.n107 a_n5934_16092.n106 0.021
R1731 a_n5934_16092.n101 a_n5934_16092.n100 0.021
R1732 a_n5934_16092.n45 a_n5934_16092.n44 0.021
R1733 a_n5934_16092.n54 a_n5934_16092.n50 0.021
R1734 a_n5934_16092.n103 a_n5934_16092.n101 0.019
R1735 a_n5934_16092.n27 a_n5934_16092.n26 0.019
R1736 a_n5934_16092.n50 a_n5934_16092.n49 0.019
R1737 a_n5934_16092.n64 a_n5934_16092.n63 0.019
R1738 a_n5934_16092.n81 a_n5934_16092.n80 0.016
R1739 a_n5934_16092.n58 a_n5934_16092.n57 0.014
R1740 a_n5934_16092.n105 a_n5934_16092.n103 0.014
R1741 a_n5934_16092.n31 a_n5934_16092.n29 0.014
R1742 a_n5934_16092.n49 a_n5934_16092.n47 0.014
R1743 a_n5934_16092.n73 a_n5934_16092.n71 0.014
C0 SS m5_n800_n3000# 4.99fF
C1 SS VIN 6.02fF
C2 S1 VOUT 19.96fF
C3 VIN D1 1.27fF
C4 VHI VOUT 1.26fF
C5 SS D1 13.20fF
C6 G_TOP VOUT 2.50fF
C7 G_TOP S1 1.40fF
C8 VHI VLO 422.33fF
C9 SS VLO 12.33fF $ **FLOATING
C10 D1 VLO 36.13fF $ **FLOATING
C11 VIN VLO 3.85fF
C12 S1 VLO 46.25fF $ **FLOATING
C13 G_TOP VLO 3.78fF
C14 a_n1934_7566# VLO 1.42fF $ **FLOATING
C15 VOUT VLO 70.01fF $ **FLOATING
C16 G4 VLO 1.28fF
C17 G8 VLO 1.10fF
C18 G1 VLO 1.06fF
C19 G2 VLO 1.29fF
C20 a_n5934_16092.n9 VLO 1.46fF $ **FLOATING
C21 a_n5934_16092.t0 VLO 9.51fF
C22 a_n6722_16092.t2 VLO 3.36fF
C23 a_n5540_16092.n88 VLO 1.54fF $ **FLOATING
C24 a_n5540_16092.t2 VLO 6.69fF
C25 a_n6328_16092.t2 VLO 2.99fF
C26 SS.n484 VLO 28.08fF $ **FLOATING
C27 D1.n0 VLO 6.27fF $ **FLOATING
C28 S1.n10 VLO 3.63fF $ **FLOATING
C29 VOUT.n59 VLO 6.00fF $ **FLOATING
C30 VOUT.n134 VLO 1.20fF $ **FLOATING
C31 VOUT.n752 VLO 61.25fF $ **FLOATING


**** end user architecture code
.ends

.GLOBAL GND
.GLOBAL GNDI
.end
