magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< nwell >>
rect -36 679 620 1471
<< poly >>
rect 114 740 144 971
rect 81 674 144 740
rect 114 443 144 674
<< locali >>
rect 0 1397 584 1431
rect 62 1162 96 1397
rect 274 1162 308 1397
rect 482 1297 516 1397
rect 64 674 98 740
rect 272 724 306 1128
rect 272 690 323 724
rect 272 286 306 690
rect 62 17 96 186
rect 274 17 308 186
rect 482 17 516 104
rect 0 -17 584 17
use sky130_sram_1r1w_24x128_8_contact_15  sky130_sram_1r1w_24x128_8_contact_15_0
timestamp 1661296025
transform 1 0 48 0 1 674
box 0 0 66 66
use sky130_sram_1r1w_24x128_8_contact_28  sky130_sram_1r1w_24x128_8_contact_28_0
timestamp 1661296025
transform 1 0 474 0 1 1256
box -59 -43 109 125
use sky130_sram_1r1w_24x128_8_contact_29  sky130_sram_1r1w_24x128_8_contact_29_0
timestamp 1661296025
transform 1 0 474 0 1 63
box -26 -26 76 108
use sky130_sram_1r1w_24x128_8_nmos_m3_w1_680_sli_dli_da_p  sky130_sram_1r1w_24x128_8_nmos_m3_w1_680_sli_dli_da_p_0
timestamp 1661296025
transform 1 0 54 0 1 51
box -26 -26 392 392
use sky130_sram_1r1w_24x128_8_pmos_m3_w1_680_sli_dli_da_p  sky130_sram_1r1w_24x128_8_pmos_m3_w1_680_sli_dli_da_p_0
timestamp 1661296025
transform 1 0 54 0 1 1027
box -59 -56 425 390
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 306 707 306 707 4 Z
port 2 nsew
rlabel locali s 292 0 292 0 4 gnd
port 3 nsew
rlabel locali s 292 1414 292 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 584 1414
<< end >>
