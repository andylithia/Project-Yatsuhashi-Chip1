magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< error_p >>
rect 4 61 70 66
rect 4 5 9 61
rect 4 0 70 5
<< metal2 >>
rect 0 5 9 61
rect 65 5 74 61
<< via2 >>
rect 9 5 65 61
<< metal3 >>
rect 4 61 70 66
rect 4 5 9 61
rect 65 5 70 61
rect 4 0 70 5
<< properties >>
string FIXED_BBOX 0 0 74 66
<< end >>
