magic
tech sky130B
magscale 1 2
timestamp 1661836362
<< metal1 >>
rect 16000 13700 20000 13900
rect -13500 13300 -11500 13400
rect -13500 13280 -13380 13300
rect -13120 13280 -12880 13300
rect -12620 13280 -12380 13300
rect -12120 13280 -11880 13300
rect -11620 13280 -11500 13300
rect -13500 13020 -13400 13280
rect -13100 13020 -12900 13280
rect -12600 13020 -12400 13280
rect -12100 13020 -11900 13280
rect -11600 13020 -11500 13280
rect -13500 13000 -13380 13020
rect -13120 13000 -12880 13020
rect -12620 13000 -12380 13020
rect -12120 13000 -11880 13020
rect -11620 13000 -11500 13020
rect -13500 12800 -11500 13000
rect -13500 12780 -13380 12800
rect -13120 12780 -12880 12800
rect -12620 12780 -12380 12800
rect -12120 12780 -11880 12800
rect -11620 12780 -11500 12800
rect -13500 12520 -13400 12780
rect -13100 12520 -12900 12780
rect -12600 12520 -12400 12780
rect -12100 12520 -11900 12780
rect -11600 12520 -11500 12780
rect -13500 12500 -13380 12520
rect -13120 12500 -12880 12520
rect -12620 12500 -12380 12520
rect -12120 12500 -11880 12520
rect -11620 12500 -11500 12520
rect -13500 12300 -11500 12500
rect -13500 12280 -13380 12300
rect -13120 12280 -12880 12300
rect -12620 12280 -12380 12300
rect -12120 12280 -11880 12300
rect -11620 12280 -11500 12300
rect -13500 12020 -13400 12280
rect -13100 12020 -12900 12280
rect -12600 12020 -12400 12280
rect -12100 12020 -11900 12280
rect -11600 12020 -11500 12280
rect -13500 12000 -13380 12020
rect -13120 12000 -12880 12020
rect -12620 12000 -12380 12020
rect -12120 12000 -11880 12020
rect -11620 12000 -11500 12020
rect -13500 11800 -11500 12000
rect -13500 11780 -13380 11800
rect -13120 11780 -12880 11800
rect -12620 11780 -12380 11800
rect -12120 11780 -11880 11800
rect -11620 11780 -11500 11800
rect -13500 11520 -13400 11780
rect -13100 11520 -12900 11780
rect -12600 11520 -12400 11780
rect -12100 11520 -11900 11780
rect -11600 11520 -11500 11780
rect -13500 11500 -13380 11520
rect -13120 11500 -12880 11520
rect -12620 11500 -12380 11520
rect -12120 11500 -11880 11520
rect -11620 11500 -11500 11520
rect -13500 11300 -11500 11500
rect -13500 11280 -13380 11300
rect -13120 11280 -12880 11300
rect -12620 11280 -12380 11300
rect -12120 11280 -11880 11300
rect -11620 11280 -11500 11300
rect -13500 11020 -13400 11280
rect -13100 11020 -12900 11280
rect -12600 11020 -12400 11280
rect -12100 11020 -11900 11280
rect -11600 11020 -11500 11280
rect -13500 11000 -13380 11020
rect -13120 11000 -12880 11020
rect -12620 11000 -12380 11020
rect -12120 11000 -11880 11020
rect -11620 11000 -11500 11020
rect -13500 10900 -11500 11000
rect -13500 10800 -3000 10900
rect -13500 10780 -13380 10800
rect -13120 10780 -12880 10800
rect -12620 10780 -12380 10800
rect -12120 10780 -11880 10800
rect -11620 10780 -11380 10800
rect -11120 10780 -10880 10800
rect -10620 10780 -10380 10800
rect -10120 10780 -9880 10800
rect -9620 10780 -9380 10800
rect -9120 10780 -8880 10800
rect -8620 10780 -8380 10800
rect -8120 10780 -7880 10800
rect -7620 10780 -7380 10800
rect -7120 10780 -6880 10800
rect -6620 10780 -6380 10800
rect -6120 10780 -5880 10800
rect -5620 10780 -5380 10800
rect -5120 10780 -4880 10800
rect -4620 10780 -4380 10800
rect -4120 10780 -3880 10800
rect -3620 10780 -3380 10800
rect -3120 10780 -3000 10800
rect -13500 10520 -13400 10780
rect -13100 10520 -12900 10780
rect -12600 10520 -12400 10780
rect -12100 10520 -11900 10780
rect -11600 10520 -11400 10780
rect -11100 10520 -10900 10780
rect -10600 10520 -10400 10780
rect -10100 10520 -9900 10780
rect -9600 10520 -9400 10780
rect -9100 10520 -8900 10780
rect -8600 10520 -8400 10780
rect -8100 10520 -7900 10780
rect -7600 10520 -7400 10780
rect -7100 10520 -6900 10780
rect -6600 10520 -6400 10780
rect -6100 10520 -5900 10780
rect -5600 10520 -5400 10780
rect -5100 10520 -4900 10780
rect -4600 10520 -4400 10780
rect -4100 10520 -3900 10780
rect -3600 10520 -3400 10780
rect -3100 10520 -3000 10780
rect -13500 10500 -13380 10520
rect -13120 10500 -12880 10520
rect -12620 10500 -12380 10520
rect -12120 10500 -11880 10520
rect -11620 10500 -11380 10520
rect -11120 10500 -10880 10520
rect -10620 10500 -10380 10520
rect -10120 10500 -9880 10520
rect -9620 10500 -9380 10520
rect -9120 10500 -8880 10520
rect -8620 10500 -8380 10520
rect -8120 10500 -7880 10520
rect -7620 10500 -7380 10520
rect -7120 10500 -6880 10520
rect -6620 10500 -6380 10520
rect -6120 10500 -5880 10520
rect -5620 10500 -5380 10520
rect -5120 10500 -4880 10520
rect -4620 10500 -4380 10520
rect -4120 10500 -3880 10520
rect -3620 10500 -3380 10520
rect -3120 10500 -3000 10520
rect -13500 10300 -3000 10500
rect -13500 10280 -13380 10300
rect -13120 10280 -12880 10300
rect -12620 10280 -12380 10300
rect -12120 10280 -11880 10300
rect -11620 10280 -11380 10300
rect -11120 10280 -10880 10300
rect -10620 10280 -10380 10300
rect -10120 10280 -9880 10300
rect -9620 10280 -9380 10300
rect -9120 10280 -8880 10300
rect -8620 10280 -8380 10300
rect -8120 10280 -7880 10300
rect -7620 10280 -7380 10300
rect -7120 10280 -6880 10300
rect -6620 10280 -6380 10300
rect -6120 10280 -5880 10300
rect -5620 10280 -5380 10300
rect -5120 10280 -4880 10300
rect -4620 10280 -4380 10300
rect -4120 10280 -3880 10300
rect -3620 10280 -3380 10300
rect -3120 10280 -3000 10300
rect -13500 10020 -13400 10280
rect -13100 10020 -12900 10280
rect -12600 10020 -12400 10280
rect -12100 10020 -11900 10280
rect -11600 10020 -11400 10280
rect -11100 10020 -10900 10280
rect -10600 10020 -10400 10280
rect -10100 10020 -9900 10280
rect -9600 10020 -9400 10280
rect -9100 10020 -8900 10280
rect -8600 10020 -8400 10280
rect -8100 10020 -7900 10280
rect -7600 10020 -7400 10280
rect -7100 10020 -6900 10280
rect -6600 10020 -6400 10280
rect -6100 10020 -5900 10280
rect -5600 10020 -5400 10280
rect -5100 10020 -4900 10280
rect -4600 10020 -4400 10280
rect -4100 10020 -3900 10280
rect -3600 10020 -3400 10280
rect -3100 10020 -3000 10280
rect -13500 10000 -13380 10020
rect -13120 10000 -12880 10020
rect -12620 10000 -12380 10020
rect -12120 10000 -11880 10020
rect -11620 10000 -11380 10020
rect -11120 10000 -10880 10020
rect -10620 10000 -10380 10020
rect -10120 10000 -9880 10020
rect -9620 10000 -9380 10020
rect -9120 10000 -8880 10020
rect -8620 10000 -8380 10020
rect -8120 10000 -7880 10020
rect -7620 10000 -7380 10020
rect -7120 10000 -6880 10020
rect -6620 10000 -6380 10020
rect -6120 10000 -5880 10020
rect -5620 10000 -5380 10020
rect -5120 10000 -4880 10020
rect -4620 10000 -4380 10020
rect -4120 10000 -3880 10020
rect -3620 10000 -3380 10020
rect -3120 10000 -3000 10020
rect -13500 9800 -3000 10000
rect -13500 9780 -13380 9800
rect -13120 9780 -12880 9800
rect -12620 9780 -12380 9800
rect -12120 9780 -11880 9800
rect -11620 9780 -11380 9800
rect -11120 9780 -10880 9800
rect -10620 9780 -10380 9800
rect -10120 9780 -9880 9800
rect -9620 9780 -9380 9800
rect -9120 9780 -8880 9800
rect -8620 9780 -8380 9800
rect -8120 9780 -7880 9800
rect -7620 9780 -7380 9800
rect -7120 9780 -6880 9800
rect -6620 9780 -6380 9800
rect -6120 9780 -5880 9800
rect -5620 9780 -5380 9800
rect -5120 9780 -4880 9800
rect -4620 9780 -4380 9800
rect -4120 9780 -3880 9800
rect -3620 9780 -3380 9800
rect -3120 9780 -3000 9800
rect -13500 9520 -13400 9780
rect -13100 9520 -12900 9780
rect -12600 9520 -12400 9780
rect -12100 9520 -11900 9780
rect -11600 9520 -11400 9780
rect -11100 9520 -10900 9780
rect -10600 9520 -10400 9780
rect -10100 9520 -9900 9780
rect -9600 9520 -9400 9780
rect -9100 9520 -8900 9780
rect -8600 9520 -8400 9780
rect -8100 9520 -7900 9780
rect -7600 9520 -7400 9780
rect -7100 9520 -6900 9780
rect -6600 9520 -6400 9780
rect -6100 9520 -5900 9780
rect -5600 9520 -5400 9780
rect -5100 9520 -4900 9780
rect -4600 9520 -4400 9780
rect -4100 9520 -3900 9780
rect -3600 9520 -3400 9780
rect -3100 9520 -3000 9780
rect -13500 9500 -13380 9520
rect -13120 9500 -12880 9520
rect -12620 9500 -12380 9520
rect -12120 9500 -11880 9520
rect -11620 9500 -11380 9520
rect -11120 9500 -10880 9520
rect -10620 9500 -10380 9520
rect -10120 9500 -9880 9520
rect -9620 9500 -9380 9520
rect -9120 9500 -8880 9520
rect -8620 9500 -8380 9520
rect -8120 9500 -7880 9520
rect -7620 9500 -7380 9520
rect -7120 9500 -6880 9520
rect -6620 9500 -6380 9520
rect -6120 9500 -5880 9520
rect -5620 9500 -5380 9520
rect -5120 9500 -4880 9520
rect -4620 9500 -4380 9520
rect -4120 9500 -3880 9520
rect -3620 9500 -3380 9520
rect -3120 9500 -3000 9520
rect -13500 9300 -3000 9500
rect -13500 9280 -13380 9300
rect -13120 9280 -12880 9300
rect -12620 9280 -12380 9300
rect -12120 9280 -11880 9300
rect -11620 9280 -11380 9300
rect -11120 9280 -10880 9300
rect -10620 9280 -10380 9300
rect -10120 9280 -9880 9300
rect -9620 9280 -9380 9300
rect -9120 9280 -8880 9300
rect -8620 9280 -8380 9300
rect -8120 9280 -7880 9300
rect -7620 9280 -7380 9300
rect -7120 9280 -6880 9300
rect -6620 9280 -6380 9300
rect -6120 9280 -5880 9300
rect -5620 9280 -5380 9300
rect -5120 9280 -4880 9300
rect -4620 9280 -4380 9300
rect -4120 9280 -3880 9300
rect -3620 9280 -3380 9300
rect -3120 9280 -3000 9300
rect -13500 9020 -13400 9280
rect -13100 9020 -12900 9280
rect -12600 9020 -12400 9280
rect -12100 9020 -11900 9280
rect -11600 9020 -11400 9280
rect -11100 9020 -10900 9280
rect -10600 9020 -10400 9280
rect -10100 9020 -9900 9280
rect -9600 9020 -9400 9280
rect -9100 9020 -8900 9280
rect -8600 9020 -8400 9280
rect -8100 9020 -7900 9280
rect -7600 9020 -7400 9280
rect -7100 9020 -6900 9280
rect -6600 9020 -6400 9280
rect -6100 9020 -5900 9280
rect -5600 9020 -5400 9280
rect -5100 9020 -4900 9280
rect -4600 9020 -4400 9280
rect -4100 9020 -3900 9280
rect -3600 9020 -3400 9280
rect -3100 9020 -3000 9280
rect -13500 9000 -13380 9020
rect -13120 9000 -12880 9020
rect -12620 9000 -12380 9020
rect -12120 9000 -11880 9020
rect -11620 9000 -11380 9020
rect -11120 9000 -10880 9020
rect -10620 9000 -10380 9020
rect -10120 9000 -9880 9020
rect -9620 9000 -9380 9020
rect -9120 9000 -8880 9020
rect -8620 9000 -8380 9020
rect -8120 9000 -7880 9020
rect -7620 9000 -7380 9020
rect -7120 9000 -6880 9020
rect -6620 9000 -6380 9020
rect -6120 9000 -5880 9020
rect -5620 9000 -5380 9020
rect -5120 9000 -4880 9020
rect -4620 9000 -4380 9020
rect -4120 9000 -3880 9020
rect -3620 9000 -3380 9020
rect -3120 9000 -3000 9020
rect -13500 8900 -3000 9000
rect -5500 8800 -3000 8900
rect -5500 8780 -5380 8800
rect -5120 8780 -4880 8800
rect -4620 8780 -4380 8800
rect -4120 8780 -3880 8800
rect -3620 8780 -3380 8800
rect -3120 8780 -3000 8800
rect -5500 8520 -5400 8780
rect -5100 8520 -4900 8780
rect -4600 8520 -4400 8780
rect -4100 8520 -3900 8780
rect -3600 8520 -3400 8780
rect -3100 8520 -3000 8780
rect -5500 8500 -5380 8520
rect -5120 8500 -4880 8520
rect -4620 8500 -4380 8520
rect -4120 8500 -3880 8520
rect -3620 8500 -3380 8520
rect -3120 8500 -3000 8520
rect -23000 8300 -15500 8400
rect -23000 8280 -22880 8300
rect -22620 8280 -22380 8300
rect -22120 8280 -21880 8300
rect -21620 8280 -21380 8300
rect -21120 8280 -20880 8300
rect -20620 8280 -20380 8300
rect -20120 8280 -19880 8300
rect -19620 8280 -19380 8300
rect -19120 8280 -18880 8300
rect -18620 8280 -18380 8300
rect -18120 8280 -17880 8300
rect -17620 8280 -17380 8300
rect -17120 8280 -16880 8300
rect -16620 8280 -16380 8300
rect -16120 8280 -15880 8300
rect -15620 8280 -15500 8300
rect -23000 8020 -22900 8280
rect -22600 8020 -22400 8280
rect -22100 8020 -21900 8280
rect -21600 8020 -21400 8280
rect -21100 8020 -20900 8280
rect -20600 8020 -20400 8280
rect -20100 8020 -19900 8280
rect -19600 8020 -19400 8280
rect -19100 8020 -18900 8280
rect -18600 8020 -18400 8280
rect -18100 8020 -17900 8280
rect -17600 8020 -17400 8280
rect -17100 8020 -16900 8280
rect -16600 8020 -16400 8280
rect -16100 8020 -15900 8280
rect -15600 8020 -15500 8280
rect -23000 8000 -22880 8020
rect -22620 8000 -22380 8020
rect -22120 8000 -21880 8020
rect -21620 8000 -21380 8020
rect -21120 8000 -20880 8020
rect -20620 8000 -20380 8020
rect -20120 8000 -19880 8020
rect -19620 8000 -19380 8020
rect -19120 8000 -18880 8020
rect -18620 8000 -18380 8020
rect -18120 8000 -17880 8020
rect -17620 8000 -17380 8020
rect -17120 8000 -16880 8020
rect -16620 8000 -16380 8020
rect -16120 8000 -15880 8020
rect -15620 8000 -15500 8020
rect -23000 7800 -15500 8000
rect -11500 8300 -7500 8400
rect -11500 8280 -11380 8300
rect -11120 8280 -10880 8300
rect -10620 8280 -10380 8300
rect -10120 8280 -9880 8300
rect -9620 8280 -9380 8300
rect -9120 8280 -8880 8300
rect -8620 8280 -8380 8300
rect -8120 8280 -7880 8300
rect -7620 8280 -7500 8300
rect -11500 8020 -11400 8280
rect -11100 8020 -10900 8280
rect -10600 8020 -10400 8280
rect -10100 8020 -9900 8280
rect -9600 8020 -9400 8280
rect -9100 8020 -8900 8280
rect -8600 8020 -8400 8280
rect -8100 8020 -7900 8280
rect -7600 8020 -7500 8280
rect -11500 8000 -11380 8020
rect -11120 8000 -10880 8020
rect -10620 8000 -10380 8020
rect -10120 8000 -9880 8020
rect -9620 8000 -9380 8020
rect -9120 8000 -8880 8020
rect -8620 8000 -8380 8020
rect -8120 8000 -7880 8020
rect -7620 8000 -7500 8020
rect -11500 7900 -7500 8000
rect -5500 8300 -3000 8500
rect -5500 8280 -5380 8300
rect -5120 8280 -4880 8300
rect -4620 8280 -4380 8300
rect -4120 8280 -3880 8300
rect -3620 8280 -3380 8300
rect -3120 8280 -3000 8300
rect -5500 8020 -5400 8280
rect -5100 8020 -4900 8280
rect -4600 8020 -4400 8280
rect -4100 8020 -3900 8280
rect -3600 8020 -3400 8280
rect -3100 8020 -3000 8280
rect -5500 8000 -5380 8020
rect -5120 8000 -4880 8020
rect -4620 8000 -4380 8020
rect -4120 8000 -3880 8020
rect -3620 8000 -3380 8020
rect -3120 8000 -3000 8020
rect -23000 7780 -22880 7800
rect -22620 7780 -22380 7800
rect -22120 7780 -21880 7800
rect -21620 7780 -21380 7800
rect -21120 7780 -20880 7800
rect -20620 7780 -20380 7800
rect -20120 7780 -19880 7800
rect -19620 7780 -19380 7800
rect -19120 7780 -18880 7800
rect -18620 7780 -18380 7800
rect -18120 7780 -17880 7800
rect -17620 7780 -17380 7800
rect -17120 7780 -16880 7800
rect -16620 7780 -16380 7800
rect -16120 7780 -15880 7800
rect -15620 7780 -15500 7800
rect -23000 7520 -22900 7780
rect -22600 7520 -22400 7780
rect -22100 7520 -21900 7780
rect -21600 7520 -21400 7780
rect -21100 7520 -20900 7780
rect -20600 7520 -20400 7780
rect -20100 7520 -19900 7780
rect -19600 7520 -19400 7780
rect -19100 7520 -18900 7780
rect -18600 7520 -18400 7780
rect -18100 7520 -17900 7780
rect -17600 7520 -17400 7780
rect -17100 7520 -16900 7780
rect -16600 7520 -16400 7780
rect -16100 7520 -15900 7780
rect -15600 7520 -15500 7780
rect -23000 7500 -22880 7520
rect -22620 7500 -22380 7520
rect -22120 7500 -21880 7520
rect -21620 7500 -21380 7520
rect -21120 7500 -20880 7520
rect -20620 7500 -20380 7520
rect -20120 7500 -19880 7520
rect -19620 7500 -19380 7520
rect -19120 7500 -18880 7520
rect -18620 7500 -18380 7520
rect -18120 7500 -17880 7520
rect -17620 7500 -17380 7520
rect -17120 7500 -16880 7520
rect -16620 7500 -16380 7520
rect -16120 7500 -15880 7520
rect -15620 7500 -15500 7520
rect -23000 7300 -15500 7500
rect -23000 7280 -22880 7300
rect -22620 7280 -22380 7300
rect -22120 7280 -21880 7300
rect -21620 7280 -21380 7300
rect -21120 7280 -20880 7300
rect -20620 7280 -20380 7300
rect -20120 7280 -19880 7300
rect -19620 7280 -19380 7300
rect -19120 7280 -18880 7300
rect -18620 7280 -18380 7300
rect -18120 7280 -17880 7300
rect -17620 7280 -17380 7300
rect -17120 7280 -16880 7300
rect -16620 7280 -16380 7300
rect -16120 7280 -15880 7300
rect -15620 7280 -15500 7300
rect -23000 7020 -22900 7280
rect -22600 7020 -22400 7280
rect -22100 7020 -21900 7280
rect -21600 7020 -21400 7280
rect -21100 7020 -20900 7280
rect -20600 7020 -20400 7280
rect -20100 7020 -19900 7280
rect -19600 7020 -19400 7280
rect -19100 7020 -18900 7280
rect -18600 7020 -18400 7280
rect -18100 7020 -17900 7280
rect -17600 7020 -17400 7280
rect -17100 7020 -16900 7280
rect -16600 7020 -16400 7280
rect -16100 7020 -15900 7280
rect -15600 7020 -15500 7280
rect -23000 7000 -22880 7020
rect -22620 7000 -22380 7020
rect -22120 7000 -21880 7020
rect -21620 7000 -21380 7020
rect -21120 7000 -20880 7020
rect -20620 7000 -20380 7020
rect -20120 7000 -19880 7020
rect -19620 7000 -19380 7020
rect -19120 7000 -18880 7020
rect -18620 7000 -18380 7020
rect -18120 7000 -17880 7020
rect -17620 7000 -17380 7020
rect -17120 7000 -16880 7020
rect -16620 7000 -16380 7020
rect -16120 7000 -15880 7020
rect -15620 7000 -15500 7020
rect -23000 6800 -15500 7000
rect -23000 6780 -22880 6800
rect -22620 6780 -22380 6800
rect -22120 6780 -21880 6800
rect -21620 6780 -21380 6800
rect -21120 6780 -20880 6800
rect -20620 6780 -20380 6800
rect -20120 6780 -19880 6800
rect -19620 6780 -19380 6800
rect -19120 6780 -18880 6800
rect -18620 6780 -18380 6800
rect -18120 6780 -17880 6800
rect -17620 6780 -17380 6800
rect -17120 6780 -16880 6800
rect -16620 6780 -16380 6800
rect -16120 6780 -15880 6800
rect -15620 6780 -15500 6800
rect -23000 6520 -22900 6780
rect -22600 6520 -22400 6780
rect -22100 6520 -21900 6780
rect -21600 6520 -21400 6780
rect -21100 6520 -20900 6780
rect -20600 6520 -20400 6780
rect -20100 6520 -19900 6780
rect -19600 6520 -19400 6780
rect -19100 6520 -18900 6780
rect -18600 6520 -18400 6780
rect -18100 6520 -17900 6780
rect -17600 6520 -17400 6780
rect -17100 6520 -16900 6780
rect -16600 6520 -16400 6780
rect -16100 6520 -15900 6780
rect -15600 6520 -15500 6780
rect -23000 6500 -22880 6520
rect -22620 6500 -22380 6520
rect -22120 6500 -21880 6520
rect -21620 6500 -21380 6520
rect -21120 6500 -20880 6520
rect -20620 6500 -20380 6520
rect -20120 6500 -19880 6520
rect -19620 6500 -19380 6520
rect -19120 6500 -18880 6520
rect -18620 6500 -18380 6520
rect -18120 6500 -17880 6520
rect -17620 6500 -17380 6520
rect -17120 6500 -16880 6520
rect -16620 6500 -16380 6520
rect -16120 6500 -15880 6520
rect -15620 6500 -15500 6520
rect -23000 6300 -15500 6500
rect -23000 6280 -22880 6300
rect -22620 6280 -22380 6300
rect -22120 6280 -21880 6300
rect -21620 6280 -21380 6300
rect -21120 6280 -20880 6300
rect -20620 6280 -20380 6300
rect -20120 6280 -19880 6300
rect -19620 6280 -19380 6300
rect -19120 6280 -18880 6300
rect -18620 6280 -18380 6300
rect -18120 6280 -17880 6300
rect -17620 6280 -17380 6300
rect -17120 6280 -16880 6300
rect -16620 6280 -16380 6300
rect -16120 6280 -15880 6300
rect -15620 6280 -15500 6300
rect -23000 6020 -22900 6280
rect -22600 6020 -22400 6280
rect -22100 6020 -21900 6280
rect -21600 6020 -21400 6280
rect -21100 6020 -20900 6280
rect -20600 6020 -20400 6280
rect -20100 6020 -19900 6280
rect -19600 6020 -19400 6280
rect -19100 6020 -18900 6280
rect -18600 6020 -18400 6280
rect -18100 6020 -17900 6280
rect -17600 6020 -17400 6280
rect -17100 6020 -16900 6280
rect -16600 6020 -16400 6280
rect -16100 6020 -15900 6280
rect -15600 6020 -15500 6280
rect -23000 6000 -22880 6020
rect -22620 6000 -22380 6020
rect -22120 6000 -21880 6020
rect -21620 6000 -21380 6020
rect -21120 6000 -20880 6020
rect -20620 6000 -20380 6020
rect -20120 6000 -19880 6020
rect -19620 6000 -19380 6020
rect -19120 6000 -18880 6020
rect -18620 6000 -18380 6020
rect -18120 6000 -17880 6020
rect -17620 6000 -17380 6020
rect -17120 6000 -16880 6020
rect -16620 6000 -16380 6020
rect -16120 6000 -15880 6020
rect -15620 6000 -15500 6020
rect -23000 5900 -15500 6000
rect -5500 7800 -3000 8000
rect -5500 7780 -5380 7800
rect -5120 7780 -4880 7800
rect -4620 7780 -4380 7800
rect -4120 7780 -3880 7800
rect -3620 7780 -3380 7800
rect -3120 7780 -3000 7800
rect -5500 7520 -5400 7780
rect -5100 7520 -4900 7780
rect -4600 7520 -4400 7780
rect -4100 7520 -3900 7780
rect -3600 7520 -3400 7780
rect -3100 7520 -3000 7780
rect -5500 7500 -5380 7520
rect -5120 7500 -4880 7520
rect -4620 7500 -4380 7520
rect -4120 7500 -3880 7520
rect -3620 7500 -3380 7520
rect -3120 7500 -3000 7520
rect -5500 7300 -3000 7500
rect -5500 7280 -5380 7300
rect -5120 7280 -4880 7300
rect -4620 7280 -4380 7300
rect -4120 7280 -3880 7300
rect -3620 7280 -3380 7300
rect -3120 7280 -3000 7300
rect -5500 7020 -5400 7280
rect -5100 7020 -4900 7280
rect -4600 7020 -4400 7280
rect -4100 7020 -3900 7280
rect -3600 7020 -3400 7280
rect -3100 7020 -3000 7280
rect -5500 7000 -5380 7020
rect -5120 7000 -4880 7020
rect -4620 7000 -4380 7020
rect -4120 7000 -3880 7020
rect -3620 7000 -3380 7020
rect -3120 7000 -3000 7020
rect -5500 6800 -3000 7000
rect -5500 6780 -5380 6800
rect -5120 6780 -4880 6800
rect -4620 6780 -4380 6800
rect -4120 6780 -3880 6800
rect -3620 6780 -3380 6800
rect -3120 6780 -3000 6800
rect -5500 6520 -5400 6780
rect -5100 6520 -4900 6780
rect -4600 6520 -4400 6780
rect -4100 6520 -3900 6780
rect -3600 6520 -3400 6780
rect -3100 6520 -3000 6780
rect -5500 6500 -5380 6520
rect -5120 6500 -4880 6520
rect -4620 6500 -4380 6520
rect -4120 6500 -3880 6520
rect -3620 6500 -3380 6520
rect -3120 6500 -3000 6520
rect -5500 6300 -3000 6500
rect -5500 6280 -5380 6300
rect -5120 6280 -4880 6300
rect -4620 6280 -4380 6300
rect -4120 6280 -3880 6300
rect -3620 6280 -3380 6300
rect -3120 6280 -3000 6300
rect -5500 6020 -5400 6280
rect -5100 6020 -4900 6280
rect -4600 6020 -4400 6280
rect -4100 6020 -3900 6280
rect -3600 6020 -3400 6280
rect -3100 6020 -3000 6280
rect -5500 6000 -5380 6020
rect -5120 6000 -4880 6020
rect -4620 6000 -4380 6020
rect -4120 6000 -3880 6020
rect -3620 6000 -3380 6020
rect -3120 6000 -3000 6020
rect -5500 5900 -3000 6000
rect -23000 5800 -21000 5900
rect -23000 5780 -22880 5800
rect -22620 5780 -22380 5800
rect -22120 5780 -21880 5800
rect -21620 5780 -21380 5800
rect -21120 5780 -21000 5800
rect -23000 5520 -22900 5780
rect -22600 5520 -22400 5780
rect -22100 5520 -21900 5780
rect -21600 5520 -21400 5780
rect -21100 5520 -21000 5780
rect -23000 5500 -22880 5520
rect -22620 5500 -22380 5520
rect -22120 5500 -21880 5520
rect -21620 5500 -21380 5520
rect -21120 5500 -21000 5520
rect -23000 5300 -21000 5500
rect -23000 5280 -22880 5300
rect -22620 5280 -22380 5300
rect -22120 5280 -21880 5300
rect -21620 5280 -21380 5300
rect -21120 5280 -21000 5300
rect -23000 5020 -22900 5280
rect -22600 5020 -22400 5280
rect -22100 5020 -21900 5280
rect -21600 5020 -21400 5280
rect -21100 5020 -21000 5280
rect -23000 5000 -22880 5020
rect -22620 5000 -22380 5020
rect -22120 5000 -21880 5020
rect -21620 5000 -21380 5020
rect -21120 5000 -21000 5020
rect -23000 4900 -21000 5000
rect -25000 4800 -21000 4900
rect -25000 4780 -24880 4800
rect -24620 4780 -24380 4800
rect -24120 4780 -23880 4800
rect -23620 4780 -23380 4800
rect -23120 4780 -22880 4800
rect -22620 4780 -22380 4800
rect -22120 4780 -21880 4800
rect -21620 4780 -21380 4800
rect -21120 4780 -21000 4800
rect -25000 4520 -24900 4780
rect -24600 4520 -24400 4780
rect -24100 4520 -23900 4780
rect -23600 4520 -23400 4780
rect -23100 4520 -22900 4780
rect -22600 4520 -22400 4780
rect -22100 4520 -21900 4780
rect -21600 4520 -21400 4780
rect -21100 4520 -21000 4780
rect -25000 4500 -24880 4520
rect -24620 4500 -24380 4520
rect -24120 4500 -23880 4520
rect -23620 4500 -23380 4520
rect -23120 4500 -22880 4520
rect -22620 4500 -22380 4520
rect -22120 4500 -21880 4520
rect -21620 4500 -21380 4520
rect -21120 4500 -21000 4520
rect -25000 4300 -21000 4500
rect -25000 4280 -24880 4300
rect -24620 4280 -24380 4300
rect -24120 4280 -23880 4300
rect -23620 4280 -23380 4300
rect -23120 4280 -22880 4300
rect -22620 4280 -22380 4300
rect -22120 4280 -21880 4300
rect -21620 4280 -21380 4300
rect -21120 4280 -21000 4300
rect -25000 4020 -24900 4280
rect -24600 4020 -24400 4280
rect -24100 4020 -23900 4280
rect -23600 4020 -23400 4280
rect -23100 4020 -22900 4280
rect -22600 4020 -22400 4280
rect -22100 4020 -21900 4280
rect -21600 4020 -21400 4280
rect -21100 4020 -21000 4280
rect -25000 4000 -24880 4020
rect -24620 4000 -24380 4020
rect -24120 4000 -23880 4020
rect -23620 4000 -23380 4020
rect -23120 4000 -22880 4020
rect -22620 4000 -22380 4020
rect -22120 4000 -21880 4020
rect -21620 4000 -21380 4020
rect -21120 4000 -21000 4020
rect -25000 3800 -21000 4000
rect -25000 3780 -24880 3800
rect -24620 3780 -24380 3800
rect -24120 3780 -23880 3800
rect -23620 3780 -23380 3800
rect -23120 3780 -22880 3800
rect -22620 3780 -22380 3800
rect -22120 3780 -21880 3800
rect -21620 3780 -21380 3800
rect -21120 3780 -21000 3800
rect -25000 3520 -24900 3780
rect -24600 3520 -24400 3780
rect -24100 3520 -23900 3780
rect -23600 3520 -23400 3780
rect -23100 3520 -22900 3780
rect -22600 3520 -22400 3780
rect -22100 3520 -21900 3780
rect -21600 3520 -21400 3780
rect -21100 3520 -21000 3780
rect -25000 3500 -24880 3520
rect -24620 3500 -24380 3520
rect -24120 3500 -23880 3520
rect -23620 3500 -23380 3520
rect -23120 3500 -22880 3520
rect -22620 3500 -22380 3520
rect -22120 3500 -21880 3520
rect -21620 3500 -21380 3520
rect -21120 3500 -21000 3520
rect -25000 3300 -21000 3500
rect -25000 3280 -24880 3300
rect -24620 3280 -24380 3300
rect -24120 3280 -23880 3300
rect -23620 3280 -23380 3300
rect -23120 3280 -22880 3300
rect -22620 3280 -22380 3300
rect -22120 3280 -21880 3300
rect -21620 3280 -21380 3300
rect -21120 3280 -21000 3300
rect -25000 3020 -24900 3280
rect -24600 3020 -24400 3280
rect -24100 3020 -23900 3280
rect -23600 3020 -23400 3280
rect -23100 3020 -22900 3280
rect -22600 3020 -22400 3280
rect -22100 3020 -21900 3280
rect -21600 3020 -21400 3280
rect -21100 3020 -21000 3280
rect -25000 3000 -24880 3020
rect -24620 3000 -24380 3020
rect -24120 3000 -23880 3020
rect -23620 3000 -23380 3020
rect -23120 3000 -22880 3020
rect -22620 3000 -22380 3020
rect -22120 3000 -21880 3020
rect -21620 3000 -21380 3020
rect -21120 3000 -21000 3020
rect -25000 2800 -21000 3000
rect -25000 2780 -24880 2800
rect -24620 2780 -24380 2800
rect -24120 2780 -23880 2800
rect -23620 2780 -23380 2800
rect -23120 2780 -22880 2800
rect -22620 2780 -22380 2800
rect -22120 2780 -21880 2800
rect -21620 2780 -21380 2800
rect -21120 2780 -21000 2800
rect -25000 2520 -24900 2780
rect -24600 2520 -24400 2780
rect -24100 2520 -23900 2780
rect -23600 2520 -23400 2780
rect -23100 2520 -22900 2780
rect -22600 2520 -22400 2780
rect -22100 2520 -21900 2780
rect -21600 2520 -21400 2780
rect -21100 2520 -21000 2780
rect -25000 2500 -24880 2520
rect -24620 2500 -24380 2520
rect -24120 2500 -23880 2520
rect -23620 2500 -23380 2520
rect -23120 2500 -22880 2520
rect -22620 2500 -22380 2520
rect -22120 2500 -21880 2520
rect -21620 2500 -21380 2520
rect -21120 2500 -21000 2520
rect -25000 2300 -21000 2500
rect -25000 2280 -24880 2300
rect -24620 2280 -24380 2300
rect -24120 2280 -23880 2300
rect -23620 2280 -23380 2300
rect -23120 2280 -22880 2300
rect -22620 2280 -22380 2300
rect -22120 2280 -21880 2300
rect -21620 2280 -21380 2300
rect -21120 2280 -21000 2300
rect -25000 2020 -24900 2280
rect -24600 2020 -24400 2280
rect -24100 2020 -23900 2280
rect -23600 2020 -23400 2280
rect -23100 2020 -22900 2280
rect -22600 2020 -22400 2280
rect -22100 2020 -21900 2280
rect -21600 2020 -21400 2280
rect -21100 2020 -21000 2280
rect -25000 2000 -24880 2020
rect -24620 2000 -24380 2020
rect -24120 2000 -23880 2020
rect -23620 2000 -23380 2020
rect -23120 2000 -22880 2020
rect -22620 2000 -22380 2020
rect -22120 2000 -21880 2020
rect -21620 2000 -21380 2020
rect -21120 2000 -21000 2020
rect -25000 1800 -21000 2000
rect -25000 1780 -24880 1800
rect -24620 1780 -24380 1800
rect -24120 1780 -23880 1800
rect -23620 1780 -23380 1800
rect -23120 1780 -22880 1800
rect -22620 1780 -22380 1800
rect -22120 1780 -21880 1800
rect -21620 1780 -21380 1800
rect -21120 1780 -21000 1800
rect -25000 1520 -24900 1780
rect -24600 1520 -24400 1780
rect -24100 1520 -23900 1780
rect -23600 1520 -23400 1780
rect -23100 1520 -22900 1780
rect -22600 1520 -22400 1780
rect -22100 1520 -21900 1780
rect -21600 1520 -21400 1780
rect -21100 1520 -21000 1780
rect -25000 1500 -24880 1520
rect -24620 1500 -24380 1520
rect -24120 1500 -23880 1520
rect -23620 1500 -23380 1520
rect -23120 1500 -22880 1520
rect -22620 1500 -22380 1520
rect -22120 1500 -21880 1520
rect -21620 1500 -21380 1520
rect -21120 1500 -21000 1520
rect -25000 1300 -21000 1500
rect -25000 1280 -24880 1300
rect -24620 1280 -24380 1300
rect -24120 1280 -23880 1300
rect -23620 1280 -23380 1300
rect -23120 1280 -22880 1300
rect -22620 1280 -22380 1300
rect -22120 1280 -21880 1300
rect -21620 1280 -21380 1300
rect -21120 1280 -21000 1300
rect -25000 1020 -24900 1280
rect -24600 1020 -24400 1280
rect -24100 1020 -23900 1280
rect -23600 1020 -23400 1280
rect -23100 1020 -22900 1280
rect -22600 1020 -22400 1280
rect -22100 1020 -21900 1280
rect -21600 1020 -21400 1280
rect -21100 1020 -21000 1280
rect -25000 1000 -24880 1020
rect -24620 1000 -24380 1020
rect -24120 1000 -23880 1020
rect -23620 1000 -23380 1020
rect -23120 1000 -22880 1020
rect -22620 1000 -22380 1020
rect -22120 1000 -21880 1020
rect -21620 1000 -21380 1020
rect -21120 1000 -21000 1020
rect -25000 800 -21000 1000
rect -25000 780 -24880 800
rect -24620 780 -24380 800
rect -24120 780 -23880 800
rect -23620 780 -23380 800
rect -23120 780 -22880 800
rect -22620 780 -22380 800
rect -22120 780 -21880 800
rect -21620 780 -21380 800
rect -21120 780 -21000 800
rect -25000 520 -24900 780
rect -24600 520 -24400 780
rect -24100 520 -23900 780
rect -23600 520 -23400 780
rect -23100 520 -22900 780
rect -22600 520 -22400 780
rect -22100 520 -21900 780
rect -21600 520 -21400 780
rect -21100 520 -21000 780
rect -25000 500 -24880 520
rect -24620 500 -24380 520
rect -24120 500 -23880 520
rect -23620 500 -23380 520
rect -23120 500 -22880 520
rect -22620 500 -22380 520
rect -22120 500 -21880 520
rect -21620 500 -21380 520
rect -21120 500 -21000 520
rect -25000 300 -21000 500
rect 13000 2300 15500 2400
rect 13000 2280 13120 2300
rect 13380 2280 13620 2300
rect 13880 2280 14120 2300
rect 14380 2280 14620 2300
rect 14880 2280 15120 2300
rect 15380 2280 15500 2300
rect 13000 2020 13100 2280
rect 13400 2020 13600 2280
rect 13900 2020 14100 2280
rect 14400 2020 14600 2280
rect 14900 2020 15100 2280
rect 15400 2020 15500 2280
rect 13000 2000 13120 2020
rect 13380 2000 13620 2020
rect 13880 2000 14120 2020
rect 14380 2000 14620 2020
rect 14880 2000 15120 2020
rect 15380 2000 15500 2020
rect 13000 1800 15500 2000
rect 13000 1780 13120 1800
rect 13380 1780 13620 1800
rect 13880 1780 14120 1800
rect 14380 1780 14620 1800
rect 14880 1780 15120 1800
rect 15380 1780 15500 1800
rect 13000 1520 13100 1780
rect 13400 1520 13600 1780
rect 13900 1520 14100 1780
rect 14400 1520 14600 1780
rect 14900 1520 15100 1780
rect 15400 1520 15500 1780
rect 13000 1500 13120 1520
rect 13380 1500 13620 1520
rect 13880 1500 14120 1520
rect 14380 1500 14620 1520
rect 14880 1500 15120 1520
rect 15380 1500 15500 1520
rect 13000 1300 15500 1500
rect 13000 1280 13120 1300
rect 13380 1280 13620 1300
rect 13880 1280 14120 1300
rect 14380 1280 14620 1300
rect 14880 1280 15120 1300
rect 15380 1280 15500 1300
rect 13000 1020 13100 1280
rect 13400 1020 13600 1280
rect 13900 1020 14100 1280
rect 14400 1020 14600 1280
rect 14900 1020 15100 1280
rect 15400 1020 15500 1280
rect 13000 1000 13120 1020
rect 13380 1000 13620 1020
rect 13880 1000 14120 1020
rect 14380 1000 14620 1020
rect 14880 1000 15120 1020
rect 15380 1000 15500 1020
rect 13000 800 15500 1000
rect 13000 780 13120 800
rect 13380 780 13620 800
rect 13880 780 14120 800
rect 14380 780 14620 800
rect 14880 780 15120 800
rect 15380 780 15500 800
rect 13000 520 13100 780
rect 13400 520 13600 780
rect 13900 520 14100 780
rect 14400 520 14600 780
rect 14900 520 15100 780
rect 15400 520 15500 780
rect 13000 500 13120 520
rect 13380 500 13620 520
rect 13880 500 14120 520
rect 14380 500 14620 520
rect 14880 500 15120 520
rect 15380 500 15500 520
rect 13000 400 15500 500
rect 17500 1300 19500 1400
rect 17500 1280 17620 1300
rect 17880 1280 18120 1300
rect 18380 1280 18620 1300
rect 18880 1280 19120 1300
rect 19380 1280 19500 1300
rect 17500 1020 17600 1280
rect 17900 1020 18100 1280
rect 18400 1020 18600 1280
rect 18900 1020 19100 1280
rect 19400 1020 19500 1280
rect 17500 1000 17620 1020
rect 17880 1000 18120 1020
rect 18380 1000 18620 1020
rect 18880 1000 19120 1020
rect 19380 1000 19500 1020
rect 17500 800 19500 1000
rect 17500 780 17620 800
rect 17880 780 18120 800
rect 18380 780 18620 800
rect 18880 780 19120 800
rect 19380 780 19500 800
rect 17500 520 17600 780
rect 17900 520 18100 780
rect 18400 520 18600 780
rect 18900 520 19100 780
rect 19400 520 19500 780
rect 17500 500 17620 520
rect 17880 500 18120 520
rect 18380 500 18620 520
rect 18880 500 19120 520
rect 19380 500 19500 520
rect -25000 280 -24880 300
rect -24620 280 -24380 300
rect -24120 280 -23880 300
rect -23620 280 -23380 300
rect -23120 280 -22880 300
rect -22620 280 -22380 300
rect -22120 280 -21880 300
rect -21620 280 -21380 300
rect -21120 280 -21000 300
rect -25000 20 -24900 280
rect -24600 20 -24400 280
rect -24100 20 -23900 280
rect -23600 20 -23400 280
rect -23100 20 -22900 280
rect -22600 20 -22400 280
rect -22100 20 -21900 280
rect -21600 20 -21400 280
rect -21100 20 -21000 280
rect -25000 0 -24880 20
rect -24620 0 -24380 20
rect -24120 0 -23880 20
rect -23620 0 -23380 20
rect -23120 0 -22880 20
rect -22620 0 -22380 20
rect -22120 0 -21880 20
rect -21620 0 -21380 20
rect -21120 0 -21000 20
rect -25000 -200 -21000 0
rect -25000 -220 -24880 -200
rect -24620 -220 -24380 -200
rect -24120 -220 -23880 -200
rect -23620 -220 -23380 -200
rect -23120 -220 -22880 -200
rect -22620 -220 -22380 -200
rect -22120 -220 -21880 -200
rect -21620 -220 -21380 -200
rect -21120 -220 -21000 -200
rect -25000 -480 -24900 -220
rect -24600 -480 -24400 -220
rect -24100 -480 -23900 -220
rect -23600 -480 -23400 -220
rect -23100 -480 -22900 -220
rect -22600 -480 -22400 -220
rect -22100 -480 -21900 -220
rect -21600 -480 -21400 -220
rect -21100 -480 -21000 -220
rect -25000 -500 -24880 -480
rect -24620 -500 -24380 -480
rect -24120 -500 -23880 -480
rect -23620 -500 -23380 -480
rect -23120 -500 -22880 -480
rect -22620 -500 -22380 -480
rect -22120 -500 -21880 -480
rect -21620 -500 -21380 -480
rect -21120 -500 -21000 -480
rect -25000 -700 -21000 -500
rect -25000 -720 -24880 -700
rect -24620 -720 -24380 -700
rect -24120 -720 -23880 -700
rect -23620 -720 -23380 -700
rect -23120 -720 -22880 -700
rect -22620 -720 -22380 -700
rect -22120 -720 -21880 -700
rect -21620 -720 -21380 -700
rect -21120 -720 -21000 -700
rect -25000 -980 -24900 -720
rect -24600 -980 -24400 -720
rect -24100 -980 -23900 -720
rect -23600 -980 -23400 -720
rect -23100 -980 -22900 -720
rect -22600 -980 -22400 -720
rect -22100 -980 -21900 -720
rect -21600 -980 -21400 -720
rect -21100 -980 -21000 -720
rect -25000 -1000 -24880 -980
rect -24620 -1000 -24380 -980
rect -24120 -1000 -23880 -980
rect -23620 -1000 -23380 -980
rect -23120 -1000 -22880 -980
rect -22620 -1000 -22380 -980
rect -22120 -1000 -21880 -980
rect -21620 -1000 -21380 -980
rect -21120 -1000 -21000 -980
rect -25000 -1200 -21000 -1000
rect -25000 -1220 -24880 -1200
rect -24620 -1220 -24380 -1200
rect -24120 -1220 -23880 -1200
rect -23620 -1220 -23380 -1200
rect -23120 -1220 -22880 -1200
rect -22620 -1220 -22380 -1200
rect -22120 -1220 -21880 -1200
rect -21620 -1220 -21380 -1200
rect -21120 -1220 -21000 -1200
rect -25000 -1480 -24900 -1220
rect -24600 -1480 -24400 -1220
rect -24100 -1480 -23900 -1220
rect -23600 -1480 -23400 -1220
rect -23100 -1480 -22900 -1220
rect -22600 -1480 -22400 -1220
rect -22100 -1480 -21900 -1220
rect -21600 -1480 -21400 -1220
rect -21100 -1480 -21000 -1220
rect -25000 -1500 -24880 -1480
rect -24620 -1500 -24380 -1480
rect -24120 -1500 -23880 -1480
rect -23620 -1500 -23380 -1480
rect -23120 -1500 -22880 -1480
rect -22620 -1500 -22380 -1480
rect -22120 -1500 -21880 -1480
rect -21620 -1500 -21380 -1480
rect -21120 -1500 -21000 -1480
rect -25000 -1700 -21000 -1500
rect -25000 -1720 -24880 -1700
rect -24620 -1720 -24380 -1700
rect -24120 -1720 -23880 -1700
rect -23620 -1720 -23380 -1700
rect -23120 -1720 -22880 -1700
rect -22620 -1720 -22380 -1700
rect -22120 -1720 -21880 -1700
rect -21620 -1720 -21380 -1700
rect -21120 -1720 -21000 -1700
rect -25000 -1980 -24900 -1720
rect -24600 -1980 -24400 -1720
rect -24100 -1980 -23900 -1720
rect -23600 -1980 -23400 -1720
rect -23100 -1980 -22900 -1720
rect -22600 -1980 -22400 -1720
rect -22100 -1980 -21900 -1720
rect -21600 -1980 -21400 -1720
rect -21100 -1980 -21000 -1720
rect -25000 -2000 -24880 -1980
rect -24620 -2000 -24380 -1980
rect -24120 -2000 -23880 -1980
rect -23620 -2000 -23380 -1980
rect -23120 -2000 -22880 -1980
rect -22620 -2000 -22380 -1980
rect -22120 -2000 -21880 -1980
rect -21620 -2000 -21380 -1980
rect -21120 -2000 -21000 -1980
rect -25000 -2200 -21000 -2000
rect -25000 -2220 -24880 -2200
rect -24620 -2220 -24380 -2200
rect -24120 -2220 -23880 -2200
rect -23620 -2220 -23380 -2200
rect -23120 -2220 -22880 -2200
rect -22620 -2220 -22380 -2200
rect -22120 -2220 -21880 -2200
rect -21620 -2220 -21380 -2200
rect -21120 -2220 -21000 -2200
rect -25000 -2480 -24900 -2220
rect -24600 -2480 -24400 -2220
rect -24100 -2480 -23900 -2220
rect -23600 -2480 -23400 -2220
rect -23100 -2480 -22900 -2220
rect -22600 -2480 -22400 -2220
rect -22100 -2480 -21900 -2220
rect -21600 -2480 -21400 -2220
rect -21100 -2480 -21000 -2220
rect -25000 -2500 -24880 -2480
rect -24620 -2500 -24380 -2480
rect -24120 -2500 -23880 -2480
rect -23620 -2500 -23380 -2480
rect -23120 -2500 -22880 -2480
rect -22620 -2500 -22380 -2480
rect -22120 -2500 -21880 -2480
rect -21620 -2500 -21380 -2480
rect -21120 -2500 -21000 -2480
rect -25000 -2700 -21000 -2500
rect -25000 -2720 -24880 -2700
rect -24620 -2720 -24380 -2700
rect -24120 -2720 -23880 -2700
rect -23620 -2720 -23380 -2700
rect -23120 -2720 -22880 -2700
rect -22620 -2720 -22380 -2700
rect -22120 -2720 -21880 -2700
rect -21620 -2720 -21380 -2700
rect -21120 -2720 -21000 -2700
rect -25000 -2980 -24900 -2720
rect -24600 -2980 -24400 -2720
rect -24100 -2980 -23900 -2720
rect -23600 -2980 -23400 -2720
rect -23100 -2980 -22900 -2720
rect -22600 -2980 -22400 -2720
rect -22100 -2980 -21900 -2720
rect -21600 -2980 -21400 -2720
rect -21100 -2980 -21000 -2720
rect -25000 -3000 -24880 -2980
rect -24620 -3000 -24380 -2980
rect -24120 -3000 -23880 -2980
rect -23620 -3000 -23380 -2980
rect -23120 -3000 -22880 -2980
rect -22620 -3000 -22380 -2980
rect -22120 -3000 -21880 -2980
rect -21620 -3000 -21380 -2980
rect -21120 -3000 -21000 -2980
rect -25000 -3100 -21000 -3000
rect 12000 300 17000 400
rect 12000 280 12120 300
rect 12380 280 12620 300
rect 12880 280 13120 300
rect 13380 280 13620 300
rect 13880 280 14120 300
rect 14380 280 14620 300
rect 14880 280 15120 300
rect 15380 280 15620 300
rect 15880 280 16120 300
rect 16380 280 16620 300
rect 16880 280 17000 300
rect 12000 20 12100 280
rect 12400 20 12600 280
rect 12900 20 13100 280
rect 13400 20 13600 280
rect 13900 20 14100 280
rect 14400 20 14600 280
rect 14900 20 15100 280
rect 15400 20 15600 280
rect 15900 20 16100 280
rect 16400 20 16600 280
rect 16900 20 17000 280
rect 12000 0 12120 20
rect 12380 0 12620 20
rect 12880 0 13120 20
rect 13380 0 13620 20
rect 13880 0 14120 20
rect 14380 0 14620 20
rect 14880 0 15120 20
rect 15380 0 15620 20
rect 15880 0 16120 20
rect 16380 0 16620 20
rect 16880 0 17000 20
rect 12000 -200 17000 0
rect 12000 -220 12120 -200
rect 12380 -220 12620 -200
rect 12880 -220 13120 -200
rect 13380 -220 13620 -200
rect 13880 -220 14120 -200
rect 14380 -220 14620 -200
rect 14880 -220 15120 -200
rect 15380 -220 15620 -200
rect 15880 -220 16120 -200
rect 16380 -220 16620 -200
rect 16880 -220 17000 -200
rect 12000 -480 12100 -220
rect 12400 -480 12600 -220
rect 12900 -480 13100 -220
rect 13400 -480 13600 -220
rect 13900 -480 14100 -220
rect 14400 -480 14600 -220
rect 14900 -480 15100 -220
rect 15400 -480 15600 -220
rect 15900 -480 16100 -220
rect 16400 -480 16600 -220
rect 16900 -480 17000 -220
rect 12000 -500 12120 -480
rect 12380 -500 12620 -480
rect 12880 -500 13120 -480
rect 13380 -500 13620 -480
rect 13880 -500 14120 -480
rect 14380 -500 14620 -480
rect 14880 -500 15120 -480
rect 15380 -500 15620 -480
rect 15880 -500 16120 -480
rect 16380 -500 16620 -480
rect 16880 -500 17000 -480
rect 12000 -700 17000 -500
rect 12000 -720 12120 -700
rect 12380 -720 12620 -700
rect 12880 -720 13120 -700
rect 13380 -720 13620 -700
rect 13880 -720 14120 -700
rect 14380 -720 14620 -700
rect 14880 -720 15120 -700
rect 15380 -720 15620 -700
rect 15880 -720 16120 -700
rect 16380 -720 16620 -700
rect 16880 -720 17000 -700
rect 12000 -980 12100 -720
rect 12400 -980 12600 -720
rect 12900 -980 13100 -720
rect 13400 -980 13600 -720
rect 13900 -980 14100 -720
rect 14400 -980 14600 -720
rect 14900 -980 15100 -720
rect 15400 -980 15600 -720
rect 15900 -980 16100 -720
rect 16400 -980 16600 -720
rect 16900 -980 17000 -720
rect 12000 -1000 12120 -980
rect 12380 -1000 12620 -980
rect 12880 -1000 13120 -980
rect 13380 -1000 13620 -980
rect 13880 -1000 14120 -980
rect 14380 -1000 14620 -980
rect 14880 -1000 15120 -980
rect 15380 -1000 15620 -980
rect 15880 -1000 16120 -980
rect 16380 -1000 16620 -980
rect 16880 -1000 17000 -980
rect 12000 -1200 17000 -1000
rect 12000 -1220 12120 -1200
rect 12380 -1220 12620 -1200
rect 12880 -1220 13120 -1200
rect 13380 -1220 13620 -1200
rect 13880 -1220 14120 -1200
rect 14380 -1220 14620 -1200
rect 14880 -1220 15120 -1200
rect 15380 -1220 15620 -1200
rect 15880 -1220 16120 -1200
rect 16380 -1220 16620 -1200
rect 16880 -1220 17000 -1200
rect 12000 -1480 12100 -1220
rect 12400 -1480 12600 -1220
rect 12900 -1480 13100 -1220
rect 13400 -1480 13600 -1220
rect 13900 -1480 14100 -1220
rect 14400 -1480 14600 -1220
rect 14900 -1480 15100 -1220
rect 15400 -1480 15600 -1220
rect 15900 -1480 16100 -1220
rect 16400 -1480 16600 -1220
rect 16900 -1480 17000 -1220
rect 12000 -1500 12120 -1480
rect 12380 -1500 12620 -1480
rect 12880 -1500 13120 -1480
rect 13380 -1500 13620 -1480
rect 13880 -1500 14120 -1480
rect 14380 -1500 14620 -1480
rect 14880 -1500 15120 -1480
rect 15380 -1500 15620 -1480
rect 15880 -1500 16120 -1480
rect 16380 -1500 16620 -1480
rect 16880 -1500 17000 -1480
rect 12000 -1700 17000 -1500
rect 12000 -1720 12120 -1700
rect 12380 -1720 12620 -1700
rect 12880 -1720 13120 -1700
rect 13380 -1720 13620 -1700
rect 13880 -1720 14120 -1700
rect 14380 -1720 14620 -1700
rect 14880 -1720 15120 -1700
rect 15380 -1720 15620 -1700
rect 15880 -1720 16120 -1700
rect 16380 -1720 16620 -1700
rect 16880 -1720 17000 -1700
rect 12000 -1980 12100 -1720
rect 12400 -1980 12600 -1720
rect 12900 -1980 13100 -1720
rect 13400 -1980 13600 -1720
rect 13900 -1980 14100 -1720
rect 14400 -1980 14600 -1720
rect 14900 -1980 15100 -1720
rect 15400 -1980 15600 -1720
rect 15900 -1980 16100 -1720
rect 16400 -1980 16600 -1720
rect 16900 -1980 17000 -1720
rect 12000 -2000 12120 -1980
rect 12380 -2000 12620 -1980
rect 12880 -2000 13120 -1980
rect 13380 -2000 13620 -1980
rect 13880 -2000 14120 -1980
rect 14380 -2000 14620 -1980
rect 14880 -2000 15120 -1980
rect 15380 -2000 15620 -1980
rect 15880 -2000 16120 -1980
rect 16380 -2000 16620 -1980
rect 16880 -2000 17000 -1980
rect 12000 -2200 17000 -2000
rect 12000 -2220 12120 -2200
rect 12380 -2220 12620 -2200
rect 12880 -2220 13120 -2200
rect 13380 -2220 13620 -2200
rect 13880 -2220 14120 -2200
rect 14380 -2220 14620 -2200
rect 14880 -2220 15120 -2200
rect 15380 -2220 15620 -2200
rect 15880 -2220 16120 -2200
rect 16380 -2220 16620 -2200
rect 16880 -2220 17000 -2200
rect 12000 -2480 12100 -2220
rect 12400 -2480 12600 -2220
rect 12900 -2480 13100 -2220
rect 13400 -2480 13600 -2220
rect 13900 -2480 14100 -2220
rect 14400 -2480 14600 -2220
rect 14900 -2480 15100 -2220
rect 15400 -2480 15600 -2220
rect 15900 -2480 16100 -2220
rect 16400 -2480 16600 -2220
rect 16900 -2480 17000 -2220
rect 12000 -2500 12120 -2480
rect 12380 -2500 12620 -2480
rect 12880 -2500 13120 -2480
rect 13380 -2500 13620 -2480
rect 13880 -2500 14120 -2480
rect 14380 -2500 14620 -2480
rect 14880 -2500 15120 -2480
rect 15380 -2500 15620 -2480
rect 15880 -2500 16120 -2480
rect 16380 -2500 16620 -2480
rect 16880 -2500 17000 -2480
rect 12000 -2700 17000 -2500
rect 12000 -2720 12120 -2700
rect 12380 -2720 12620 -2700
rect 12880 -2720 13120 -2700
rect 13380 -2720 13620 -2700
rect 13880 -2720 14120 -2700
rect 14380 -2720 14620 -2700
rect 14880 -2720 15120 -2700
rect 15380 -2720 15620 -2700
rect 15880 -2720 16120 -2700
rect 16380 -2720 16620 -2700
rect 16880 -2720 17000 -2700
rect 12000 -2980 12100 -2720
rect 12400 -2980 12600 -2720
rect 12900 -2980 13100 -2720
rect 13400 -2980 13600 -2720
rect 13900 -2980 14100 -2720
rect 14400 -2980 14600 -2720
rect 14900 -2980 15100 -2720
rect 15400 -2980 15600 -2720
rect 15900 -2980 16100 -2720
rect 16400 -2980 16600 -2720
rect 16900 -2980 17000 -2720
rect 12000 -3000 12120 -2980
rect 12380 -3000 12620 -2980
rect 12880 -3000 13120 -2980
rect 13380 -3000 13620 -2980
rect 13880 -3000 14120 -2980
rect 14380 -3000 14620 -2980
rect 14880 -3000 15120 -2980
rect 15380 -3000 15620 -2980
rect 15880 -3000 16120 -2980
rect 16380 -3000 16620 -2980
rect 16880 -3000 17000 -2980
rect -23500 -3200 -14500 -3100
rect -23500 -3220 -23380 -3200
rect -23120 -3220 -22880 -3200
rect -22620 -3220 -22380 -3200
rect -22120 -3220 -21880 -3200
rect -21620 -3220 -21380 -3200
rect -21120 -3220 -20880 -3200
rect -20620 -3220 -20380 -3200
rect -20120 -3220 -19880 -3200
rect -19620 -3220 -19380 -3200
rect -19120 -3220 -18880 -3200
rect -18620 -3220 -18380 -3200
rect -18120 -3220 -17880 -3200
rect -17620 -3220 -17380 -3200
rect -17120 -3220 -16880 -3200
rect -16620 -3220 -16380 -3200
rect -16120 -3220 -15880 -3200
rect -15620 -3220 -15380 -3200
rect -15120 -3220 -14880 -3200
rect -14620 -3220 -14500 -3200
rect -23500 -3480 -23400 -3220
rect -23100 -3480 -22900 -3220
rect -22600 -3480 -22400 -3220
rect -22100 -3480 -21900 -3220
rect -21600 -3480 -21400 -3220
rect -21100 -3480 -20900 -3220
rect -20600 -3480 -20400 -3220
rect -20100 -3480 -19900 -3220
rect -19600 -3480 -19400 -3220
rect -19100 -3480 -18900 -3220
rect -18600 -3480 -18400 -3220
rect -18100 -3480 -17900 -3220
rect -17600 -3480 -17400 -3220
rect -17100 -3480 -16900 -3220
rect -16600 -3480 -16400 -3220
rect -16100 -3480 -15900 -3220
rect -15600 -3480 -15400 -3220
rect -15100 -3480 -14900 -3220
rect -14600 -3480 -14500 -3220
rect -23500 -3500 -23380 -3480
rect -23120 -3500 -22880 -3480
rect -22620 -3500 -22380 -3480
rect -22120 -3500 -21880 -3480
rect -21620 -3500 -21380 -3480
rect -21120 -3500 -20880 -3480
rect -20620 -3500 -20380 -3480
rect -20120 -3500 -19880 -3480
rect -19620 -3500 -19380 -3480
rect -19120 -3500 -18880 -3480
rect -18620 -3500 -18380 -3480
rect -18120 -3500 -17880 -3480
rect -17620 -3500 -17380 -3480
rect -17120 -3500 -16880 -3480
rect -16620 -3500 -16380 -3480
rect -16120 -3500 -15880 -3480
rect -15620 -3500 -15380 -3480
rect -15120 -3500 -14880 -3480
rect -14620 -3500 -14500 -3480
rect -23500 -3600 -14500 -3500
rect 12000 -3200 17000 -3000
rect 12000 -3220 12120 -3200
rect 12380 -3220 12620 -3200
rect 12880 -3220 13120 -3200
rect 13380 -3220 13620 -3200
rect 13880 -3220 14120 -3200
rect 14380 -3220 14620 -3200
rect 14880 -3220 15120 -3200
rect 15380 -3220 15620 -3200
rect 15880 -3220 16120 -3200
rect 16380 -3220 16620 -3200
rect 16880 -3220 17000 -3200
rect 12000 -3480 12100 -3220
rect 12400 -3480 12600 -3220
rect 12900 -3480 13100 -3220
rect 13400 -3480 13600 -3220
rect 13900 -3480 14100 -3220
rect 14400 -3480 14600 -3220
rect 14900 -3480 15100 -3220
rect 15400 -3480 15600 -3220
rect 15900 -3480 16100 -3220
rect 16400 -3480 16600 -3220
rect 16900 -3480 17000 -3220
rect 12000 -3500 12120 -3480
rect 12380 -3500 12620 -3480
rect 12880 -3500 13120 -3480
rect 13380 -3500 13620 -3480
rect 13880 -3500 14120 -3480
rect 14380 -3500 14620 -3480
rect 14880 -3500 15120 -3480
rect 15380 -3500 15620 -3480
rect 15880 -3500 16120 -3480
rect 16380 -3500 16620 -3480
rect 16880 -3500 17000 -3480
rect 12000 -3600 17000 -3500
rect 17500 300 19500 500
rect 17500 280 17620 300
rect 17880 280 18120 300
rect 18380 280 18620 300
rect 18880 280 19120 300
rect 19380 280 19500 300
rect 17500 20 17600 280
rect 17900 20 18100 280
rect 18400 20 18600 280
rect 18900 20 19100 280
rect 19400 20 19500 280
rect 17500 0 17620 20
rect 17880 0 18120 20
rect 18380 0 18620 20
rect 18880 0 19120 20
rect 19380 0 19500 20
rect 17500 -200 19500 0
rect 17500 -220 17620 -200
rect 17880 -220 18120 -200
rect 18380 -220 18620 -200
rect 18880 -220 19120 -200
rect 19380 -220 19500 -200
rect 17500 -480 17600 -220
rect 17900 -480 18100 -220
rect 18400 -480 18600 -220
rect 18900 -480 19100 -220
rect 19400 -480 19500 -220
rect 17500 -500 17620 -480
rect 17880 -500 18120 -480
rect 18380 -500 18620 -480
rect 18880 -500 19120 -480
rect 19380 -500 19500 -480
rect 17500 -700 19500 -500
rect 17500 -720 17620 -700
rect 17880 -720 18120 -700
rect 18380 -720 18620 -700
rect 18880 -720 19120 -700
rect 19380 -720 19500 -700
rect 17500 -980 17600 -720
rect 17900 -980 18100 -720
rect 18400 -980 18600 -720
rect 18900 -980 19100 -720
rect 19400 -980 19500 -720
rect 17500 -1000 17620 -980
rect 17880 -1000 18120 -980
rect 18380 -1000 18620 -980
rect 18880 -1000 19120 -980
rect 19380 -1000 19500 -980
rect 17500 -1200 19500 -1000
rect 17500 -1220 17620 -1200
rect 17880 -1220 18120 -1200
rect 18380 -1220 18620 -1200
rect 18880 -1220 19120 -1200
rect 19380 -1220 19500 -1200
rect 17500 -1480 17600 -1220
rect 17900 -1480 18100 -1220
rect 18400 -1480 18600 -1220
rect 18900 -1480 19100 -1220
rect 19400 -1480 19500 -1220
rect 17500 -1500 17620 -1480
rect 17880 -1500 18120 -1480
rect 18380 -1500 18620 -1480
rect 18880 -1500 19120 -1480
rect 19380 -1500 19500 -1480
rect 17500 -1700 19500 -1500
rect 17500 -1720 17620 -1700
rect 17880 -1720 18120 -1700
rect 18380 -1720 18620 -1700
rect 18880 -1720 19120 -1700
rect 19380 -1720 19500 -1700
rect 17500 -1980 17600 -1720
rect 17900 -1980 18100 -1720
rect 18400 -1980 18600 -1720
rect 18900 -1980 19100 -1720
rect 19400 -1980 19500 -1720
rect 17500 -2000 17620 -1980
rect 17880 -2000 18120 -1980
rect 18380 -2000 18620 -1980
rect 18880 -2000 19120 -1980
rect 19380 -2000 19500 -1980
rect 17500 -2200 19500 -2000
rect 17500 -2220 17620 -2200
rect 17880 -2220 18120 -2200
rect 18380 -2220 18620 -2200
rect 18880 -2220 19120 -2200
rect 19380 -2220 19500 -2200
rect 17500 -2480 17600 -2220
rect 17900 -2480 18100 -2220
rect 18400 -2480 18600 -2220
rect 18900 -2480 19100 -2220
rect 19400 -2480 19500 -2220
rect 17500 -2500 17620 -2480
rect 17880 -2500 18120 -2480
rect 18380 -2500 18620 -2480
rect 18880 -2500 19120 -2480
rect 19380 -2500 19500 -2480
rect 17500 -2700 19500 -2500
rect 17500 -2720 17620 -2700
rect 17880 -2720 18120 -2700
rect 18380 -2720 18620 -2700
rect 18880 -2720 19120 -2700
rect 19380 -2720 19500 -2700
rect 17500 -2980 17600 -2720
rect 17900 -2980 18100 -2720
rect 18400 -2980 18600 -2720
rect 18900 -2980 19100 -2720
rect 19400 -2980 19500 -2720
rect 17500 -3000 17620 -2980
rect 17880 -3000 18120 -2980
rect 18380 -3000 18620 -2980
rect 18880 -3000 19120 -2980
rect 19380 -3000 19500 -2980
rect 17500 -3200 19500 -3000
rect 17500 -3220 17620 -3200
rect 17880 -3220 18120 -3200
rect 18380 -3220 18620 -3200
rect 18880 -3220 19120 -3200
rect 19380 -3220 19500 -3200
rect 17500 -3480 17600 -3220
rect 17900 -3480 18100 -3220
rect 18400 -3480 18600 -3220
rect 18900 -3480 19100 -3220
rect 19400 -3480 19500 -3220
rect 17500 -3500 17620 -3480
rect 17880 -3500 18120 -3480
rect 18380 -3500 18620 -3480
rect 18880 -3500 19120 -3480
rect 19380 -3500 19500 -3480
rect 17500 -3600 19500 -3500
rect 32500 1300 33500 1400
rect 32500 1280 32620 1300
rect 32880 1280 33120 1300
rect 33380 1280 33500 1300
rect 32500 1020 32600 1280
rect 32900 1020 33100 1280
rect 33400 1020 33500 1280
rect 32500 1000 32620 1020
rect 32880 1000 33120 1020
rect 33380 1000 33500 1020
rect 32500 800 33500 1000
rect 32500 780 32620 800
rect 32880 780 33120 800
rect 33380 780 33500 800
rect 32500 520 32600 780
rect 32900 520 33100 780
rect 33400 520 33500 780
rect 32500 500 32620 520
rect 32880 500 33120 520
rect 33380 500 33500 520
rect 32500 300 33500 500
rect 32500 280 32620 300
rect 32880 280 33120 300
rect 33380 280 33500 300
rect 32500 20 32600 280
rect 32900 20 33100 280
rect 33400 20 33500 280
rect 32500 0 32620 20
rect 32880 0 33120 20
rect 33380 0 33500 20
rect 32500 -200 33500 0
rect 32500 -220 32620 -200
rect 32880 -220 33120 -200
rect 33380 -220 33500 -200
rect 32500 -480 32600 -220
rect 32900 -480 33100 -220
rect 33400 -480 33500 -220
rect 32500 -500 32620 -480
rect 32880 -500 33120 -480
rect 33380 -500 33500 -480
rect 32500 -700 33500 -500
rect 32500 -720 32620 -700
rect 32880 -720 33120 -700
rect 33380 -720 33500 -700
rect 32500 -980 32600 -720
rect 32900 -980 33100 -720
rect 33400 -980 33500 -720
rect 32500 -1000 32620 -980
rect 32880 -1000 33120 -980
rect 33380 -1000 33500 -980
rect 32500 -1200 33500 -1000
rect 32500 -1220 32620 -1200
rect 32880 -1220 33120 -1200
rect 33380 -1220 33500 -1200
rect 32500 -1480 32600 -1220
rect 32900 -1480 33100 -1220
rect 33400 -1480 33500 -1220
rect 32500 -1500 32620 -1480
rect 32880 -1500 33120 -1480
rect 33380 -1500 33500 -1480
rect 32500 -1700 33500 -1500
rect 32500 -1720 32620 -1700
rect 32880 -1720 33120 -1700
rect 33380 -1720 33500 -1700
rect 32500 -1980 32600 -1720
rect 32900 -1980 33100 -1720
rect 33400 -1980 33500 -1720
rect 32500 -2000 32620 -1980
rect 32880 -2000 33120 -1980
rect 33380 -2000 33500 -1980
rect 32500 -2200 33500 -2000
rect 32500 -2220 32620 -2200
rect 32880 -2220 33120 -2200
rect 33380 -2220 33500 -2200
rect 32500 -2480 32600 -2220
rect 32900 -2480 33100 -2220
rect 33400 -2480 33500 -2220
rect 32500 -2500 32620 -2480
rect 32880 -2500 33120 -2480
rect 33380 -2500 33500 -2480
rect 32500 -2700 33500 -2500
rect 32500 -2720 32620 -2700
rect 32880 -2720 33120 -2700
rect 33380 -2720 33500 -2700
rect 32500 -2980 32600 -2720
rect 32900 -2980 33100 -2720
rect 33400 -2980 33500 -2720
rect 32500 -3000 32620 -2980
rect 32880 -3000 33120 -2980
rect 33380 -3000 33500 -2980
rect 32500 -3200 33500 -3000
rect 32500 -3220 32620 -3200
rect 32880 -3220 33120 -3200
rect 33380 -3220 33500 -3200
rect 32500 -3480 32600 -3220
rect 32900 -3480 33100 -3220
rect 33400 -3480 33500 -3220
rect 32500 -3500 32620 -3480
rect 32880 -3500 33120 -3480
rect 33380 -3500 33500 -3480
rect 32500 -3600 33500 -3500
rect -23500 -3700 -15000 -3600
rect -23500 -3720 -23380 -3700
rect -23120 -3720 -22880 -3700
rect -22620 -3720 -22380 -3700
rect -22120 -3720 -21880 -3700
rect -21620 -3720 -21380 -3700
rect -21120 -3720 -20880 -3700
rect -20620 -3720 -20380 -3700
rect -20120 -3720 -19880 -3700
rect -19620 -3720 -19380 -3700
rect -19120 -3720 -18880 -3700
rect -18620 -3720 -18380 -3700
rect -18120 -3720 -17880 -3700
rect -17620 -3720 -17380 -3700
rect -17120 -3720 -16880 -3700
rect -16620 -3720 -16380 -3700
rect -16120 -3720 -15880 -3700
rect -15620 -3720 -15380 -3700
rect -15120 -3720 -15000 -3700
rect -23500 -3980 -23400 -3720
rect -23100 -3980 -22900 -3720
rect -22600 -3980 -22400 -3720
rect -22100 -3980 -21900 -3720
rect -21600 -3980 -21400 -3720
rect -21100 -3980 -20900 -3720
rect -20600 -3980 -20400 -3720
rect -20100 -3980 -19900 -3720
rect -19600 -3980 -19400 -3720
rect -19100 -3980 -18900 -3720
rect -18600 -3980 -18400 -3720
rect -18100 -3980 -17900 -3720
rect -17600 -3980 -17400 -3720
rect -17100 -3980 -16900 -3720
rect -16600 -3980 -16400 -3720
rect -16100 -3980 -15900 -3720
rect -15600 -3980 -15400 -3720
rect -15100 -3980 -15000 -3720
rect -23500 -4000 -23380 -3980
rect -23120 -4000 -22880 -3980
rect -22620 -4000 -22380 -3980
rect -22120 -4000 -21880 -3980
rect -21620 -4000 -21380 -3980
rect -21120 -4000 -20880 -3980
rect -20620 -4000 -20380 -3980
rect -20120 -4000 -19880 -3980
rect -19620 -4000 -19380 -3980
rect -19120 -4000 -18880 -3980
rect -18620 -4000 -18380 -3980
rect -18120 -4000 -17880 -3980
rect -17620 -4000 -17380 -3980
rect -17120 -4000 -16880 -3980
rect -16620 -4000 -16380 -3980
rect -16120 -4000 -15880 -3980
rect -15620 -4000 -15380 -3980
rect -15120 -4000 -15000 -3980
rect -23500 -4200 -15000 -4000
rect -23500 -4220 -23380 -4200
rect -23120 -4220 -22880 -4200
rect -22620 -4220 -22380 -4200
rect -22120 -4220 -21880 -4200
rect -21620 -4220 -21380 -4200
rect -21120 -4220 -20880 -4200
rect -20620 -4220 -20380 -4200
rect -20120 -4220 -19880 -4200
rect -19620 -4220 -19380 -4200
rect -19120 -4220 -18880 -4200
rect -18620 -4220 -18380 -4200
rect -18120 -4220 -17880 -4200
rect -17620 -4220 -17380 -4200
rect -17120 -4220 -16880 -4200
rect -16620 -4220 -16380 -4200
rect -16120 -4220 -15880 -4200
rect -15620 -4220 -15380 -4200
rect -15120 -4220 -15000 -4200
rect -23500 -4480 -23400 -4220
rect -23100 -4480 -22900 -4220
rect -22600 -4480 -22400 -4220
rect -22100 -4480 -21900 -4220
rect -21600 -4480 -21400 -4220
rect -21100 -4480 -20900 -4220
rect -20600 -4480 -20400 -4220
rect -20100 -4480 -19900 -4220
rect -19600 -4480 -19400 -4220
rect -19100 -4480 -18900 -4220
rect -18600 -4480 -18400 -4220
rect -18100 -4480 -17900 -4220
rect -17600 -4480 -17400 -4220
rect -17100 -4480 -16900 -4220
rect -16600 -4480 -16400 -4220
rect -16100 -4480 -15900 -4220
rect -15600 -4480 -15400 -4220
rect -15100 -4480 -15000 -4220
rect -23500 -4500 -23380 -4480
rect -23120 -4500 -22880 -4480
rect -22620 -4500 -22380 -4480
rect -22120 -4500 -21880 -4480
rect -21620 -4500 -21380 -4480
rect -21120 -4500 -20880 -4480
rect -20620 -4500 -20380 -4480
rect -20120 -4500 -19880 -4480
rect -19620 -4500 -19380 -4480
rect -19120 -4500 -18880 -4480
rect -18620 -4500 -18380 -4480
rect -18120 -4500 -17880 -4480
rect -17620 -4500 -17380 -4480
rect -17120 -4500 -16880 -4480
rect -16620 -4500 -16380 -4480
rect -16120 -4500 -15880 -4480
rect -15620 -4500 -15380 -4480
rect -15120 -4500 -15000 -4480
rect -23500 -4700 -15000 -4500
rect -23500 -4720 -23380 -4700
rect -23120 -4720 -22880 -4700
rect -22620 -4720 -22380 -4700
rect -22120 -4720 -21880 -4700
rect -21620 -4720 -21380 -4700
rect -21120 -4720 -20880 -4700
rect -20620 -4720 -20380 -4700
rect -20120 -4720 -19880 -4700
rect -19620 -4720 -19380 -4700
rect -19120 -4720 -18880 -4700
rect -18620 -4720 -18380 -4700
rect -18120 -4720 -17880 -4700
rect -17620 -4720 -17380 -4700
rect -17120 -4720 -16880 -4700
rect -16620 -4720 -16380 -4700
rect -16120 -4720 -15880 -4700
rect -15620 -4720 -15380 -4700
rect -15120 -4720 -15000 -4700
rect -23500 -4980 -23400 -4720
rect -23100 -4980 -22900 -4720
rect -22600 -4980 -22400 -4720
rect -22100 -4980 -21900 -4720
rect -21600 -4980 -21400 -4720
rect -21100 -4980 -20900 -4720
rect -20600 -4980 -20400 -4720
rect -20100 -4980 -19900 -4720
rect -19600 -4980 -19400 -4720
rect -19100 -4980 -18900 -4720
rect -18600 -4980 -18400 -4720
rect -18100 -4980 -17900 -4720
rect -17600 -4980 -17400 -4720
rect -17100 -4980 -16900 -4720
rect -16600 -4980 -16400 -4720
rect -16100 -4980 -15900 -4720
rect -15600 -4980 -15400 -4720
rect -15100 -4980 -15000 -4720
rect -23500 -5000 -23380 -4980
rect -23120 -5000 -22880 -4980
rect -22620 -5000 -22380 -4980
rect -22120 -5000 -21880 -4980
rect -21620 -5000 -21380 -4980
rect -21120 -5000 -20880 -4980
rect -20620 -5000 -20380 -4980
rect -20120 -5000 -19880 -4980
rect -19620 -5000 -19380 -4980
rect -19120 -5000 -18880 -4980
rect -18620 -5000 -18380 -4980
rect -18120 -5000 -17880 -4980
rect -17620 -5000 -17380 -4980
rect -17120 -5000 -16880 -4980
rect -16620 -5000 -16380 -4980
rect -16120 -5000 -15880 -4980
rect -15620 -5000 -15380 -4980
rect -15120 -5000 -15000 -4980
rect -23500 -5200 -15000 -5000
rect -23500 -5220 -23380 -5200
rect -23120 -5220 -22880 -5200
rect -22620 -5220 -22380 -5200
rect -22120 -5220 -21880 -5200
rect -21620 -5220 -21380 -5200
rect -21120 -5220 -20880 -5200
rect -20620 -5220 -20380 -5200
rect -20120 -5220 -19880 -5200
rect -19620 -5220 -19380 -5200
rect -19120 -5220 -18880 -5200
rect -18620 -5220 -18380 -5200
rect -18120 -5220 -17880 -5200
rect -17620 -5220 -17380 -5200
rect -17120 -5220 -16880 -5200
rect -16620 -5220 -16380 -5200
rect -16120 -5220 -15880 -5200
rect -15620 -5220 -15380 -5200
rect -15120 -5220 -15000 -5200
rect -23500 -5480 -23400 -5220
rect -23100 -5480 -22900 -5220
rect -22600 -5480 -22400 -5220
rect -22100 -5480 -21900 -5220
rect -21600 -5480 -21400 -5220
rect -21100 -5480 -20900 -5220
rect -20600 -5480 -20400 -5220
rect -20100 -5480 -19900 -5220
rect -19600 -5480 -19400 -5220
rect -19100 -5480 -18900 -5220
rect -18600 -5480 -18400 -5220
rect -18100 -5480 -17900 -5220
rect -17600 -5480 -17400 -5220
rect -17100 -5480 -16900 -5220
rect -16600 -5480 -16400 -5220
rect -16100 -5480 -15900 -5220
rect -15600 -5480 -15400 -5220
rect -15100 -5480 -15000 -5220
rect -23500 -5500 -23380 -5480
rect -23120 -5500 -22880 -5480
rect -22620 -5500 -22380 -5480
rect -22120 -5500 -21880 -5480
rect -21620 -5500 -21380 -5480
rect -21120 -5500 -20880 -5480
rect -20620 -5500 -20380 -5480
rect -20120 -5500 -19880 -5480
rect -19620 -5500 -19380 -5480
rect -19120 -5500 -18880 -5480
rect -18620 -5500 -18380 -5480
rect -18120 -5500 -17880 -5480
rect -17620 -5500 -17380 -5480
rect -17120 -5500 -16880 -5480
rect -16620 -5500 -16380 -5480
rect -16120 -5500 -15880 -5480
rect -15620 -5500 -15380 -5480
rect -15120 -5500 -15000 -5480
rect -23500 -5700 -15000 -5500
rect -23500 -5720 -23380 -5700
rect -23120 -5720 -22880 -5700
rect -22620 -5720 -22380 -5700
rect -22120 -5720 -21880 -5700
rect -21620 -5720 -21380 -5700
rect -21120 -5720 -20880 -5700
rect -20620 -5720 -20380 -5700
rect -20120 -5720 -19880 -5700
rect -19620 -5720 -19380 -5700
rect -19120 -5720 -18880 -5700
rect -18620 -5720 -18380 -5700
rect -18120 -5720 -17880 -5700
rect -17620 -5720 -17380 -5700
rect -17120 -5720 -16880 -5700
rect -16620 -5720 -16380 -5700
rect -16120 -5720 -15880 -5700
rect -15620 -5720 -15380 -5700
rect -15120 -5720 -15000 -5700
rect -23500 -5980 -23400 -5720
rect -23100 -5980 -22900 -5720
rect -22600 -5980 -22400 -5720
rect -22100 -5980 -21900 -5720
rect -21600 -5980 -21400 -5720
rect -21100 -5980 -20900 -5720
rect -20600 -5980 -20400 -5720
rect -20100 -5980 -19900 -5720
rect -19600 -5980 -19400 -5720
rect -19100 -5980 -18900 -5720
rect -18600 -5980 -18400 -5720
rect -18100 -5980 -17900 -5720
rect -17600 -5980 -17400 -5720
rect -17100 -5980 -16900 -5720
rect -16600 -5980 -16400 -5720
rect -16100 -5980 -15900 -5720
rect -15600 -5980 -15400 -5720
rect -15100 -5980 -15000 -5720
rect -23500 -6000 -23380 -5980
rect -23120 -6000 -22880 -5980
rect -22620 -6000 -22380 -5980
rect -22120 -6000 -21880 -5980
rect -21620 -6000 -21380 -5980
rect -21120 -6000 -20880 -5980
rect -20620 -6000 -20380 -5980
rect -20120 -6000 -19880 -5980
rect -19620 -6000 -19380 -5980
rect -19120 -6000 -18880 -5980
rect -18620 -6000 -18380 -5980
rect -18120 -6000 -17880 -5980
rect -17620 -6000 -17380 -5980
rect -17120 -6000 -16880 -5980
rect -16620 -6000 -16380 -5980
rect -16120 -6000 -15880 -5980
rect -15620 -6000 -15380 -5980
rect -15120 -6000 -15000 -5980
rect -23500 -6200 -15000 -6000
rect -23500 -6220 -23380 -6200
rect -23120 -6220 -22880 -6200
rect -22620 -6220 -22380 -6200
rect -22120 -6220 -21880 -6200
rect -21620 -6220 -21380 -6200
rect -21120 -6220 -20880 -6200
rect -20620 -6220 -20380 -6200
rect -20120 -6220 -19880 -6200
rect -19620 -6220 -19380 -6200
rect -19120 -6220 -18880 -6200
rect -18620 -6220 -18380 -6200
rect -18120 -6220 -17880 -6200
rect -17620 -6220 -17380 -6200
rect -17120 -6220 -16880 -6200
rect -16620 -6220 -16380 -6200
rect -16120 -6220 -15880 -6200
rect -15620 -6220 -15380 -6200
rect -15120 -6220 -15000 -6200
rect -23500 -6480 -23400 -6220
rect -23100 -6480 -22900 -6220
rect -22600 -6480 -22400 -6220
rect -22100 -6480 -21900 -6220
rect -21600 -6480 -21400 -6220
rect -21100 -6480 -20900 -6220
rect -20600 -6480 -20400 -6220
rect -20100 -6480 -19900 -6220
rect -19600 -6480 -19400 -6220
rect -19100 -6480 -18900 -6220
rect -18600 -6480 -18400 -6220
rect -18100 -6480 -17900 -6220
rect -17600 -6480 -17400 -6220
rect -17100 -6480 -16900 -6220
rect -16600 -6480 -16400 -6220
rect -16100 -6480 -15900 -6220
rect -15600 -6480 -15400 -6220
rect -15100 -6480 -15000 -6220
rect -23500 -6500 -23380 -6480
rect -23120 -6500 -22880 -6480
rect -22620 -6500 -22380 -6480
rect -22120 -6500 -21880 -6480
rect -21620 -6500 -21380 -6480
rect -21120 -6500 -20880 -6480
rect -20620 -6500 -20380 -6480
rect -20120 -6500 -19880 -6480
rect -19620 -6500 -19380 -6480
rect -19120 -6500 -18880 -6480
rect -18620 -6500 -18380 -6480
rect -18120 -6500 -17880 -6480
rect -17620 -6500 -17380 -6480
rect -17120 -6500 -16880 -6480
rect -16620 -6500 -16380 -6480
rect -16120 -6500 -15880 -6480
rect -15620 -6500 -15380 -6480
rect -15120 -6500 -15000 -6480
rect -23500 -6700 -15000 -6500
rect -23500 -6720 -23380 -6700
rect -23120 -6720 -22880 -6700
rect -22620 -6720 -22380 -6700
rect -22120 -6720 -21880 -6700
rect -21620 -6720 -21380 -6700
rect -21120 -6720 -20880 -6700
rect -20620 -6720 -20380 -6700
rect -20120 -6720 -19880 -6700
rect -19620 -6720 -19380 -6700
rect -19120 -6720 -18880 -6700
rect -18620 -6720 -18380 -6700
rect -18120 -6720 -17880 -6700
rect -17620 -6720 -17380 -6700
rect -17120 -6720 -16880 -6700
rect -16620 -6720 -16380 -6700
rect -16120 -6720 -15880 -6700
rect -15620 -6720 -15380 -6700
rect -15120 -6720 -15000 -6700
rect -23500 -6980 -23400 -6720
rect -23100 -6980 -22900 -6720
rect -22600 -6980 -22400 -6720
rect -22100 -6980 -21900 -6720
rect -21600 -6980 -21400 -6720
rect -21100 -6980 -20900 -6720
rect -20600 -6980 -20400 -6720
rect -20100 -6980 -19900 -6720
rect -19600 -6980 -19400 -6720
rect -19100 -6980 -18900 -6720
rect -18600 -6980 -18400 -6720
rect -18100 -6980 -17900 -6720
rect -17600 -6980 -17400 -6720
rect -17100 -6980 -16900 -6720
rect -16600 -6980 -16400 -6720
rect -16100 -6980 -15900 -6720
rect -15600 -6980 -15400 -6720
rect -15100 -6980 -15000 -6720
rect -23500 -7000 -23380 -6980
rect -23120 -7000 -22880 -6980
rect -22620 -7000 -22380 -6980
rect -22120 -7000 -21880 -6980
rect -21620 -7000 -21380 -6980
rect -21120 -7000 -20880 -6980
rect -20620 -7000 -20380 -6980
rect -20120 -7000 -19880 -6980
rect -19620 -7000 -19380 -6980
rect -19120 -7000 -18880 -6980
rect -18620 -7000 -18380 -6980
rect -18120 -7000 -17880 -6980
rect -17620 -7000 -17380 -6980
rect -17120 -7000 -16880 -6980
rect -16620 -7000 -16380 -6980
rect -16120 -7000 -15880 -6980
rect -15620 -7000 -15380 -6980
rect -15120 -7000 -15000 -6980
rect -23500 -7200 -15000 -7000
rect -23500 -7220 -23380 -7200
rect -23120 -7220 -22880 -7200
rect -22620 -7220 -22380 -7200
rect -22120 -7220 -21880 -7200
rect -21620 -7220 -21380 -7200
rect -21120 -7220 -20880 -7200
rect -20620 -7220 -20380 -7200
rect -20120 -7220 -19880 -7200
rect -19620 -7220 -19380 -7200
rect -19120 -7220 -18880 -7200
rect -18620 -7220 -18380 -7200
rect -18120 -7220 -17880 -7200
rect -17620 -7220 -17380 -7200
rect -17120 -7220 -16880 -7200
rect -16620 -7220 -16380 -7200
rect -16120 -7220 -15880 -7200
rect -15620 -7220 -15380 -7200
rect -15120 -7220 -15000 -7200
rect -23500 -7480 -23400 -7220
rect -23100 -7480 -22900 -7220
rect -22600 -7480 -22400 -7220
rect -22100 -7480 -21900 -7220
rect -21600 -7480 -21400 -7220
rect -21100 -7480 -20900 -7220
rect -20600 -7480 -20400 -7220
rect -20100 -7480 -19900 -7220
rect -19600 -7480 -19400 -7220
rect -19100 -7480 -18900 -7220
rect -18600 -7480 -18400 -7220
rect -18100 -7480 -17900 -7220
rect -17600 -7480 -17400 -7220
rect -17100 -7480 -16900 -7220
rect -16600 -7480 -16400 -7220
rect -16100 -7480 -15900 -7220
rect -15600 -7480 -15400 -7220
rect -15100 -7480 -15000 -7220
rect -23500 -7500 -23380 -7480
rect -23120 -7500 -22880 -7480
rect -22620 -7500 -22380 -7480
rect -22120 -7500 -21880 -7480
rect -21620 -7500 -21380 -7480
rect -21120 -7500 -20880 -7480
rect -20620 -7500 -20380 -7480
rect -20120 -7500 -19880 -7480
rect -19620 -7500 -19380 -7480
rect -19120 -7500 -18880 -7480
rect -18620 -7500 -18380 -7480
rect -18120 -7500 -17880 -7480
rect -17620 -7500 -17380 -7480
rect -17120 -7500 -16880 -7480
rect -16620 -7500 -16380 -7480
rect -16120 -7500 -15880 -7480
rect -15620 -7500 -15380 -7480
rect -15120 -7500 -15000 -7480
rect -28000 -8100 -27500 -7600
rect -23500 -7700 -15000 -7500
rect -23500 -7720 -23380 -7700
rect -23120 -7720 -22880 -7700
rect -22620 -7720 -22380 -7700
rect -22120 -7720 -21880 -7700
rect -21620 -7720 -21380 -7700
rect -21120 -7720 -20880 -7700
rect -20620 -7720 -20380 -7700
rect -20120 -7720 -19880 -7700
rect -19620 -7720 -19380 -7700
rect -19120 -7720 -18880 -7700
rect -18620 -7720 -18380 -7700
rect -18120 -7720 -17880 -7700
rect -17620 -7720 -17380 -7700
rect -17120 -7720 -16880 -7700
rect -16620 -7720 -16380 -7700
rect -16120 -7720 -15880 -7700
rect -15620 -7720 -15380 -7700
rect -15120 -7720 -15000 -7700
rect -23500 -7980 -23400 -7720
rect -23100 -7980 -22900 -7720
rect -22600 -7980 -22400 -7720
rect -22100 -7980 -21900 -7720
rect -21600 -7980 -21400 -7720
rect -21100 -7980 -20900 -7720
rect -20600 -7980 -20400 -7720
rect -20100 -7980 -19900 -7720
rect -19600 -7980 -19400 -7720
rect -19100 -7980 -18900 -7720
rect -18600 -7980 -18400 -7720
rect -18100 -7980 -17900 -7720
rect -17600 -7980 -17400 -7720
rect -17100 -7980 -16900 -7720
rect -16600 -7980 -16400 -7720
rect -16100 -7980 -15900 -7720
rect -15600 -7980 -15400 -7720
rect -15100 -7980 -15000 -7720
rect -23500 -8000 -23380 -7980
rect -23120 -8000 -22880 -7980
rect -22620 -8000 -22380 -7980
rect -22120 -8000 -21880 -7980
rect -21620 -8000 -21380 -7980
rect -21120 -8000 -20880 -7980
rect -20620 -8000 -20380 -7980
rect -20120 -8000 -19880 -7980
rect -19620 -8000 -19380 -7980
rect -19120 -8000 -18880 -7980
rect -18620 -8000 -18380 -7980
rect -18120 -8000 -17880 -7980
rect -17620 -8000 -17380 -7980
rect -17120 -8000 -16880 -7980
rect -16620 -8000 -16380 -7980
rect -16120 -8000 -15880 -7980
rect -15620 -8000 -15380 -7980
rect -15120 -8000 -15000 -7980
rect -23500 -8100 -15000 -8000
rect -27500 -8200 -15000 -8100
rect -27500 -8220 -27380 -8200
rect -27120 -8220 -26880 -8200
rect -26620 -8220 -26380 -8200
rect -26120 -8220 -25880 -8200
rect -25620 -8220 -25380 -8200
rect -25120 -8220 -24880 -8200
rect -24620 -8220 -24380 -8200
rect -24120 -8220 -23880 -8200
rect -23620 -8220 -23380 -8200
rect -23120 -8220 -22880 -8200
rect -22620 -8220 -22380 -8200
rect -22120 -8220 -21880 -8200
rect -21620 -8220 -21380 -8200
rect -21120 -8220 -20880 -8200
rect -20620 -8220 -20380 -8200
rect -20120 -8220 -19880 -8200
rect -19620 -8220 -19380 -8200
rect -19120 -8220 -18880 -8200
rect -18620 -8220 -18380 -8200
rect -18120 -8220 -17880 -8200
rect -17620 -8220 -17380 -8200
rect -17120 -8220 -16880 -8200
rect -16620 -8220 -16380 -8200
rect -16120 -8220 -15880 -8200
rect -15620 -8220 -15380 -8200
rect -15120 -8220 -15000 -8200
rect -27500 -8480 -27400 -8220
rect -27100 -8480 -26900 -8220
rect -26600 -8480 -26400 -8220
rect -26100 -8480 -25900 -8220
rect -25600 -8480 -25400 -8220
rect -25100 -8480 -24900 -8220
rect -24600 -8480 -24400 -8220
rect -24100 -8480 -23900 -8220
rect -23600 -8480 -23400 -8220
rect -23100 -8480 -22900 -8220
rect -22600 -8480 -22400 -8220
rect -22100 -8480 -21900 -8220
rect -21600 -8480 -21400 -8220
rect -21100 -8480 -20900 -8220
rect -20600 -8480 -20400 -8220
rect -20100 -8480 -19900 -8220
rect -19600 -8480 -19400 -8220
rect -19100 -8480 -18900 -8220
rect -18600 -8480 -18400 -8220
rect -18100 -8480 -17900 -8220
rect -17600 -8480 -17400 -8220
rect -17100 -8480 -16900 -8220
rect -16600 -8480 -16400 -8220
rect -16100 -8480 -15900 -8220
rect -15600 -8480 -15400 -8220
rect -15100 -8480 -15000 -8220
rect -27500 -8500 -27380 -8480
rect -27120 -8500 -26880 -8480
rect -26620 -8500 -26380 -8480
rect -26120 -8500 -25880 -8480
rect -25620 -8500 -25380 -8480
rect -25120 -8500 -24880 -8480
rect -24620 -8500 -24380 -8480
rect -24120 -8500 -23880 -8480
rect -23620 -8500 -23380 -8480
rect -23120 -8500 -22880 -8480
rect -22620 -8500 -22380 -8480
rect -22120 -8500 -21880 -8480
rect -21620 -8500 -21380 -8480
rect -21120 -8500 -20880 -8480
rect -20620 -8500 -20380 -8480
rect -20120 -8500 -19880 -8480
rect -19620 -8500 -19380 -8480
rect -19120 -8500 -18880 -8480
rect -18620 -8500 -18380 -8480
rect -18120 -8500 -17880 -8480
rect -17620 -8500 -17380 -8480
rect -17120 -8500 -16880 -8480
rect -16620 -8500 -16380 -8480
rect -16120 -8500 -15880 -8480
rect -15620 -8500 -15380 -8480
rect -15120 -8500 -15000 -8480
rect -27500 -8700 -15000 -8500
rect -27500 -8720 -27380 -8700
rect -27120 -8720 -26880 -8700
rect -26620 -8720 -26380 -8700
rect -26120 -8720 -25880 -8700
rect -25620 -8720 -25380 -8700
rect -25120 -8720 -24880 -8700
rect -24620 -8720 -24380 -8700
rect -24120 -8720 -23880 -8700
rect -23620 -8720 -23380 -8700
rect -23120 -8720 -22880 -8700
rect -22620 -8720 -22380 -8700
rect -22120 -8720 -21880 -8700
rect -21620 -8720 -21380 -8700
rect -21120 -8720 -20880 -8700
rect -20620 -8720 -20380 -8700
rect -20120 -8720 -19880 -8700
rect -19620 -8720 -19380 -8700
rect -19120 -8720 -18880 -8700
rect -18620 -8720 -18380 -8700
rect -18120 -8720 -17880 -8700
rect -17620 -8720 -17380 -8700
rect -17120 -8720 -16880 -8700
rect -16620 -8720 -16380 -8700
rect -16120 -8720 -15880 -8700
rect -15620 -8720 -15380 -8700
rect -15120 -8720 -15000 -8700
rect -27500 -8980 -27400 -8720
rect -27100 -8980 -26900 -8720
rect -26600 -8980 -26400 -8720
rect -26100 -8980 -25900 -8720
rect -25600 -8980 -25400 -8720
rect -25100 -8980 -24900 -8720
rect -24600 -8980 -24400 -8720
rect -24100 -8980 -23900 -8720
rect -23600 -8980 -23400 -8720
rect -23100 -8980 -22900 -8720
rect -22600 -8980 -22400 -8720
rect -22100 -8980 -21900 -8720
rect -21600 -8980 -21400 -8720
rect -21100 -8980 -20900 -8720
rect -20600 -8980 -20400 -8720
rect -20100 -8980 -19900 -8720
rect -19600 -8980 -19400 -8720
rect -19100 -8980 -18900 -8720
rect -18600 -8980 -18400 -8720
rect -18100 -8980 -17900 -8720
rect -17600 -8980 -17400 -8720
rect -17100 -8980 -16900 -8720
rect -16600 -8980 -16400 -8720
rect -16100 -8980 -15900 -8720
rect -15600 -8980 -15400 -8720
rect -15100 -8980 -15000 -8720
rect -27500 -9000 -27380 -8980
rect -27120 -9000 -26880 -8980
rect -26620 -9000 -26380 -8980
rect -26120 -9000 -25880 -8980
rect -25620 -9000 -25380 -8980
rect -25120 -9000 -24880 -8980
rect -24620 -9000 -24380 -8980
rect -24120 -9000 -23880 -8980
rect -23620 -9000 -23380 -8980
rect -23120 -9000 -22880 -8980
rect -22620 -9000 -22380 -8980
rect -22120 -9000 -21880 -8980
rect -21620 -9000 -21380 -8980
rect -21120 -9000 -20880 -8980
rect -20620 -9000 -20380 -8980
rect -20120 -9000 -19880 -8980
rect -19620 -9000 -19380 -8980
rect -19120 -9000 -18880 -8980
rect -18620 -9000 -18380 -8980
rect -18120 -9000 -17880 -8980
rect -17620 -9000 -17380 -8980
rect -17120 -9000 -16880 -8980
rect -16620 -9000 -16380 -8980
rect -16120 -9000 -15880 -8980
rect -15620 -9000 -15380 -8980
rect -15120 -9000 -15000 -8980
rect -27500 -9200 -15000 -9000
rect -27500 -9220 -27380 -9200
rect -27120 -9220 -26880 -9200
rect -26620 -9220 -26380 -9200
rect -26120 -9220 -25880 -9200
rect -25620 -9220 -25380 -9200
rect -25120 -9220 -24880 -9200
rect -24620 -9220 -24380 -9200
rect -24120 -9220 -23880 -9200
rect -23620 -9220 -23380 -9200
rect -23120 -9220 -22880 -9200
rect -22620 -9220 -22380 -9200
rect -22120 -9220 -21880 -9200
rect -21620 -9220 -21380 -9200
rect -21120 -9220 -20880 -9200
rect -20620 -9220 -20380 -9200
rect -20120 -9220 -19880 -9200
rect -19620 -9220 -19380 -9200
rect -19120 -9220 -18880 -9200
rect -18620 -9220 -18380 -9200
rect -18120 -9220 -17880 -9200
rect -17620 -9220 -17380 -9200
rect -17120 -9220 -16880 -9200
rect -16620 -9220 -16380 -9200
rect -16120 -9220 -15880 -9200
rect -15620 -9220 -15380 -9200
rect -15120 -9220 -15000 -9200
rect -27500 -9480 -27400 -9220
rect -27100 -9480 -26900 -9220
rect -26600 -9480 -26400 -9220
rect -26100 -9480 -25900 -9220
rect -25600 -9480 -25400 -9220
rect -25100 -9480 -24900 -9220
rect -24600 -9480 -24400 -9220
rect -24100 -9480 -23900 -9220
rect -23600 -9480 -23400 -9220
rect -23100 -9480 -22900 -9220
rect -22600 -9480 -22400 -9220
rect -22100 -9480 -21900 -9220
rect -21600 -9480 -21400 -9220
rect -21100 -9480 -20900 -9220
rect -20600 -9480 -20400 -9220
rect -20100 -9480 -19900 -9220
rect -19600 -9480 -19400 -9220
rect -19100 -9480 -18900 -9220
rect -18600 -9480 -18400 -9220
rect -18100 -9480 -17900 -9220
rect -17600 -9480 -17400 -9220
rect -17100 -9480 -16900 -9220
rect -16600 -9480 -16400 -9220
rect -16100 -9480 -15900 -9220
rect -15600 -9480 -15400 -9220
rect -15100 -9480 -15000 -9220
rect -27500 -9500 -27380 -9480
rect -27120 -9500 -26880 -9480
rect -26620 -9500 -26380 -9480
rect -26120 -9500 -25880 -9480
rect -25620 -9500 -25380 -9480
rect -25120 -9500 -24880 -9480
rect -24620 -9500 -24380 -9480
rect -24120 -9500 -23880 -9480
rect -23620 -9500 -23380 -9480
rect -23120 -9500 -22880 -9480
rect -22620 -9500 -22380 -9480
rect -22120 -9500 -21880 -9480
rect -21620 -9500 -21380 -9480
rect -21120 -9500 -20880 -9480
rect -20620 -9500 -20380 -9480
rect -20120 -9500 -19880 -9480
rect -19620 -9500 -19380 -9480
rect -19120 -9500 -18880 -9480
rect -18620 -9500 -18380 -9480
rect -18120 -9500 -17880 -9480
rect -17620 -9500 -17380 -9480
rect -17120 -9500 -16880 -9480
rect -16620 -9500 -16380 -9480
rect -16120 -9500 -15880 -9480
rect -15620 -9500 -15380 -9480
rect -15120 -9500 -15000 -9480
rect -27500 -9700 -15000 -9500
rect -27500 -9720 -27380 -9700
rect -27120 -9720 -26880 -9700
rect -26620 -9720 -26380 -9700
rect -26120 -9720 -25880 -9700
rect -25620 -9720 -25380 -9700
rect -25120 -9720 -24880 -9700
rect -24620 -9720 -24380 -9700
rect -24120 -9720 -23880 -9700
rect -23620 -9720 -23380 -9700
rect -23120 -9720 -22880 -9700
rect -22620 -9720 -22380 -9700
rect -22120 -9720 -21880 -9700
rect -21620 -9720 -21380 -9700
rect -21120 -9720 -20880 -9700
rect -20620 -9720 -20380 -9700
rect -20120 -9720 -19880 -9700
rect -19620 -9720 -19380 -9700
rect -19120 -9720 -18880 -9700
rect -18620 -9720 -18380 -9700
rect -18120 -9720 -17880 -9700
rect -17620 -9720 -17380 -9700
rect -17120 -9720 -16880 -9700
rect -16620 -9720 -16380 -9700
rect -16120 -9720 -15880 -9700
rect -15620 -9720 -15380 -9700
rect -15120 -9720 -15000 -9700
rect -27500 -9980 -27400 -9720
rect -27100 -9980 -26900 -9720
rect -26600 -9980 -26400 -9720
rect -26100 -9980 -25900 -9720
rect -25600 -9980 -25400 -9720
rect -25100 -9980 -24900 -9720
rect -24600 -9980 -24400 -9720
rect -24100 -9980 -23900 -9720
rect -23600 -9980 -23400 -9720
rect -23100 -9980 -22900 -9720
rect -22600 -9980 -22400 -9720
rect -22100 -9980 -21900 -9720
rect -21600 -9980 -21400 -9720
rect -21100 -9980 -20900 -9720
rect -20600 -9980 -20400 -9720
rect -20100 -9980 -19900 -9720
rect -19600 -9980 -19400 -9720
rect -19100 -9980 -18900 -9720
rect -18600 -9980 -18400 -9720
rect -18100 -9980 -17900 -9720
rect -17600 -9980 -17400 -9720
rect -17100 -9980 -16900 -9720
rect -16600 -9980 -16400 -9720
rect -16100 -9980 -15900 -9720
rect -15600 -9980 -15400 -9720
rect -15100 -9980 -15000 -9720
rect -27500 -10000 -27380 -9980
rect -27120 -10000 -26880 -9980
rect -26620 -10000 -26380 -9980
rect -26120 -10000 -25880 -9980
rect -25620 -10000 -25380 -9980
rect -25120 -10000 -24880 -9980
rect -24620 -10000 -24380 -9980
rect -24120 -10000 -23880 -9980
rect -23620 -10000 -23380 -9980
rect -23120 -10000 -22880 -9980
rect -22620 -10000 -22380 -9980
rect -22120 -10000 -21880 -9980
rect -21620 -10000 -21380 -9980
rect -21120 -10000 -20880 -9980
rect -20620 -10000 -20380 -9980
rect -20120 -10000 -19880 -9980
rect -19620 -10000 -19380 -9980
rect -19120 -10000 -18880 -9980
rect -18620 -10000 -18380 -9980
rect -18120 -10000 -17880 -9980
rect -17620 -10000 -17380 -9980
rect -17120 -10000 -16880 -9980
rect -16620 -10000 -16380 -9980
rect -16120 -10000 -15880 -9980
rect -15620 -10000 -15380 -9980
rect -15120 -10000 -15000 -9980
rect -27500 -10200 -15000 -10000
rect -27500 -10220 -27380 -10200
rect -27120 -10220 -26880 -10200
rect -26620 -10220 -26380 -10200
rect -26120 -10220 -25880 -10200
rect -25620 -10220 -25380 -10200
rect -25120 -10220 -24880 -10200
rect -24620 -10220 -24380 -10200
rect -24120 -10220 -23880 -10200
rect -23620 -10220 -23380 -10200
rect -23120 -10220 -22880 -10200
rect -22620 -10220 -22380 -10200
rect -22120 -10220 -21880 -10200
rect -21620 -10220 -21380 -10200
rect -21120 -10220 -20880 -10200
rect -20620 -10220 -20380 -10200
rect -20120 -10220 -19880 -10200
rect -19620 -10220 -19380 -10200
rect -19120 -10220 -18880 -10200
rect -18620 -10220 -18380 -10200
rect -18120 -10220 -17880 -10200
rect -17620 -10220 -17380 -10200
rect -17120 -10220 -16880 -10200
rect -16620 -10220 -16380 -10200
rect -16120 -10220 -15880 -10200
rect -15620 -10220 -15380 -10200
rect -15120 -10220 -15000 -10200
rect -27500 -10480 -27400 -10220
rect -27100 -10480 -26900 -10220
rect -26600 -10480 -26400 -10220
rect -26100 -10480 -25900 -10220
rect -25600 -10480 -25400 -10220
rect -25100 -10480 -24900 -10220
rect -24600 -10480 -24400 -10220
rect -24100 -10480 -23900 -10220
rect -23600 -10480 -23400 -10220
rect -23100 -10480 -22900 -10220
rect -22600 -10480 -22400 -10220
rect -22100 -10480 -21900 -10220
rect -21600 -10480 -21400 -10220
rect -21100 -10480 -20900 -10220
rect -20600 -10480 -20400 -10220
rect -20100 -10480 -19900 -10220
rect -19600 -10480 -19400 -10220
rect -19100 -10480 -18900 -10220
rect -18600 -10480 -18400 -10220
rect -18100 -10480 -17900 -10220
rect -17600 -10480 -17400 -10220
rect -17100 -10480 -16900 -10220
rect -16600 -10480 -16400 -10220
rect -16100 -10480 -15900 -10220
rect -15600 -10480 -15400 -10220
rect -15100 -10480 -15000 -10220
rect -27500 -10500 -27380 -10480
rect -27120 -10500 -26880 -10480
rect -26620 -10500 -26380 -10480
rect -26120 -10500 -25880 -10480
rect -25620 -10500 -25380 -10480
rect -25120 -10500 -24880 -10480
rect -24620 -10500 -24380 -10480
rect -24120 -10500 -23880 -10480
rect -23620 -10500 -23380 -10480
rect -23120 -10500 -22880 -10480
rect -22620 -10500 -22380 -10480
rect -22120 -10500 -21880 -10480
rect -21620 -10500 -21380 -10480
rect -21120 -10500 -20880 -10480
rect -20620 -10500 -20380 -10480
rect -20120 -10500 -19880 -10480
rect -19620 -10500 -19380 -10480
rect -19120 -10500 -18880 -10480
rect -18620 -10500 -18380 -10480
rect -18120 -10500 -17880 -10480
rect -17620 -10500 -17380 -10480
rect -17120 -10500 -16880 -10480
rect -16620 -10500 -16380 -10480
rect -16120 -10500 -15880 -10480
rect -15620 -10500 -15380 -10480
rect -15120 -10500 -15000 -10480
rect -27500 -10700 -15000 -10500
rect -27500 -10720 -27380 -10700
rect -27120 -10720 -26880 -10700
rect -26620 -10720 -26380 -10700
rect -26120 -10720 -25880 -10700
rect -25620 -10720 -25380 -10700
rect -25120 -10720 -24880 -10700
rect -24620 -10720 -24380 -10700
rect -24120 -10720 -23880 -10700
rect -23620 -10720 -23380 -10700
rect -23120 -10720 -22880 -10700
rect -22620 -10720 -22380 -10700
rect -22120 -10720 -21880 -10700
rect -21620 -10720 -21380 -10700
rect -21120 -10720 -20880 -10700
rect -20620 -10720 -20380 -10700
rect -20120 -10720 -19880 -10700
rect -19620 -10720 -19380 -10700
rect -19120 -10720 -18880 -10700
rect -18620 -10720 -18380 -10700
rect -18120 -10720 -17880 -10700
rect -17620 -10720 -17380 -10700
rect -17120 -10720 -16880 -10700
rect -16620 -10720 -16380 -10700
rect -16120 -10720 -15880 -10700
rect -15620 -10720 -15380 -10700
rect -15120 -10720 -15000 -10700
rect -27500 -10980 -27400 -10720
rect -27100 -10980 -26900 -10720
rect -26600 -10980 -26400 -10720
rect -26100 -10980 -25900 -10720
rect -25600 -10980 -25400 -10720
rect -25100 -10980 -24900 -10720
rect -24600 -10980 -24400 -10720
rect -24100 -10980 -23900 -10720
rect -23600 -10980 -23400 -10720
rect -23100 -10980 -22900 -10720
rect -22600 -10980 -22400 -10720
rect -22100 -10980 -21900 -10720
rect -21600 -10980 -21400 -10720
rect -21100 -10980 -20900 -10720
rect -20600 -10980 -20400 -10720
rect -20100 -10980 -19900 -10720
rect -19600 -10980 -19400 -10720
rect -19100 -10980 -18900 -10720
rect -18600 -10980 -18400 -10720
rect -18100 -10980 -17900 -10720
rect -17600 -10980 -17400 -10720
rect -17100 -10980 -16900 -10720
rect -16600 -10980 -16400 -10720
rect -16100 -10980 -15900 -10720
rect -15600 -10980 -15400 -10720
rect -15100 -10980 -15000 -10720
rect -27500 -11000 -27380 -10980
rect -27120 -11000 -26880 -10980
rect -26620 -11000 -26380 -10980
rect -26120 -11000 -25880 -10980
rect -25620 -11000 -25380 -10980
rect -25120 -11000 -24880 -10980
rect -24620 -11000 -24380 -10980
rect -24120 -11000 -23880 -10980
rect -23620 -11000 -23380 -10980
rect -23120 -11000 -22880 -10980
rect -22620 -11000 -22380 -10980
rect -22120 -11000 -21880 -10980
rect -21620 -11000 -21380 -10980
rect -21120 -11000 -20880 -10980
rect -20620 -11000 -20380 -10980
rect -20120 -11000 -19880 -10980
rect -19620 -11000 -19380 -10980
rect -19120 -11000 -18880 -10980
rect -18620 -11000 -18380 -10980
rect -18120 -11000 -17880 -10980
rect -17620 -11000 -17380 -10980
rect -17120 -11000 -16880 -10980
rect -16620 -11000 -16380 -10980
rect -16120 -11000 -15880 -10980
rect -15620 -11000 -15380 -10980
rect -15120 -11000 -15000 -10980
rect -27500 -11200 -15000 -11000
rect -27500 -11220 -27380 -11200
rect -27120 -11220 -26880 -11200
rect -26620 -11220 -26380 -11200
rect -26120 -11220 -25880 -11200
rect -25620 -11220 -25380 -11200
rect -25120 -11220 -24880 -11200
rect -24620 -11220 -24380 -11200
rect -24120 -11220 -23880 -11200
rect -23620 -11220 -23380 -11200
rect -23120 -11220 -22880 -11200
rect -22620 -11220 -22380 -11200
rect -22120 -11220 -21880 -11200
rect -21620 -11220 -21380 -11200
rect -21120 -11220 -20880 -11200
rect -20620 -11220 -20380 -11200
rect -20120 -11220 -19880 -11200
rect -19620 -11220 -19380 -11200
rect -19120 -11220 -18880 -11200
rect -18620 -11220 -18380 -11200
rect -18120 -11220 -17880 -11200
rect -17620 -11220 -17380 -11200
rect -17120 -11220 -16880 -11200
rect -16620 -11220 -16380 -11200
rect -16120 -11220 -15880 -11200
rect -15620 -11220 -15380 -11200
rect -15120 -11220 -15000 -11200
rect -27500 -11480 -27400 -11220
rect -27100 -11480 -26900 -11220
rect -26600 -11480 -26400 -11220
rect -26100 -11480 -25900 -11220
rect -25600 -11480 -25400 -11220
rect -25100 -11480 -24900 -11220
rect -24600 -11480 -24400 -11220
rect -24100 -11480 -23900 -11220
rect -23600 -11480 -23400 -11220
rect -23100 -11480 -22900 -11220
rect -22600 -11480 -22400 -11220
rect -22100 -11480 -21900 -11220
rect -21600 -11480 -21400 -11220
rect -21100 -11480 -20900 -11220
rect -20600 -11480 -20400 -11220
rect -20100 -11480 -19900 -11220
rect -19600 -11480 -19400 -11220
rect -19100 -11480 -18900 -11220
rect -18600 -11480 -18400 -11220
rect -18100 -11480 -17900 -11220
rect -17600 -11480 -17400 -11220
rect -17100 -11480 -16900 -11220
rect -16600 -11480 -16400 -11220
rect -16100 -11480 -15900 -11220
rect -15600 -11480 -15400 -11220
rect -15100 -11480 -15000 -11220
rect -27500 -11500 -27380 -11480
rect -27120 -11500 -26880 -11480
rect -26620 -11500 -26380 -11480
rect -26120 -11500 -25880 -11480
rect -25620 -11500 -25380 -11480
rect -25120 -11500 -24880 -11480
rect -24620 -11500 -24380 -11480
rect -24120 -11500 -23880 -11480
rect -23620 -11500 -23380 -11480
rect -23120 -11500 -22880 -11480
rect -22620 -11500 -22380 -11480
rect -22120 -11500 -21880 -11480
rect -21620 -11500 -21380 -11480
rect -21120 -11500 -20880 -11480
rect -20620 -11500 -20380 -11480
rect -20120 -11500 -19880 -11480
rect -19620 -11500 -19380 -11480
rect -19120 -11500 -18880 -11480
rect -18620 -11500 -18380 -11480
rect -18120 -11500 -17880 -11480
rect -17620 -11500 -17380 -11480
rect -17120 -11500 -16880 -11480
rect -16620 -11500 -16380 -11480
rect -16120 -11500 -15880 -11480
rect -15620 -11500 -15380 -11480
rect -15120 -11500 -15000 -11480
rect -27500 -11600 -15000 -11500
rect -27500 -11700 -18200 -11600
rect -18000 -11700 -15000 -11600
rect -27500 -11720 -27380 -11700
rect -27120 -11720 -26880 -11700
rect -26620 -11720 -26380 -11700
rect -26120 -11720 -25880 -11700
rect -25620 -11720 -25380 -11700
rect -25120 -11720 -24880 -11700
rect -24620 -11720 -24380 -11700
rect -24120 -11720 -23880 -11700
rect -23620 -11720 -23380 -11700
rect -23120 -11720 -22880 -11700
rect -22620 -11720 -22380 -11700
rect -22120 -11720 -21880 -11700
rect -21620 -11720 -21380 -11700
rect -21120 -11720 -20880 -11700
rect -20620 -11720 -20380 -11700
rect -20120 -11720 -19880 -11700
rect -19620 -11720 -19380 -11700
rect -19120 -11720 -18880 -11700
rect -18620 -11720 -18380 -11700
rect -18000 -11720 -17880 -11700
rect -17620 -11720 -17380 -11700
rect -17120 -11720 -16880 -11700
rect -16620 -11720 -16380 -11700
rect -16120 -11720 -15880 -11700
rect -15620 -11720 -15380 -11700
rect -15120 -11720 -15000 -11700
rect -27500 -11980 -27400 -11720
rect -27100 -11980 -26900 -11720
rect -26600 -11980 -26400 -11720
rect -26100 -11980 -25900 -11720
rect -25600 -11980 -25400 -11720
rect -25100 -11980 -24900 -11720
rect -24600 -11980 -24400 -11720
rect -24100 -11980 -23900 -11720
rect -23600 -11980 -23400 -11720
rect -23100 -11980 -22900 -11720
rect -22600 -11980 -22400 -11720
rect -22100 -11980 -21900 -11720
rect -21600 -11980 -21400 -11720
rect -21100 -11980 -20900 -11720
rect -20600 -11980 -20400 -11720
rect -20100 -11980 -19900 -11720
rect -19600 -11980 -19400 -11720
rect -19100 -11980 -18900 -11720
rect -18600 -11980 -18400 -11720
rect -18000 -11900 -17900 -11720
rect -18100 -11980 -17900 -11900
rect -17600 -11980 -17400 -11720
rect -17100 -11980 -16900 -11720
rect -16600 -11980 -16400 -11720
rect -16100 -11980 -15900 -11720
rect -15600 -11980 -15400 -11720
rect -15100 -11980 -15000 -11720
rect -27500 -12000 -27380 -11980
rect -27120 -12000 -26880 -11980
rect -26620 -12000 -26380 -11980
rect -26120 -12000 -25880 -11980
rect -25620 -12000 -25380 -11980
rect -25120 -12000 -24880 -11980
rect -24620 -12000 -24380 -11980
rect -24120 -12000 -23880 -11980
rect -23620 -12000 -23380 -11980
rect -23120 -12000 -22880 -11980
rect -22620 -12000 -22380 -11980
rect -22120 -12000 -21880 -11980
rect -21620 -12000 -21380 -11980
rect -21120 -12000 -20880 -11980
rect -20620 -12000 -20380 -11980
rect -20120 -12000 -19880 -11980
rect -19620 -12000 -19380 -11980
rect -19120 -12000 -18880 -11980
rect -18620 -12000 -18380 -11980
rect -18120 -12000 -17880 -11980
rect -17620 -12000 -17380 -11980
rect -17120 -12000 -16880 -11980
rect -16620 -12000 -16380 -11980
rect -16120 -12000 -15880 -11980
rect -15620 -12000 -15380 -11980
rect -15120 -12000 -15000 -11980
rect -27500 -12200 -15000 -12000
rect -27500 -12220 -27380 -12200
rect -27120 -12220 -26880 -12200
rect -26620 -12220 -26380 -12200
rect -26120 -12220 -25880 -12200
rect -25620 -12220 -25380 -12200
rect -25120 -12220 -24880 -12200
rect -24620 -12220 -24380 -12200
rect -24120 -12220 -23880 -12200
rect -23620 -12220 -23380 -12200
rect -23120 -12220 -22880 -12200
rect -22620 -12220 -22380 -12200
rect -22120 -12220 -21880 -12200
rect -21620 -12220 -21380 -12200
rect -21120 -12220 -20880 -12200
rect -20620 -12220 -20380 -12200
rect -20120 -12220 -19880 -12200
rect -19620 -12220 -19380 -12200
rect -19120 -12220 -18880 -12200
rect -18620 -12220 -18380 -12200
rect -18120 -12220 -17880 -12200
rect -17620 -12220 -17380 -12200
rect -17120 -12220 -16880 -12200
rect -16620 -12220 -16380 -12200
rect -16120 -12220 -15880 -12200
rect -15620 -12220 -15380 -12200
rect -15120 -12220 -15000 -12200
rect -27500 -12480 -27400 -12220
rect -27100 -12480 -26900 -12220
rect -26600 -12480 -26400 -12220
rect -26100 -12480 -25900 -12220
rect -25600 -12480 -25400 -12220
rect -25100 -12480 -24900 -12220
rect -24600 -12480 -24400 -12220
rect -24100 -12480 -23900 -12220
rect -23600 -12480 -23400 -12220
rect -23100 -12480 -22900 -12220
rect -22600 -12480 -22400 -12220
rect -22100 -12480 -21900 -12220
rect -21600 -12480 -21400 -12220
rect -21100 -12480 -20900 -12220
rect -20600 -12480 -20400 -12220
rect -20100 -12480 -19900 -12220
rect -19600 -12480 -19400 -12220
rect -19100 -12480 -18900 -12220
rect -18600 -12480 -18400 -12220
rect -18100 -12480 -17900 -12220
rect -17600 -12480 -17400 -12220
rect -17100 -12480 -16900 -12220
rect -16600 -12480 -16400 -12220
rect -16100 -12480 -15900 -12220
rect -15600 -12480 -15400 -12220
rect -15100 -12480 -15000 -12220
rect -27500 -12500 -27380 -12480
rect -27120 -12500 -26880 -12480
rect -26620 -12500 -26380 -12480
rect -26120 -12500 -25880 -12480
rect -25620 -12500 -25380 -12480
rect -25120 -12500 -24880 -12480
rect -24620 -12500 -24380 -12480
rect -24120 -12500 -23880 -12480
rect -23620 -12500 -23380 -12480
rect -23120 -12500 -22880 -12480
rect -22620 -12500 -22380 -12480
rect -22120 -12500 -21880 -12480
rect -21620 -12500 -21380 -12480
rect -21120 -12500 -20880 -12480
rect -20620 -12500 -20380 -12480
rect -20120 -12500 -19880 -12480
rect -19620 -12500 -19380 -12480
rect -19120 -12500 -18880 -12480
rect -18620 -12500 -18380 -12480
rect -18120 -12500 -17880 -12480
rect -17620 -12500 -17380 -12480
rect -17120 -12500 -16880 -12480
rect -16620 -12500 -16380 -12480
rect -16120 -12500 -15880 -12480
rect -15620 -12500 -15380 -12480
rect -15120 -12500 -15000 -12480
rect -27500 -12700 -15000 -12500
rect -27500 -12720 -27380 -12700
rect -27120 -12720 -26880 -12700
rect -26620 -12720 -26380 -12700
rect -26120 -12720 -25880 -12700
rect -25620 -12720 -25380 -12700
rect -25120 -12720 -24880 -12700
rect -24620 -12720 -24380 -12700
rect -24120 -12720 -23880 -12700
rect -23620 -12720 -23380 -12700
rect -23120 -12720 -22880 -12700
rect -22620 -12720 -22380 -12700
rect -22120 -12720 -21880 -12700
rect -21620 -12720 -21380 -12700
rect -21120 -12720 -20880 -12700
rect -20620 -12720 -20380 -12700
rect -20120 -12720 -19880 -12700
rect -19620 -12720 -19380 -12700
rect -19120 -12720 -18880 -12700
rect -18620 -12720 -18380 -12700
rect -18120 -12720 -17880 -12700
rect -17620 -12720 -17380 -12700
rect -17120 -12720 -16880 -12700
rect -16620 -12720 -16380 -12700
rect -16120 -12720 -15880 -12700
rect -15620 -12720 -15380 -12700
rect -15120 -12720 -15000 -12700
rect -27500 -12980 -27400 -12720
rect -27100 -12980 -26900 -12720
rect -26600 -12980 -26400 -12720
rect -26100 -12980 -25900 -12720
rect -25600 -12980 -25400 -12720
rect -25100 -12980 -24900 -12720
rect -24600 -12980 -24400 -12720
rect -24100 -12980 -23900 -12720
rect -23600 -12980 -23400 -12720
rect -23100 -12980 -22900 -12720
rect -22600 -12980 -22400 -12720
rect -22100 -12980 -21900 -12720
rect -21600 -12980 -21400 -12720
rect -21100 -12980 -20900 -12720
rect -20600 -12980 -20400 -12720
rect -20100 -12980 -19900 -12720
rect -19600 -12980 -19400 -12720
rect -19100 -12980 -18900 -12720
rect -18600 -12980 -18400 -12720
rect -18100 -12980 -17900 -12720
rect -17600 -12980 -17400 -12720
rect -17100 -12980 -16900 -12720
rect -16600 -12980 -16400 -12720
rect -16100 -12980 -15900 -12720
rect -15600 -12980 -15400 -12720
rect -15100 -12980 -15000 -12720
rect -27500 -13000 -27380 -12980
rect -27120 -13000 -26880 -12980
rect -26620 -13000 -26380 -12980
rect -26120 -13000 -25880 -12980
rect -25620 -13000 -25380 -12980
rect -25120 -13000 -24880 -12980
rect -24620 -13000 -24380 -12980
rect -24120 -13000 -23880 -12980
rect -23620 -13000 -23380 -12980
rect -23120 -13000 -22880 -12980
rect -22620 -13000 -22380 -12980
rect -22120 -13000 -21880 -12980
rect -21620 -13000 -21380 -12980
rect -21120 -13000 -20880 -12980
rect -20620 -13000 -20380 -12980
rect -20120 -13000 -19880 -12980
rect -19620 -13000 -19380 -12980
rect -19120 -13000 -18880 -12980
rect -18620 -13000 -18380 -12980
rect -18120 -13000 -17880 -12980
rect -17620 -13000 -17380 -12980
rect -17120 -13000 -16880 -12980
rect -16620 -13000 -16380 -12980
rect -16120 -13000 -15880 -12980
rect -15620 -13000 -15380 -12980
rect -15120 -13000 -15000 -12980
rect -27500 -13200 -15000 -13000
rect 14500 -3700 33500 -3600
rect 14500 -3720 14620 -3700
rect 14880 -3720 15120 -3700
rect 15380 -3720 15620 -3700
rect 15880 -3720 16120 -3700
rect 16380 -3720 16620 -3700
rect 16880 -3720 17120 -3700
rect 17380 -3720 17620 -3700
rect 17880 -3720 18120 -3700
rect 18380 -3720 18620 -3700
rect 18880 -3720 19120 -3700
rect 19380 -3720 19620 -3700
rect 19880 -3720 20120 -3700
rect 20380 -3720 20620 -3700
rect 20880 -3720 21120 -3700
rect 21380 -3720 21620 -3700
rect 21880 -3720 22120 -3700
rect 22380 -3720 22620 -3700
rect 22880 -3720 23120 -3700
rect 23380 -3720 23620 -3700
rect 23880 -3720 24120 -3700
rect 24380 -3720 24620 -3700
rect 24880 -3720 25120 -3700
rect 25380 -3720 25620 -3700
rect 25880 -3720 26120 -3700
rect 26380 -3720 26620 -3700
rect 26880 -3720 27120 -3700
rect 27380 -3720 27620 -3700
rect 27880 -3720 28120 -3700
rect 28380 -3720 28620 -3700
rect 28880 -3720 29120 -3700
rect 29380 -3720 29620 -3700
rect 29880 -3720 30120 -3700
rect 30380 -3720 30620 -3700
rect 30880 -3720 31120 -3700
rect 31380 -3720 31620 -3700
rect 31880 -3720 32120 -3700
rect 32380 -3720 32620 -3700
rect 32880 -3720 33120 -3700
rect 33380 -3720 33500 -3700
rect 14500 -3980 14600 -3720
rect 14900 -3980 15100 -3720
rect 15400 -3980 15600 -3720
rect 15900 -3980 16100 -3720
rect 16400 -3980 16600 -3720
rect 16900 -3980 17100 -3720
rect 17400 -3980 17600 -3720
rect 17900 -3980 18100 -3720
rect 18400 -3980 18600 -3720
rect 18900 -3980 19100 -3720
rect 19400 -3980 19600 -3720
rect 19900 -3980 20100 -3720
rect 20400 -3980 20600 -3720
rect 20900 -3980 21100 -3720
rect 21400 -3980 21600 -3720
rect 21900 -3980 22100 -3720
rect 22400 -3980 22600 -3720
rect 22900 -3980 23100 -3720
rect 23400 -3980 23600 -3720
rect 23900 -3980 24100 -3720
rect 24400 -3980 24600 -3720
rect 24900 -3980 25100 -3720
rect 25400 -3980 25600 -3720
rect 25900 -3980 26100 -3720
rect 26400 -3980 26600 -3720
rect 26900 -3980 27100 -3720
rect 27400 -3980 27600 -3720
rect 27900 -3980 28100 -3720
rect 28400 -3980 28600 -3720
rect 28900 -3980 29100 -3720
rect 29400 -3980 29600 -3720
rect 29900 -3980 30100 -3720
rect 30400 -3980 30600 -3720
rect 30900 -3980 31100 -3720
rect 31400 -3980 31600 -3720
rect 31900 -3980 32100 -3720
rect 32400 -3980 32600 -3720
rect 32900 -3980 33100 -3720
rect 33400 -3980 33500 -3720
rect 14500 -4000 14620 -3980
rect 14880 -4000 15120 -3980
rect 15380 -4000 15620 -3980
rect 15880 -4000 16120 -3980
rect 16380 -4000 16620 -3980
rect 16880 -4000 17120 -3980
rect 17380 -4000 17620 -3980
rect 17880 -4000 18120 -3980
rect 18380 -4000 18620 -3980
rect 18880 -4000 19120 -3980
rect 19380 -4000 19620 -3980
rect 19880 -4000 20120 -3980
rect 20380 -4000 20620 -3980
rect 20880 -4000 21120 -3980
rect 21380 -4000 21620 -3980
rect 21880 -4000 22120 -3980
rect 22380 -4000 22620 -3980
rect 22880 -4000 23120 -3980
rect 23380 -4000 23620 -3980
rect 23880 -4000 24120 -3980
rect 24380 -4000 24620 -3980
rect 24880 -4000 25120 -3980
rect 25380 -4000 25620 -3980
rect 25880 -4000 26120 -3980
rect 26380 -4000 26620 -3980
rect 26880 -4000 27120 -3980
rect 27380 -4000 27620 -3980
rect 27880 -4000 28120 -3980
rect 28380 -4000 28620 -3980
rect 28880 -4000 29120 -3980
rect 29380 -4000 29620 -3980
rect 29880 -4000 30120 -3980
rect 30380 -4000 30620 -3980
rect 30880 -4000 31120 -3980
rect 31380 -4000 31620 -3980
rect 31880 -4000 32120 -3980
rect 32380 -4000 32620 -3980
rect 32880 -4000 33120 -3980
rect 33380 -4000 33500 -3980
rect 14500 -4200 33500 -4000
rect 14500 -4220 14620 -4200
rect 14880 -4220 15120 -4200
rect 15380 -4220 15620 -4200
rect 15880 -4220 16120 -4200
rect 16380 -4220 16620 -4200
rect 16880 -4220 17120 -4200
rect 17380 -4220 17620 -4200
rect 17880 -4220 18120 -4200
rect 18380 -4220 18620 -4200
rect 18880 -4220 19120 -4200
rect 19380 -4220 19620 -4200
rect 19880 -4220 20120 -4200
rect 20380 -4220 20620 -4200
rect 20880 -4220 21120 -4200
rect 21380 -4220 21620 -4200
rect 21880 -4220 22120 -4200
rect 22380 -4220 22620 -4200
rect 22880 -4220 23120 -4200
rect 23380 -4220 23620 -4200
rect 23880 -4220 24120 -4200
rect 24380 -4220 24620 -4200
rect 24880 -4220 25120 -4200
rect 25380 -4220 25620 -4200
rect 25880 -4220 26120 -4200
rect 26380 -4220 26620 -4200
rect 26880 -4220 27120 -4200
rect 27380 -4220 27620 -4200
rect 27880 -4220 28120 -4200
rect 28380 -4220 28620 -4200
rect 28880 -4220 29120 -4200
rect 29380 -4220 29620 -4200
rect 29880 -4220 30120 -4200
rect 30380 -4220 30620 -4200
rect 30880 -4220 31120 -4200
rect 31380 -4220 31620 -4200
rect 31880 -4220 32120 -4200
rect 32380 -4220 32620 -4200
rect 32880 -4220 33120 -4200
rect 33380 -4220 33500 -4200
rect 14500 -4480 14600 -4220
rect 14900 -4480 15100 -4220
rect 15400 -4480 15600 -4220
rect 15900 -4480 16100 -4220
rect 16400 -4480 16600 -4220
rect 16900 -4480 17100 -4220
rect 17400 -4480 17600 -4220
rect 17900 -4480 18100 -4220
rect 18400 -4480 18600 -4220
rect 18900 -4480 19100 -4220
rect 19400 -4480 19600 -4220
rect 19900 -4480 20100 -4220
rect 20400 -4480 20600 -4220
rect 20900 -4480 21100 -4220
rect 21400 -4480 21600 -4220
rect 21900 -4480 22100 -4220
rect 22400 -4480 22600 -4220
rect 22900 -4480 23100 -4220
rect 23400 -4480 23600 -4220
rect 23900 -4480 24100 -4220
rect 24400 -4480 24600 -4220
rect 24900 -4480 25100 -4220
rect 25400 -4480 25600 -4220
rect 25900 -4480 26100 -4220
rect 26400 -4480 26600 -4220
rect 26900 -4480 27100 -4220
rect 27400 -4480 27600 -4220
rect 27900 -4480 28100 -4220
rect 28400 -4480 28600 -4220
rect 28900 -4480 29100 -4220
rect 29400 -4480 29600 -4220
rect 29900 -4480 30100 -4220
rect 30400 -4480 30600 -4220
rect 30900 -4480 31100 -4220
rect 31400 -4480 31600 -4220
rect 31900 -4480 32100 -4220
rect 32400 -4480 32600 -4220
rect 32900 -4480 33100 -4220
rect 33400 -4480 33500 -4220
rect 14500 -4500 14620 -4480
rect 14880 -4500 15120 -4480
rect 15380 -4500 15620 -4480
rect 15880 -4500 16120 -4480
rect 16380 -4500 16620 -4480
rect 16880 -4500 17120 -4480
rect 17380 -4500 17620 -4480
rect 17880 -4500 18120 -4480
rect 18380 -4500 18620 -4480
rect 18880 -4500 19120 -4480
rect 19380 -4500 19620 -4480
rect 19880 -4500 20120 -4480
rect 20380 -4500 20620 -4480
rect 20880 -4500 21120 -4480
rect 21380 -4500 21620 -4480
rect 21880 -4500 22120 -4480
rect 22380 -4500 22620 -4480
rect 22880 -4500 23120 -4480
rect 23380 -4500 23620 -4480
rect 23880 -4500 24120 -4480
rect 24380 -4500 24620 -4480
rect 24880 -4500 25120 -4480
rect 25380 -4500 25620 -4480
rect 25880 -4500 26120 -4480
rect 26380 -4500 26620 -4480
rect 26880 -4500 27120 -4480
rect 27380 -4500 27620 -4480
rect 27880 -4500 28120 -4480
rect 28380 -4500 28620 -4480
rect 28880 -4500 29120 -4480
rect 29380 -4500 29620 -4480
rect 29880 -4500 30120 -4480
rect 30380 -4500 30620 -4480
rect 30880 -4500 31120 -4480
rect 31380 -4500 31620 -4480
rect 31880 -4500 32120 -4480
rect 32380 -4500 32620 -4480
rect 32880 -4500 33120 -4480
rect 33380 -4500 33500 -4480
rect 14500 -4700 33500 -4500
rect 14500 -4720 14620 -4700
rect 14880 -4720 15120 -4700
rect 15380 -4720 15620 -4700
rect 15880 -4720 16120 -4700
rect 16380 -4720 16620 -4700
rect 16880 -4720 17120 -4700
rect 17380 -4720 17620 -4700
rect 17880 -4720 18120 -4700
rect 18380 -4720 18620 -4700
rect 18880 -4720 19120 -4700
rect 19380 -4720 19620 -4700
rect 19880 -4720 20120 -4700
rect 20380 -4720 20620 -4700
rect 20880 -4720 21120 -4700
rect 21380 -4720 21620 -4700
rect 21880 -4720 22120 -4700
rect 22380 -4720 22620 -4700
rect 22880 -4720 23120 -4700
rect 23380 -4720 23620 -4700
rect 23880 -4720 24120 -4700
rect 24380 -4720 24620 -4700
rect 24880 -4720 25120 -4700
rect 25380 -4720 25620 -4700
rect 25880 -4720 26120 -4700
rect 26380 -4720 26620 -4700
rect 26880 -4720 27120 -4700
rect 27380 -4720 27620 -4700
rect 27880 -4720 28120 -4700
rect 28380 -4720 28620 -4700
rect 28880 -4720 29120 -4700
rect 29380 -4720 29620 -4700
rect 29880 -4720 30120 -4700
rect 30380 -4720 30620 -4700
rect 30880 -4720 31120 -4700
rect 31380 -4720 31620 -4700
rect 31880 -4720 32120 -4700
rect 32380 -4720 32620 -4700
rect 32880 -4720 33120 -4700
rect 33380 -4720 33500 -4700
rect 14500 -4980 14600 -4720
rect 14900 -4980 15100 -4720
rect 15400 -4980 15600 -4720
rect 15900 -4980 16100 -4720
rect 16400 -4980 16600 -4720
rect 16900 -4980 17100 -4720
rect 17400 -4980 17600 -4720
rect 17900 -4980 18100 -4720
rect 18400 -4980 18600 -4720
rect 18900 -4980 19100 -4720
rect 19400 -4980 19600 -4720
rect 19900 -4980 20100 -4720
rect 20400 -4980 20600 -4720
rect 20900 -4980 21100 -4720
rect 21400 -4980 21600 -4720
rect 21900 -4980 22100 -4720
rect 22400 -4980 22600 -4720
rect 22900 -4980 23100 -4720
rect 23400 -4980 23600 -4720
rect 23900 -4980 24100 -4720
rect 24400 -4980 24600 -4720
rect 24900 -4980 25100 -4720
rect 25400 -4980 25600 -4720
rect 25900 -4980 26100 -4720
rect 26400 -4980 26600 -4720
rect 26900 -4980 27100 -4720
rect 27400 -4980 27600 -4720
rect 27900 -4980 28100 -4720
rect 28400 -4980 28600 -4720
rect 28900 -4980 29100 -4720
rect 29400 -4980 29600 -4720
rect 29900 -4980 30100 -4720
rect 30400 -4980 30600 -4720
rect 30900 -4980 31100 -4720
rect 31400 -4980 31600 -4720
rect 31900 -4980 32100 -4720
rect 32400 -4980 32600 -4720
rect 32900 -4980 33100 -4720
rect 33400 -4980 33500 -4720
rect 14500 -5000 14620 -4980
rect 14880 -5000 15120 -4980
rect 15380 -5000 15620 -4980
rect 15880 -5000 16120 -4980
rect 16380 -5000 16620 -4980
rect 16880 -5000 17120 -4980
rect 17380 -5000 17620 -4980
rect 17880 -5000 18120 -4980
rect 18380 -5000 18620 -4980
rect 18880 -5000 19120 -4980
rect 19380 -5000 19620 -4980
rect 19880 -5000 20120 -4980
rect 20380 -5000 20620 -4980
rect 20880 -5000 21120 -4980
rect 21380 -5000 21620 -4980
rect 21880 -5000 22120 -4980
rect 22380 -5000 22620 -4980
rect 22880 -5000 23120 -4980
rect 23380 -5000 23620 -4980
rect 23880 -5000 24120 -4980
rect 24380 -5000 24620 -4980
rect 24880 -5000 25120 -4980
rect 25380 -5000 25620 -4980
rect 25880 -5000 26120 -4980
rect 26380 -5000 26620 -4980
rect 26880 -5000 27120 -4980
rect 27380 -5000 27620 -4980
rect 27880 -5000 28120 -4980
rect 28380 -5000 28620 -4980
rect 28880 -5000 29120 -4980
rect 29380 -5000 29620 -4980
rect 29880 -5000 30120 -4980
rect 30380 -5000 30620 -4980
rect 30880 -5000 31120 -4980
rect 31380 -5000 31620 -4980
rect 31880 -5000 32120 -4980
rect 32380 -5000 32620 -4980
rect 32880 -5000 33120 -4980
rect 33380 -5000 33500 -4980
rect 14500 -5200 33500 -5000
rect 14500 -5220 14620 -5200
rect 14880 -5220 15120 -5200
rect 15380 -5220 15620 -5200
rect 15880 -5220 16120 -5200
rect 16380 -5220 16620 -5200
rect 16880 -5220 17120 -5200
rect 17380 -5220 17620 -5200
rect 17880 -5220 18120 -5200
rect 18380 -5220 18620 -5200
rect 18880 -5220 19120 -5200
rect 19380 -5220 19620 -5200
rect 19880 -5220 20120 -5200
rect 20380 -5220 20620 -5200
rect 20880 -5220 21120 -5200
rect 21380 -5220 21620 -5200
rect 21880 -5220 22120 -5200
rect 22380 -5220 22620 -5200
rect 22880 -5220 23120 -5200
rect 23380 -5220 23620 -5200
rect 23880 -5220 24120 -5200
rect 24380 -5220 24620 -5200
rect 24880 -5220 25120 -5200
rect 25380 -5220 25620 -5200
rect 25880 -5220 26120 -5200
rect 26380 -5220 26620 -5200
rect 26880 -5220 27120 -5200
rect 27380 -5220 27620 -5200
rect 27880 -5220 28120 -5200
rect 28380 -5220 28620 -5200
rect 28880 -5220 29120 -5200
rect 29380 -5220 29620 -5200
rect 29880 -5220 30120 -5200
rect 30380 -5220 30620 -5200
rect 30880 -5220 31120 -5200
rect 31380 -5220 31620 -5200
rect 31880 -5220 32120 -5200
rect 32380 -5220 32620 -5200
rect 32880 -5220 33120 -5200
rect 33380 -5220 33500 -5200
rect 14500 -5480 14600 -5220
rect 14900 -5480 15100 -5220
rect 15400 -5480 15600 -5220
rect 15900 -5480 16100 -5220
rect 16400 -5480 16600 -5220
rect 16900 -5480 17100 -5220
rect 17400 -5480 17600 -5220
rect 17900 -5480 18100 -5220
rect 18400 -5480 18600 -5220
rect 18900 -5480 19100 -5220
rect 19400 -5480 19600 -5220
rect 19900 -5480 20100 -5220
rect 20400 -5480 20600 -5220
rect 20900 -5480 21100 -5220
rect 21400 -5480 21600 -5220
rect 21900 -5480 22100 -5220
rect 22400 -5480 22600 -5220
rect 22900 -5480 23100 -5220
rect 23400 -5480 23600 -5220
rect 23900 -5480 24100 -5220
rect 24400 -5480 24600 -5220
rect 24900 -5480 25100 -5220
rect 25400 -5480 25600 -5220
rect 25900 -5480 26100 -5220
rect 26400 -5480 26600 -5220
rect 26900 -5480 27100 -5220
rect 27400 -5480 27600 -5220
rect 27900 -5480 28100 -5220
rect 28400 -5480 28600 -5220
rect 28900 -5480 29100 -5220
rect 29400 -5480 29600 -5220
rect 29900 -5480 30100 -5220
rect 30400 -5480 30600 -5220
rect 30900 -5480 31100 -5220
rect 31400 -5480 31600 -5220
rect 31900 -5480 32100 -5220
rect 32400 -5480 32600 -5220
rect 32900 -5480 33100 -5220
rect 33400 -5480 33500 -5220
rect 14500 -5500 14620 -5480
rect 14880 -5500 15120 -5480
rect 15380 -5500 15620 -5480
rect 15880 -5500 16120 -5480
rect 16380 -5500 16620 -5480
rect 16880 -5500 17120 -5480
rect 17380 -5500 17620 -5480
rect 17880 -5500 18120 -5480
rect 18380 -5500 18620 -5480
rect 18880 -5500 19120 -5480
rect 19380 -5500 19620 -5480
rect 19880 -5500 20120 -5480
rect 20380 -5500 20620 -5480
rect 20880 -5500 21120 -5480
rect 21380 -5500 21620 -5480
rect 21880 -5500 22120 -5480
rect 22380 -5500 22620 -5480
rect 22880 -5500 23120 -5480
rect 23380 -5500 23620 -5480
rect 23880 -5500 24120 -5480
rect 24380 -5500 24620 -5480
rect 24880 -5500 25120 -5480
rect 25380 -5500 25620 -5480
rect 25880 -5500 26120 -5480
rect 26380 -5500 26620 -5480
rect 26880 -5500 27120 -5480
rect 27380 -5500 27620 -5480
rect 27880 -5500 28120 -5480
rect 28380 -5500 28620 -5480
rect 28880 -5500 29120 -5480
rect 29380 -5500 29620 -5480
rect 29880 -5500 30120 -5480
rect 30380 -5500 30620 -5480
rect 30880 -5500 31120 -5480
rect 31380 -5500 31620 -5480
rect 31880 -5500 32120 -5480
rect 32380 -5500 32620 -5480
rect 32880 -5500 33120 -5480
rect 33380 -5500 33500 -5480
rect 14500 -5600 33500 -5500
rect 14500 -5700 24000 -5600
rect 14500 -5720 14620 -5700
rect 14880 -5720 15120 -5700
rect 15380 -5720 15620 -5700
rect 15880 -5720 16120 -5700
rect 16380 -5720 16620 -5700
rect 16880 -5720 17120 -5700
rect 17380 -5720 17620 -5700
rect 17880 -5720 18120 -5700
rect 18380 -5720 18620 -5700
rect 18880 -5720 19120 -5700
rect 19380 -5720 19620 -5700
rect 19880 -5720 20120 -5700
rect 20380 -5720 20620 -5700
rect 20880 -5720 21120 -5700
rect 21380 -5720 21620 -5700
rect 21880 -5720 22120 -5700
rect 22380 -5720 22620 -5700
rect 22880 -5720 23120 -5700
rect 23380 -5720 23620 -5700
rect 23880 -5720 24000 -5700
rect 14500 -5980 14600 -5720
rect 14900 -5980 15100 -5720
rect 15400 -5980 15600 -5720
rect 15900 -5980 16100 -5720
rect 16400 -5980 16600 -5720
rect 16900 -5980 17100 -5720
rect 17400 -5980 17600 -5720
rect 17900 -5980 18100 -5720
rect 18400 -5980 18600 -5720
rect 18900 -5980 19100 -5720
rect 19400 -5980 19600 -5720
rect 19900 -5980 20100 -5720
rect 20400 -5980 20600 -5720
rect 20900 -5980 21100 -5720
rect 21400 -5980 21600 -5720
rect 21900 -5980 22100 -5720
rect 22400 -5980 22600 -5720
rect 22900 -5980 23100 -5720
rect 23400 -5980 23600 -5720
rect 23900 -5980 24000 -5720
rect 14500 -6000 14620 -5980
rect 14880 -6000 15120 -5980
rect 15380 -6000 15620 -5980
rect 15880 -6000 16120 -5980
rect 16380 -6000 16620 -5980
rect 16880 -6000 17120 -5980
rect 17380 -6000 17620 -5980
rect 17880 -6000 18120 -5980
rect 18380 -6000 18620 -5980
rect 18880 -6000 19120 -5980
rect 19380 -6000 19620 -5980
rect 19880 -6000 20120 -5980
rect 20380 -6000 20620 -5980
rect 20880 -6000 21120 -5980
rect 21380 -6000 21620 -5980
rect 21880 -6000 22120 -5980
rect 22380 -6000 22620 -5980
rect 22880 -6000 23120 -5980
rect 23380 -6000 23620 -5980
rect 23880 -6000 24000 -5980
rect 14500 -6200 24000 -6000
rect 14500 -6220 14620 -6200
rect 14880 -6220 15120 -6200
rect 15380 -6220 15620 -6200
rect 15880 -6220 16120 -6200
rect 16380 -6220 16620 -6200
rect 16880 -6220 17120 -6200
rect 17380 -6220 17620 -6200
rect 17880 -6220 18120 -6200
rect 18380 -6220 18620 -6200
rect 18880 -6220 19120 -6200
rect 19380 -6220 19620 -6200
rect 19880 -6220 20120 -6200
rect 20380 -6220 20620 -6200
rect 20880 -6220 21120 -6200
rect 21380 -6220 21620 -6200
rect 21880 -6220 22120 -6200
rect 22380 -6220 22620 -6200
rect 22880 -6220 23120 -6200
rect 23380 -6220 23620 -6200
rect 23880 -6220 24000 -6200
rect 14500 -6480 14600 -6220
rect 14900 -6480 15100 -6220
rect 15400 -6480 15600 -6220
rect 15900 -6480 16100 -6220
rect 16400 -6480 16600 -6220
rect 16900 -6480 17100 -6220
rect 17400 -6480 17600 -6220
rect 17900 -6480 18100 -6220
rect 18400 -6480 18600 -6220
rect 18900 -6480 19100 -6220
rect 19400 -6480 19600 -6220
rect 19900 -6480 20100 -6220
rect 20400 -6480 20600 -6220
rect 20900 -6480 21100 -6220
rect 21400 -6480 21600 -6220
rect 21900 -6480 22100 -6220
rect 22400 -6480 22600 -6220
rect 22900 -6480 23100 -6220
rect 23400 -6480 23600 -6220
rect 23900 -6480 24000 -6220
rect 14500 -6500 14620 -6480
rect 14880 -6500 15120 -6480
rect 15380 -6500 15620 -6480
rect 15880 -6500 16120 -6480
rect 16380 -6500 16620 -6480
rect 16880 -6500 17120 -6480
rect 17380 -6500 17620 -6480
rect 17880 -6500 18120 -6480
rect 18380 -6500 18620 -6480
rect 18880 -6500 19120 -6480
rect 19380 -6500 19620 -6480
rect 19880 -6500 20120 -6480
rect 20380 -6500 20620 -6480
rect 20880 -6500 21120 -6480
rect 21380 -6500 21620 -6480
rect 21880 -6500 22120 -6480
rect 22380 -6500 22620 -6480
rect 22880 -6500 23120 -6480
rect 23380 -6500 23620 -6480
rect 23880 -6500 24000 -6480
rect 14500 -6700 24000 -6500
rect 14500 -6720 14620 -6700
rect 14880 -6720 15120 -6700
rect 15380 -6720 15620 -6700
rect 15880 -6720 16120 -6700
rect 16380 -6720 16620 -6700
rect 16880 -6720 17120 -6700
rect 17380 -6720 17620 -6700
rect 17880 -6720 18120 -6700
rect 18380 -6720 18620 -6700
rect 18880 -6720 19120 -6700
rect 19380 -6720 19620 -6700
rect 19880 -6720 20120 -6700
rect 20380 -6720 20620 -6700
rect 20880 -6720 21120 -6700
rect 21380 -6720 21620 -6700
rect 21880 -6720 22120 -6700
rect 22380 -6720 22620 -6700
rect 22880 -6720 23120 -6700
rect 23380 -6720 23620 -6700
rect 23880 -6720 24000 -6700
rect 14500 -6980 14600 -6720
rect 14900 -6980 15100 -6720
rect 15400 -6980 15600 -6720
rect 15900 -6980 16100 -6720
rect 16400 -6980 16600 -6720
rect 16900 -6980 17100 -6720
rect 17400 -6980 17600 -6720
rect 17900 -6980 18100 -6720
rect 18400 -6980 18600 -6720
rect 18900 -6980 19100 -6720
rect 19400 -6980 19600 -6720
rect 19900 -6980 20100 -6720
rect 20400 -6980 20600 -6720
rect 20900 -6980 21100 -6720
rect 21400 -6980 21600 -6720
rect 21900 -6980 22100 -6720
rect 22400 -6980 22600 -6720
rect 22900 -6980 23100 -6720
rect 23400 -6980 23600 -6720
rect 23900 -6980 24000 -6720
rect 14500 -7000 14620 -6980
rect 14880 -7000 15120 -6980
rect 15380 -7000 15620 -6980
rect 15880 -7000 16120 -6980
rect 16380 -7000 16620 -6980
rect 16880 -7000 17120 -6980
rect 17380 -7000 17620 -6980
rect 17880 -7000 18120 -6980
rect 18380 -7000 18620 -6980
rect 18880 -7000 19120 -6980
rect 19380 -7000 19620 -6980
rect 19880 -7000 20120 -6980
rect 20380 -7000 20620 -6980
rect 20880 -7000 21120 -6980
rect 21380 -7000 21620 -6980
rect 21880 -7000 22120 -6980
rect 22380 -7000 22620 -6980
rect 22880 -7000 23120 -6980
rect 23380 -7000 23620 -6980
rect 23880 -7000 24000 -6980
rect 14500 -7200 24000 -7000
rect 14500 -7220 14620 -7200
rect 14880 -7220 15120 -7200
rect 15380 -7220 15620 -7200
rect 15880 -7220 16120 -7200
rect 16380 -7220 16620 -7200
rect 16880 -7220 17120 -7200
rect 17380 -7220 17620 -7200
rect 17880 -7220 18120 -7200
rect 18380 -7220 18620 -7200
rect 18880 -7220 19120 -7200
rect 19380 -7220 19620 -7200
rect 19880 -7220 20120 -7200
rect 20380 -7220 20620 -7200
rect 20880 -7220 21120 -7200
rect 21380 -7220 21620 -7200
rect 21880 -7220 22120 -7200
rect 22380 -7220 22620 -7200
rect 22880 -7220 23120 -7200
rect 23380 -7220 23620 -7200
rect 23880 -7220 24000 -7200
rect 14500 -7480 14600 -7220
rect 14900 -7480 15100 -7220
rect 15400 -7480 15600 -7220
rect 15900 -7480 16100 -7220
rect 16400 -7480 16600 -7220
rect 16900 -7480 17100 -7220
rect 17400 -7480 17600 -7220
rect 17900 -7480 18100 -7220
rect 18400 -7480 18600 -7220
rect 18900 -7480 19100 -7220
rect 19400 -7480 19600 -7220
rect 19900 -7480 20100 -7220
rect 20400 -7480 20600 -7220
rect 20900 -7480 21100 -7220
rect 21400 -7480 21600 -7220
rect 21900 -7480 22100 -7220
rect 22400 -7480 22600 -7220
rect 22900 -7480 23100 -7220
rect 23400 -7480 23600 -7220
rect 23900 -7480 24000 -7220
rect 14500 -7500 14620 -7480
rect 14880 -7500 15120 -7480
rect 15380 -7500 15620 -7480
rect 15880 -7500 16120 -7480
rect 16380 -7500 16620 -7480
rect 16880 -7500 17120 -7480
rect 17380 -7500 17620 -7480
rect 17880 -7500 18120 -7480
rect 18380 -7500 18620 -7480
rect 18880 -7500 19120 -7480
rect 19380 -7500 19620 -7480
rect 19880 -7500 20120 -7480
rect 20380 -7500 20620 -7480
rect 20880 -7500 21120 -7480
rect 21380 -7500 21620 -7480
rect 21880 -7500 22120 -7480
rect 22380 -7500 22620 -7480
rect 22880 -7500 23120 -7480
rect 23380 -7500 23620 -7480
rect 23880 -7500 24000 -7480
rect 14500 -7700 24000 -7500
rect 14500 -7720 14620 -7700
rect 14880 -7720 15120 -7700
rect 15380 -7720 15620 -7700
rect 15880 -7720 16120 -7700
rect 16380 -7720 16620 -7700
rect 16880 -7720 17120 -7700
rect 17380 -7720 17620 -7700
rect 17880 -7720 18120 -7700
rect 18380 -7720 18620 -7700
rect 18880 -7720 19120 -7700
rect 19380 -7720 19620 -7700
rect 19880 -7720 20120 -7700
rect 20380 -7720 20620 -7700
rect 20880 -7720 21120 -7700
rect 21380 -7720 21620 -7700
rect 21880 -7720 22120 -7700
rect 22380 -7720 22620 -7700
rect 22880 -7720 23120 -7700
rect 23380 -7720 23620 -7700
rect 23880 -7720 24000 -7700
rect 14500 -7980 14600 -7720
rect 14900 -7980 15100 -7720
rect 15400 -7980 15600 -7720
rect 15900 -7980 16100 -7720
rect 16400 -7980 16600 -7720
rect 16900 -7980 17100 -7720
rect 17400 -7980 17600 -7720
rect 17900 -7980 18100 -7720
rect 18400 -7980 18600 -7720
rect 18900 -7980 19100 -7720
rect 19400 -7980 19600 -7720
rect 19900 -7980 20100 -7720
rect 20400 -7980 20600 -7720
rect 20900 -7980 21100 -7720
rect 21400 -7980 21600 -7720
rect 21900 -7980 22100 -7720
rect 22400 -7980 22600 -7720
rect 22900 -7980 23100 -7720
rect 23400 -7980 23600 -7720
rect 23900 -7980 24000 -7720
rect 14500 -8000 14620 -7980
rect 14880 -8000 15120 -7980
rect 15380 -8000 15620 -7980
rect 15880 -8000 16120 -7980
rect 16380 -8000 16620 -7980
rect 16880 -8000 17120 -7980
rect 17380 -8000 17620 -7980
rect 17880 -8000 18120 -7980
rect 18380 -8000 18620 -7980
rect 18880 -8000 19120 -7980
rect 19380 -8000 19620 -7980
rect 19880 -8000 20120 -7980
rect 20380 -8000 20620 -7980
rect 20880 -8000 21120 -7980
rect 21380 -8000 21620 -7980
rect 21880 -8000 22120 -7980
rect 22380 -8000 22620 -7980
rect 22880 -8000 23120 -7980
rect 23380 -8000 23620 -7980
rect 23880 -8000 24000 -7980
rect 14500 -8200 24000 -8000
rect 14500 -8220 14620 -8200
rect 14880 -8220 15120 -8200
rect 15380 -8220 15620 -8200
rect 15880 -8220 16120 -8200
rect 16380 -8220 16620 -8200
rect 16880 -8220 17120 -8200
rect 17380 -8220 17620 -8200
rect 17880 -8220 18120 -8200
rect 18380 -8220 18620 -8200
rect 18880 -8220 19120 -8200
rect 19380 -8220 19620 -8200
rect 19880 -8220 20120 -8200
rect 20380 -8220 20620 -8200
rect 20880 -8220 21120 -8200
rect 21380 -8220 21620 -8200
rect 21880 -8220 22120 -8200
rect 22380 -8220 22620 -8200
rect 22880 -8220 23120 -8200
rect 23380 -8220 23620 -8200
rect 23880 -8220 24000 -8200
rect 14500 -8480 14600 -8220
rect 14900 -8480 15100 -8220
rect 15400 -8480 15600 -8220
rect 15900 -8480 16100 -8220
rect 16400 -8480 16600 -8220
rect 16900 -8480 17100 -8220
rect 17400 -8480 17600 -8220
rect 17900 -8480 18100 -8220
rect 18400 -8480 18600 -8220
rect 18900 -8480 19100 -8220
rect 19400 -8480 19600 -8220
rect 19900 -8480 20100 -8220
rect 20400 -8480 20600 -8220
rect 20900 -8480 21100 -8220
rect 21400 -8480 21600 -8220
rect 21900 -8480 22100 -8220
rect 22400 -8480 22600 -8220
rect 22900 -8480 23100 -8220
rect 23400 -8480 23600 -8220
rect 23900 -8480 24000 -8220
rect 14500 -8500 14620 -8480
rect 14880 -8500 15120 -8480
rect 15380 -8500 15620 -8480
rect 15880 -8500 16120 -8480
rect 16380 -8500 16620 -8480
rect 16880 -8500 17120 -8480
rect 17380 -8500 17620 -8480
rect 17880 -8500 18120 -8480
rect 18380 -8500 18620 -8480
rect 18880 -8500 19120 -8480
rect 19380 -8500 19620 -8480
rect 19880 -8500 20120 -8480
rect 20380 -8500 20620 -8480
rect 20880 -8500 21120 -8480
rect 21380 -8500 21620 -8480
rect 21880 -8500 22120 -8480
rect 22380 -8500 22620 -8480
rect 22880 -8500 23120 -8480
rect 23380 -8500 23620 -8480
rect 23880 -8500 24000 -8480
rect 14500 -8600 24000 -8500
rect 14500 -8700 17000 -8600
rect 14500 -8720 14620 -8700
rect 14880 -8720 15120 -8700
rect 15380 -8720 15620 -8700
rect 15880 -8720 16120 -8700
rect 16380 -8720 16620 -8700
rect 16880 -8720 17000 -8700
rect 14500 -8980 14600 -8720
rect 14900 -8980 15100 -8720
rect 15400 -8980 15600 -8720
rect 15900 -8980 16100 -8720
rect 16400 -8980 16600 -8720
rect 16900 -8980 17000 -8720
rect 14500 -9000 14620 -8980
rect 14880 -9000 15120 -8980
rect 15380 -9000 15620 -8980
rect 15880 -9000 16120 -8980
rect 16380 -9000 16620 -8980
rect 16880 -9000 17000 -8980
rect 14500 -9200 17000 -9000
rect 14500 -9220 14620 -9200
rect 14880 -9220 15120 -9200
rect 15380 -9220 15620 -9200
rect 15880 -9220 16120 -9200
rect 16380 -9220 16620 -9200
rect 16880 -9220 17000 -9200
rect 14500 -9480 14600 -9220
rect 14900 -9480 15100 -9220
rect 15400 -9480 15600 -9220
rect 15900 -9480 16100 -9220
rect 16400 -9480 16600 -9220
rect 16900 -9480 17000 -9220
rect 14500 -9500 14620 -9480
rect 14880 -9500 15120 -9480
rect 15380 -9500 15620 -9480
rect 15880 -9500 16120 -9480
rect 16380 -9500 16620 -9480
rect 16880 -9500 17000 -9480
rect 14500 -9700 17000 -9500
rect 14500 -9720 14620 -9700
rect 14880 -9720 15120 -9700
rect 15380 -9720 15620 -9700
rect 15880 -9720 16120 -9700
rect 16380 -9720 16620 -9700
rect 16880 -9720 17000 -9700
rect 14500 -9980 14600 -9720
rect 14900 -9980 15100 -9720
rect 15400 -9980 15600 -9720
rect 15900 -9980 16100 -9720
rect 16400 -9980 16600 -9720
rect 16900 -9980 17000 -9720
rect 14500 -10000 14620 -9980
rect 14880 -10000 15120 -9980
rect 15380 -10000 15620 -9980
rect 15880 -10000 16120 -9980
rect 16380 -10000 16620 -9980
rect 16880 -10000 17000 -9980
rect 14500 -10200 17000 -10000
rect 14500 -10220 14620 -10200
rect 14880 -10220 15120 -10200
rect 15380 -10220 15620 -10200
rect 15880 -10220 16120 -10200
rect 16380 -10220 16620 -10200
rect 16880 -10220 17000 -10200
rect 14500 -10480 14600 -10220
rect 14900 -10480 15100 -10220
rect 15400 -10480 15600 -10220
rect 15900 -10480 16100 -10220
rect 16400 -10480 16600 -10220
rect 16900 -10480 17000 -10220
rect 14500 -10500 14620 -10480
rect 14880 -10500 15120 -10480
rect 15380 -10500 15620 -10480
rect 15880 -10500 16120 -10480
rect 16380 -10500 16620 -10480
rect 16880 -10500 17000 -10480
rect 14500 -10700 17000 -10500
rect 14500 -10720 14620 -10700
rect 14880 -10720 15120 -10700
rect 15380 -10720 15620 -10700
rect 15880 -10720 16120 -10700
rect 16380 -10720 16620 -10700
rect 16880 -10720 17000 -10700
rect 14500 -10980 14600 -10720
rect 14900 -10980 15100 -10720
rect 15400 -10980 15600 -10720
rect 15900 -10980 16100 -10720
rect 16400 -10980 16600 -10720
rect 16900 -10980 17000 -10720
rect 14500 -11000 14620 -10980
rect 14880 -11000 15120 -10980
rect 15380 -11000 15620 -10980
rect 15880 -11000 16120 -10980
rect 16380 -11000 16620 -10980
rect 16880 -11000 17000 -10980
rect 14500 -11200 17000 -11000
rect 14500 -11220 14620 -11200
rect 14880 -11220 15120 -11200
rect 15380 -11220 15620 -11200
rect 15880 -11220 16120 -11200
rect 16380 -11220 16620 -11200
rect 16880 -11220 17000 -11200
rect 14500 -11480 14600 -11220
rect 14900 -11480 15100 -11220
rect 15400 -11480 15600 -11220
rect 15900 -11480 16100 -11220
rect 16400 -11480 16600 -11220
rect 16900 -11480 17000 -11220
rect 14500 -11500 14620 -11480
rect 14880 -11500 15120 -11480
rect 15380 -11500 15620 -11480
rect 15880 -11500 16120 -11480
rect 16380 -11500 16620 -11480
rect 16880 -11500 17000 -11480
rect 14500 -11700 17000 -11500
rect 14500 -11720 14620 -11700
rect 14880 -11720 15120 -11700
rect 15380 -11720 15620 -11700
rect 15880 -11720 16120 -11700
rect 16380 -11720 16620 -11700
rect 16880 -11720 17000 -11700
rect 14500 -11980 14600 -11720
rect 14900 -11980 15100 -11720
rect 15400 -11980 15600 -11720
rect 15900 -11980 16100 -11720
rect 16400 -11980 16600 -11720
rect 16900 -11980 17000 -11720
rect 14500 -12000 14620 -11980
rect 14880 -12000 15120 -11980
rect 15380 -12000 15620 -11980
rect 15880 -12000 16120 -11980
rect 16380 -12000 16620 -11980
rect 16880 -12000 17000 -11980
rect 14500 -12200 17000 -12000
rect 14500 -12220 14620 -12200
rect 14880 -12220 15120 -12200
rect 15380 -12220 15620 -12200
rect 15880 -12220 16120 -12200
rect 16380 -12220 16620 -12200
rect 16880 -12220 17000 -12200
rect 14500 -12480 14600 -12220
rect 14900 -12480 15100 -12220
rect 15400 -12480 15600 -12220
rect 15900 -12480 16100 -12220
rect 16400 -12480 16600 -12220
rect 16900 -12480 17000 -12220
rect 14500 -12500 14620 -12480
rect 14880 -12500 15120 -12480
rect 15380 -12500 15620 -12480
rect 15880 -12500 16120 -12480
rect 16380 -12500 16620 -12480
rect 16880 -12500 17000 -12480
rect 14500 -12700 17000 -12500
rect 14500 -12720 14620 -12700
rect 14880 -12720 15120 -12700
rect 15380 -12720 15620 -12700
rect 15880 -12720 16120 -12700
rect 16380 -12720 16620 -12700
rect 16880 -12720 17000 -12700
rect 14500 -12980 14600 -12720
rect 14900 -12980 15100 -12720
rect 15400 -12980 15600 -12720
rect 15900 -12980 16100 -12720
rect 16400 -12980 16600 -12720
rect 16900 -12980 17000 -12720
rect 14500 -13000 14620 -12980
rect 14880 -13000 15120 -12980
rect 15380 -13000 15620 -12980
rect 15880 -13000 16120 -12980
rect 16380 -13000 16620 -12980
rect 16880 -13000 17000 -12980
rect 14500 -13100 17000 -13000
rect 23500 -8700 24000 -8600
rect 23500 -8720 23620 -8700
rect 23880 -8720 24000 -8700
rect 23500 -8980 23600 -8720
rect 23900 -8980 24000 -8720
rect 23500 -9000 23620 -8980
rect 23880 -9000 24000 -8980
rect 23500 -9200 24000 -9000
rect 23500 -9220 23620 -9200
rect 23880 -9220 24000 -9200
rect 23500 -9480 23600 -9220
rect 23900 -9480 24000 -9220
rect 23500 -9500 23620 -9480
rect 23880 -9500 24000 -9480
rect 23500 -9700 24000 -9500
rect 23500 -9720 23620 -9700
rect 23880 -9720 24000 -9700
rect 23500 -9980 23600 -9720
rect 23900 -9980 24000 -9720
rect 23500 -10000 23620 -9980
rect 23880 -10000 24000 -9980
rect 23500 -10200 24000 -10000
rect 23500 -10220 23620 -10200
rect 23880 -10220 24000 -10200
rect 23500 -10480 23600 -10220
rect 23900 -10480 24000 -10220
rect 23500 -10500 23620 -10480
rect 23880 -10500 24000 -10480
rect 23500 -10700 24000 -10500
rect 23500 -10720 23620 -10700
rect 23880 -10720 24000 -10700
rect 23500 -10980 23600 -10720
rect 23900 -10980 24000 -10720
rect 23500 -11000 23620 -10980
rect 23880 -11000 24000 -10980
rect 23500 -11200 24000 -11000
rect 23500 -11220 23620 -11200
rect 23880 -11220 24000 -11200
rect 23500 -11480 23600 -11220
rect 23900 -11480 24000 -11220
rect 23500 -11500 23620 -11480
rect 23880 -11500 24000 -11480
rect 23500 -11700 24000 -11500
rect 23500 -11720 23620 -11700
rect 23880 -11720 24000 -11700
rect 23500 -11980 23600 -11720
rect 23900 -11980 24000 -11720
rect 23500 -12000 23620 -11980
rect 23880 -12000 24000 -11980
rect 23500 -12200 24000 -12000
rect 23500 -12220 23620 -12200
rect 23880 -12220 24000 -12200
rect 23500 -12480 23600 -12220
rect 23900 -12480 24000 -12220
rect 23500 -12500 23620 -12480
rect 23880 -12500 24000 -12480
rect 23500 -12700 24000 -12500
rect 23500 -12720 23620 -12700
rect 23880 -12720 24000 -12700
rect 23500 -12980 23600 -12720
rect 23900 -12980 24000 -12720
rect 23500 -13000 23620 -12980
rect 23880 -13000 24000 -12980
rect -27500 -13220 -27380 -13200
rect -27120 -13220 -26880 -13200
rect -26620 -13220 -26380 -13200
rect -26120 -13220 -25880 -13200
rect -25620 -13220 -25380 -13200
rect -25120 -13220 -24880 -13200
rect -24620 -13220 -24380 -13200
rect -24120 -13220 -23880 -13200
rect -23620 -13220 -23380 -13200
rect -23120 -13220 -22880 -13200
rect -22620 -13220 -22380 -13200
rect -22120 -13220 -21880 -13200
rect -21620 -13220 -21380 -13200
rect -21120 -13220 -20880 -13200
rect -20620 -13220 -20380 -13200
rect -20120 -13220 -19880 -13200
rect -19620 -13220 -19380 -13200
rect -19120 -13220 -18880 -13200
rect -18620 -13220 -18380 -13200
rect -18120 -13220 -17880 -13200
rect -17620 -13220 -17380 -13200
rect -17120 -13220 -16880 -13200
rect -16620 -13220 -16380 -13200
rect -16120 -13220 -15880 -13200
rect -15620 -13220 -15380 -13200
rect -15120 -13220 -15000 -13200
rect -27500 -13480 -27400 -13220
rect -27100 -13480 -26900 -13220
rect -26600 -13480 -26400 -13220
rect -26100 -13480 -25900 -13220
rect -25600 -13480 -25400 -13220
rect -25100 -13480 -24900 -13220
rect -24600 -13480 -24400 -13220
rect -24100 -13480 -23900 -13220
rect -23600 -13480 -23400 -13220
rect -23100 -13480 -22900 -13220
rect -22600 -13480 -22400 -13220
rect -22100 -13480 -21900 -13220
rect -21600 -13480 -21400 -13220
rect -21100 -13480 -20900 -13220
rect -20600 -13480 -20400 -13220
rect -20100 -13480 -19900 -13220
rect -19600 -13480 -19400 -13220
rect -19100 -13480 -18900 -13220
rect -18600 -13480 -18400 -13220
rect -18100 -13480 -17900 -13220
rect -17600 -13480 -17400 -13220
rect -17100 -13480 -16900 -13220
rect -16600 -13480 -16400 -13220
rect -16100 -13480 -15900 -13220
rect -15600 -13480 -15400 -13220
rect -15100 -13480 -15000 -13220
rect -27500 -13500 -27380 -13480
rect -27120 -13500 -26880 -13480
rect -26620 -13500 -26380 -13480
rect -26120 -13500 -25880 -13480
rect -25620 -13500 -25380 -13480
rect -25120 -13500 -24880 -13480
rect -24620 -13500 -24380 -13480
rect -24120 -13500 -23880 -13480
rect -23620 -13500 -23380 -13480
rect -23120 -13500 -22880 -13480
rect -22620 -13500 -22380 -13480
rect -22120 -13500 -21880 -13480
rect -21620 -13500 -21380 -13480
rect -21120 -13500 -20880 -13480
rect -20620 -13500 -20380 -13480
rect -20120 -13500 -19880 -13480
rect -19620 -13500 -19380 -13480
rect -19120 -13500 -18880 -13480
rect -18620 -13500 -18380 -13480
rect -18120 -13500 -17880 -13480
rect -17620 -13500 -17380 -13480
rect -17120 -13500 -16880 -13480
rect -16620 -13500 -16380 -13480
rect -16120 -13500 -15880 -13480
rect -15620 -13500 -15380 -13480
rect -15120 -13500 -15000 -13480
rect -27500 -13600 -15000 -13500
rect -29500 -13700 -15000 -13600
rect -29500 -13720 -29380 -13700
rect -29120 -13720 -28880 -13700
rect -28620 -13720 -28380 -13700
rect -28120 -13720 -27880 -13700
rect -27620 -13720 -27380 -13700
rect -27120 -13720 -26880 -13700
rect -26620 -13720 -26380 -13700
rect -26120 -13720 -25880 -13700
rect -25620 -13720 -25380 -13700
rect -25120 -13720 -24880 -13700
rect -24620 -13720 -24380 -13700
rect -24120 -13720 -23880 -13700
rect -23620 -13720 -23380 -13700
rect -23120 -13720 -22880 -13700
rect -22620 -13720 -22380 -13700
rect -22120 -13720 -21880 -13700
rect -21620 -13720 -21380 -13700
rect -21120 -13720 -20880 -13700
rect -20620 -13720 -20380 -13700
rect -20120 -13720 -19880 -13700
rect -19620 -13720 -19380 -13700
rect -19120 -13720 -18880 -13700
rect -18620 -13720 -18380 -13700
rect -18120 -13720 -17880 -13700
rect -17620 -13720 -17380 -13700
rect -17120 -13720 -16880 -13700
rect -16620 -13720 -16380 -13700
rect -16120 -13720 -15880 -13700
rect -15620 -13720 -15380 -13700
rect -15120 -13720 -15000 -13700
rect -29500 -13980 -29400 -13720
rect -29100 -13980 -28900 -13720
rect -28600 -13980 -28400 -13720
rect -28100 -13980 -27900 -13720
rect -27600 -13980 -27400 -13720
rect -27100 -13980 -26900 -13720
rect -26600 -13980 -26400 -13720
rect -26100 -13980 -25900 -13720
rect -25600 -13980 -25400 -13720
rect -25100 -13980 -24900 -13720
rect -24600 -13980 -24400 -13720
rect -24100 -13980 -23900 -13720
rect -23600 -13980 -23400 -13720
rect -23100 -13980 -22900 -13720
rect -22600 -13980 -22400 -13720
rect -22100 -13980 -21900 -13720
rect -21600 -13980 -21400 -13720
rect -21100 -13980 -20900 -13720
rect -20600 -13980 -20400 -13720
rect -20100 -13980 -19900 -13720
rect -19600 -13980 -19400 -13720
rect -19100 -13980 -18900 -13720
rect -18600 -13980 -18400 -13720
rect -18100 -13980 -17900 -13720
rect -17600 -13980 -17400 -13720
rect -17100 -13980 -16900 -13720
rect -16600 -13980 -16400 -13720
rect -16100 -13980 -15900 -13720
rect -15600 -13980 -15400 -13720
rect -15100 -13980 -15000 -13720
rect -29500 -14000 -29380 -13980
rect -29120 -14000 -28880 -13980
rect -28620 -14000 -28380 -13980
rect -28120 -14000 -27880 -13980
rect -27620 -14000 -27380 -13980
rect -27120 -14000 -26880 -13980
rect -26620 -14000 -26380 -13980
rect -26120 -14000 -25880 -13980
rect -25620 -14000 -25380 -13980
rect -25120 -14000 -24880 -13980
rect -24620 -14000 -24380 -13980
rect -24120 -14000 -23880 -13980
rect -23620 -14000 -23380 -13980
rect -23120 -14000 -22880 -13980
rect -22620 -14000 -22380 -13980
rect -22120 -14000 -21880 -13980
rect -21620 -14000 -21380 -13980
rect -21120 -14000 -20880 -13980
rect -20620 -14000 -20380 -13980
rect -20120 -14000 -19880 -13980
rect -19620 -14000 -19380 -13980
rect -19120 -14000 -18880 -13980
rect -18620 -14000 -18380 -13980
rect -18120 -14000 -17880 -13980
rect -17620 -14000 -17380 -13980
rect -17120 -14000 -16880 -13980
rect -16620 -14000 -16380 -13980
rect -16120 -14000 -15880 -13980
rect -15620 -14000 -15380 -13980
rect -15120 -14000 -15000 -13980
rect -29500 -14200 -15000 -14000
rect -29500 -14220 -29380 -14200
rect -29120 -14220 -28880 -14200
rect -28620 -14220 -28380 -14200
rect -28120 -14220 -27880 -14200
rect -27620 -14220 -27380 -14200
rect -27120 -14220 -26880 -14200
rect -26620 -14220 -26380 -14200
rect -26120 -14220 -25880 -14200
rect -25620 -14220 -25380 -14200
rect -25120 -14220 -24880 -14200
rect -24620 -14220 -24380 -14200
rect -24120 -14220 -23880 -14200
rect -23620 -14220 -23380 -14200
rect -23120 -14220 -22880 -14200
rect -22620 -14220 -22380 -14200
rect -22120 -14220 -21880 -14200
rect -21620 -14220 -21380 -14200
rect -21120 -14220 -20880 -14200
rect -20620 -14220 -20380 -14200
rect -20120 -14220 -19880 -14200
rect -19620 -14220 -19380 -14200
rect -19120 -14220 -18880 -14200
rect -18620 -14220 -18380 -14200
rect -18120 -14220 -17880 -14200
rect -17620 -14220 -17380 -14200
rect -17120 -14220 -16880 -14200
rect -16620 -14220 -16380 -14200
rect -16120 -14220 -15880 -14200
rect -15620 -14220 -15380 -14200
rect -15120 -14220 -15000 -14200
rect -29500 -14480 -29400 -14220
rect -29100 -14480 -28900 -14220
rect -28600 -14480 -28400 -14220
rect -28100 -14480 -27900 -14220
rect -27600 -14480 -27400 -14220
rect -27100 -14480 -26900 -14220
rect -26600 -14480 -26400 -14220
rect -26100 -14480 -25900 -14220
rect -25600 -14480 -25400 -14220
rect -25100 -14480 -24900 -14220
rect -24600 -14480 -24400 -14220
rect -24100 -14480 -23900 -14220
rect -23600 -14480 -23400 -14220
rect -23100 -14480 -22900 -14220
rect -22600 -14480 -22400 -14220
rect -22100 -14480 -21900 -14220
rect -21600 -14480 -21400 -14220
rect -21100 -14480 -20900 -14220
rect -20600 -14480 -20400 -14220
rect -20100 -14480 -19900 -14220
rect -19600 -14480 -19400 -14220
rect -19100 -14480 -18900 -14220
rect -18600 -14480 -18400 -14220
rect -18100 -14480 -17900 -14220
rect -17600 -14480 -17400 -14220
rect -17100 -14480 -16900 -14220
rect -16600 -14480 -16400 -14220
rect -16100 -14480 -15900 -14220
rect -15600 -14480 -15400 -14220
rect -15100 -14480 -15000 -14220
rect -29500 -14500 -29380 -14480
rect -29120 -14500 -28880 -14480
rect -28620 -14500 -28380 -14480
rect -28120 -14500 -27880 -14480
rect -27620 -14500 -27380 -14480
rect -27120 -14500 -26880 -14480
rect -26620 -14500 -26380 -14480
rect -26120 -14500 -25880 -14480
rect -25620 -14500 -25380 -14480
rect -25120 -14500 -24880 -14480
rect -24620 -14500 -24380 -14480
rect -24120 -14500 -23880 -14480
rect -23620 -14500 -23380 -14480
rect -23120 -14500 -22880 -14480
rect -22620 -14500 -22380 -14480
rect -22120 -14500 -21880 -14480
rect -21620 -14500 -21380 -14480
rect -21120 -14500 -20880 -14480
rect -20620 -14500 -20380 -14480
rect -20120 -14500 -19880 -14480
rect -19620 -14500 -19380 -14480
rect -19120 -14500 -18880 -14480
rect -18620 -14500 -18380 -14480
rect -18120 -14500 -17880 -14480
rect -17620 -14500 -17380 -14480
rect -17120 -14500 -16880 -14480
rect -16620 -14500 -16380 -14480
rect -16120 -14500 -15880 -14480
rect -15620 -14500 -15380 -14480
rect -15120 -14500 -15000 -14480
rect -29500 -14700 -15000 -14500
rect -29500 -14720 -29380 -14700
rect -29120 -14720 -28880 -14700
rect -28620 -14720 -28380 -14700
rect -28120 -14720 -27880 -14700
rect -27620 -14720 -27380 -14700
rect -27120 -14720 -26880 -14700
rect -26620 -14720 -26380 -14700
rect -26120 -14720 -25880 -14700
rect -25620 -14720 -25380 -14700
rect -25120 -14720 -24880 -14700
rect -24620 -14720 -24380 -14700
rect -24120 -14720 -23880 -14700
rect -23620 -14720 -23380 -14700
rect -23120 -14720 -22880 -14700
rect -22620 -14720 -22380 -14700
rect -22120 -14720 -21880 -14700
rect -21620 -14720 -21380 -14700
rect -21120 -14720 -20880 -14700
rect -20620 -14720 -20380 -14700
rect -20120 -14720 -19880 -14700
rect -19620 -14720 -19380 -14700
rect -19120 -14720 -18880 -14700
rect -18620 -14720 -18380 -14700
rect -18120 -14720 -17880 -14700
rect -17620 -14720 -17380 -14700
rect -17120 -14720 -16880 -14700
rect -16620 -14720 -16380 -14700
rect -16120 -14720 -15880 -14700
rect -15620 -14720 -15380 -14700
rect -15120 -14720 -15000 -14700
rect -29500 -14980 -29400 -14720
rect -29100 -14980 -28900 -14720
rect -28600 -14980 -28400 -14720
rect -28100 -14980 -27900 -14720
rect -27600 -14980 -27400 -14720
rect -27100 -14980 -26900 -14720
rect -26600 -14980 -26400 -14720
rect -26100 -14980 -25900 -14720
rect -25600 -14980 -25400 -14720
rect -25100 -14980 -24900 -14720
rect -24600 -14980 -24400 -14720
rect -24100 -14980 -23900 -14720
rect -23600 -14980 -23400 -14720
rect -23100 -14980 -22900 -14720
rect -22600 -14980 -22400 -14720
rect -22100 -14980 -21900 -14720
rect -21600 -14980 -21400 -14720
rect -21100 -14980 -20900 -14720
rect -20600 -14980 -20400 -14720
rect -20100 -14980 -19900 -14720
rect -19600 -14980 -19400 -14720
rect -19100 -14980 -18900 -14720
rect -18600 -14980 -18400 -14720
rect -18100 -14980 -17900 -14720
rect -17600 -14980 -17400 -14720
rect -17100 -14980 -16900 -14720
rect -16600 -14980 -16400 -14720
rect -16100 -14980 -15900 -14720
rect -15600 -14980 -15400 -14720
rect -15100 -14980 -15000 -14720
rect -29500 -15000 -29380 -14980
rect -29120 -15000 -28880 -14980
rect -28620 -15000 -28380 -14980
rect -28120 -15000 -27880 -14980
rect -27620 -15000 -27380 -14980
rect -27120 -15000 -26880 -14980
rect -26620 -15000 -26380 -14980
rect -26120 -15000 -25880 -14980
rect -25620 -15000 -25380 -14980
rect -25120 -15000 -24880 -14980
rect -24620 -15000 -24380 -14980
rect -24120 -15000 -23880 -14980
rect -23620 -15000 -23380 -14980
rect -23120 -15000 -22880 -14980
rect -22620 -15000 -22380 -14980
rect -22120 -15000 -21880 -14980
rect -21620 -15000 -21380 -14980
rect -21120 -15000 -20880 -14980
rect -20620 -15000 -20380 -14980
rect -20120 -15000 -19880 -14980
rect -19620 -15000 -19380 -14980
rect -19120 -15000 -18880 -14980
rect -18620 -15000 -18380 -14980
rect -18120 -15000 -17880 -14980
rect -17620 -15000 -17380 -14980
rect -17120 -15000 -16880 -14980
rect -16620 -15000 -16380 -14980
rect -16120 -15000 -15880 -14980
rect -15620 -15000 -15380 -14980
rect -15120 -15000 -15000 -14980
rect -29500 -15200 -15000 -15000
rect -29500 -15220 -29380 -15200
rect -29120 -15220 -28880 -15200
rect -28620 -15220 -28380 -15200
rect -28120 -15220 -27880 -15200
rect -27620 -15220 -27380 -15200
rect -27120 -15220 -26880 -15200
rect -26620 -15220 -26380 -15200
rect -26120 -15220 -25880 -15200
rect -25620 -15220 -25380 -15200
rect -25120 -15220 -24880 -15200
rect -24620 -15220 -24380 -15200
rect -24120 -15220 -23880 -15200
rect -23620 -15220 -23380 -15200
rect -23120 -15220 -22880 -15200
rect -22620 -15220 -22380 -15200
rect -22120 -15220 -21880 -15200
rect -21620 -15220 -21380 -15200
rect -21120 -15220 -20880 -15200
rect -20620 -15220 -20380 -15200
rect -20120 -15220 -19880 -15200
rect -19620 -15220 -19380 -15200
rect -19120 -15220 -18880 -15200
rect -18620 -15220 -18380 -15200
rect -18120 -15220 -17880 -15200
rect -17620 -15220 -17380 -15200
rect -17120 -15220 -16880 -15200
rect -16620 -15220 -16380 -15200
rect -16120 -15220 -15880 -15200
rect -15620 -15220 -15380 -15200
rect -15120 -15220 -15000 -15200
rect -29500 -15480 -29400 -15220
rect -29100 -15480 -28900 -15220
rect -28600 -15480 -28400 -15220
rect -28100 -15480 -27900 -15220
rect -27600 -15480 -27400 -15220
rect -27100 -15480 -26900 -15220
rect -26600 -15480 -26400 -15220
rect -26100 -15480 -25900 -15220
rect -25600 -15480 -25400 -15220
rect -25100 -15480 -24900 -15220
rect -24600 -15480 -24400 -15220
rect -24100 -15480 -23900 -15220
rect -23600 -15480 -23400 -15220
rect -23100 -15480 -22900 -15220
rect -22600 -15480 -22400 -15220
rect -22100 -15480 -21900 -15220
rect -21600 -15480 -21400 -15220
rect -21100 -15480 -20900 -15220
rect -20600 -15480 -20400 -15220
rect -20100 -15480 -19900 -15220
rect -19600 -15480 -19400 -15220
rect -19100 -15480 -18900 -15220
rect -18600 -15480 -18400 -15220
rect -18100 -15480 -17900 -15220
rect -17600 -15480 -17400 -15220
rect -17100 -15480 -16900 -15220
rect -16600 -15480 -16400 -15220
rect -16100 -15480 -15900 -15220
rect -15600 -15480 -15400 -15220
rect -15100 -15480 -15000 -15220
rect -29500 -15500 -29380 -15480
rect -29120 -15500 -28880 -15480
rect -28620 -15500 -28380 -15480
rect -28120 -15500 -27880 -15480
rect -27620 -15500 -27380 -15480
rect -27120 -15500 -26880 -15480
rect -26620 -15500 -26380 -15480
rect -26120 -15500 -25880 -15480
rect -25620 -15500 -25380 -15480
rect -25120 -15500 -24880 -15480
rect -24620 -15500 -24380 -15480
rect -24120 -15500 -23880 -15480
rect -23620 -15500 -23380 -15480
rect -23120 -15500 -22880 -15480
rect -22620 -15500 -22380 -15480
rect -22120 -15500 -21880 -15480
rect -21620 -15500 -21380 -15480
rect -21120 -15500 -20880 -15480
rect -20620 -15500 -20380 -15480
rect -20120 -15500 -19880 -15480
rect -19620 -15500 -19380 -15480
rect -19120 -15500 -18880 -15480
rect -18620 -15500 -18380 -15480
rect -18120 -15500 -17880 -15480
rect -17620 -15500 -17380 -15480
rect -17120 -15500 -16880 -15480
rect -16620 -15500 -16380 -15480
rect -16120 -15500 -15880 -15480
rect -15620 -15500 -15380 -15480
rect -15120 -15500 -15000 -15480
rect -29500 -15700 -15000 -15500
rect -29500 -15720 -29380 -15700
rect -29120 -15720 -28880 -15700
rect -28620 -15720 -28380 -15700
rect -28120 -15720 -27880 -15700
rect -27620 -15720 -27380 -15700
rect -27120 -15720 -26880 -15700
rect -26620 -15720 -26380 -15700
rect -26120 -15720 -25880 -15700
rect -25620 -15720 -25380 -15700
rect -25120 -15720 -24880 -15700
rect -24620 -15720 -24380 -15700
rect -24120 -15720 -23880 -15700
rect -23620 -15720 -23380 -15700
rect -23120 -15720 -22880 -15700
rect -22620 -15720 -22380 -15700
rect -22120 -15720 -21880 -15700
rect -21620 -15720 -21380 -15700
rect -21120 -15720 -20880 -15700
rect -20620 -15720 -20380 -15700
rect -20120 -15720 -19880 -15700
rect -19620 -15720 -19380 -15700
rect -19120 -15720 -18880 -15700
rect -18620 -15720 -18380 -15700
rect -18120 -15720 -17880 -15700
rect -17620 -15720 -17380 -15700
rect -17120 -15720 -16880 -15700
rect -16620 -15720 -16380 -15700
rect -16120 -15720 -15880 -15700
rect -15620 -15720 -15380 -15700
rect -15120 -15720 -15000 -15700
rect -29500 -15980 -29400 -15720
rect -29100 -15980 -28900 -15720
rect -28600 -15980 -28400 -15720
rect -28100 -15980 -27900 -15720
rect -27600 -15980 -27400 -15720
rect -27100 -15980 -26900 -15720
rect -26600 -15980 -26400 -15720
rect -26100 -15980 -25900 -15720
rect -25600 -15980 -25400 -15720
rect -25100 -15980 -24900 -15720
rect -24600 -15980 -24400 -15720
rect -24100 -15980 -23900 -15720
rect -23600 -15980 -23400 -15720
rect -23100 -15980 -22900 -15720
rect -22600 -15980 -22400 -15720
rect -22100 -15980 -21900 -15720
rect -21600 -15980 -21400 -15720
rect -21100 -15980 -20900 -15720
rect -20600 -15980 -20400 -15720
rect -20100 -15980 -19900 -15720
rect -19600 -15980 -19400 -15720
rect -19100 -15980 -18900 -15720
rect -18600 -15980 -18400 -15720
rect -18100 -15980 -17900 -15720
rect -17600 -15980 -17400 -15720
rect -17100 -15980 -16900 -15720
rect -16600 -15980 -16400 -15720
rect -16100 -15980 -15900 -15720
rect -15600 -15980 -15400 -15720
rect -15100 -15980 -15000 -15720
rect -29500 -16000 -29380 -15980
rect -29120 -16000 -28880 -15980
rect -28620 -16000 -28380 -15980
rect -28120 -16000 -27880 -15980
rect -27620 -16000 -27380 -15980
rect -27120 -16000 -26880 -15980
rect -26620 -16000 -26380 -15980
rect -26120 -16000 -25880 -15980
rect -25620 -16000 -25380 -15980
rect -25120 -16000 -24880 -15980
rect -24620 -16000 -24380 -15980
rect -24120 -16000 -23880 -15980
rect -23620 -16000 -23380 -15980
rect -23120 -16000 -22880 -15980
rect -22620 -16000 -22380 -15980
rect -22120 -16000 -21880 -15980
rect -21620 -16000 -21380 -15980
rect -21120 -16000 -20880 -15980
rect -20620 -16000 -20380 -15980
rect -20120 -16000 -19880 -15980
rect -19620 -16000 -19380 -15980
rect -19120 -16000 -18880 -15980
rect -18620 -16000 -18380 -15980
rect -18120 -16000 -17880 -15980
rect -17620 -16000 -17380 -15980
rect -17120 -16000 -16880 -15980
rect -16620 -16000 -16380 -15980
rect -16120 -16000 -15880 -15980
rect -15620 -16000 -15380 -15980
rect -15120 -16000 -15000 -15980
rect -29500 -16100 -15000 -16000
rect -31500 -16200 -15000 -16100
rect -31500 -16220 -31380 -16200
rect -31120 -16220 -30880 -16200
rect -30620 -16220 -30380 -16200
rect -30120 -16220 -29880 -16200
rect -29620 -16220 -29380 -16200
rect -29120 -16220 -28880 -16200
rect -28620 -16220 -28380 -16200
rect -28120 -16220 -27880 -16200
rect -27620 -16220 -27380 -16200
rect -27120 -16220 -26880 -16200
rect -26620 -16220 -26380 -16200
rect -26120 -16220 -25880 -16200
rect -25620 -16220 -25380 -16200
rect -25120 -16220 -24880 -16200
rect -24620 -16220 -24380 -16200
rect -24120 -16220 -23880 -16200
rect -23620 -16220 -23380 -16200
rect -23120 -16220 -22880 -16200
rect -22620 -16220 -22380 -16200
rect -22120 -16220 -21880 -16200
rect -21620 -16220 -21380 -16200
rect -21120 -16220 -20880 -16200
rect -20620 -16220 -20380 -16200
rect -20120 -16220 -19880 -16200
rect -19620 -16220 -19380 -16200
rect -19120 -16220 -18880 -16200
rect -18620 -16220 -18380 -16200
rect -18120 -16220 -17880 -16200
rect -17620 -16220 -17380 -16200
rect -17120 -16220 -16880 -16200
rect -16620 -16220 -16380 -16200
rect -16120 -16220 -15880 -16200
rect -15620 -16220 -15380 -16200
rect -15120 -16220 -15000 -16200
rect -31500 -16480 -31400 -16220
rect -31100 -16480 -30900 -16220
rect -30600 -16480 -30400 -16220
rect -30100 -16480 -29900 -16220
rect -29600 -16480 -29400 -16220
rect -29100 -16480 -28900 -16220
rect -28600 -16480 -28400 -16220
rect -28100 -16480 -27900 -16220
rect -27600 -16480 -27400 -16220
rect -27100 -16480 -26900 -16220
rect -26600 -16480 -26400 -16220
rect -26100 -16480 -25900 -16220
rect -25600 -16480 -25400 -16220
rect -25100 -16480 -24900 -16220
rect -24600 -16480 -24400 -16220
rect -24100 -16480 -23900 -16220
rect -23600 -16480 -23400 -16220
rect -23100 -16480 -22900 -16220
rect -22600 -16480 -22400 -16220
rect -22100 -16480 -21900 -16220
rect -21600 -16480 -21400 -16220
rect -21100 -16480 -20900 -16220
rect -20600 -16480 -20400 -16220
rect -20100 -16480 -19900 -16220
rect -19600 -16480 -19400 -16220
rect -19100 -16480 -18900 -16220
rect -18600 -16480 -18400 -16220
rect -18100 -16480 -17900 -16220
rect -17600 -16480 -17400 -16220
rect -17100 -16480 -16900 -16220
rect -16600 -16480 -16400 -16220
rect -16100 -16480 -15900 -16220
rect -15600 -16480 -15400 -16220
rect -15100 -16480 -15000 -16220
rect -31500 -16500 -31380 -16480
rect -31120 -16500 -30880 -16480
rect -30620 -16500 -30380 -16480
rect -30120 -16500 -29880 -16480
rect -29620 -16500 -29380 -16480
rect -29120 -16500 -28880 -16480
rect -28620 -16500 -28380 -16480
rect -28120 -16500 -27880 -16480
rect -27620 -16500 -27380 -16480
rect -27120 -16500 -26880 -16480
rect -26620 -16500 -26380 -16480
rect -26120 -16500 -25880 -16480
rect -25620 -16500 -25380 -16480
rect -25120 -16500 -24880 -16480
rect -24620 -16500 -24380 -16480
rect -24120 -16500 -23880 -16480
rect -23620 -16500 -23380 -16480
rect -23120 -16500 -22880 -16480
rect -22620 -16500 -22380 -16480
rect -22120 -16500 -21880 -16480
rect -21620 -16500 -21380 -16480
rect -21120 -16500 -20880 -16480
rect -20620 -16500 -20380 -16480
rect -20120 -16500 -19880 -16480
rect -19620 -16500 -19380 -16480
rect -19120 -16500 -18880 -16480
rect -18620 -16500 -18380 -16480
rect -18120 -16500 -17880 -16480
rect -17620 -16500 -17380 -16480
rect -17120 -16500 -16880 -16480
rect -16620 -16500 -16380 -16480
rect -16120 -16500 -15880 -16480
rect -15620 -16500 -15380 -16480
rect -15120 -16500 -15000 -16480
rect -31500 -16600 -15000 -16500
rect -31500 -16700 -23000 -16600
rect -31500 -16720 -31380 -16700
rect -31120 -16720 -30880 -16700
rect -30620 -16720 -30380 -16700
rect -30120 -16720 -29880 -16700
rect -29620 -16720 -29380 -16700
rect -29120 -16720 -28880 -16700
rect -28620 -16720 -28380 -16700
rect -28120 -16720 -27880 -16700
rect -27620 -16720 -27380 -16700
rect -27120 -16720 -26880 -16700
rect -26620 -16720 -26380 -16700
rect -26120 -16720 -25880 -16700
rect -25620 -16720 -25380 -16700
rect -25120 -16720 -24880 -16700
rect -24620 -16720 -24380 -16700
rect -24120 -16720 -23880 -16700
rect -23620 -16720 -23380 -16700
rect -23120 -16720 -23000 -16700
rect -31500 -16980 -31400 -16720
rect -31100 -16980 -30900 -16720
rect -30600 -16980 -30400 -16720
rect -30100 -16980 -29900 -16720
rect -29600 -16980 -29400 -16720
rect -29100 -16980 -28900 -16720
rect -28600 -16980 -28400 -16720
rect -28100 -16980 -27900 -16720
rect -27600 -16980 -27400 -16720
rect -27100 -16980 -26900 -16720
rect -26600 -16980 -26400 -16720
rect -26100 -16980 -25900 -16720
rect -25600 -16980 -25400 -16720
rect -25100 -16980 -24900 -16720
rect -24600 -16980 -24400 -16720
rect -24100 -16980 -23900 -16720
rect -23600 -16980 -23400 -16720
rect -23100 -16980 -23000 -16720
rect -31500 -17000 -31380 -16980
rect -31120 -17000 -30880 -16980
rect -30620 -17000 -30380 -16980
rect -30120 -17000 -29880 -16980
rect -29620 -17000 -29380 -16980
rect -29120 -17000 -28880 -16980
rect -28620 -17000 -28380 -16980
rect -28120 -17000 -27880 -16980
rect -27620 -17000 -27380 -16980
rect -27120 -17000 -26880 -16980
rect -26620 -17000 -26380 -16980
rect -26120 -17000 -25880 -16980
rect -25620 -17000 -25380 -16980
rect -25120 -17000 -24880 -16980
rect -24620 -17000 -24380 -16980
rect -24120 -17000 -23880 -16980
rect -23620 -17000 -23380 -16980
rect -23120 -17000 -23000 -16980
rect -31500 -17200 -23000 -17000
rect -31500 -17220 -31380 -17200
rect -31120 -17220 -30880 -17200
rect -30620 -17220 -30380 -17200
rect -30120 -17220 -29880 -17200
rect -29620 -17220 -29380 -17200
rect -29120 -17220 -28880 -17200
rect -28620 -17220 -28380 -17200
rect -28120 -17220 -27880 -17200
rect -27620 -17220 -27380 -17200
rect -27120 -17220 -26880 -17200
rect -26620 -17220 -26380 -17200
rect -26120 -17220 -25880 -17200
rect -25620 -17220 -25380 -17200
rect -25120 -17220 -24880 -17200
rect -24620 -17220 -24380 -17200
rect -24120 -17220 -23880 -17200
rect -23620 -17220 -23380 -17200
rect -23120 -17220 -23000 -17200
rect -31500 -17480 -31400 -17220
rect -31100 -17480 -30900 -17220
rect -30600 -17480 -30400 -17220
rect -30100 -17480 -29900 -17220
rect -29600 -17480 -29400 -17220
rect -29100 -17480 -28900 -17220
rect -28600 -17480 -28400 -17220
rect -28100 -17480 -27900 -17220
rect -27600 -17480 -27400 -17220
rect -27100 -17480 -26900 -17220
rect -26600 -17480 -26400 -17220
rect -26100 -17480 -25900 -17220
rect -25600 -17480 -25400 -17220
rect -25100 -17480 -24900 -17220
rect -24600 -17480 -24400 -17220
rect -24100 -17480 -23900 -17220
rect -23600 -17480 -23400 -17220
rect -23100 -17480 -23000 -17220
rect -31500 -17500 -31380 -17480
rect -31120 -17500 -30880 -17480
rect -30620 -17500 -30380 -17480
rect -30120 -17500 -29880 -17480
rect -29620 -17500 -29380 -17480
rect -29120 -17500 -28880 -17480
rect -28620 -17500 -28380 -17480
rect -28120 -17500 -27880 -17480
rect -27620 -17500 -27380 -17480
rect -27120 -17500 -26880 -17480
rect -26620 -17500 -26380 -17480
rect -26120 -17500 -25880 -17480
rect -25620 -17500 -25380 -17480
rect -25120 -17500 -24880 -17480
rect -24620 -17500 -24380 -17480
rect -24120 -17500 -23880 -17480
rect -23620 -17500 -23380 -17480
rect -23120 -17500 -23000 -17480
rect -31500 -17600 -23000 -17500
rect -31500 -17700 -27500 -17600
rect -31500 -17720 -31380 -17700
rect -31120 -17720 -30880 -17700
rect -30620 -17720 -30380 -17700
rect -30120 -17720 -29880 -17700
rect -29620 -17720 -29380 -17700
rect -29120 -17720 -28880 -17700
rect -28620 -17720 -28380 -17700
rect -28120 -17720 -27880 -17700
rect -27620 -17720 -27500 -17700
rect -31500 -17980 -31400 -17720
rect -31100 -17980 -30900 -17720
rect -30600 -17980 -30400 -17720
rect -30100 -17980 -29900 -17720
rect -29600 -17980 -29400 -17720
rect -29100 -17980 -28900 -17720
rect -28600 -17980 -28400 -17720
rect -28100 -17980 -27900 -17720
rect -27600 -17980 -27500 -17720
rect -31500 -18000 -31380 -17980
rect -31120 -18000 -30880 -17980
rect -30620 -18000 -30380 -17980
rect -30120 -18000 -29880 -17980
rect -29620 -18000 -29380 -17980
rect -29120 -18000 -28880 -17980
rect -28620 -18000 -28380 -17980
rect -28120 -18000 -27880 -17980
rect -27620 -18000 -27500 -17980
rect -31500 -18100 -27500 -18000
rect -26500 -17700 -23000 -17600
rect -26500 -17720 -26380 -17700
rect -26120 -17720 -25880 -17700
rect -25620 -17720 -25380 -17700
rect -25120 -17720 -24880 -17700
rect -24620 -17720 -24380 -17700
rect -24120 -17720 -23880 -17700
rect -23620 -17720 -23380 -17700
rect -23120 -17720 -23000 -17700
rect -26500 -17980 -26400 -17720
rect -26100 -17980 -25900 -17720
rect -25600 -17980 -25400 -17720
rect -25100 -17980 -24900 -17720
rect -24600 -17980 -24400 -17720
rect -24100 -17980 -23900 -17720
rect -23600 -17980 -23400 -17720
rect -23100 -17980 -23000 -17720
rect -26500 -18000 -26380 -17980
rect -26120 -18000 -25880 -17980
rect -25620 -18000 -25380 -17980
rect -25120 -18000 -24880 -17980
rect -24620 -18000 -24380 -17980
rect -24120 -18000 -23880 -17980
rect -23620 -18000 -23380 -17980
rect -23120 -18000 -23000 -17980
rect -31500 -18200 -29500 -18100
rect -31500 -18220 -31380 -18200
rect -31120 -18220 -30880 -18200
rect -30620 -18220 -30380 -18200
rect -30120 -18220 -29880 -18200
rect -29620 -18220 -29500 -18200
rect -31500 -18480 -31400 -18220
rect -31100 -18480 -30900 -18220
rect -30600 -18480 -30400 -18220
rect -30100 -18480 -29900 -18220
rect -29600 -18480 -29500 -18220
rect -31500 -18500 -31380 -18480
rect -31120 -18500 -30880 -18480
rect -30620 -18500 -30380 -18480
rect -30120 -18500 -29880 -18480
rect -29620 -18500 -29500 -18480
rect -31500 -18700 -29500 -18500
rect -31500 -18720 -31380 -18700
rect -31120 -18720 -30880 -18700
rect -30620 -18720 -30380 -18700
rect -30120 -18720 -29880 -18700
rect -29620 -18720 -29500 -18700
rect -31500 -18980 -31400 -18720
rect -31100 -18980 -30900 -18720
rect -30600 -18980 -30400 -18720
rect -30100 -18980 -29900 -18720
rect -29600 -18980 -29500 -18720
rect -31500 -19000 -31380 -18980
rect -31120 -19000 -30880 -18980
rect -30620 -19000 -30380 -18980
rect -30120 -19000 -29880 -18980
rect -29620 -19000 -29500 -18980
rect -31500 -19200 -29500 -19000
rect -31500 -19220 -31380 -19200
rect -31120 -19220 -30880 -19200
rect -30620 -19220 -30380 -19200
rect -30120 -19220 -29880 -19200
rect -29620 -19220 -29500 -19200
rect -31500 -19480 -31400 -19220
rect -31100 -19480 -30900 -19220
rect -30600 -19480 -30400 -19220
rect -30100 -19480 -29900 -19220
rect -29600 -19480 -29500 -19220
rect -31500 -19500 -31380 -19480
rect -31120 -19500 -30880 -19480
rect -30620 -19500 -30380 -19480
rect -30120 -19500 -29880 -19480
rect -29620 -19500 -29500 -19480
rect -31500 -19700 -29500 -19500
rect -31500 -19720 -31380 -19700
rect -31120 -19720 -30880 -19700
rect -30620 -19720 -30380 -19700
rect -30120 -19720 -29880 -19700
rect -29620 -19720 -29500 -19700
rect -31500 -19980 -31400 -19720
rect -31100 -19980 -30900 -19720
rect -30600 -19980 -30400 -19720
rect -30100 -19980 -29900 -19720
rect -29600 -19980 -29500 -19720
rect -31500 -20000 -31380 -19980
rect -31120 -20000 -30880 -19980
rect -30620 -20000 -30380 -19980
rect -30120 -20000 -29880 -19980
rect -29620 -20000 -29500 -19980
rect -31500 -20200 -29500 -20000
rect -31500 -20220 -31380 -20200
rect -31120 -20220 -30880 -20200
rect -30620 -20220 -30380 -20200
rect -30120 -20220 -29880 -20200
rect -29620 -20220 -29500 -20200
rect -31500 -20480 -31400 -20220
rect -31100 -20480 -30900 -20220
rect -30600 -20480 -30400 -20220
rect -30100 -20480 -29900 -20220
rect -29600 -20480 -29500 -20220
rect -31500 -20500 -31380 -20480
rect -31120 -20500 -30880 -20480
rect -30620 -20500 -30380 -20480
rect -30120 -20500 -29880 -20480
rect -29620 -20500 -29500 -20480
rect -31500 -20700 -29500 -20500
rect -31500 -20720 -31380 -20700
rect -31120 -20720 -30880 -20700
rect -30620 -20720 -30380 -20700
rect -30120 -20720 -29880 -20700
rect -29620 -20720 -29500 -20700
rect -31500 -20980 -31400 -20720
rect -31100 -20980 -30900 -20720
rect -30600 -20980 -30400 -20720
rect -30100 -20980 -29900 -20720
rect -29600 -20980 -29500 -20720
rect -31500 -21000 -31380 -20980
rect -31120 -21000 -30880 -20980
rect -30620 -21000 -30380 -20980
rect -30120 -21000 -29880 -20980
rect -29620 -21000 -29500 -20980
rect -31500 -21200 -29500 -21000
rect -31500 -21220 -31380 -21200
rect -31120 -21220 -30880 -21200
rect -30620 -21220 -30380 -21200
rect -30120 -21220 -29880 -21200
rect -29620 -21220 -29500 -21200
rect -31500 -21480 -31400 -21220
rect -31100 -21480 -30900 -21220
rect -30600 -21480 -30400 -21220
rect -30100 -21480 -29900 -21220
rect -29600 -21480 -29500 -21220
rect -31500 -21500 -31380 -21480
rect -31120 -21500 -30880 -21480
rect -30620 -21500 -30380 -21480
rect -30120 -21500 -29880 -21480
rect -29620 -21500 -29500 -21480
rect -31500 -21700 -29500 -21500
rect -31500 -21720 -31380 -21700
rect -31120 -21720 -30880 -21700
rect -30620 -21720 -30380 -21700
rect -30120 -21720 -29880 -21700
rect -29620 -21720 -29500 -21700
rect -31500 -21980 -31400 -21720
rect -31100 -21980 -30900 -21720
rect -30600 -21980 -30400 -21720
rect -30100 -21980 -29900 -21720
rect -29600 -21980 -29500 -21720
rect -31500 -22000 -31380 -21980
rect -31120 -22000 -30880 -21980
rect -30620 -22000 -30380 -21980
rect -30120 -22000 -29880 -21980
rect -29620 -22000 -29500 -21980
rect -31500 -22200 -29500 -22000
rect -31500 -22220 -31380 -22200
rect -31120 -22220 -30880 -22200
rect -30620 -22220 -30380 -22200
rect -30120 -22220 -29880 -22200
rect -29620 -22220 -29500 -22200
rect -31500 -22480 -31400 -22220
rect -31100 -22480 -30900 -22220
rect -30600 -22480 -30400 -22220
rect -30100 -22480 -29900 -22220
rect -29600 -22480 -29500 -22220
rect -31500 -22500 -31380 -22480
rect -31120 -22500 -30880 -22480
rect -30620 -22500 -30380 -22480
rect -30120 -22500 -29880 -22480
rect -29620 -22500 -29500 -22480
rect -31500 -22700 -29500 -22500
rect -31500 -22720 -31380 -22700
rect -31120 -22720 -30880 -22700
rect -30620 -22720 -30380 -22700
rect -30120 -22720 -29880 -22700
rect -29620 -22720 -29500 -22700
rect -31500 -22980 -31400 -22720
rect -31100 -22980 -30900 -22720
rect -30600 -22980 -30400 -22720
rect -30100 -22980 -29900 -22720
rect -29600 -22980 -29500 -22720
rect -31500 -23000 -31380 -22980
rect -31120 -23000 -30880 -22980
rect -30620 -23000 -30380 -22980
rect -30120 -23000 -29880 -22980
rect -29620 -23000 -29500 -22980
rect -31500 -23200 -29500 -23000
rect -31500 -23220 -31380 -23200
rect -31120 -23220 -30880 -23200
rect -30620 -23220 -30380 -23200
rect -30120 -23220 -29880 -23200
rect -29620 -23220 -29500 -23200
rect -31500 -23480 -31400 -23220
rect -31100 -23480 -30900 -23220
rect -30600 -23480 -30400 -23220
rect -30100 -23480 -29900 -23220
rect -29600 -23480 -29500 -23220
rect -31500 -23500 -31380 -23480
rect -31120 -23500 -30880 -23480
rect -30620 -23500 -30380 -23480
rect -30120 -23500 -29880 -23480
rect -29620 -23500 -29500 -23480
rect -31500 -23700 -29500 -23500
rect -31500 -23720 -31380 -23700
rect -31120 -23720 -30880 -23700
rect -30620 -23720 -30380 -23700
rect -30120 -23720 -29880 -23700
rect -29620 -23720 -29500 -23700
rect -31500 -23980 -31400 -23720
rect -31100 -23980 -30900 -23720
rect -30600 -23980 -30400 -23720
rect -30100 -23980 -29900 -23720
rect -29600 -23980 -29500 -23720
rect -31500 -24000 -31380 -23980
rect -31120 -24000 -30880 -23980
rect -30620 -24000 -30380 -23980
rect -30120 -24000 -29880 -23980
rect -29620 -24000 -29500 -23980
rect -31500 -24200 -29500 -24000
rect -31500 -24220 -31380 -24200
rect -31120 -24220 -30880 -24200
rect -30620 -24220 -30380 -24200
rect -30120 -24220 -29880 -24200
rect -29620 -24220 -29500 -24200
rect -31500 -24480 -31400 -24220
rect -31100 -24480 -30900 -24220
rect -30600 -24480 -30400 -24220
rect -30100 -24480 -29900 -24220
rect -29600 -24480 -29500 -24220
rect -31500 -24500 -31380 -24480
rect -31120 -24500 -30880 -24480
rect -30620 -24500 -30380 -24480
rect -30120 -24500 -29880 -24480
rect -29620 -24500 -29500 -24480
rect -31500 -24700 -29500 -24500
rect -31500 -24720 -31380 -24700
rect -31120 -24720 -30880 -24700
rect -30620 -24720 -30380 -24700
rect -30120 -24720 -29880 -24700
rect -29620 -24720 -29500 -24700
rect -31500 -24980 -31400 -24720
rect -31100 -24980 -30900 -24720
rect -30600 -24980 -30400 -24720
rect -30100 -24980 -29900 -24720
rect -29600 -24980 -29500 -24720
rect -31500 -25000 -31380 -24980
rect -31120 -25000 -30880 -24980
rect -30620 -25000 -30380 -24980
rect -30120 -25000 -29880 -24980
rect -29620 -25000 -29500 -24980
rect -31500 -25200 -29500 -25000
rect -31500 -25220 -31380 -25200
rect -31120 -25220 -30880 -25200
rect -30620 -25220 -30380 -25200
rect -30120 -25220 -29880 -25200
rect -29620 -25220 -29500 -25200
rect -31500 -25480 -31400 -25220
rect -31100 -25480 -30900 -25220
rect -30600 -25480 -30400 -25220
rect -30100 -25480 -29900 -25220
rect -29600 -25480 -29500 -25220
rect -31500 -25500 -31380 -25480
rect -31120 -25500 -30880 -25480
rect -30620 -25500 -30380 -25480
rect -30120 -25500 -29880 -25480
rect -29620 -25500 -29500 -25480
rect -31500 -25700 -29500 -25500
rect -31500 -25720 -31380 -25700
rect -31120 -25720 -30880 -25700
rect -30620 -25720 -30380 -25700
rect -30120 -25720 -29880 -25700
rect -29620 -25720 -29500 -25700
rect -31500 -25980 -31400 -25720
rect -31100 -25980 -30900 -25720
rect -30600 -25980 -30400 -25720
rect -30100 -25980 -29900 -25720
rect -29600 -25980 -29500 -25720
rect -31500 -26000 -31380 -25980
rect -31120 -26000 -30880 -25980
rect -30620 -26000 -30380 -25980
rect -30120 -26000 -29880 -25980
rect -29620 -26000 -29500 -25980
rect -31500 -26200 -29500 -26000
rect -31500 -26220 -31380 -26200
rect -31120 -26220 -30880 -26200
rect -30620 -26220 -30380 -26200
rect -30120 -26220 -29880 -26200
rect -29620 -26220 -29500 -26200
rect -31500 -26480 -31400 -26220
rect -31100 -26480 -30900 -26220
rect -30600 -26480 -30400 -26220
rect -30100 -26480 -29900 -26220
rect -29600 -26480 -29500 -26220
rect -31500 -26500 -31380 -26480
rect -31120 -26500 -30880 -26480
rect -30620 -26500 -30380 -26480
rect -30120 -26500 -29880 -26480
rect -29620 -26500 -29500 -26480
rect -31500 -26700 -29500 -26500
rect -31500 -26720 -31380 -26700
rect -31120 -26720 -30880 -26700
rect -30620 -26720 -30380 -26700
rect -30120 -26720 -29880 -26700
rect -29620 -26720 -29500 -26700
rect -31500 -26980 -31400 -26720
rect -31100 -26980 -30900 -26720
rect -30600 -26980 -30400 -26720
rect -30100 -26980 -29900 -26720
rect -29600 -26980 -29500 -26720
rect -31500 -27000 -31380 -26980
rect -31120 -27000 -30880 -26980
rect -30620 -27000 -30380 -26980
rect -30120 -27000 -29880 -26980
rect -29620 -27000 -29500 -26980
rect -31500 -27200 -29500 -27000
rect -31500 -27220 -31380 -27200
rect -31120 -27220 -30880 -27200
rect -30620 -27220 -30380 -27200
rect -30120 -27220 -29880 -27200
rect -29620 -27220 -29500 -27200
rect -31500 -27480 -31400 -27220
rect -31100 -27480 -30900 -27220
rect -30600 -27480 -30400 -27220
rect -30100 -27480 -29900 -27220
rect -29600 -27480 -29500 -27220
rect -31500 -27500 -31380 -27480
rect -31120 -27500 -30880 -27480
rect -30620 -27500 -30380 -27480
rect -30120 -27500 -29880 -27480
rect -29620 -27500 -29500 -27480
rect -31500 -27700 -29500 -27500
rect -31500 -27720 -31380 -27700
rect -31120 -27720 -30880 -27700
rect -30620 -27720 -30380 -27700
rect -30120 -27720 -29880 -27700
rect -29620 -27720 -29500 -27700
rect -31500 -27980 -31400 -27720
rect -31100 -27980 -30900 -27720
rect -30600 -27980 -30400 -27720
rect -30100 -27980 -29900 -27720
rect -29600 -27980 -29500 -27720
rect -31500 -28000 -31380 -27980
rect -31120 -28000 -30880 -27980
rect -30620 -28000 -30380 -27980
rect -30120 -28000 -29880 -27980
rect -29620 -28000 -29500 -27980
rect -31500 -28200 -29500 -28000
rect -31500 -28220 -31380 -28200
rect -31120 -28220 -30880 -28200
rect -30620 -28220 -30380 -28200
rect -30120 -28220 -29880 -28200
rect -29620 -28220 -29500 -28200
rect -31500 -28480 -31400 -28220
rect -31100 -28480 -30900 -28220
rect -30600 -28480 -30400 -28220
rect -30100 -28480 -29900 -28220
rect -29600 -28480 -29500 -28220
rect -31500 -28500 -31380 -28480
rect -31120 -28500 -30880 -28480
rect -30620 -28500 -30380 -28480
rect -30120 -28500 -29880 -28480
rect -29620 -28500 -29500 -28480
rect -31500 -28700 -29500 -28500
rect -31500 -28720 -31380 -28700
rect -31120 -28720 -30880 -28700
rect -30620 -28720 -30380 -28700
rect -30120 -28720 -29880 -28700
rect -29620 -28720 -29500 -28700
rect -31500 -28980 -31400 -28720
rect -31100 -28980 -30900 -28720
rect -30600 -28980 -30400 -28720
rect -30100 -28980 -29900 -28720
rect -29600 -28980 -29500 -28720
rect -31500 -29000 -31380 -28980
rect -31120 -29000 -30880 -28980
rect -30620 -29000 -30380 -28980
rect -30120 -29000 -29880 -28980
rect -29620 -29000 -29500 -28980
rect -31500 -29200 -29500 -29000
rect -31500 -29220 -31380 -29200
rect -31120 -29220 -30880 -29200
rect -30620 -29220 -30380 -29200
rect -30120 -29220 -29880 -29200
rect -29620 -29220 -29500 -29200
rect -31500 -29480 -31400 -29220
rect -31100 -29480 -30900 -29220
rect -30600 -29480 -30400 -29220
rect -30100 -29480 -29900 -29220
rect -29600 -29480 -29500 -29220
rect -31500 -29500 -31380 -29480
rect -31120 -29500 -30880 -29480
rect -30620 -29500 -30380 -29480
rect -30120 -29500 -29880 -29480
rect -29620 -29500 -29500 -29480
rect -31500 -29600 -29500 -29500
rect -26500 -18200 -23000 -18000
rect -26500 -18220 -26380 -18200
rect -26120 -18220 -25880 -18200
rect -25620 -18220 -25380 -18200
rect -25120 -18220 -24880 -18200
rect -24620 -18220 -24380 -18200
rect -24120 -18220 -23880 -18200
rect -23620 -18220 -23380 -18200
rect -23120 -18220 -23000 -18200
rect -26500 -18480 -26400 -18220
rect -26100 -18480 -25900 -18220
rect -25600 -18480 -25400 -18220
rect -25100 -18480 -24900 -18220
rect -24600 -18480 -24400 -18220
rect -24100 -18480 -23900 -18220
rect -23600 -18480 -23400 -18220
rect -23100 -18480 -23000 -18220
rect -26500 -18500 -26380 -18480
rect -26120 -18500 -25880 -18480
rect -25620 -18500 -25380 -18480
rect -25120 -18500 -24880 -18480
rect -24620 -18500 -24380 -18480
rect -24120 -18500 -23880 -18480
rect -23620 -18500 -23380 -18480
rect -23120 -18500 -23000 -18480
rect -26500 -18700 -23000 -18500
rect -26500 -18720 -26380 -18700
rect -26120 -18720 -25880 -18700
rect -25620 -18720 -25380 -18700
rect -25120 -18720 -24880 -18700
rect -24620 -18720 -24380 -18700
rect -24120 -18720 -23880 -18700
rect -23620 -18720 -23380 -18700
rect -23120 -18720 -23000 -18700
rect -26500 -18980 -26400 -18720
rect -26100 -18980 -25900 -18720
rect -25600 -18980 -25400 -18720
rect -25100 -18980 -24900 -18720
rect -24600 -18980 -24400 -18720
rect -24100 -18980 -23900 -18720
rect -23600 -18980 -23400 -18720
rect -23100 -18980 -23000 -18720
rect -26500 -19000 -26380 -18980
rect -26120 -19000 -25880 -18980
rect -25620 -19000 -25380 -18980
rect -25120 -19000 -24880 -18980
rect -24620 -19000 -24380 -18980
rect -24120 -19000 -23880 -18980
rect -23620 -19000 -23380 -18980
rect -23120 -19000 -23000 -18980
rect -26500 -19200 -23000 -19000
rect -26500 -19220 -26380 -19200
rect -26120 -19220 -25880 -19200
rect -25620 -19220 -25380 -19200
rect -25120 -19220 -24880 -19200
rect -24620 -19220 -24380 -19200
rect -24120 -19220 -23880 -19200
rect -23620 -19220 -23380 -19200
rect -23120 -19220 -23000 -19200
rect -26500 -19480 -26400 -19220
rect -26100 -19480 -25900 -19220
rect -25600 -19480 -25400 -19220
rect -25100 -19480 -24900 -19220
rect -24600 -19480 -24400 -19220
rect -24100 -19480 -23900 -19220
rect -23600 -19480 -23400 -19220
rect -23100 -19480 -23000 -19220
rect -26500 -19500 -26380 -19480
rect -26120 -19500 -25880 -19480
rect -25620 -19500 -25380 -19480
rect -25120 -19500 -24880 -19480
rect -24620 -19500 -24380 -19480
rect -24120 -19500 -23880 -19480
rect -23620 -19500 -23380 -19480
rect -23120 -19500 -23000 -19480
rect -26500 -19700 -23000 -19500
rect -26500 -19720 -26380 -19700
rect -26120 -19720 -25880 -19700
rect -25620 -19720 -25380 -19700
rect -25120 -19720 -24880 -19700
rect -24620 -19720 -24380 -19700
rect -24120 -19720 -23880 -19700
rect -23620 -19720 -23380 -19700
rect -23120 -19720 -23000 -19700
rect -26500 -19980 -26400 -19720
rect -26100 -19980 -25900 -19720
rect -25600 -19980 -25400 -19720
rect -25100 -19980 -24900 -19720
rect -24600 -19980 -24400 -19720
rect -24100 -19980 -23900 -19720
rect -23600 -19980 -23400 -19720
rect -23100 -19980 -23000 -19720
rect -26500 -20000 -26380 -19980
rect -26120 -20000 -25880 -19980
rect -25620 -20000 -25380 -19980
rect -25120 -20000 -24880 -19980
rect -24620 -20000 -24380 -19980
rect -24120 -20000 -23880 -19980
rect -23620 -20000 -23380 -19980
rect -23120 -20000 -23000 -19980
rect -26500 -20200 -23000 -20000
rect -26500 -20220 -26380 -20200
rect -26120 -20220 -25880 -20200
rect -25620 -20220 -25380 -20200
rect -25120 -20220 -24880 -20200
rect -24620 -20220 -24380 -20200
rect -24120 -20220 -23880 -20200
rect -23620 -20220 -23380 -20200
rect -23120 -20220 -23000 -20200
rect -26500 -20480 -26400 -20220
rect -26100 -20480 -25900 -20220
rect -25600 -20480 -25400 -20220
rect -25100 -20480 -24900 -20220
rect -24600 -20480 -24400 -20220
rect -24100 -20480 -23900 -20220
rect -23600 -20480 -23400 -20220
rect -23100 -20480 -23000 -20220
rect -26500 -20500 -26380 -20480
rect -26120 -20500 -25880 -20480
rect -25620 -20500 -25380 -20480
rect -25120 -20500 -24880 -20480
rect -24620 -20500 -24380 -20480
rect -24120 -20500 -23880 -20480
rect -23620 -20500 -23380 -20480
rect -23120 -20500 -23000 -20480
rect -26500 -20700 -23000 -20500
rect -26500 -20720 -26380 -20700
rect -26120 -20720 -25880 -20700
rect -25620 -20720 -25380 -20700
rect -25120 -20720 -24880 -20700
rect -24620 -20720 -24380 -20700
rect -24120 -20720 -23880 -20700
rect -23620 -20720 -23380 -20700
rect -23120 -20720 -23000 -20700
rect -26500 -20980 -26400 -20720
rect -26100 -20980 -25900 -20720
rect -25600 -20980 -25400 -20720
rect -25100 -20980 -24900 -20720
rect -24600 -20980 -24400 -20720
rect -24100 -20980 -23900 -20720
rect -23600 -20980 -23400 -20720
rect -23100 -20980 -23000 -20720
rect -26500 -21000 -26380 -20980
rect -26120 -21000 -25880 -20980
rect -25620 -21000 -25380 -20980
rect -25120 -21000 -24880 -20980
rect -24620 -21000 -24380 -20980
rect -24120 -21000 -23880 -20980
rect -23620 -21000 -23380 -20980
rect -23120 -21000 -23000 -20980
rect -26500 -21100 -23000 -21000
rect -19000 -16700 -15000 -16600
rect -19000 -16720 -18880 -16700
rect -18620 -16720 -18380 -16700
rect -18120 -16720 -17880 -16700
rect -17620 -16720 -17380 -16700
rect -17120 -16720 -16880 -16700
rect -16620 -16720 -16380 -16700
rect -16120 -16720 -15880 -16700
rect -15620 -16720 -15380 -16700
rect -15120 -16720 -15000 -16700
rect -19000 -16980 -18900 -16720
rect -18600 -16980 -18400 -16720
rect -18100 -16980 -17900 -16720
rect -17600 -16980 -17400 -16720
rect -17100 -16980 -16900 -16720
rect -16600 -16980 -16400 -16720
rect -16100 -16980 -15900 -16720
rect -15600 -16980 -15400 -16720
rect -15100 -16980 -15000 -16720
rect -19000 -17000 -18880 -16980
rect -18620 -17000 -18380 -16980
rect -18120 -17000 -17880 -16980
rect -17620 -17000 -17380 -16980
rect -17120 -17000 -16880 -16980
rect -16620 -17000 -16380 -16980
rect -16120 -17000 -15880 -16980
rect -15620 -17000 -15380 -16980
rect -15120 -17000 -15000 -16980
rect -19000 -17200 -15000 -17000
rect -19000 -17220 -18880 -17200
rect -18620 -17220 -18380 -17200
rect -18120 -17220 -17880 -17200
rect -17620 -17220 -17380 -17200
rect -17120 -17220 -16880 -17200
rect -16620 -17220 -16380 -17200
rect -16120 -17220 -15880 -17200
rect -15620 -17220 -15380 -17200
rect -15120 -17220 -15000 -17200
rect -19000 -17480 -18900 -17220
rect -18600 -17480 -18400 -17220
rect -18100 -17480 -17900 -17220
rect -17600 -17480 -17400 -17220
rect -17100 -17480 -16900 -17220
rect -16600 -17480 -16400 -17220
rect -16100 -17480 -15900 -17220
rect -15600 -17480 -15400 -17220
rect -15100 -17480 -15000 -17220
rect -19000 -17500 -18880 -17480
rect -18620 -17500 -18380 -17480
rect -18120 -17500 -17880 -17480
rect -17620 -17500 -17380 -17480
rect -17120 -17500 -16880 -17480
rect -16620 -17500 -16380 -17480
rect -16120 -17500 -15880 -17480
rect -15620 -17500 -15380 -17480
rect -15120 -17500 -15000 -17480
rect -19000 -17700 -15000 -17500
rect -19000 -17720 -18880 -17700
rect -18620 -17720 -18380 -17700
rect -18120 -17720 -17880 -17700
rect -17620 -17720 -17380 -17700
rect -17120 -17720 -16880 -17700
rect -16620 -17720 -16380 -17700
rect -16120 -17720 -15880 -17700
rect -15620 -17720 -15380 -17700
rect -15120 -17720 -15000 -17700
rect -19000 -17980 -18900 -17720
rect -18600 -17980 -18400 -17720
rect -18100 -17980 -17900 -17720
rect -17600 -17980 -17400 -17720
rect -17100 -17980 -16900 -17720
rect -16600 -17980 -16400 -17720
rect -16100 -17980 -15900 -17720
rect -15600 -17980 -15400 -17720
rect -15100 -17980 -15000 -17720
rect -19000 -18000 -18880 -17980
rect -18620 -18000 -18380 -17980
rect -18120 -18000 -17880 -17980
rect -17620 -18000 -17380 -17980
rect -17120 -18000 -16880 -17980
rect -16620 -18000 -16380 -17980
rect -16120 -18000 -15880 -17980
rect -15620 -18000 -15380 -17980
rect -15120 -18000 -15000 -17980
rect -19000 -18200 -15000 -18000
rect -19000 -18220 -18880 -18200
rect -18620 -18220 -18380 -18200
rect -18120 -18220 -17880 -18200
rect -17620 -18220 -17380 -18200
rect -17120 -18220 -16880 -18200
rect -16620 -18220 -16380 -18200
rect -16120 -18220 -15880 -18200
rect -15620 -18220 -15380 -18200
rect -15120 -18220 -15000 -18200
rect -19000 -18480 -18900 -18220
rect -18600 -18480 -18400 -18220
rect -18100 -18480 -17900 -18220
rect -17600 -18480 -17400 -18220
rect -17100 -18480 -16900 -18220
rect -16600 -18480 -16400 -18220
rect -16100 -18480 -15900 -18220
rect -15600 -18480 -15400 -18220
rect -15100 -18480 -15000 -18220
rect -19000 -18500 -18880 -18480
rect -18620 -18500 -18380 -18480
rect -18120 -18500 -17880 -18480
rect -17620 -18500 -17380 -18480
rect -17120 -18500 -16880 -18480
rect -16620 -18500 -16380 -18480
rect -16120 -18500 -15880 -18480
rect -15620 -18500 -15380 -18480
rect -15120 -18500 -15000 -18480
rect -19000 -18700 -15000 -18500
rect -19000 -18720 -18880 -18700
rect -18620 -18720 -18380 -18700
rect -18120 -18720 -17880 -18700
rect -17620 -18720 -17380 -18700
rect -17120 -18720 -16880 -18700
rect -16620 -18720 -16380 -18700
rect -16120 -18720 -15880 -18700
rect -15620 -18720 -15380 -18700
rect -15120 -18720 -15000 -18700
rect -19000 -18980 -18900 -18720
rect -18600 -18980 -18400 -18720
rect -18100 -18980 -17900 -18720
rect -17600 -18980 -17400 -18720
rect -17100 -18980 -16900 -18720
rect -16600 -18980 -16400 -18720
rect -16100 -18980 -15900 -18720
rect -15600 -18980 -15400 -18720
rect -15100 -18980 -15000 -18720
rect -19000 -19000 -18880 -18980
rect -18620 -19000 -18380 -18980
rect -18120 -19000 -17880 -18980
rect -17620 -19000 -17380 -18980
rect -17120 -19000 -16880 -18980
rect -16620 -19000 -16380 -18980
rect -16120 -19000 -15880 -18980
rect -15620 -19000 -15380 -18980
rect -15120 -19000 -15000 -18980
rect -19000 -19200 -15000 -19000
rect -19000 -19220 -18880 -19200
rect -18620 -19220 -18380 -19200
rect -18120 -19220 -17880 -19200
rect -17620 -19220 -17380 -19200
rect -17120 -19220 -16880 -19200
rect -16620 -19220 -16380 -19200
rect -16120 -19220 -15880 -19200
rect -15620 -19220 -15380 -19200
rect -15120 -19220 -15000 -19200
rect -19000 -19480 -18900 -19220
rect -18600 -19480 -18400 -19220
rect -18100 -19480 -17900 -19220
rect -17600 -19480 -17400 -19220
rect -17100 -19480 -16900 -19220
rect -16600 -19480 -16400 -19220
rect -16100 -19480 -15900 -19220
rect -15600 -19480 -15400 -19220
rect -15100 -19480 -15000 -19220
rect -19000 -19500 -18880 -19480
rect -18620 -19500 -18380 -19480
rect -18120 -19500 -17880 -19480
rect -17620 -19500 -17380 -19480
rect -17120 -19500 -16880 -19480
rect -16620 -19500 -16380 -19480
rect -16120 -19500 -15880 -19480
rect -15620 -19500 -15380 -19480
rect -15120 -19500 -15000 -19480
rect -19000 -19700 -15000 -19500
rect -19000 -19720 -18880 -19700
rect -18620 -19720 -18380 -19700
rect -18120 -19720 -17880 -19700
rect -17620 -19720 -17380 -19700
rect -17120 -19720 -16880 -19700
rect -16620 -19720 -16380 -19700
rect -16120 -19720 -15880 -19700
rect -15620 -19720 -15380 -19700
rect -15120 -19720 -15000 -19700
rect -19000 -19980 -18900 -19720
rect -18600 -19980 -18400 -19720
rect -18100 -19980 -17900 -19720
rect -17600 -19980 -17400 -19720
rect -17100 -19980 -16900 -19720
rect -16600 -19980 -16400 -19720
rect -16100 -19980 -15900 -19720
rect -15600 -19980 -15400 -19720
rect -15100 -19980 -15000 -19720
rect -19000 -20000 -18880 -19980
rect -18620 -20000 -18380 -19980
rect -18120 -20000 -17880 -19980
rect -17620 -20000 -17380 -19980
rect -17120 -20000 -16880 -19980
rect -16620 -20000 -16380 -19980
rect -16120 -20000 -15880 -19980
rect -15620 -20000 -15380 -19980
rect -15120 -20000 -15000 -19980
rect -19000 -20200 -15000 -20000
rect -19000 -20220 -18880 -20200
rect -18620 -20220 -18380 -20200
rect -18120 -20220 -17880 -20200
rect -17620 -20220 -17380 -20200
rect -17120 -20220 -16880 -20200
rect -16620 -20220 -16380 -20200
rect -16120 -20220 -15880 -20200
rect -15620 -20220 -15380 -20200
rect -15120 -20220 -15000 -20200
rect -19000 -20480 -18900 -20220
rect -18600 -20480 -18400 -20220
rect -18100 -20480 -17900 -20220
rect -17600 -20480 -17400 -20220
rect -17100 -20480 -16900 -20220
rect -16600 -20480 -16400 -20220
rect -16100 -20480 -15900 -20220
rect -15600 -20480 -15400 -20220
rect -15100 -20480 -15000 -20220
rect -19000 -20500 -18880 -20480
rect -18620 -20500 -18380 -20480
rect -18120 -20500 -17880 -20480
rect -17620 -20500 -17380 -20480
rect -17120 -20500 -16880 -20480
rect -16620 -20500 -16380 -20480
rect -16120 -20500 -15880 -20480
rect -15620 -20500 -15380 -20480
rect -15120 -20500 -15000 -20480
rect -19000 -20700 -15000 -20500
rect -19000 -20720 -18880 -20700
rect -18620 -20720 -18380 -20700
rect -18120 -20720 -17880 -20700
rect -17620 -20720 -17380 -20700
rect -17120 -20720 -16880 -20700
rect -16620 -20720 -16380 -20700
rect -16120 -20720 -15880 -20700
rect -15620 -20720 -15380 -20700
rect -15120 -20720 -15000 -20700
rect -19000 -20980 -18900 -20720
rect -18600 -20980 -18400 -20720
rect -18100 -20980 -17900 -20720
rect -17600 -20980 -17400 -20720
rect -17100 -20980 -16900 -20720
rect -16600 -20980 -16400 -20720
rect -16100 -20980 -15900 -20720
rect -15600 -20980 -15400 -20720
rect -15100 -20980 -15000 -20720
rect -19000 -21000 -18880 -20980
rect -18620 -21000 -18380 -20980
rect -18120 -21000 -17880 -20980
rect -17620 -21000 -17380 -20980
rect -17120 -21000 -16880 -20980
rect -16620 -21000 -16380 -20980
rect -16120 -21000 -15880 -20980
rect -15620 -21000 -15380 -20980
rect -15120 -21000 -15000 -20980
rect -19000 -21100 -15000 -21000
rect -26500 -21200 -15000 -21100
rect -26500 -21220 -26380 -21200
rect -26120 -21220 -25880 -21200
rect -25620 -21220 -25380 -21200
rect -25120 -21220 -24880 -21200
rect -24620 -21220 -24380 -21200
rect -24120 -21220 -23880 -21200
rect -23620 -21220 -23380 -21200
rect -23120 -21220 -22880 -21200
rect -22620 -21220 -22380 -21200
rect -22120 -21220 -21880 -21200
rect -21620 -21220 -21380 -21200
rect -21120 -21220 -20880 -21200
rect -20620 -21220 -20380 -21200
rect -20120 -21220 -19880 -21200
rect -19620 -21220 -19380 -21200
rect -19120 -21220 -18880 -21200
rect -18620 -21220 -18380 -21200
rect -18120 -21220 -17880 -21200
rect -17620 -21220 -17380 -21200
rect -17120 -21220 -16880 -21200
rect -16620 -21220 -16380 -21200
rect -16120 -21220 -15880 -21200
rect -15620 -21220 -15380 -21200
rect -15120 -21220 -15000 -21200
rect -26500 -21480 -26400 -21220
rect -26100 -21480 -25900 -21220
rect -25600 -21480 -25400 -21220
rect -25100 -21480 -24900 -21220
rect -24600 -21480 -24400 -21220
rect -24100 -21480 -23900 -21220
rect -23600 -21480 -23400 -21220
rect -23100 -21480 -22900 -21220
rect -22600 -21480 -22400 -21220
rect -22100 -21480 -21900 -21220
rect -21600 -21480 -21400 -21220
rect -21100 -21480 -20900 -21220
rect -20600 -21480 -20400 -21220
rect -20100 -21480 -19900 -21220
rect -19600 -21480 -19400 -21220
rect -19100 -21480 -18900 -21220
rect -18600 -21480 -18400 -21220
rect -18100 -21480 -17900 -21220
rect -17600 -21480 -17400 -21220
rect -17100 -21480 -16900 -21220
rect -16600 -21480 -16400 -21220
rect -16100 -21480 -15900 -21220
rect -15600 -21480 -15400 -21220
rect -15100 -21480 -15000 -21220
rect -26500 -21500 -26380 -21480
rect -26120 -21500 -25880 -21480
rect -25620 -21500 -25380 -21480
rect -25120 -21500 -24880 -21480
rect -24620 -21500 -24380 -21480
rect -24120 -21500 -23880 -21480
rect -23620 -21500 -23380 -21480
rect -23120 -21500 -22880 -21480
rect -22620 -21500 -22380 -21480
rect -22120 -21500 -21880 -21480
rect -21620 -21500 -21380 -21480
rect -21120 -21500 -20880 -21480
rect -20620 -21500 -20380 -21480
rect -20120 -21500 -19880 -21480
rect -19620 -21500 -19380 -21480
rect -19120 -21500 -18880 -21480
rect -18620 -21500 -18380 -21480
rect -18120 -21500 -17880 -21480
rect -17620 -21500 -17380 -21480
rect -17120 -21500 -16880 -21480
rect -16620 -21500 -16380 -21480
rect -16120 -21500 -15880 -21480
rect -15620 -21500 -15380 -21480
rect -15120 -21500 -15000 -21480
rect -26500 -21700 -15000 -21500
rect -26500 -21720 -26380 -21700
rect -26120 -21720 -25880 -21700
rect -25620 -21720 -25380 -21700
rect -25120 -21720 -24880 -21700
rect -24620 -21720 -24380 -21700
rect -24120 -21720 -23880 -21700
rect -23620 -21720 -23380 -21700
rect -23120 -21720 -22880 -21700
rect -22620 -21720 -22380 -21700
rect -22120 -21720 -21880 -21700
rect -21620 -21720 -21380 -21700
rect -21120 -21720 -20880 -21700
rect -20620 -21720 -20380 -21700
rect -20120 -21720 -19880 -21700
rect -19620 -21720 -19380 -21700
rect -19120 -21720 -18880 -21700
rect -18620 -21720 -18380 -21700
rect -18120 -21720 -17880 -21700
rect -17620 -21720 -17380 -21700
rect -17120 -21720 -16880 -21700
rect -16620 -21720 -16380 -21700
rect -16120 -21720 -15880 -21700
rect -15620 -21720 -15380 -21700
rect -15120 -21720 -15000 -21700
rect -26500 -21980 -26400 -21720
rect -26100 -21980 -25900 -21720
rect -25600 -21980 -25400 -21720
rect -25100 -21980 -24900 -21720
rect -24600 -21980 -24400 -21720
rect -24100 -21980 -23900 -21720
rect -23600 -21980 -23400 -21720
rect -23100 -21980 -22900 -21720
rect -22600 -21980 -22400 -21720
rect -22100 -21980 -21900 -21720
rect -21600 -21980 -21400 -21720
rect -21100 -21980 -20900 -21720
rect -20600 -21980 -20400 -21720
rect -20100 -21980 -19900 -21720
rect -19600 -21980 -19400 -21720
rect -19100 -21980 -18900 -21720
rect -18600 -21980 -18400 -21720
rect -18100 -21980 -17900 -21720
rect -17600 -21980 -17400 -21720
rect -17100 -21980 -16900 -21720
rect -16600 -21980 -16400 -21720
rect -16100 -21980 -15900 -21720
rect -15600 -21980 -15400 -21720
rect -15100 -21980 -15000 -21720
rect -26500 -22000 -26380 -21980
rect -26120 -22000 -25880 -21980
rect -25620 -22000 -25380 -21980
rect -25120 -22000 -24880 -21980
rect -24620 -22000 -24380 -21980
rect -24120 -22000 -23880 -21980
rect -23620 -22000 -23380 -21980
rect -23120 -22000 -22880 -21980
rect -22620 -22000 -22380 -21980
rect -22120 -22000 -21880 -21980
rect -21620 -22000 -21380 -21980
rect -21120 -22000 -20880 -21980
rect -20620 -22000 -20380 -21980
rect -20120 -22000 -19880 -21980
rect -19620 -22000 -19380 -21980
rect -19120 -22000 -18880 -21980
rect -18620 -22000 -18380 -21980
rect -18120 -22000 -17880 -21980
rect -17620 -22000 -17380 -21980
rect -17120 -22000 -16880 -21980
rect -16620 -22000 -16380 -21980
rect -16120 -22000 -15880 -21980
rect -15620 -22000 -15380 -21980
rect -15120 -22000 -15000 -21980
rect -26500 -22200 -15000 -22000
rect -26500 -22220 -26380 -22200
rect -26120 -22220 -25880 -22200
rect -25620 -22220 -25380 -22200
rect -25120 -22220 -24880 -22200
rect -24620 -22220 -24380 -22200
rect -24120 -22220 -23880 -22200
rect -23620 -22220 -23380 -22200
rect -23120 -22220 -22880 -22200
rect -22620 -22220 -22380 -22200
rect -22120 -22220 -21880 -22200
rect -21620 -22220 -21380 -22200
rect -21120 -22220 -20880 -22200
rect -20620 -22220 -20380 -22200
rect -20120 -22220 -19880 -22200
rect -19620 -22220 -19380 -22200
rect -19120 -22220 -18880 -22200
rect -18620 -22220 -18380 -22200
rect -18120 -22220 -17880 -22200
rect -17620 -22220 -17380 -22200
rect -17120 -22220 -16880 -22200
rect -16620 -22220 -16380 -22200
rect -16120 -22220 -15880 -22200
rect -15620 -22220 -15380 -22200
rect -15120 -22220 -15000 -22200
rect -26500 -22480 -26400 -22220
rect -26100 -22480 -25900 -22220
rect -25600 -22480 -25400 -22220
rect -25100 -22480 -24900 -22220
rect -24600 -22480 -24400 -22220
rect -24100 -22480 -23900 -22220
rect -23600 -22480 -23400 -22220
rect -23100 -22480 -22900 -22220
rect -22600 -22480 -22400 -22220
rect -22100 -22480 -21900 -22220
rect -21600 -22480 -21400 -22220
rect -21100 -22480 -20900 -22220
rect -20600 -22480 -20400 -22220
rect -20100 -22480 -19900 -22220
rect -19600 -22480 -19400 -22220
rect -19100 -22480 -18900 -22220
rect -18600 -22480 -18400 -22220
rect -18100 -22480 -17900 -22220
rect -17600 -22480 -17400 -22220
rect -17100 -22480 -16900 -22220
rect -16600 -22480 -16400 -22220
rect -16100 -22480 -15900 -22220
rect -15600 -22480 -15400 -22220
rect -15100 -22480 -15000 -22220
rect -26500 -22500 -26380 -22480
rect -26120 -22500 -25880 -22480
rect -25620 -22500 -25380 -22480
rect -25120 -22500 -24880 -22480
rect -24620 -22500 -24380 -22480
rect -24120 -22500 -23880 -22480
rect -23620 -22500 -23380 -22480
rect -23120 -22500 -22880 -22480
rect -22620 -22500 -22380 -22480
rect -22120 -22500 -21880 -22480
rect -21620 -22500 -21380 -22480
rect -21120 -22500 -20880 -22480
rect -20620 -22500 -20380 -22480
rect -20120 -22500 -19880 -22480
rect -19620 -22500 -19380 -22480
rect -19120 -22500 -18880 -22480
rect -18620 -22500 -18380 -22480
rect -18120 -22500 -17880 -22480
rect -17620 -22500 -17380 -22480
rect -17120 -22500 -16880 -22480
rect -16620 -22500 -16380 -22480
rect -16120 -22500 -15880 -22480
rect -15620 -22500 -15380 -22480
rect -15120 -22500 -15000 -22480
rect -26500 -22700 -15000 -22500
rect -26500 -22720 -26380 -22700
rect -26120 -22720 -25880 -22700
rect -25620 -22720 -25380 -22700
rect -25120 -22720 -24880 -22700
rect -24620 -22720 -24380 -22700
rect -24120 -22720 -23880 -22700
rect -23620 -22720 -23380 -22700
rect -23120 -22720 -22880 -22700
rect -22620 -22720 -22380 -22700
rect -22120 -22720 -21880 -22700
rect -21620 -22720 -21380 -22700
rect -21120 -22720 -20880 -22700
rect -20620 -22720 -20380 -22700
rect -20120 -22720 -19880 -22700
rect -19620 -22720 -19380 -22700
rect -19120 -22720 -18880 -22700
rect -18620 -22720 -18380 -22700
rect -18120 -22720 -17880 -22700
rect -17620 -22720 -17380 -22700
rect -17120 -22720 -16880 -22700
rect -16620 -22720 -16380 -22700
rect -16120 -22720 -15880 -22700
rect -15620 -22720 -15380 -22700
rect -15120 -22720 -15000 -22700
rect -26500 -22980 -26400 -22720
rect -26100 -22980 -25900 -22720
rect -25600 -22980 -25400 -22720
rect -25100 -22980 -24900 -22720
rect -24600 -22980 -24400 -22720
rect -24100 -22980 -23900 -22720
rect -23600 -22980 -23400 -22720
rect -23100 -22980 -22900 -22720
rect -22600 -22980 -22400 -22720
rect -22100 -22980 -21900 -22720
rect -21600 -22980 -21400 -22720
rect -21100 -22980 -20900 -22720
rect -20600 -22980 -20400 -22720
rect -20100 -22980 -19900 -22720
rect -19600 -22980 -19400 -22720
rect -19100 -22980 -18900 -22720
rect -18600 -22980 -18400 -22720
rect -18100 -22980 -17900 -22720
rect -17600 -22980 -17400 -22720
rect -17100 -22980 -16900 -22720
rect -16600 -22980 -16400 -22720
rect -16100 -22980 -15900 -22720
rect -15600 -22980 -15400 -22720
rect -15100 -22980 -15000 -22720
rect -26500 -23000 -26380 -22980
rect -26120 -23000 -25880 -22980
rect -25620 -23000 -25380 -22980
rect -25120 -23000 -24880 -22980
rect -24620 -23000 -24380 -22980
rect -24120 -23000 -23880 -22980
rect -23620 -23000 -23380 -22980
rect -23120 -23000 -22880 -22980
rect -22620 -23000 -22380 -22980
rect -22120 -23000 -21880 -22980
rect -21620 -23000 -21380 -22980
rect -21120 -23000 -20880 -22980
rect -20620 -23000 -20380 -22980
rect -20120 -23000 -19880 -22980
rect -19620 -23000 -19380 -22980
rect -19120 -23000 -18880 -22980
rect -18620 -23000 -18380 -22980
rect -18120 -23000 -17880 -22980
rect -17620 -23000 -17380 -22980
rect -17120 -23000 -16880 -22980
rect -16620 -23000 -16380 -22980
rect -16120 -23000 -15880 -22980
rect -15620 -23000 -15380 -22980
rect -15120 -23000 -15000 -22980
rect -26500 -23200 -15000 -23000
rect -26500 -23220 -26380 -23200
rect -26120 -23220 -25880 -23200
rect -25620 -23220 -25380 -23200
rect -25120 -23220 -24880 -23200
rect -24620 -23220 -24380 -23200
rect -24120 -23220 -23880 -23200
rect -23620 -23220 -23380 -23200
rect -23120 -23220 -22880 -23200
rect -22620 -23220 -22380 -23200
rect -22120 -23220 -21880 -23200
rect -21620 -23220 -21380 -23200
rect -21120 -23220 -20880 -23200
rect -20620 -23220 -20380 -23200
rect -20120 -23220 -19880 -23200
rect -19620 -23220 -19380 -23200
rect -19120 -23220 -18880 -23200
rect -18620 -23220 -18380 -23200
rect -18120 -23220 -17880 -23200
rect -17620 -23220 -17380 -23200
rect -17120 -23220 -16880 -23200
rect -16620 -23220 -16380 -23200
rect -16120 -23220 -15880 -23200
rect -15620 -23220 -15380 -23200
rect -15120 -23220 -15000 -23200
rect -26500 -23480 -26400 -23220
rect -26100 -23480 -25900 -23220
rect -25600 -23480 -25400 -23220
rect -25100 -23480 -24900 -23220
rect -24600 -23480 -24400 -23220
rect -24100 -23480 -23900 -23220
rect -23600 -23480 -23400 -23220
rect -23100 -23480 -22900 -23220
rect -22600 -23480 -22400 -23220
rect -22100 -23480 -21900 -23220
rect -21600 -23480 -21400 -23220
rect -21100 -23480 -20900 -23220
rect -20600 -23480 -20400 -23220
rect -20100 -23480 -19900 -23220
rect -19600 -23480 -19400 -23220
rect -19100 -23480 -18900 -23220
rect -18600 -23480 -18400 -23220
rect -18100 -23480 -17900 -23220
rect -17600 -23480 -17400 -23220
rect -17100 -23480 -16900 -23220
rect -16600 -23480 -16400 -23220
rect -16100 -23480 -15900 -23220
rect -15600 -23480 -15400 -23220
rect -15100 -23480 -15000 -23220
rect -26500 -23500 -26380 -23480
rect -26120 -23500 -25880 -23480
rect -25620 -23500 -25380 -23480
rect -25120 -23500 -24880 -23480
rect -24620 -23500 -24380 -23480
rect -24120 -23500 -23880 -23480
rect -23620 -23500 -23380 -23480
rect -23120 -23500 -22880 -23480
rect -22620 -23500 -22380 -23480
rect -22120 -23500 -21880 -23480
rect -21620 -23500 -21380 -23480
rect -21120 -23500 -20880 -23480
rect -20620 -23500 -20380 -23480
rect -20120 -23500 -19880 -23480
rect -19620 -23500 -19380 -23480
rect -19120 -23500 -18880 -23480
rect -18620 -23500 -18380 -23480
rect -18120 -23500 -17880 -23480
rect -17620 -23500 -17380 -23480
rect -17120 -23500 -16880 -23480
rect -16620 -23500 -16380 -23480
rect -16120 -23500 -15880 -23480
rect -15620 -23500 -15380 -23480
rect -15120 -23500 -15000 -23480
rect -26500 -23700 -15000 -23500
rect -26500 -23720 -26380 -23700
rect -26120 -23720 -25880 -23700
rect -25620 -23720 -25380 -23700
rect -25120 -23720 -24880 -23700
rect -24620 -23720 -24380 -23700
rect -24120 -23720 -23880 -23700
rect -23620 -23720 -23380 -23700
rect -23120 -23720 -22880 -23700
rect -22620 -23720 -22380 -23700
rect -22120 -23720 -21880 -23700
rect -21620 -23720 -21380 -23700
rect -21120 -23720 -20880 -23700
rect -20620 -23720 -20380 -23700
rect -20120 -23720 -19880 -23700
rect -19620 -23720 -19380 -23700
rect -19120 -23720 -18880 -23700
rect -18620 -23720 -18380 -23700
rect -18120 -23720 -17880 -23700
rect -17620 -23720 -17380 -23700
rect -17120 -23720 -16880 -23700
rect -16620 -23720 -16380 -23700
rect -16120 -23720 -15880 -23700
rect -15620 -23720 -15380 -23700
rect -15120 -23720 -15000 -23700
rect -26500 -23980 -26400 -23720
rect -26100 -23980 -25900 -23720
rect -25600 -23980 -25400 -23720
rect -25100 -23980 -24900 -23720
rect -24600 -23980 -24400 -23720
rect -24100 -23980 -23900 -23720
rect -23600 -23980 -23400 -23720
rect -23100 -23980 -22900 -23720
rect -22600 -23980 -22400 -23720
rect -22100 -23980 -21900 -23720
rect -21600 -23980 -21400 -23720
rect -21100 -23980 -20900 -23720
rect -20600 -23980 -20400 -23720
rect -20100 -23980 -19900 -23720
rect -19600 -23980 -19400 -23720
rect -19100 -23980 -18900 -23720
rect -18600 -23980 -18400 -23720
rect -18100 -23980 -17900 -23720
rect -17600 -23980 -17400 -23720
rect -17100 -23980 -16900 -23720
rect -16600 -23980 -16400 -23720
rect -16100 -23980 -15900 -23720
rect -15600 -23980 -15400 -23720
rect -15100 -23980 -15000 -23720
rect -26500 -24000 -26380 -23980
rect -26120 -24000 -25880 -23980
rect -25620 -24000 -25380 -23980
rect -25120 -24000 -24880 -23980
rect -24620 -24000 -24380 -23980
rect -24120 -24000 -23880 -23980
rect -23620 -24000 -23380 -23980
rect -23120 -24000 -22880 -23980
rect -22620 -24000 -22380 -23980
rect -22120 -24000 -21880 -23980
rect -21620 -24000 -21380 -23980
rect -21120 -24000 -20880 -23980
rect -20620 -24000 -20380 -23980
rect -20120 -24000 -19880 -23980
rect -19620 -24000 -19380 -23980
rect -19120 -24000 -18880 -23980
rect -18620 -24000 -18380 -23980
rect -18120 -24000 -17880 -23980
rect -17620 -24000 -17380 -23980
rect -17120 -24000 -16880 -23980
rect -16620 -24000 -16380 -23980
rect -16120 -24000 -15880 -23980
rect -15620 -24000 -15380 -23980
rect -15120 -24000 -15000 -23980
rect -26500 -24100 -15000 -24000
rect 23500 -13200 24000 -13000
rect 23500 -13220 23620 -13200
rect 23880 -13220 24000 -13200
rect 23500 -13480 23600 -13220
rect 23900 -13480 24000 -13220
rect 23500 -13500 23620 -13480
rect 23880 -13500 24000 -13480
rect 23500 -13700 24000 -13500
rect 23500 -13720 23620 -13700
rect 23880 -13720 24000 -13700
rect 23500 -13980 23600 -13720
rect 23900 -13980 24000 -13720
rect 23500 -14000 23620 -13980
rect 23880 -14000 24000 -13980
rect 23500 -14200 24000 -14000
rect 23500 -14220 23620 -14200
rect 23880 -14220 24000 -14200
rect 23500 -14480 23600 -14220
rect 23900 -14480 24000 -14220
rect 23500 -14500 23620 -14480
rect 23880 -14500 24000 -14480
rect 23500 -14700 24000 -14500
rect 23500 -14720 23620 -14700
rect 23880 -14720 24000 -14700
rect 23500 -14980 23600 -14720
rect 23900 -14980 24000 -14720
rect 23500 -15000 23620 -14980
rect 23880 -15000 24000 -14980
rect 23500 -15200 24000 -15000
rect 23500 -15220 23620 -15200
rect 23880 -15220 24000 -15200
rect 23500 -15480 23600 -15220
rect 23900 -15480 24000 -15220
rect 23500 -15500 23620 -15480
rect 23880 -15500 24000 -15480
rect 23500 -15700 24000 -15500
rect 23500 -15720 23620 -15700
rect 23880 -15720 24000 -15700
rect 23500 -15980 23600 -15720
rect 23900 -15980 24000 -15720
rect 23500 -16000 23620 -15980
rect 23880 -16000 24000 -15980
rect 23500 -16200 24000 -16000
rect 23500 -16220 23620 -16200
rect 23880 -16220 24000 -16200
rect 23500 -16480 23600 -16220
rect 23900 -16480 24000 -16220
rect 23500 -16500 23620 -16480
rect 23880 -16500 24000 -16480
rect 23500 -16700 24000 -16500
rect 23500 -16720 23620 -16700
rect 23880 -16720 24000 -16700
rect 23500 -16980 23600 -16720
rect 23900 -16980 24000 -16720
rect 23500 -17000 23620 -16980
rect 23880 -17000 24000 -16980
rect 23500 -17200 24000 -17000
rect 23500 -17220 23620 -17200
rect 23880 -17220 24000 -17200
rect 23500 -17480 23600 -17220
rect 23900 -17480 24000 -17220
rect 23500 -17500 23620 -17480
rect 23880 -17500 24000 -17480
rect 23500 -17700 24000 -17500
rect 23500 -17720 23620 -17700
rect 23880 -17720 24000 -17700
rect 23500 -17980 23600 -17720
rect 23900 -17980 24000 -17720
rect 23500 -18000 23620 -17980
rect 23880 -18000 24000 -17980
rect 23500 -18200 24000 -18000
rect 23500 -18220 23620 -18200
rect 23880 -18220 24000 -18200
rect 23500 -18480 23600 -18220
rect 23900 -18480 24000 -18220
rect 23500 -18500 23620 -18480
rect 23880 -18500 24000 -18480
rect 23500 -18700 24000 -18500
rect 23500 -18720 23620 -18700
rect 23880 -18720 24000 -18700
rect 23500 -18980 23600 -18720
rect 23900 -18980 24000 -18720
rect 23500 -19000 23620 -18980
rect 23880 -19000 24000 -18980
rect 23500 -19200 24000 -19000
rect 23500 -19220 23620 -19200
rect 23880 -19220 24000 -19200
rect 23500 -19480 23600 -19220
rect 23900 -19480 24000 -19220
rect 23500 -19500 23620 -19480
rect 23880 -19500 24000 -19480
rect 23500 -19700 24000 -19500
rect 23500 -19720 23620 -19700
rect 23880 -19720 24000 -19700
rect 23500 -19980 23600 -19720
rect 23900 -19980 24000 -19720
rect 23500 -20000 23620 -19980
rect 23880 -20000 24000 -19980
rect 23500 -20200 24000 -20000
rect 23500 -20220 23620 -20200
rect 23880 -20220 24000 -20200
rect 23500 -20480 23600 -20220
rect 23900 -20480 24000 -20220
rect 23500 -20500 23620 -20480
rect 23880 -20500 24000 -20480
rect 23500 -20700 24000 -20500
rect 23500 -20720 23620 -20700
rect 23880 -20720 24000 -20700
rect 23500 -20980 23600 -20720
rect 23900 -20980 24000 -20720
rect 23500 -21000 23620 -20980
rect 23880 -21000 24000 -20980
rect 23500 -21200 24000 -21000
rect 23500 -21220 23620 -21200
rect 23880 -21220 24000 -21200
rect 23500 -21480 23600 -21220
rect 23900 -21480 24000 -21220
rect 23500 -21500 23620 -21480
rect 23880 -21500 24000 -21480
rect 23500 -21700 24000 -21500
rect 23500 -21720 23620 -21700
rect 23880 -21720 24000 -21700
rect 23500 -21980 23600 -21720
rect 23900 -21980 24000 -21720
rect 23500 -22000 23620 -21980
rect 23880 -22000 24000 -21980
rect 23500 -22200 24000 -22000
rect 23500 -22220 23620 -22200
rect 23880 -22220 24000 -22200
rect 23500 -22480 23600 -22220
rect 23900 -22480 24000 -22220
rect 23500 -22500 23620 -22480
rect 23880 -22500 24000 -22480
rect 23500 -22700 24000 -22500
rect 23500 -22720 23620 -22700
rect 23880 -22720 24000 -22700
rect 23500 -22980 23600 -22720
rect 23900 -22980 24000 -22720
rect 23500 -23000 23620 -22980
rect 23880 -23000 24000 -22980
rect 23500 -23200 24000 -23000
rect 23500 -23220 23620 -23200
rect 23880 -23220 24000 -23200
rect 23500 -23480 23600 -23220
rect 23900 -23480 24000 -23220
rect 23500 -23500 23620 -23480
rect 23880 -23500 24000 -23480
rect 23500 -23700 24000 -23500
rect 23500 -23720 23620 -23700
rect 23880 -23720 24000 -23700
rect 23500 -23980 23600 -23720
rect 23900 -23980 24000 -23720
rect 23500 -24000 23620 -23980
rect 23880 -24000 24000 -23980
rect -26500 -24200 -17000 -24100
rect -26500 -24220 -26380 -24200
rect -26120 -24220 -25880 -24200
rect -25620 -24220 -25380 -24200
rect -25120 -24220 -24880 -24200
rect -24620 -24220 -24380 -24200
rect -24120 -24220 -23880 -24200
rect -23620 -24220 -23380 -24200
rect -23120 -24220 -22880 -24200
rect -22620 -24220 -22380 -24200
rect -22120 -24220 -21880 -24200
rect -21620 -24220 -21380 -24200
rect -21120 -24220 -20880 -24200
rect -20620 -24220 -20380 -24200
rect -20120 -24220 -19880 -24200
rect -19620 -24220 -19380 -24200
rect -19120 -24220 -18880 -24200
rect -18620 -24220 -18380 -24200
rect -18120 -24220 -17880 -24200
rect -17620 -24220 -17380 -24200
rect -17120 -24220 -17000 -24200
rect -26500 -24480 -26400 -24220
rect -26100 -24480 -25900 -24220
rect -25600 -24480 -25400 -24220
rect -25100 -24480 -24900 -24220
rect -24600 -24480 -24400 -24220
rect -24100 -24480 -23900 -24220
rect -23600 -24480 -23400 -24220
rect -23100 -24480 -22900 -24220
rect -22600 -24480 -22400 -24220
rect -22100 -24480 -21900 -24220
rect -21600 -24480 -21400 -24220
rect -21100 -24480 -20900 -24220
rect -20600 -24480 -20400 -24220
rect -20100 -24480 -19900 -24220
rect -19600 -24480 -19400 -24220
rect -19100 -24480 -18900 -24220
rect -18600 -24480 -18400 -24220
rect -18100 -24480 -17900 -24220
rect -17600 -24480 -17400 -24220
rect -17100 -24480 -17000 -24220
rect -26500 -24500 -26380 -24480
rect -26120 -24500 -25880 -24480
rect -25620 -24500 -25380 -24480
rect -25120 -24500 -24880 -24480
rect -24620 -24500 -24380 -24480
rect -24120 -24500 -23880 -24480
rect -23620 -24500 -23380 -24480
rect -23120 -24500 -22880 -24480
rect -22620 -24500 -22380 -24480
rect -22120 -24500 -21880 -24480
rect -21620 -24500 -21380 -24480
rect -21120 -24500 -20880 -24480
rect -20620 -24500 -20380 -24480
rect -20120 -24500 -19880 -24480
rect -19620 -24500 -19380 -24480
rect -19120 -24500 -18880 -24480
rect -18620 -24500 -18380 -24480
rect -18120 -24500 -17880 -24480
rect -17620 -24500 -17380 -24480
rect -17120 -24500 -17000 -24480
rect -26500 -24600 -17000 -24500
rect 23500 -24200 24000 -24000
rect 23500 -24220 23620 -24200
rect 23880 -24220 24000 -24200
rect 23500 -24480 23600 -24220
rect 23900 -24480 24000 -24220
rect 23500 -24500 23620 -24480
rect 23880 -24500 24000 -24480
rect -26500 -24700 -19000 -24600
rect -26500 -24720 -26380 -24700
rect -26120 -24720 -25880 -24700
rect -25620 -24720 -25380 -24700
rect -25120 -24720 -24880 -24700
rect -24620 -24720 -24380 -24700
rect -24120 -24720 -23880 -24700
rect -23620 -24720 -23380 -24700
rect -23120 -24720 -22880 -24700
rect -22620 -24720 -22380 -24700
rect -22120 -24720 -21880 -24700
rect -21620 -24720 -21380 -24700
rect -21120 -24720 -20880 -24700
rect -20620 -24720 -20380 -24700
rect -20120 -24720 -19880 -24700
rect -19620 -24720 -19380 -24700
rect -19120 -24720 -19000 -24700
rect -26500 -24980 -26400 -24720
rect -26100 -24980 -25900 -24720
rect -25600 -24980 -25400 -24720
rect -25100 -24980 -24900 -24720
rect -24600 -24980 -24400 -24720
rect -24100 -24980 -23900 -24720
rect -23600 -24980 -23400 -24720
rect -23100 -24980 -22900 -24720
rect -22600 -24980 -22400 -24720
rect -22100 -24980 -21900 -24720
rect -21600 -24980 -21400 -24720
rect -21100 -24980 -20900 -24720
rect -20600 -24980 -20400 -24720
rect -20100 -24980 -19900 -24720
rect -19600 -24980 -19400 -24720
rect -19100 -24980 -19000 -24720
rect -26500 -25000 -26380 -24980
rect -26120 -25000 -25880 -24980
rect -25620 -25000 -25380 -24980
rect -25120 -25000 -24880 -24980
rect -24620 -25000 -24380 -24980
rect -24120 -25000 -23880 -24980
rect -23620 -25000 -23380 -24980
rect -23120 -25000 -22880 -24980
rect -22620 -25000 -22380 -24980
rect -22120 -25000 -21880 -24980
rect -21620 -25000 -21380 -24980
rect -21120 -25000 -20880 -24980
rect -20620 -25000 -20380 -24980
rect -20120 -25000 -19880 -24980
rect -19620 -25000 -19380 -24980
rect -19120 -25000 -19000 -24980
rect -26500 -25100 -19000 -25000
rect 23500 -24700 24000 -24500
rect 23500 -24720 23620 -24700
rect 23880 -24720 24000 -24700
rect 23500 -24980 23600 -24720
rect 23900 -24980 24000 -24720
rect 23500 -25000 23620 -24980
rect 23880 -25000 24000 -24980
rect -26500 -25200 -21500 -25100
rect -26500 -25220 -26380 -25200
rect -26120 -25220 -25880 -25200
rect -25620 -25220 -25380 -25200
rect -25120 -25220 -24880 -25200
rect -24620 -25220 -24380 -25200
rect -24120 -25220 -23880 -25200
rect -23620 -25220 -23380 -25200
rect -23120 -25220 -22880 -25200
rect -22620 -25220 -22380 -25200
rect -22120 -25220 -21880 -25200
rect -21620 -25220 -21500 -25200
rect -26500 -25480 -26400 -25220
rect -26100 -25480 -25900 -25220
rect -25600 -25480 -25400 -25220
rect -25100 -25480 -24900 -25220
rect -24600 -25480 -24400 -25220
rect -24100 -25480 -23900 -25220
rect -23600 -25480 -23400 -25220
rect -23100 -25480 -22900 -25220
rect -22600 -25480 -22400 -25220
rect -22100 -25480 -21900 -25220
rect -21600 -25480 -21500 -25220
rect -26500 -25500 -26380 -25480
rect -26120 -25500 -25880 -25480
rect -25620 -25500 -25380 -25480
rect -25120 -25500 -24880 -25480
rect -24620 -25500 -24380 -25480
rect -24120 -25500 -23880 -25480
rect -23620 -25500 -23380 -25480
rect -23120 -25500 -22880 -25480
rect -22620 -25500 -22380 -25480
rect -22120 -25500 -21880 -25480
rect -21620 -25500 -21500 -25480
rect -26500 -25700 -21500 -25500
rect -26500 -25720 -26380 -25700
rect -26120 -25720 -25880 -25700
rect -25620 -25720 -25380 -25700
rect -25120 -25720 -24880 -25700
rect -24620 -25720 -24380 -25700
rect -24120 -25720 -23880 -25700
rect -23620 -25720 -23380 -25700
rect -23120 -25720 -22880 -25700
rect -22620 -25720 -22380 -25700
rect -22120 -25720 -21880 -25700
rect -21620 -25720 -21500 -25700
rect -26500 -25980 -26400 -25720
rect -26100 -25980 -25900 -25720
rect -25600 -25980 -25400 -25720
rect -25100 -25980 -24900 -25720
rect -24600 -25980 -24400 -25720
rect -24100 -25980 -23900 -25720
rect -23600 -25980 -23400 -25720
rect -23100 -25980 -22900 -25720
rect -22600 -25980 -22400 -25720
rect -22100 -25980 -21900 -25720
rect -21600 -25980 -21500 -25720
rect -26500 -26000 -26380 -25980
rect -26120 -26000 -25880 -25980
rect -25620 -26000 -25380 -25980
rect -25120 -26000 -24880 -25980
rect -24620 -26000 -24380 -25980
rect -24120 -26000 -23880 -25980
rect -23620 -26000 -23380 -25980
rect -23120 -26000 -22880 -25980
rect -22620 -26000 -22380 -25980
rect -22120 -26000 -21880 -25980
rect -21620 -26000 -21500 -25980
rect -26500 -26200 -21500 -26000
rect -26500 -26220 -26380 -26200
rect -26120 -26220 -25880 -26200
rect -25620 -26220 -25380 -26200
rect -25120 -26220 -24880 -26200
rect -24620 -26220 -24380 -26200
rect -24120 -26220 -23880 -26200
rect -23620 -26220 -23380 -26200
rect -23120 -26220 -22880 -26200
rect -22620 -26220 -22380 -26200
rect -22120 -26220 -21880 -26200
rect -21620 -26220 -21500 -26200
rect -26500 -26480 -26400 -26220
rect -26100 -26480 -25900 -26220
rect -25600 -26480 -25400 -26220
rect -25100 -26480 -24900 -26220
rect -24600 -26480 -24400 -26220
rect -24100 -26480 -23900 -26220
rect -23600 -26480 -23400 -26220
rect -23100 -26480 -22900 -26220
rect -22600 -26480 -22400 -26220
rect -22100 -26480 -21900 -26220
rect -21600 -26480 -21500 -26220
rect -26500 -26500 -26380 -26480
rect -26120 -26500 -25880 -26480
rect -25620 -26500 -25380 -26480
rect -25120 -26500 -24880 -26480
rect -24620 -26500 -24380 -26480
rect -24120 -26500 -23880 -26480
rect -23620 -26500 -23380 -26480
rect -23120 -26500 -22880 -26480
rect -22620 -26500 -22380 -26480
rect -22120 -26500 -21880 -26480
rect -21620 -26500 -21500 -26480
rect -26500 -26700 -21500 -26500
rect -26500 -26720 -26380 -26700
rect -26120 -26720 -25880 -26700
rect -25620 -26720 -25380 -26700
rect -25120 -26720 -24880 -26700
rect -24620 -26720 -24380 -26700
rect -24120 -26720 -23880 -26700
rect -23620 -26720 -23380 -26700
rect -23120 -26720 -22880 -26700
rect -22620 -26720 -22380 -26700
rect -22120 -26720 -21880 -26700
rect -21620 -26720 -21500 -26700
rect -26500 -26980 -26400 -26720
rect -26100 -26980 -25900 -26720
rect -25600 -26980 -25400 -26720
rect -25100 -26980 -24900 -26720
rect -24600 -26980 -24400 -26720
rect -24100 -26980 -23900 -26720
rect -23600 -26980 -23400 -26720
rect -23100 -26980 -22900 -26720
rect -22600 -26980 -22400 -26720
rect -22100 -26980 -21900 -26720
rect -21600 -26980 -21500 -26720
rect -26500 -27000 -26380 -26980
rect -26120 -27000 -25880 -26980
rect -25620 -27000 -25380 -26980
rect -25120 -27000 -24880 -26980
rect -24620 -27000 -24380 -26980
rect -24120 -27000 -23880 -26980
rect -23620 -27000 -23380 -26980
rect -23120 -27000 -22880 -26980
rect -22620 -27000 -22380 -26980
rect -22120 -27000 -21880 -26980
rect -21620 -27000 -21500 -26980
rect -26500 -27200 -21500 -27000
rect -26500 -27220 -26380 -27200
rect -26120 -27220 -25880 -27200
rect -25620 -27220 -25380 -27200
rect -25120 -27220 -24880 -27200
rect -24620 -27220 -24380 -27200
rect -24120 -27220 -23880 -27200
rect -23620 -27220 -23380 -27200
rect -23120 -27220 -22880 -27200
rect -22620 -27220 -22380 -27200
rect -22120 -27220 -21880 -27200
rect -21620 -27220 -21500 -27200
rect -26500 -27480 -26400 -27220
rect -26100 -27480 -25900 -27220
rect -25600 -27480 -25400 -27220
rect -25100 -27480 -24900 -27220
rect -24600 -27480 -24400 -27220
rect -24100 -27480 -23900 -27220
rect -23600 -27480 -23400 -27220
rect -23100 -27480 -22900 -27220
rect -22600 -27480 -22400 -27220
rect -22100 -27480 -21900 -27220
rect -21600 -27480 -21500 -27220
rect -26500 -27500 -26380 -27480
rect -26120 -27500 -25880 -27480
rect -25620 -27500 -25380 -27480
rect -25120 -27500 -24880 -27480
rect -24620 -27500 -24380 -27480
rect -24120 -27500 -23880 -27480
rect -23620 -27500 -23380 -27480
rect -23120 -27500 -22880 -27480
rect -22620 -27500 -22380 -27480
rect -22120 -27500 -21880 -27480
rect -21620 -27500 -21500 -27480
rect -26500 -27700 -21500 -27500
rect -26500 -27720 -26380 -27700
rect -26120 -27720 -25880 -27700
rect -25620 -27720 -25380 -27700
rect -25120 -27720 -24880 -27700
rect -24620 -27720 -24380 -27700
rect -24120 -27720 -23880 -27700
rect -23620 -27720 -23380 -27700
rect -23120 -27720 -22880 -27700
rect -22620 -27720 -22380 -27700
rect -22120 -27720 -21880 -27700
rect -21620 -27720 -21500 -27700
rect -26500 -27980 -26400 -27720
rect -26100 -27980 -25900 -27720
rect -25600 -27980 -25400 -27720
rect -25100 -27980 -24900 -27720
rect -24600 -27980 -24400 -27720
rect -24100 -27980 -23900 -27720
rect -23600 -27980 -23400 -27720
rect -23100 -27980 -22900 -27720
rect -22600 -27980 -22400 -27720
rect -22100 -27980 -21900 -27720
rect -21600 -27980 -21500 -27720
rect -26500 -28000 -26380 -27980
rect -26120 -28000 -25880 -27980
rect -25620 -28000 -25380 -27980
rect -25120 -28000 -24880 -27980
rect -24620 -28000 -24380 -27980
rect -24120 -28000 -23880 -27980
rect -23620 -28000 -23380 -27980
rect -23120 -28000 -22880 -27980
rect -22620 -28000 -22380 -27980
rect -22120 -28000 -21880 -27980
rect -21620 -28000 -21500 -27980
rect -26500 -28200 -21500 -28000
rect -26500 -28220 -26380 -28200
rect -26120 -28220 -25880 -28200
rect -25620 -28220 -25380 -28200
rect -25120 -28220 -24880 -28200
rect -24620 -28220 -24380 -28200
rect -24120 -28220 -23880 -28200
rect -23620 -28220 -23380 -28200
rect -23120 -28220 -22880 -28200
rect -22620 -28220 -22380 -28200
rect -22120 -28220 -21880 -28200
rect -21620 -28220 -21500 -28200
rect -26500 -28480 -26400 -28220
rect -26100 -28480 -25900 -28220
rect -25600 -28480 -25400 -28220
rect -25100 -28480 -24900 -28220
rect -24600 -28480 -24400 -28220
rect -24100 -28480 -23900 -28220
rect -23600 -28480 -23400 -28220
rect -23100 -28480 -22900 -28220
rect -22600 -28480 -22400 -28220
rect -22100 -28480 -21900 -28220
rect -21600 -28480 -21500 -28220
rect -26500 -28500 -26380 -28480
rect -26120 -28500 -25880 -28480
rect -25620 -28500 -25380 -28480
rect -25120 -28500 -24880 -28480
rect -24620 -28500 -24380 -28480
rect -24120 -28500 -23880 -28480
rect -23620 -28500 -23380 -28480
rect -23120 -28500 -22880 -28480
rect -22620 -28500 -22380 -28480
rect -22120 -28500 -21880 -28480
rect -21620 -28500 -21500 -28480
rect -26500 -28700 -21500 -28500
rect -26500 -28720 -26380 -28700
rect -26120 -28720 -25880 -28700
rect -25620 -28720 -25380 -28700
rect -25120 -28720 -24880 -28700
rect -24620 -28720 -24380 -28700
rect -24120 -28720 -23880 -28700
rect -23620 -28720 -23380 -28700
rect -23120 -28720 -22880 -28700
rect -22620 -28720 -22380 -28700
rect -22120 -28720 -21880 -28700
rect -21620 -28720 -21500 -28700
rect -26500 -28980 -26400 -28720
rect -26100 -28980 -25900 -28720
rect -25600 -28980 -25400 -28720
rect -25100 -28980 -24900 -28720
rect -24600 -28980 -24400 -28720
rect -24100 -28980 -23900 -28720
rect -23600 -28980 -23400 -28720
rect -23100 -28980 -22900 -28720
rect -22600 -28980 -22400 -28720
rect -22100 -28980 -21900 -28720
rect -21600 -28980 -21500 -28720
rect -26500 -29000 -26380 -28980
rect -26120 -29000 -25880 -28980
rect -25620 -29000 -25380 -28980
rect -25120 -29000 -24880 -28980
rect -24620 -29000 -24380 -28980
rect -24120 -29000 -23880 -28980
rect -23620 -29000 -23380 -28980
rect -23120 -29000 -22880 -28980
rect -22620 -29000 -22380 -28980
rect -22120 -29000 -21880 -28980
rect -21620 -29000 -21500 -28980
rect -26500 -29200 -21500 -29000
rect -26500 -29220 -26380 -29200
rect -26120 -29220 -25880 -29200
rect -25620 -29220 -25380 -29200
rect -25120 -29220 -24880 -29200
rect -24620 -29220 -24380 -29200
rect -24120 -29220 -23880 -29200
rect -23620 -29220 -23380 -29200
rect -23120 -29220 -22880 -29200
rect -22620 -29220 -22380 -29200
rect -22120 -29220 -21880 -29200
rect -21620 -29220 -21500 -29200
rect -26500 -29480 -26400 -29220
rect -26100 -29480 -25900 -29220
rect -25600 -29480 -25400 -29220
rect -25100 -29480 -24900 -29220
rect -24600 -29480 -24400 -29220
rect -24100 -29480 -23900 -29220
rect -23600 -29480 -23400 -29220
rect -23100 -29480 -22900 -29220
rect -22600 -29480 -22400 -29220
rect -22100 -29480 -21900 -29220
rect -21600 -29480 -21500 -29220
rect -26500 -29500 -26380 -29480
rect -26120 -29500 -25880 -29480
rect -25620 -29500 -25380 -29480
rect -25120 -29500 -24880 -29480
rect -24620 -29500 -24380 -29480
rect -24120 -29500 -23880 -29480
rect -23620 -29500 -23380 -29480
rect -23120 -29500 -22880 -29480
rect -22620 -29500 -22380 -29480
rect -22120 -29500 -21880 -29480
rect -21620 -29500 -21500 -29480
rect -26500 -29600 -21500 -29500
rect 23500 -25200 24000 -25000
rect 23500 -25220 23620 -25200
rect 23880 -25220 24000 -25200
rect 23500 -25480 23600 -25220
rect 23900 -25480 24000 -25220
rect 23500 -25500 23620 -25480
rect 23880 -25500 24000 -25480
rect 23500 -25700 24000 -25500
rect 23500 -25720 23620 -25700
rect 23880 -25720 24000 -25700
rect 23500 -25980 23600 -25720
rect 23900 -25980 24000 -25720
rect 23500 -26000 23620 -25980
rect 23880 -26000 24000 -25980
rect 23500 -26200 24000 -26000
rect 23500 -26220 23620 -26200
rect 23880 -26220 24000 -26200
rect 23500 -26480 23600 -26220
rect 23900 -26480 24000 -26220
rect 23500 -26500 23620 -26480
rect 23880 -26500 24000 -26480
rect 23500 -26700 24000 -26500
rect 23500 -26720 23620 -26700
rect 23880 -26720 24000 -26700
rect 23500 -26980 23600 -26720
rect 23900 -26980 24000 -26720
rect 23500 -27000 23620 -26980
rect 23880 -27000 24000 -26980
rect 23500 -27200 24000 -27000
rect 23500 -27220 23620 -27200
rect 23880 -27220 24000 -27200
rect 23500 -27480 23600 -27220
rect 23900 -27480 24000 -27220
rect 23500 -27500 23620 -27480
rect 23880 -27500 24000 -27480
rect 23500 -27700 24000 -27500
rect 23500 -27720 23620 -27700
rect 23880 -27720 24000 -27700
rect 23500 -27980 23600 -27720
rect 23900 -27980 24000 -27720
rect 23500 -28000 23620 -27980
rect 23880 -28000 24000 -27980
rect 23500 -28200 24000 -28000
rect 23500 -28220 23620 -28200
rect 23880 -28220 24000 -28200
rect 23500 -28480 23600 -28220
rect 23900 -28480 24000 -28220
rect 23500 -28500 23620 -28480
rect 23880 -28500 24000 -28480
rect 23500 -28700 24000 -28500
rect 23500 -28720 23620 -28700
rect 23880 -28720 24000 -28700
rect 23500 -28980 23600 -28720
rect 23900 -28980 24000 -28720
rect 23500 -29000 23620 -28980
rect 23880 -29000 24000 -28980
rect 23500 -29200 24000 -29000
rect 23500 -29220 23620 -29200
rect 23880 -29220 24000 -29200
rect 23500 -29480 23600 -29220
rect 23900 -29480 24000 -29220
rect 23500 -29500 23620 -29480
rect 23880 -29500 24000 -29480
rect 23500 -29700 24000 -29500
rect 23500 -29720 23620 -29700
rect 23880 -29720 24000 -29700
rect 23500 -29980 23600 -29720
rect 23900 -29980 24000 -29720
rect 23500 -30000 23620 -29980
rect 23880 -30000 24000 -29980
rect 23500 -30200 24000 -30000
rect 23500 -30220 23620 -30200
rect 23880 -30220 24000 -30200
rect 23500 -30480 23600 -30220
rect 23900 -30480 24000 -30220
rect 23500 -30500 23620 -30480
rect 23880 -30500 24000 -30480
rect 23500 -30700 24000 -30500
rect 23500 -30720 23620 -30700
rect 23880 -30720 24000 -30700
rect 23500 -30980 23600 -30720
rect 23900 -30980 24000 -30720
rect 23500 -31000 23620 -30980
rect 23880 -31000 24000 -30980
rect 23500 -31200 24000 -31000
rect 23500 -31220 23620 -31200
rect 23880 -31220 24000 -31200
rect 23500 -31480 23600 -31220
rect 23900 -31480 24000 -31220
rect 23500 -31500 23620 -31480
rect 23880 -31500 24000 -31480
rect 23500 -31700 24000 -31500
rect 23500 -31720 23620 -31700
rect 23880 -31720 24000 -31700
rect 23500 -31980 23600 -31720
rect 23900 -31980 24000 -31720
rect 23500 -32000 23620 -31980
rect 23880 -32000 24000 -31980
rect 23500 -32200 24000 -32000
rect 23500 -32220 23620 -32200
rect 23880 -32220 24000 -32200
rect 23500 -32480 23600 -32220
rect 23900 -32480 24000 -32220
rect 23500 -32500 23620 -32480
rect 23880 -32500 24000 -32480
rect 23500 -32700 24000 -32500
rect 23500 -32720 23620 -32700
rect 23880 -32720 24000 -32700
rect 23500 -32980 23600 -32720
rect 23900 -32980 24000 -32720
rect 23500 -33000 23620 -32980
rect 23880 -33000 24000 -32980
rect 23500 -33200 24000 -33000
rect 23500 -33220 23620 -33200
rect 23880 -33220 24000 -33200
rect 23500 -33480 23600 -33220
rect 23900 -33480 24000 -33220
rect 23500 -33500 23620 -33480
rect 23880 -33500 24000 -33480
rect 23500 -33600 24000 -33500
rect 32800 -5700 33500 -5600
rect 32800 -5720 33120 -5700
rect 33380 -5720 33500 -5700
rect 32800 -5980 33100 -5720
rect 33400 -5980 33500 -5720
rect 32800 -6000 33120 -5980
rect 33380 -6000 33500 -5980
rect 32800 -6200 33500 -6000
rect 32800 -6220 33120 -6200
rect 33380 -6220 33500 -6200
rect 32800 -6480 33100 -6220
rect 33400 -6480 33500 -6220
rect 32800 -6500 33120 -6480
rect 33380 -6500 33500 -6480
rect 32800 -6700 33500 -6500
rect 32800 -6720 33120 -6700
rect 33380 -6720 33500 -6700
rect 32800 -6980 33100 -6720
rect 33400 -6980 33500 -6720
rect 32800 -7000 33120 -6980
rect 33380 -7000 33500 -6980
rect 32800 -7200 33500 -7000
rect 32800 -7220 33120 -7200
rect 33380 -7220 33500 -7200
rect 32800 -7480 33100 -7220
rect 33400 -7480 33500 -7220
rect 32800 -7500 33120 -7480
rect 33380 -7500 33500 -7480
rect 32800 -7700 33500 -7500
rect 32800 -7720 33120 -7700
rect 33380 -7720 33500 -7700
rect 32800 -7980 33100 -7720
rect 33400 -7980 33500 -7720
rect 32800 -8000 33120 -7980
rect 33380 -8000 33500 -7980
rect 32800 -8200 33500 -8000
rect 32800 -8220 33120 -8200
rect 33380 -8220 33500 -8200
rect 32800 -8480 33100 -8220
rect 33400 -8480 33500 -8220
rect 32800 -8500 33120 -8480
rect 33380 -8500 33500 -8480
rect 32800 -8700 33500 -8500
rect 32800 -8720 33120 -8700
rect 33380 -8720 33500 -8700
rect 32800 -8980 33100 -8720
rect 33400 -8980 33500 -8720
rect 32800 -9000 33120 -8980
rect 33380 -9000 33500 -8980
rect 32800 -9200 33500 -9000
rect 32800 -9220 33120 -9200
rect 33380 -9220 33500 -9200
rect 32800 -9480 33100 -9220
rect 33400 -9480 33500 -9220
rect 32800 -9500 33120 -9480
rect 33380 -9500 33500 -9480
rect 32800 -9700 33500 -9500
rect 32800 -9720 33120 -9700
rect 33380 -9720 33500 -9700
rect 32800 -9980 33100 -9720
rect 33400 -9980 33500 -9720
rect 32800 -10000 33120 -9980
rect 33380 -10000 33500 -9980
rect 32800 -10200 33500 -10000
rect 32800 -10220 33120 -10200
rect 33380 -10220 33500 -10200
rect 32800 -10480 33100 -10220
rect 33400 -10480 33500 -10220
rect 32800 -10500 33120 -10480
rect 33380 -10500 33500 -10480
rect 32800 -10700 33500 -10500
rect 32800 -10720 33120 -10700
rect 33380 -10720 33500 -10700
rect 32800 -10980 33100 -10720
rect 33400 -10980 33500 -10720
rect 32800 -11000 33120 -10980
rect 33380 -11000 33500 -10980
rect 32800 -11200 33500 -11000
rect 32800 -11220 33120 -11200
rect 33380 -11220 33500 -11200
rect 32800 -11480 33100 -11220
rect 33400 -11480 33500 -11220
rect 32800 -11500 33120 -11480
rect 33380 -11500 33500 -11480
rect 32800 -11700 33500 -11500
rect 32800 -11720 33120 -11700
rect 33380 -11720 33500 -11700
rect 32800 -11980 33100 -11720
rect 33400 -11980 33500 -11720
rect 32800 -12000 33120 -11980
rect 33380 -12000 33500 -11980
rect 32800 -12200 33500 -12000
rect 32800 -12220 33120 -12200
rect 33380 -12220 33500 -12200
rect 32800 -12480 33100 -12220
rect 33400 -12480 33500 -12220
rect 32800 -12500 33120 -12480
rect 33380 -12500 33500 -12480
rect 32800 -12700 33500 -12500
rect 32800 -12720 33120 -12700
rect 33380 -12720 33500 -12700
rect 32800 -12980 33100 -12720
rect 33400 -12980 33500 -12720
rect 32800 -13000 33120 -12980
rect 33380 -13000 33500 -12980
rect 32800 -13200 33500 -13000
rect 32800 -13220 33120 -13200
rect 33380 -13220 33500 -13200
rect 32800 -13480 33100 -13220
rect 33400 -13480 33500 -13220
rect 32800 -13500 33120 -13480
rect 33380 -13500 33500 -13480
rect 32800 -13700 33500 -13500
rect 32800 -13720 33120 -13700
rect 33380 -13720 33500 -13700
rect 32800 -13980 33100 -13720
rect 33400 -13980 33500 -13720
rect 32800 -14000 33120 -13980
rect 33380 -14000 33500 -13980
rect 32800 -14200 33500 -14000
rect 32800 -14220 33120 -14200
rect 33380 -14220 33500 -14200
rect 32800 -14480 33100 -14220
rect 33400 -14480 33500 -14220
rect 32800 -14500 33120 -14480
rect 33380 -14500 33500 -14480
rect 32800 -14700 33500 -14500
rect 32800 -14720 33120 -14700
rect 33380 -14720 33500 -14700
rect 32800 -14980 33100 -14720
rect 33400 -14980 33500 -14720
rect 32800 -15000 33120 -14980
rect 33380 -15000 33500 -14980
rect 32800 -15200 33500 -15000
rect 32800 -15220 33120 -15200
rect 33380 -15220 33500 -15200
rect 32800 -15480 33100 -15220
rect 33400 -15480 33500 -15220
rect 32800 -15500 33120 -15480
rect 33380 -15500 33500 -15480
rect 32800 -15700 33500 -15500
rect 32800 -15720 33120 -15700
rect 33380 -15720 33500 -15700
rect 32800 -15980 33100 -15720
rect 33400 -15980 33500 -15720
rect 32800 -16000 33120 -15980
rect 33380 -16000 33500 -15980
rect 32800 -16200 33500 -16000
rect 32800 -16220 33120 -16200
rect 33380 -16220 33500 -16200
rect 32800 -16480 33100 -16220
rect 33400 -16480 33500 -16220
rect 32800 -16500 33120 -16480
rect 33380 -16500 33500 -16480
rect 32800 -16700 33500 -16500
rect 32800 -16720 33120 -16700
rect 33380 -16720 33500 -16700
rect 32800 -16980 33100 -16720
rect 33400 -16980 33500 -16720
rect 32800 -17000 33120 -16980
rect 33380 -17000 33500 -16980
rect 32800 -17200 33500 -17000
rect 32800 -17220 33120 -17200
rect 33380 -17220 33500 -17200
rect 32800 -17480 33100 -17220
rect 33400 -17480 33500 -17220
rect 32800 -17500 33120 -17480
rect 33380 -17500 33500 -17480
rect 32800 -17700 33500 -17500
rect 32800 -17720 33120 -17700
rect 33380 -17720 33500 -17700
rect 32800 -17980 33100 -17720
rect 33400 -17980 33500 -17720
rect 32800 -18000 33120 -17980
rect 33380 -18000 33500 -17980
rect 32800 -18200 33500 -18000
rect 32800 -18220 33120 -18200
rect 33380 -18220 33500 -18200
rect 32800 -18480 33100 -18220
rect 33400 -18480 33500 -18220
rect 32800 -18500 33120 -18480
rect 33380 -18500 33500 -18480
rect 32800 -18700 33500 -18500
rect 32800 -18720 33120 -18700
rect 33380 -18720 33500 -18700
rect 32800 -18980 33100 -18720
rect 33400 -18980 33500 -18720
rect 32800 -19000 33120 -18980
rect 33380 -19000 33500 -18980
rect 32800 -19200 33500 -19000
rect 32800 -19220 33120 -19200
rect 33380 -19220 33500 -19200
rect 32800 -19480 33100 -19220
rect 33400 -19480 33500 -19220
rect 32800 -19500 33120 -19480
rect 33380 -19500 33500 -19480
rect 32800 -19700 33500 -19500
rect 32800 -19720 33120 -19700
rect 33380 -19720 33500 -19700
rect 32800 -19980 33100 -19720
rect 33400 -19980 33500 -19720
rect 32800 -20000 33120 -19980
rect 33380 -20000 33500 -19980
rect 32800 -20100 33500 -20000
rect 32800 -20200 34500 -20100
rect 32800 -20220 33120 -20200
rect 33380 -20220 33620 -20200
rect 33880 -20220 34120 -20200
rect 34380 -20220 34500 -20200
rect 32800 -20480 33100 -20220
rect 33400 -20480 33600 -20220
rect 33900 -20480 34100 -20220
rect 34400 -20480 34500 -20220
rect 32800 -20500 33120 -20480
rect 33380 -20500 33620 -20480
rect 33880 -20500 34120 -20480
rect 34380 -20500 34500 -20480
rect 32800 -20700 34500 -20500
rect 32800 -20720 33120 -20700
rect 33380 -20720 33620 -20700
rect 33880 -20720 34120 -20700
rect 34380 -20720 34500 -20700
rect 32800 -20980 33100 -20720
rect 33400 -20980 33600 -20720
rect 33900 -20980 34100 -20720
rect 34400 -20980 34500 -20720
rect 32800 -21000 33120 -20980
rect 33380 -21000 33620 -20980
rect 33880 -21000 34120 -20980
rect 34380 -21000 34500 -20980
rect 32800 -21200 34500 -21000
rect 32800 -21220 33120 -21200
rect 33380 -21220 33620 -21200
rect 33880 -21220 34120 -21200
rect 34380 -21220 34500 -21200
rect 32800 -21480 33100 -21220
rect 33400 -21480 33600 -21220
rect 33900 -21480 34100 -21220
rect 34400 -21480 34500 -21220
rect 32800 -21500 33120 -21480
rect 33380 -21500 33620 -21480
rect 33880 -21500 34120 -21480
rect 34380 -21500 34500 -21480
rect 32800 -21700 34500 -21500
rect 32800 -21720 33120 -21700
rect 33380 -21720 33620 -21700
rect 33880 -21720 34120 -21700
rect 34380 -21720 34500 -21700
rect 32800 -21980 33100 -21720
rect 33400 -21980 33600 -21720
rect 33900 -21980 34100 -21720
rect 34400 -21980 34500 -21720
rect 32800 -22000 33120 -21980
rect 33380 -22000 33620 -21980
rect 33880 -22000 34120 -21980
rect 34380 -22000 34500 -21980
rect 32800 -22200 34500 -22000
rect 32800 -22220 33120 -22200
rect 33380 -22220 33620 -22200
rect 33880 -22220 34120 -22200
rect 34380 -22220 34500 -22200
rect 32800 -22480 33100 -22220
rect 33400 -22480 33600 -22220
rect 33900 -22480 34100 -22220
rect 34400 -22480 34500 -22220
rect 32800 -22500 33120 -22480
rect 33380 -22500 33620 -22480
rect 33880 -22500 34120 -22480
rect 34380 -22500 34500 -22480
rect 32800 -22700 34500 -22500
rect 32800 -22720 33120 -22700
rect 33380 -22720 33620 -22700
rect 33880 -22720 34120 -22700
rect 34380 -22720 34500 -22700
rect 32800 -22980 33100 -22720
rect 33400 -22980 33600 -22720
rect 33900 -22980 34100 -22720
rect 34400 -22980 34500 -22720
rect 32800 -23000 33120 -22980
rect 33380 -23000 33620 -22980
rect 33880 -23000 34120 -22980
rect 34380 -23000 34500 -22980
rect 32800 -23200 34500 -23000
rect 32800 -23220 33120 -23200
rect 33380 -23220 33620 -23200
rect 33880 -23220 34120 -23200
rect 34380 -23220 34500 -23200
rect 32800 -23480 33100 -23220
rect 33400 -23480 33600 -23220
rect 33900 -23480 34100 -23220
rect 34400 -23480 34500 -23220
rect 32800 -23500 33120 -23480
rect 33380 -23500 33620 -23480
rect 33880 -23500 34120 -23480
rect 34380 -23500 34500 -23480
rect 32800 -23700 34500 -23500
rect 32800 -23720 33120 -23700
rect 33380 -23720 33620 -23700
rect 33880 -23720 34120 -23700
rect 34380 -23720 34500 -23700
rect 32800 -23980 33100 -23720
rect 33400 -23980 33600 -23720
rect 33900 -23980 34100 -23720
rect 34400 -23980 34500 -23720
rect 32800 -24000 33120 -23980
rect 33380 -24000 33620 -23980
rect 33880 -24000 34120 -23980
rect 34380 -24000 34500 -23980
rect 32800 -24200 34500 -24000
rect 32800 -24220 33120 -24200
rect 33380 -24220 33620 -24200
rect 33880 -24220 34120 -24200
rect 34380 -24220 34500 -24200
rect 32800 -24480 33100 -24220
rect 33400 -24480 33600 -24220
rect 33900 -24480 34100 -24220
rect 34400 -24480 34500 -24220
rect 32800 -24500 33120 -24480
rect 33380 -24500 33620 -24480
rect 33880 -24500 34120 -24480
rect 34380 -24500 34500 -24480
rect 32800 -24700 34500 -24500
rect 32800 -24720 33120 -24700
rect 33380 -24720 33620 -24700
rect 33880 -24720 34120 -24700
rect 34380 -24720 34500 -24700
rect 32800 -24980 33100 -24720
rect 33400 -24980 33600 -24720
rect 33900 -24980 34100 -24720
rect 34400 -24980 34500 -24720
rect 32800 -25000 33120 -24980
rect 33380 -25000 33620 -24980
rect 33880 -25000 34120 -24980
rect 34380 -25000 34500 -24980
rect 32800 -25200 34500 -25000
rect 32800 -25220 33120 -25200
rect 33380 -25220 33620 -25200
rect 33880 -25220 34120 -25200
rect 34380 -25220 34500 -25200
rect 32800 -25480 33100 -25220
rect 33400 -25480 33600 -25220
rect 33900 -25480 34100 -25220
rect 34400 -25480 34500 -25220
rect 32800 -25500 33120 -25480
rect 33380 -25500 33620 -25480
rect 33880 -25500 34120 -25480
rect 34380 -25500 34500 -25480
rect 32800 -25700 34500 -25500
rect 32800 -25720 33120 -25700
rect 33380 -25720 33620 -25700
rect 33880 -25720 34120 -25700
rect 34380 -25720 34500 -25700
rect 32800 -25980 33100 -25720
rect 33400 -25980 33600 -25720
rect 33900 -25980 34100 -25720
rect 34400 -25980 34500 -25720
rect 32800 -26000 33120 -25980
rect 33380 -26000 33620 -25980
rect 33880 -26000 34120 -25980
rect 34380 -26000 34500 -25980
rect 32800 -26200 34500 -26000
rect 32800 -26220 33120 -26200
rect 33380 -26220 33620 -26200
rect 33880 -26220 34120 -26200
rect 34380 -26220 34500 -26200
rect 32800 -26480 33100 -26220
rect 33400 -26480 33600 -26220
rect 33900 -26480 34100 -26220
rect 34400 -26480 34500 -26220
rect 32800 -26500 33120 -26480
rect 33380 -26500 33620 -26480
rect 33880 -26500 34120 -26480
rect 34380 -26500 34500 -26480
rect 32800 -26700 34500 -26500
rect 32800 -26720 33120 -26700
rect 33380 -26720 33620 -26700
rect 33880 -26720 34120 -26700
rect 34380 -26720 34500 -26700
rect 32800 -26980 33100 -26720
rect 33400 -26980 33600 -26720
rect 33900 -26980 34100 -26720
rect 34400 -26980 34500 -26720
rect 32800 -27000 33120 -26980
rect 33380 -27000 33620 -26980
rect 33880 -27000 34120 -26980
rect 34380 -27000 34500 -26980
rect 32800 -27200 34500 -27000
rect 32800 -27220 33120 -27200
rect 33380 -27220 33620 -27200
rect 33880 -27220 34120 -27200
rect 34380 -27220 34500 -27200
rect 32800 -27480 33100 -27220
rect 33400 -27480 33600 -27220
rect 33900 -27480 34100 -27220
rect 34400 -27480 34500 -27220
rect 32800 -27500 33120 -27480
rect 33380 -27500 33620 -27480
rect 33880 -27500 34120 -27480
rect 34380 -27500 34500 -27480
rect 32800 -27700 34500 -27500
rect 32800 -27720 33120 -27700
rect 33380 -27720 33620 -27700
rect 33880 -27720 34120 -27700
rect 34380 -27720 34500 -27700
rect 32800 -27980 33100 -27720
rect 33400 -27980 33600 -27720
rect 33900 -27980 34100 -27720
rect 34400 -27980 34500 -27720
rect 32800 -28000 33120 -27980
rect 33380 -28000 33620 -27980
rect 33880 -28000 34120 -27980
rect 34380 -28000 34500 -27980
rect 32800 -28200 34500 -28000
rect 32800 -28220 33120 -28200
rect 33380 -28220 33620 -28200
rect 33880 -28220 34120 -28200
rect 34380 -28220 34500 -28200
rect 32800 -28480 33100 -28220
rect 33400 -28480 33600 -28220
rect 33900 -28480 34100 -28220
rect 34400 -28480 34500 -28220
rect 32800 -28500 33120 -28480
rect 33380 -28500 33620 -28480
rect 33880 -28500 34120 -28480
rect 34380 -28500 34500 -28480
rect 32800 -28700 34500 -28500
rect 32800 -28720 33120 -28700
rect 33380 -28720 33620 -28700
rect 33880 -28720 34120 -28700
rect 34380 -28720 34500 -28700
rect 32800 -28980 33100 -28720
rect 33400 -28980 33600 -28720
rect 33900 -28980 34100 -28720
rect 34400 -28980 34500 -28720
rect 32800 -29000 33120 -28980
rect 33380 -29000 33620 -28980
rect 33880 -29000 34120 -28980
rect 34380 -29000 34500 -28980
rect 32800 -29200 34500 -29000
rect 32800 -29220 33120 -29200
rect 33380 -29220 33620 -29200
rect 33880 -29220 34120 -29200
rect 34380 -29220 34500 -29200
rect 32800 -29480 33100 -29220
rect 33400 -29480 33600 -29220
rect 33900 -29480 34100 -29220
rect 34400 -29480 34500 -29220
rect 32800 -29500 33120 -29480
rect 33380 -29500 33620 -29480
rect 33880 -29500 34120 -29480
rect 34380 -29500 34500 -29480
rect 32800 -29700 34500 -29500
rect 32800 -29720 33120 -29700
rect 33380 -29720 33620 -29700
rect 33880 -29720 34120 -29700
rect 34380 -29720 34500 -29700
rect 32800 -29980 33100 -29720
rect 33400 -29980 33600 -29720
rect 33900 -29980 34100 -29720
rect 34400 -29980 34500 -29720
rect 32800 -30000 33120 -29980
rect 33380 -30000 33620 -29980
rect 33880 -30000 34120 -29980
rect 34380 -30000 34500 -29980
rect 32800 -30200 34500 -30000
rect 32800 -30220 33120 -30200
rect 33380 -30220 33620 -30200
rect 33880 -30220 34120 -30200
rect 34380 -30220 34500 -30200
rect 32800 -30480 33100 -30220
rect 33400 -30480 33600 -30220
rect 33900 -30480 34100 -30220
rect 34400 -30480 34500 -30220
rect 32800 -30500 33120 -30480
rect 33380 -30500 33620 -30480
rect 33880 -30500 34120 -30480
rect 34380 -30500 34500 -30480
rect 32800 -30700 34500 -30500
rect 32800 -30720 33120 -30700
rect 33380 -30720 33620 -30700
rect 33880 -30720 34120 -30700
rect 34380 -30720 34500 -30700
rect 32800 -30980 33100 -30720
rect 33400 -30980 33600 -30720
rect 33900 -30980 34100 -30720
rect 34400 -30980 34500 -30720
rect 32800 -31000 33120 -30980
rect 33380 -31000 33620 -30980
rect 33880 -31000 34120 -30980
rect 34380 -31000 34500 -30980
rect 32800 -31200 34500 -31000
rect 32800 -31220 33120 -31200
rect 33380 -31220 33620 -31200
rect 33880 -31220 34120 -31200
rect 34380 -31220 34500 -31200
rect 32800 -31480 33100 -31220
rect 33400 -31480 33600 -31220
rect 33900 -31480 34100 -31220
rect 34400 -31480 34500 -31220
rect 32800 -31500 33120 -31480
rect 33380 -31500 33620 -31480
rect 33880 -31500 34120 -31480
rect 34380 -31500 34500 -31480
rect 32800 -31700 34500 -31500
rect 32800 -31720 33120 -31700
rect 33380 -31720 33620 -31700
rect 33880 -31720 34120 -31700
rect 34380 -31720 34500 -31700
rect 32800 -31980 33100 -31720
rect 33400 -31980 33600 -31720
rect 33900 -31980 34100 -31720
rect 34400 -31980 34500 -31720
rect 32800 -32000 33120 -31980
rect 33380 -32000 33620 -31980
rect 33880 -32000 34120 -31980
rect 34380 -32000 34500 -31980
rect 32800 -32200 34500 -32000
rect 32800 -32220 33120 -32200
rect 33380 -32220 33620 -32200
rect 33880 -32220 34120 -32200
rect 34380 -32220 34500 -32200
rect 32800 -32480 33100 -32220
rect 33400 -32480 33600 -32220
rect 33900 -32480 34100 -32220
rect 34400 -32480 34500 -32220
rect 32800 -32500 33120 -32480
rect 33380 -32500 33620 -32480
rect 33880 -32500 34120 -32480
rect 34380 -32500 34500 -32480
rect 32800 -32700 34500 -32500
rect 32800 -32720 33120 -32700
rect 33380 -32720 33620 -32700
rect 33880 -32720 34120 -32700
rect 34380 -32720 34500 -32700
rect 32800 -32980 33100 -32720
rect 33400 -32980 33600 -32720
rect 33900 -32980 34100 -32720
rect 34400 -32980 34500 -32720
rect 32800 -33000 33120 -32980
rect 33380 -33000 33620 -32980
rect 33880 -33000 34120 -32980
rect 34380 -33000 34500 -32980
rect 32800 -33200 34500 -33000
rect 32800 -33220 33120 -33200
rect 33380 -33220 33620 -33200
rect 33880 -33220 34120 -33200
rect 34380 -33220 34500 -33200
rect 32800 -33480 33100 -33220
rect 33400 -33480 33600 -33220
rect 33900 -33480 34100 -33220
rect 34400 -33480 34500 -33220
rect 32800 -33500 33120 -33480
rect 33380 -33500 33620 -33480
rect 33880 -33500 34120 -33480
rect 34380 -33500 34500 -33480
rect 32800 -33600 34500 -33500
<< metal2 >>
rect 16000 13700 20000 13900
rect 13400 10200 14200 10220
rect 13400 9900 13560 10200
rect 14180 9900 14200 10200
rect 13400 9160 14200 9900
rect 13400 1800 13700 9160
rect 13400 1400 15300 1800
rect 14700 -10800 15300 1400
rect -18000 -11400 15300 -10800
rect -23500 -12000 -22700 -11950
rect -23700 -16300 -23450 -12000
rect -22750 -16300 -22700 -12000
rect -23700 -16350 -22700 -16300
rect -23700 -17000 -23000 -16350
rect -23700 -17200 -22700 -17000
rect -18000 -17200 -17200 -11400
rect -23700 -17400 -23000 -17200
rect -19500 -17300 -17200 -17200
rect -23700 -17600 -22700 -17400
rect -19500 -17500 -19300 -17300
rect -18900 -17500 -17200 -17300
rect -23700 -17800 -23000 -17600
rect -19500 -17700 -17200 -17500
rect -23700 -18000 -22700 -17800
rect -19500 -17900 -19300 -17700
rect -18900 -17900 -17200 -17700
rect -23700 -18200 -23000 -18000
rect -19500 -18100 -17200 -17900
rect -23700 -18400 -22700 -18200
rect -19500 -18300 -19300 -18100
rect -18900 -18300 -17200 -18100
rect -23700 -18600 -23000 -18400
rect -19500 -18500 -17200 -18300
rect -23700 -18800 -22700 -18600
rect -19500 -18700 -19300 -18500
rect -18900 -18700 -17200 -18500
rect -23700 -19000 -23000 -18800
rect -23700 -19200 -22700 -19000
rect -23700 -19400 -23000 -19200
rect -23700 -19600 -22700 -19400
rect -23700 -19800 -23000 -19600
rect -23700 -20000 -22700 -19800
rect -23700 -20200 -23000 -20000
rect -23700 -20400 -22700 -20200
rect -23700 -20600 -23000 -20400
rect -23700 -20800 -22700 -20600
rect 23500 -33600 24000 -5600
rect 32800 -32100 34000 -20100
<< via2 >>
rect 13560 9900 14180 10200
rect -23450 -16300 -22750 -12000
<< metal3 >>
rect -14700 13850 -14300 13900
rect -14700 12650 -14650 13850
rect -14350 13000 -14300 13850
rect 16000 13700 20000 13900
rect -14350 12650 -12000 13000
rect -14700 12600 -12000 12650
rect -13200 11850 -12800 12000
rect -14850 11550 -12800 11850
rect -13200 9600 -12800 11550
rect -12400 10400 -12000 12600
rect -12400 10000 -3800 10400
rect -13200 9200 -4600 9600
rect -18300 8200 -18100 8800
rect -22600 8000 -18100 8200
rect -22600 -1300 -22400 8000
rect -17600 7900 -17400 8800
rect -23400 -1400 -22400 -1300
rect -22300 7700 -17400 7900
rect -28000 -8100 -27500 -7600
rect -23400 -8300 -23200 -1400
rect -22300 -1500 -22100 7700
rect -17200 7600 -17000 8800
rect -27200 -8400 -23200 -8300
rect -23100 -1600 -22100 -1500
rect -22000 7400 -17000 7600
rect -27200 -16400 -27000 -8400
rect -23100 -8500 -22900 -1600
rect -22000 -1700 -21800 7400
rect -16400 7300 -16200 8800
rect -31300 -16500 -27000 -16400
rect -26900 -8600 -22900 -8500
rect -22800 -1800 -21800 -1700
rect -21700 7100 -16200 7300
rect -31300 -30000 -31100 -16500
rect -26900 -16600 -26700 -8600
rect -22800 -8700 -22600 -1800
rect -21700 -1900 -21500 7100
rect -16000 7000 -15800 8800
rect -31000 -16700 -26700 -16600
rect -26600 -8800 -22600 -8700
rect -22500 -2000 -21500 -1900
rect -21400 6800 -15800 7000
rect -31000 -30000 -30800 -16700
rect -26600 -16800 -26400 -8800
rect -22500 -8900 -22300 -2000
rect -21400 -2100 -21200 6800
rect -21000 5900 -15800 6500
rect -5000 6000 -4600 9200
rect -4200 6000 -3800 10000
rect 10700 700 12400 8600
rect -13100 -1300 -13000 400
rect -30700 -16900 -26400 -16800
rect -26300 -9000 -22300 -8900
rect -22200 -2200 -21200 -2100
rect -21000 -1400 -13000 -1300
rect -30700 -30000 -30500 -16900
rect -26300 -17000 -26100 -9000
rect -22200 -9100 -22000 -2200
rect -21000 -2400 -20800 -1400
rect -12900 -1500 -12800 400
rect -30400 -17100 -26100 -17000
rect -26000 -9200 -22000 -9100
rect -21900 -2500 -20800 -2400
rect -20700 -1600 -12800 -1500
rect -30400 -30000 -30200 -17100
rect -26000 -17200 -25800 -9200
rect -21900 -9400 -21700 -2500
rect -20700 -2600 -20500 -1600
rect -12700 -1700 -12600 400
rect -30100 -17300 -25800 -17200
rect -25300 -9500 -21700 -9400
rect -21600 -2700 -20500 -2600
rect -20400 -1800 -12600 -1700
rect -30100 -30000 -29900 -17300
rect -25300 -30000 -25100 -9500
rect -21600 -9600 -21400 -2700
rect -20400 -2800 -20200 -1800
rect -12500 -1900 -12400 400
rect -25000 -9700 -21400 -9600
rect -21300 -2900 -20200 -2800
rect -20100 -2000 -12400 -1900
rect -25000 -30000 -24800 -9700
rect -21300 -9800 -21100 -2900
rect -20100 -3000 -19900 -2000
rect -12300 -2100 -12200 400
rect -24700 -9900 -21100 -9800
rect -21000 -3100 -19900 -3000
rect -19800 -2200 -12200 -2100
rect -24700 -30000 -24500 -9900
rect -21000 -10000 -20800 -3100
rect -19800 -3200 -19600 -2200
rect -24400 -10100 -20800 -10000
rect -20700 -3300 -19600 -3200
rect -24400 -30000 -24200 -10100
rect -20700 -10200 -20500 -3300
rect -24100 -10300 -20500 -10200
rect -24100 -30000 -23900 -10300
rect -23500 -12000 -22700 -11950
rect -23500 -16300 -23450 -12000
rect -22750 -16300 -22700 -12000
rect -23500 -16350 -22700 -16300
rect -22500 -16400 -18000 -11900
rect -23600 -19600 -22400 -19400
rect -21350 -19570 -21160 -19560
rect -23600 -21400 -23500 -19600
rect -21350 -19690 -21330 -19570
rect -21170 -19690 -21160 -19570
rect -21350 -19700 -21160 -19690
rect -23800 -21600 -23500 -21400
rect -23400 -19900 -22400 -19700
rect -23800 -30000 -23600 -21600
rect -23400 -21700 -23300 -19900
rect -23500 -30000 -23300 -21700
rect -23200 -20200 -22400 -20000
rect -23200 -21900 -23100 -20200
rect -23000 -20500 -22400 -20300
rect -23000 -21700 -22900 -20500
rect -22800 -20800 -22400 -20600
rect -22800 -21400 -22700 -20800
rect -22800 -21600 -22400 -21400
rect -23000 -21800 -22700 -21700
rect -23200 -30000 -23000 -21900
rect -22900 -30000 -22700 -21800
rect -22600 -30000 -22400 -21600
rect 23500 -33600 24000 -5600
rect 32800 -32100 34000 -20100
<< via3 >>
rect -14650 12650 -14350 13850
rect -23450 -16300 -22750 -12000
rect -21330 -19690 -21170 -19570
<< mimcap >>
rect -22400 -12100 -18300 -12000
rect -22400 -16200 -22300 -12100
rect -18400 -16200 -18300 -12100
rect -22400 -16300 -18300 -16200
<< mimcapcontact >>
rect -22300 -16200 -18400 -12100
<< metal4 >>
rect 24600 21300 26100 25900
rect 24600 19900 26400 21300
rect 24500 13900 26300 19900
rect -14700 13850 -14300 13900
rect -14700 12650 -14650 13850
rect -14350 12650 -14300 13850
rect 16000 13700 20000 13900
rect -14700 12600 -14300 12650
rect 25900 8000 30500 8100
rect -21800 7700 -18800 7800
rect -21800 4700 -21700 7700
rect -18900 4700 -18800 7700
rect -21800 4600 -18800 4700
rect 17500 -1300 17900 2400
rect 25900 -1800 26000 8000
rect 30400 -1800 30500 8000
rect 25900 -1900 30500 -1800
rect -22700 -11950 -18100 -11900
rect -23600 -12000 -18100 -11950
rect -23600 -16300 -23450 -12000
rect -22750 -12100 -18100 -12000
rect -22750 -16200 -22300 -12100
rect -18400 -16200 -18100 -12100
rect -22750 -16300 -18100 -16200
rect -23600 -16400 -18100 -16300
rect -21370 -19570 -21130 -19560
rect -21134 -19810 -21130 -19570
rect -21370 -19820 -21130 -19810
rect 23500 -33600 24000 -5600
rect 32800 -32100 34000 -20100
<< via4 >>
rect -21700 4700 -18900 7700
rect 26000 -1800 30400 8000
rect -21370 -19690 -21330 -19570
rect -21330 -19690 -21170 -19570
rect -21170 -19690 -21134 -19570
rect -21370 -19810 -21134 -19690
<< mimcap2 >>
rect -22400 -12100 -18300 -12000
rect -22400 -16200 -22300 -12100
rect -18400 -16200 -18300 -12100
rect -22400 -16300 -18300 -16200
<< mimcap2contact >>
rect -22300 -16200 -18400 -12100
<< metal5 >>
rect 25900 8000 30500 8100
rect -21800 7700 -18800 7800
rect -21800 4700 -21700 7700
rect -18900 4700 -18800 7700
rect -21800 4600 -18800 4700
rect -21800 800 -19800 4600
rect -17500 1500 -10500 2100
rect -25100 -2300 -23100 -2200
rect -21800 -2300 -18800 800
rect -25100 -4100 -18800 -2300
rect -25100 -7100 -23100 -4100
rect -21800 -7100 -18800 -4100
rect -25100 -8900 -18800 -7100
rect -25100 -11900 -23100 -8900
rect -21800 -11900 -18800 -8900
rect -26900 -12000 -18100 -11900
rect -27200 -12100 -18100 -12000
rect -27200 -13700 -22300 -12100
rect -27200 -15600 -25800 -13700
rect -25200 -15600 -22300 -13700
rect -27200 -16200 -22300 -15600
rect -18400 -16200 -18100 -12100
rect -27200 -16400 -18100 -16200
rect -17500 -19400 -16800 1500
rect 25900 -1600 26000 8000
rect 25800 -1800 26000 -1600
rect 30400 -1600 30500 8000
rect 30400 -1800 30600 -1600
rect 25800 -2000 30600 -1800
rect 26600 -4200 30200 -2000
rect -21700 -19570 -16800 -19400
rect -21700 -19810 -21370 -19570
rect -21134 -19810 -16800 -19570
rect -21700 -20000 -16800 -19810
rect -21700 -20050 -20900 -20000
use CPW_chunk_1_W20  CPW_chunk_1_W20_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660959839
transform 1 0 26000 0 1 -11600
box -2000 -600 6800 7400
use CPW_chunk_1_W20  CPW_chunk_1_W20_1
timestamp 1660959839
transform 1 0 26000 0 1 -19600
box -2000 -600 6800 7400
use CPW_chunk_1_W20  CPW_chunk_1_W20_2
timestamp 1660959839
transform 1 0 26000 0 1 -27600
box -2000 -600 6800 7400
use CPW_chunk_1_W20  CPW_chunk_1_W20_3
timestamp 1660959839
transform 1 0 26000 0 1 -35600
box -2000 -600 6800 7400
use OSC_5GHz_1  OSC_5GHz_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/OSC
timestamp 1661649873
transform -1 0 -3300 0 1 5900
box 10000 -21000 68022 34000
use PA_complete  PA_complete_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/PA
timestamp 1661127237
transform 1 0 14099 0 1 2080
box -18800 -26000 70600 43800
use VGA_complete_1  VGA_complete_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/PA
timestamp 1661836362
transform 1 0 500 0 1 -15300
box -21500 -7100 11600 21400
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660275339
transform 1 0 -24600 0 1 4500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_1
timestamp 1660275339
transform 1 0 -24100 0 1 4500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_2
timestamp 1660275339
transform 1 0 -23600 0 1 4500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_3
timestamp 1660275339
transform 1 0 -24600 0 1 4000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_4
timestamp 1660275339
transform 1 0 -24100 0 1 4000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_5
timestamp 1660275339
transform 1 0 -23600 0 1 4000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_6
timestamp 1660275339
transform 1 0 -24600 0 1 3500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_7
timestamp 1660275339
transform 1 0 -24100 0 1 3500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_8
timestamp 1660275339
transform 1 0 -23600 0 1 3500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_9
timestamp 1660275339
transform 1 0 -24600 0 1 3000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_10
timestamp 1660275339
transform 1 0 -24100 0 1 3000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_11
timestamp 1660275339
transform 1 0 -23600 0 1 3000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_12
timestamp 1660275339
transform 1 0 -24600 0 1 2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_13
timestamp 1660275339
transform 1 0 -24100 0 1 2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_14
timestamp 1660275339
transform 1 0 -23600 0 1 2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_15
timestamp 1660275339
transform 1 0 -24600 0 1 2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_16
timestamp 1660275339
transform 1 0 -24100 0 1 2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_17
timestamp 1660275339
transform 1 0 -23600 0 1 2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_18
timestamp 1660275339
transform 1 0 -24600 0 1 1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_19
timestamp 1660275339
transform 1 0 -24100 0 1 1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_20
timestamp 1660275339
transform 1 0 -23600 0 1 1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_21
timestamp 1660275339
transform 1 0 -24600 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_22
timestamp 1660275339
transform 1 0 -24100 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_23
timestamp 1660275339
transform 1 0 -23600 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_24
timestamp 1660275339
transform 1 0 -24600 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_25
timestamp 1660275339
transform 1 0 -24100 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_26
timestamp 1660275339
transform 1 0 -23600 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_27
timestamp 1660275339
transform 1 0 -24600 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_28
timestamp 1660275339
transform 1 0 -24100 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_29
timestamp 1660275339
transform 1 0 -23600 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_30
timestamp 1660275339
transform 1 0 -12100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_31
timestamp 1660275339
transform 1 0 -10600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_32
timestamp 1660275339
transform 1 0 -10100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_33
timestamp 1660275339
transform 1 0 -10600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_34
timestamp 1660275339
transform 1 0 -10100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_35
timestamp 1660275339
transform 1 0 -11600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_36
timestamp 1660275339
transform 1 0 -11100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_37
timestamp 1660275339
transform 1 0 -11600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_38
timestamp 1660275339
transform 1 0 -15600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_39
timestamp 1660275339
transform 1 0 -15100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_40
timestamp 1660275339
transform 1 0 -15600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_41
timestamp 1660275339
transform 1 0 -15100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_42
timestamp 1660275339
transform 1 0 -14600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_43
timestamp 1660275339
transform 1 0 -14600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_44
timestamp 1660275339
transform 1 0 -14100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_45
timestamp 1660275339
transform 1 0 -14100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_46
timestamp 1660275339
transform 1 0 -11100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_47
timestamp 1660275339
transform 1 0 -12600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_48
timestamp 1660275339
transform 1 0 -13100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_49
timestamp 1660275339
transform 1 0 -13600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_50
timestamp 1660275339
transform 1 0 -8600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_51
timestamp 1660275339
transform 1 0 -8100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_52
timestamp 1660275339
transform 1 0 -9600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_53
timestamp 1660275339
transform 1 0 -9100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_54
timestamp 1660275339
transform 1 0 -8600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_55
timestamp 1660275339
transform 1 0 -13600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_56
timestamp 1660275339
transform 1 0 -8100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_57
timestamp 1660275339
transform 1 0 -9600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_58
timestamp 1660275339
transform 1 0 -9100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_59
timestamp 1660275339
transform 1 0 -6100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_60
timestamp 1660275339
transform 1 0 -6600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_61
timestamp 1660275339
transform 1 0 -7600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_62
timestamp 1660275339
transform 1 0 -7100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_63
timestamp 1660275339
transform 1 0 -6100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_64
timestamp 1660275339
transform 1 0 -6600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_65
timestamp 1660275339
transform 1 0 -7600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_66
timestamp 1660275339
transform 1 0 -7100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_67
timestamp 1660275339
transform 1 0 -8600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_68
timestamp 1660275339
transform 1 0 -8100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_69
timestamp 1660275339
transform 1 0 -12100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_70
timestamp 1660275339
transform 1 0 -8600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_71
timestamp 1660275339
transform 1 0 -12600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_72
timestamp 1660275339
transform 1 0 -13100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_73
timestamp 1660275339
transform 1 0 -8100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_74
timestamp 1660275339
transform 1 0 -9100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_75
timestamp 1660275339
transform 1 0 -9600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_76
timestamp 1660275339
transform 1 0 -9600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_77
timestamp 1660275339
transform 1 0 -9100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_78
timestamp 1660275339
transform 1 0 -6100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_79
timestamp 1660275339
transform 1 0 -6100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_80
timestamp 1660275339
transform 1 0 -6600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_81
timestamp 1660275339
transform 1 0 -6600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_82
timestamp 1660275339
transform 1 0 -7100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_83
timestamp 1660275339
transform 1 0 -7600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_84
timestamp 1660275339
transform 1 0 -7600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_85
timestamp 1660275339
transform 1 0 -7100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_86
timestamp 1660275339
transform 1 0 -10100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_87
timestamp 1660275339
transform 1 0 -10100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_88
timestamp 1660275339
transform 1 0 -10600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_89
timestamp 1660275339
transform 1 0 -10600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_90
timestamp 1660275339
transform 1 0 -11100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_91
timestamp 1660275339
transform 1 0 -11600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_92
timestamp 1660275339
transform 1 0 -11600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_93
timestamp 1660275339
transform 1 0 -11100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_94
timestamp 1660275339
transform 1 0 -10100 0 1 13500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_95
timestamp 1660275339
transform 1 0 -10100 0 1 13000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_96
timestamp 1660275339
transform 1 0 -10600 0 1 13500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_97
timestamp 1660275339
transform 1 0 -10600 0 1 13000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_98
timestamp 1660275339
transform 1 0 -11100 0 1 13500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_99
timestamp 1660275339
transform 1 0 -11600 0 1 13500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_100
timestamp 1660275339
transform 1 0 -11600 0 1 13000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_101
timestamp 1660275339
transform 1 0 -11100 0 1 13000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_102
timestamp 1660275339
transform 1 0 -10100 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_103
timestamp 1660275339
transform 1 0 -10100 0 1 14000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_104
timestamp 1660275339
transform 1 0 -10600 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_105
timestamp 1660275339
transform 1 0 -10600 0 1 14000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_106
timestamp 1660275339
transform 1 0 -11100 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_107
timestamp 1660275339
transform 1 0 -11600 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_108
timestamp 1660275339
transform 1 0 -11600 0 1 14000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_109
timestamp 1660275339
transform 1 0 -11100 0 1 14000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_110
timestamp 1660275339
transform 1 0 -11600 0 1 15000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_111
timestamp 1660275339
transform 1 0 -12100 0 1 15000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_112
timestamp 1660275339
transform 1 0 -12100 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_113
timestamp 1660275339
transform 1 0 -12600 0 1 15000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_114
timestamp 1660275339
transform 1 0 -13100 0 1 15000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_115
timestamp 1660275339
transform 1 0 -13100 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_116
timestamp 1660275339
transform 1 0 -12600 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_117
timestamp 1660275339
transform 1 0 -5600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_118
timestamp 1660275339
transform 1 0 -5100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_119
timestamp 1660275339
transform 1 0 -4600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_120
timestamp 1660275339
transform 1 0 -4100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_121
timestamp 1660275339
transform 1 0 -3600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_122
timestamp 1660275339
transform 1 0 -3100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_123
timestamp 1660275339
transform 1 0 -5600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_124
timestamp 1660275339
transform 1 0 -5100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_125
timestamp 1660275339
transform 1 0 -4600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_126
timestamp 1660275339
transform 1 0 -4100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_127
timestamp 1660275339
transform 1 0 -3600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_128
timestamp 1660275339
transform 1 0 -3100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_129
timestamp 1660275339
transform 1 0 -2600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_130
timestamp 1660275339
transform 1 0 -2100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_131
timestamp 1660275339
transform 1 0 -2600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_132
timestamp 1660275339
transform 1 0 -2100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_133
timestamp 1660275339
transform 1 0 -2600 0 1 11500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_134
timestamp 1660275339
transform 1 0 -2100 0 1 11500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_135
timestamp 1660275339
transform 1 0 -2600 0 1 11000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_136
timestamp 1660275339
transform 1 0 -2100 0 1 11000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_137
timestamp 1660275339
transform 1 0 -2600 0 1 10500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_138
timestamp 1660275339
transform 1 0 -2100 0 1 10500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_139
timestamp 1660275339
transform 1 0 -2600 0 1 10000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_140
timestamp 1660275339
transform 1 0 -2100 0 1 10000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_141
timestamp 1660275339
transform 1 0 -2600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_142
timestamp 1660275339
transform 1 0 -2100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_143
timestamp 1660275339
transform 1 0 -2600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_144
timestamp 1660275339
transform 1 0 -2100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_145
timestamp 1660275339
transform 1 0 -2600 0 1 8500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_146
timestamp 1660275339
transform 1 0 -2100 0 1 8500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_147
timestamp 1660275339
transform 1 0 -2600 0 1 8000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_148
timestamp 1660275339
transform 1 0 -2100 0 1 8000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_149
timestamp 1660275339
transform 1 0 -2600 0 1 7500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_150
timestamp 1660275339
transform 1 0 -2100 0 1 7500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_151
timestamp 1660275339
transform 1 0 -2600 0 1 7000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_152
timestamp 1660275339
transform 1 0 -2100 0 1 7000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_153
timestamp 1660275339
transform 1 0 -3100 0 1 11500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_154
timestamp 1660275339
transform 1 0 -3100 0 1 11000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_155
timestamp 1660275339
transform 1 0 -3100 0 1 10500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_156
timestamp 1660275339
transform 1 0 -24100 0 1 5000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_157
timestamp 1660275339
transform 1 0 -24600 0 1 5000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_158
timestamp 1660275339
transform 1 0 -24600 0 1 5500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_159
timestamp 1660275339
transform 1 0 -24100 0 1 5500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_160
timestamp 1660275339
transform 1 0 -3100 0 1 10000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_161
timestamp 1660275339
transform 1 0 -23600 0 1 5000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_162
timestamp 1660275339
transform 1 0 -23600 0 1 5500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_163
timestamp 1660275339
transform 1 0 -3100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_164
timestamp 1660275339
transform 1 0 -3100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_165
timestamp 1660275339
transform 1 0 -3100 0 1 8500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_166
timestamp 1660275339
transform 1 0 -3100 0 1 8000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_167
timestamp 1660275339
transform 1 0 -3100 0 1 7000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_168
timestamp 1660275339
transform 1 0 -3100 0 1 7500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_169
timestamp 1660275339
transform 1 0 13400 0 1 -1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_170
timestamp 1660275339
transform 1 0 13400 0 1 -1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_171
timestamp 1660275339
transform 1 0 13400 0 1 -2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_172
timestamp 1660275339
transform 1 0 13400 0 1 -2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_173
timestamp 1660275339
transform 1 0 13400 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_174
timestamp 1660275339
transform 1 0 13400 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_175
timestamp 1660275339
transform 1 0 13400 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_176
timestamp 1660275339
transform 1 0 13400 0 1 -500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_177
timestamp 1660275339
transform 1 0 13900 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_178
timestamp 1660275339
transform 1 0 13900 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_179
timestamp 1660275339
transform 1 0 13900 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_180
timestamp 1660275339
transform 1 0 13900 0 1 -500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_181
timestamp 1660275339
transform 1 0 13900 0 1 -1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_182
timestamp 1660275339
transform 1 0 13900 0 1 -1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_183
timestamp 1660275339
transform 1 0 13900 0 1 -2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_184
timestamp 1660275339
transform 1 0 13900 0 1 -2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_185
timestamp 1660275339
transform 1 0 15400 0 1 -3500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_186
timestamp 1660275339
transform 1 0 15400 0 1 -3000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_187
timestamp 1660275339
transform 1 0 15400 0 1 -4000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5#0  hash_m1m2m3_W2p5L2p5_188
timestamp 1660275339
transform 1 0 15400 0 1 -4500
box 100 -1100 600 -600
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660789662
transform 1 0 22500 0 1 -8900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_1
timestamp 1660789662
transform 1 0 22500 0 1 -9900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_2
timestamp 1660789662
transform 1 0 22500 0 1 -10900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_3
timestamp 1660789662
transform 1 0 22500 0 1 -11900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_4
timestamp 1660789662
transform 1 0 22500 0 1 -14900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_5
timestamp 1660789662
transform 1 0 22500 0 1 -13900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_6
timestamp 1660789662
transform 1 0 22500 0 1 -12900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_7
timestamp 1660789662
transform 1 0 22500 0 1 -17900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_8
timestamp 1660789662
transform 1 0 22500 0 1 -16900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_9
timestamp 1660789662
transform 1 0 22500 0 1 -15900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_10
timestamp 1660789662
transform 1 0 22500 0 1 -20900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_11
timestamp 1660789662
transform 1 0 22500 0 1 -19900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_12
timestamp 1660789662
transform 1 0 22500 0 1 -18900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_13
timestamp 1660789662
transform 1 0 22500 0 1 -23900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_14
timestamp 1660789662
transform 1 0 22500 0 1 -22900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_15
timestamp 1660789662
transform 1 0 22500 0 1 -21900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_16
timestamp 1660789662
transform 1 0 22500 0 1 -26900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_17
timestamp 1660789662
transform 1 0 22500 0 1 -25900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_18
timestamp 1660789662
transform 1 0 22500 0 1 -24900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_19
timestamp 1660789662
transform 1 0 22500 0 1 -29900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_20
timestamp 1660789662
transform 1 0 22500 0 1 -28900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_21
timestamp 1660789662
transform 1 0 22500 0 1 -27900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_22
timestamp 1660789662
transform 1 0 -17000 0 1 -2400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_23
timestamp 1660789662
transform 1 0 22500 0 1 -31900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_24
timestamp 1660789662
transform 1 0 22500 0 1 -30900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_25
timestamp 1660789662
transform 1 0 -16000 0 1 -2400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_26
timestamp 1660789662
transform 1 0 -16500 0 1 -18400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5#0  hash_m1m2m3_W5L5_27
timestamp 1660789662
transform 1 0 -16500 0 1 -17400
box 0 -1700 1000 -700
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660789662
transform 1 0 -11500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_1
timestamp 1660789662
transform 1 0 -15500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_2
timestamp 1660789662
transform 1 0 -13500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_3
timestamp 1660789662
transform 1 0 -9500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_4
timestamp 1660789662
transform 1 0 -7500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_5
timestamp 1660789662
transform 1 0 -7500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_6
timestamp 1660789662
transform 1 0 -9500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_7
timestamp 1660789662
transform 1 0 500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_8
timestamp 1660789662
transform 1 0 500 0 1 9600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_9
timestamp 1660789662
transform 1 0 -3500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_10
timestamp 1660789662
transform 1 0 -5500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_11
timestamp 1660789662
transform 1 0 500 0 1 11600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_12
timestamp 1660789662
transform 1 0 -1500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_13
timestamp 1660789662
transform 1 0 2500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_14
timestamp 1660789662
transform 1 0 -1500 0 1 11600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_15
timestamp 1660789662
transform 1 0 2500 0 1 9600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_16
timestamp 1660789662
transform 1 0 -1500 0 1 9600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_17
timestamp 1660789662
transform 1 0 2500 0 1 11600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_18
timestamp 1660789662
transform 1 0 -1500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_19
timestamp 1660789662
transform 1 0 16000 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_20
timestamp 1660789662
transform 1 0 -3500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_21
timestamp 1660789662
transform 1 0 -5500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_22
timestamp 1660789662
transform 1 0 -7500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_23
timestamp 1660789662
transform 1 0 -9500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_24
timestamp 1660789662
transform 1 0 -11500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_25
timestamp 1660789662
transform 1 0 -11500 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_26
timestamp 1660789662
transform 1 0 -9500 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_27
timestamp 1660789662
transform 1 0 -7500 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_28
timestamp 1660789662
transform 1 0 -5500 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_29
timestamp 1660789662
transform 1 0 18000 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_30
timestamp 1660789662
transform 1 0 -11500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_31
timestamp 1660789662
transform 1 0 -9500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_32
timestamp 1660789662
transform 1 0 -7500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_33
timestamp 1660789662
transform 1 0 20000 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_34
timestamp 1660789662
transform 1 0 26000 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_35
timestamp 1660789662
transform 1 0 9500 0 1 100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_36
timestamp 1660789662
transform 1 0 11500 0 1 100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_37
timestamp 1660789662
transform 1 0 11500 0 1 -1900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_38
timestamp 1660789662
transform 1 0 19500 0 1 -3900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_39
timestamp 1660789662
transform 1 0 15500 0 1 100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_40
timestamp 1660789662
transform 1 0 15500 0 1 -1900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_41
timestamp 1660789662
transform 1 0 15500 0 1 2100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_42
timestamp 1660789662
transform 1 0 21500 0 1 -3900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_43
timestamp 1660789662
transform 1 0 28000 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_44
timestamp 1660789662
transform 1 0 24000 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_45
timestamp 1660789662
transform 1 0 22000 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_46
timestamp 1660789662
transform 1 0 20000 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_47
timestamp 1660789662
transform 1 0 30000 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_48
timestamp 1660789662
transform 1 0 32000 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_49
timestamp 1660789662
transform 1 0 26000 0 1 29600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_50
timestamp 1660789662
transform 1 0 26000 0 1 31600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_51
timestamp 1660789662
transform 1 0 26000 0 1 33600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_52
timestamp 1660789662
transform 1 0 26000 0 1 35600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_53
timestamp 1660789662
transform 1 0 26000 0 1 37600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_54
timestamp 1660789662
transform 1 0 26000 0 1 39600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_55
timestamp 1660789662
transform 1 0 34500 0 1 -24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_56
timestamp 1660789662
transform 1 0 34500 0 1 -26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_57
timestamp 1660789662
transform 1 0 34500 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_58
timestamp 1660789662
transform 1 0 34500 0 1 -28400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_59
timestamp 1660789662
transform 1 0 26000 0 1 41600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_60
timestamp 1660789662
transform 1 0 26000 0 1 43600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_61
timestamp 1660789662
transform 1 0 34000 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_62
timestamp 1660789662
transform 1 0 34000 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_63
timestamp 1660789662
transform 1 0 34000 0 1 -24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_64
timestamp 1660789662
transform 1 0 34000 0 1 -26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_65
timestamp 1660789662
transform 1 0 34000 0 1 -28400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_66
timestamp 1660789662
transform 1 0 34000 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_67
timestamp 1660789662
transform 1 0 34000 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_68
timestamp 1660789662
transform 1 0 -15500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_69
timestamp 1660789662
transform 1 0 -13500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_70
timestamp 1660789662
transform 1 0 -19500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_71
timestamp 1660789662
transform 1 0 -17500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_72
timestamp 1660789662
transform 1 0 22000 0 1 47600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_73
timestamp 1660789662
transform 1 0 -3500 0 1 47600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_74
timestamp 1660789662
transform 1 0 -7500 0 1 43600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_75
timestamp 1660789662
transform 1 0 22000 0 1 45600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_76
timestamp 1660789662
transform 1 0 24000 0 1 43600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_77
timestamp 1660789662
transform 1 0 20000 0 1 47600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_78
timestamp 1660789662
transform 1 0 36000 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_79
timestamp 1660789662
transform 1 0 38000 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_80
timestamp 1660789662
transform 1 0 -17500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_81
timestamp 1660789662
transform 1 0 -17500 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_82
timestamp 1660789662
transform 1 0 -19500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_83
timestamp 1660789662
transform 1 0 -21500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_84
timestamp 1660789662
transform 1 0 -21500 0 1 -24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_85
timestamp 1660789662
transform 1 0 -21500 0 1 -26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_86
timestamp 1660789662
transform 1 0 -21500 0 1 -28400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_87
timestamp 1660789662
transform 1 0 -21500 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_160
timestamp 1660789662
transform 1 0 34500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_168
timestamp 1660789662
transform 1 0 34500 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_183
timestamp 1660789662
transform 1 0 12500 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_185
timestamp 1660789662
transform 1 0 12500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_186
timestamp 1660789662
transform 1 0 10500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_255
timestamp 1660789662
transform 1 0 -11500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_256
timestamp 1660789662
transform 1 0 -15500 0 1 -18400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_258
timestamp 1660789662
transform 1 0 -17000 0 1 -16400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_259
timestamp 1660789662
transform 1 0 -17000 0 1 -14400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_260
timestamp 1660789662
transform 1 0 -17000 0 1 -12400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_261
timestamp 1660789662
transform 1 0 -17000 0 1 -4400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_262
timestamp 1660789662
transform 1 0 -17000 0 1 -8400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_263
timestamp 1660789662
transform 1 0 -17000 0 1 -6400
box 0 -1700 2000 300
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501637
transform 1 0 -11500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_1
timestamp 1659501637
transform 1 0 -7500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_2
timestamp 1659501637
transform 1 0 24000 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_3
timestamp 1659501637
transform 1 0 -27500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_4
timestamp 1659501637
transform 1 0 -83500 0 1 31900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_5
timestamp 1659501637
transform 1 0 -15500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_6
timestamp 1659501637
transform 1 0 -19500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_7
timestamp 1659501637
transform 1 0 -27500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_8
timestamp 1659501637
transform 1 0 -23500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_9
timestamp 1659501637
transform 1 0 28000 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_10
timestamp 1659501637
transform 1 0 22000 0 1 13900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_11
timestamp 1659501637
transform 1 0 32000 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_12
timestamp 1659501637
transform 1 0 36000 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_13
timestamp 1659501637
transform 1 0 -31500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_14
timestamp 1659501637
transform 1 0 -19500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_15
timestamp 1659501637
transform 1 0 -29500 0 1 -21600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_16
timestamp 1659501637
transform 1 0 -19500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_17
timestamp 1659501637
transform 1 0 -29500 0 1 -25600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_18
timestamp 1659501637
transform 1 0 15500 0 1 -5600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_19
timestamp 1659501637
transform 1 0 15500 0 1 -9600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_20
timestamp 1659501637
transform 1 0 19500 0 1 -9600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_21
timestamp 1659501637
transform 1 0 -83500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_22
timestamp 1659501637
transform 1 0 -71500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_23
timestamp 1659501637
transform 1 0 -83500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_24
timestamp 1659501637
transform 1 0 -83500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_25
timestamp 1659501637
transform 1 0 -83500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_26
timestamp 1659501637
transform 1 0 -83500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_27
timestamp 1659501637
transform 1 0 -29500 0 1 -29600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_28
timestamp 1659501637
transform 1 0 -83500 0 1 51900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_29
timestamp 1659501637
transform 1 0 -83500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_30
timestamp 1659501637
transform 1 0 -83500 0 1 -20100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_31
timestamp 1659501637
transform 1 0 -83500 0 1 -24100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_32
timestamp 1659501637
transform 1 0 -35500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_33
timestamp 1659501637
transform 1 0 -83500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_34
timestamp 1659501637
transform 1 0 -27500 0 1 23900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_35
timestamp 1659501637
transform 1 0 -31500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_36
timestamp 1659501637
transform 1 0 -63500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_37
timestamp 1659501637
transform 1 0 -27500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_38
timestamp 1659501637
transform 1 0 -27500 0 1 -8100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_39
timestamp 1659501637
transform 1 0 -59500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_40
timestamp 1659501637
transform 1 0 -27500 0 1 -4100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_41
timestamp 1659501637
transform 1 0 -55500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_42
timestamp 1659501637
transform 1 0 -51500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_43
timestamp 1659501637
transform 1 0 -47500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_44
timestamp 1659501637
transform 1 0 -43500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_45
timestamp 1659501637
transform 1 0 -71500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_46
timestamp 1659501637
transform 1 0 -31500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_47
timestamp 1659501637
transform 1 0 -39500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_48
timestamp 1659501637
transform 1 0 -27500 0 1 -100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_49
timestamp 1659501637
transform 1 0 76500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_50
timestamp 1659501637
transform 1 0 -35500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_51
timestamp 1659501637
transform 1 0 84500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_52
timestamp 1659501637
transform 1 0 -35500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_53
timestamp 1659501637
transform 1 0 -27500 0 1 31900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_55
timestamp 1659501637
transform 1 0 76500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_56
timestamp 1659501637
transform 1 0 -15500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_57
timestamp 1659501637
transform 1 0 -3500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_58
timestamp 1659501637
transform 1 0 -7500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_59
timestamp 1659501637
transform 1 0 12500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_60
timestamp 1659501637
transform 1 0 8500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_61
timestamp 1659501637
transform 1 0 88500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_62
timestamp 1659501637
transform 1 0 4500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_63
timestamp 1659501637
transform 1 0 500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_64
timestamp 1659501637
transform 1 0 92500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_65
timestamp 1659501637
transform 1 0 -11500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_66
timestamp 1659501637
transform 1 0 14500 0 1 -24100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_67
timestamp 1659501637
transform 1 0 84500 0 1 -20100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_68
timestamp 1659501637
transform 1 0 18500 0 1 -24100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_69
timestamp 1659501637
transform 1 0 18500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_70
timestamp 1659501637
transform 1 0 16500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_71
timestamp 1659501637
transform 1 0 36500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_73
timestamp 1659501637
transform 1 0 14500 0 1 -20100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_74
timestamp 1659501637
transform 1 0 18500 0 1 -20100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_75
timestamp 1659501637
transform 1 0 84500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_76
timestamp 1659501637
transform 1 0 88500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_77
timestamp 1659501637
transform 1 0 92500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_78
timestamp 1659501637
transform 1 0 80500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_79
timestamp 1659501637
transform 1 0 76500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_80
timestamp 1659501637
transform 1 0 72500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_81
timestamp 1659501637
transform 1 0 68500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_82
timestamp 1659501637
transform 1 0 64500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_83
timestamp 1659501637
transform 1 0 60500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_84
timestamp 1659501637
transform 1 0 56500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_85
timestamp 1659501637
transform 1 0 52500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_87
timestamp 1659501637
transform 1 0 36500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_88
timestamp 1659501637
transform 1 0 40500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_89
timestamp 1659501637
transform 1 0 44500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_90
timestamp 1659501637
transform 1 0 48500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_91
timestamp 1659501637
transform 1 0 14500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_92
timestamp 1659501637
transform 1 0 16500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_93
timestamp 1659501637
transform 1 0 18500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_94
timestamp 1659501637
transform 1 0 18500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_95
timestamp 1659501637
transform 1 0 8500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_96
timestamp 1659501637
transform 1 0 12500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_98
timestamp 1659501637
transform 1 0 16500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_99
timestamp 1659501637
transform 1 0 18500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_102
timestamp 1659501637
transform 1 0 -39500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_103
timestamp 1659501637
transform 1 0 -35500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_110
timestamp 1659501637
transform 1 0 -71500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_111
timestamp 1659501637
transform 1 0 -67500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_112
timestamp 1659501637
transform 1 0 -79500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_113
timestamp 1659501637
transform 1 0 -75500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_116
timestamp 1659501637
transform 1 0 -11500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_117
timestamp 1659501637
transform 1 0 -15500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_118
timestamp 1659501637
transform 1 0 -15500 0 1 -24100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_119
timestamp 1659501637
transform 1 0 -7500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_120
timestamp 1659501637
transform 1 0 -3500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_121
timestamp 1659501637
transform 1 0 500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_122
timestamp 1659501637
transform 1 0 4500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660792292
transform 1 0 -15500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_1
timestamp 1660792292
transform 1 0 -15500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_2
timestamp 1660792292
transform 1 0 -23500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_3
timestamp 1660792292
transform 1 0 -15500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_4
timestamp 1660792292
transform 1 0 -23500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_5
timestamp 1660792292
transform 1 0 -31500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_6
timestamp 1660792292
transform 1 0 -15500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_7
timestamp 1660792292
transform 1 0 -23500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_8
timestamp 1660792292
transform 1 0 -31500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_9
timestamp 1660792292
transform 1 0 -39500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_10
timestamp 1660792292
transform 1 0 -7500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_11
timestamp 1660792292
transform 1 0 500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_12
timestamp 1660792292
transform 1 0 8500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_13
timestamp 1660792292
transform 1 0 16500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_14
timestamp 1660792292
transform 1 0 24500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_15
timestamp 1660792292
transform 1 0 -63500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_16
timestamp 1660792292
transform 1 0 -47500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_17
timestamp 1660792292
transform 1 0 -55500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_18
timestamp 1660792292
transform 1 0 -55500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_19
timestamp 1660792292
transform 1 0 -47500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_20
timestamp 1660792292
transform 1 0 -63500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_21
timestamp 1660792292
transform 1 0 -23500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_22
timestamp 1660792292
transform 1 0 -71500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_23
timestamp 1660792292
transform 1 0 -71500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_24
timestamp 1660792292
transform 1 0 -79500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_25
timestamp 1660792292
transform 1 0 -79500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_27
timestamp 1660792292
transform 1 0 -83500 0 1 -8100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_28
timestamp 1660792292
transform 1 0 -83500 0 1 -100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_29
timestamp 1660792292
transform 1 0 -83500 0 1 7900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_30
timestamp 1660792292
transform 1 0 -83500 0 1 15900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_31
timestamp 1660792292
transform 1 0 -83500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_32
timestamp 1660792292
transform 1 0 -79500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_36
timestamp 1660792292
transform 1 0 -79500 0 1 -16100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_37
timestamp 1660792292
transform 1 0 -79500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_38
timestamp 1660792292
transform 1 0 -71500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_42
timestamp 1660792292
transform 1 0 -39500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_44
timestamp 1660792292
transform 1 0 32500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_45
timestamp 1660792292
transform 1 0 40500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_46
timestamp 1660792292
transform 1 0 48500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_47
timestamp 1660792292
transform 1 0 56500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_48
timestamp 1660792292
transform 1 0 64500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_49
timestamp 1660792292
transform 1 0 72500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_50
timestamp 1660792292
transform 1 0 80500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_51
timestamp 1660792292
transform 1 0 88500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_52
timestamp 1660792292
transform 1 0 28000 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_53
timestamp 1660792292
transform 1 0 36000 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_54
timestamp 1660792292
transform 1 0 44000 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_55
timestamp 1660792292
transform 1 0 52000 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_56
timestamp 1660792292
transform 1 0 60000 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_57
timestamp 1660792292
transform 1 0 68000 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_58
timestamp 1660792292
transform 1 0 76000 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_59
timestamp 1660792292
transform 1 0 88500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_60
timestamp 1660792292
transform 1 0 88500 0 1 27900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_61
timestamp 1660792292
transform 1 0 88500 0 1 19900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_62
timestamp 1660792292
transform 1 0 88500 0 1 11900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_63
timestamp 1660792292
transform 1 0 88500 0 1 3900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_64
timestamp 1660792292
transform 1 0 88500 0 1 -4100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_65
timestamp 1660792292
transform 1 0 88500 0 1 -12100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_66
timestamp 1660792292
transform 1 0 88500 0 1 -20100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_67
timestamp 1660792292
transform 1 0 84000 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_68
timestamp 1660792292
transform 1 0 88500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_69
timestamp 1660792292
transform 1 0 84000 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_70
timestamp 1660792292
transform 1 0 76000 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_71
timestamp 1660792292
transform 1 0 68000 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_72
timestamp 1660792292
transform 1 0 60000 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_73
timestamp 1660792292
transform 1 0 52000 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_74
timestamp 1660792292
transform 1 0 44000 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_75
timestamp 1660792292
transform 1 0 36000 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_76
timestamp 1660792292
transform 1 0 28000 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_77
timestamp 1660792292
transform 1 0 80500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_78
timestamp 1660792292
transform 1 0 80500 0 1 23900
box 0 0 8000 8000
use pmirror_pfet_64x_complete  pmirror_pfet_64x_complete_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660185098
transform 0 1 -22800 -1 0 -16650
box 0 0 4280 3344
<< labels >>
rlabel metal4 -23600 -16400 -22500 -16300 1 VHI
rlabel metal3 -23600 -21300 -23500 -21100 1 G32
rlabel metal3 -23400 -21300 -23300 -21100 1 G16
rlabel metal3 -23200 -21300 -23100 -21100 1 G2
rlabel metal3 -23000 -21300 -22900 -21100 1 G4
rlabel metal3 -22800 -21300 -22700 -21100 1 G8
rlabel metal5 -21700 -20050 -20900 -19450 3 IREF
<< end >>
