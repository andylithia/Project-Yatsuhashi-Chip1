magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< error_s >>
rect 38 26482 80 26491
rect 38 26465 113 26482
rect 42 26448 76 26465
rect 79 26448 113 26465
rect 42 26369 46 26403
rect 72 26369 76 26403
rect -25 26332 25 26334
rect 0 26324 14 26325
rect 0 26323 17 26324
rect 25 26323 27 26332
rect 0 26316 38 26323
rect 0 26315 34 26316
rect 0 26299 8 26315
rect 14 26299 34 26315
rect 0 26298 34 26299
rect 0 26291 38 26298
rect 14 26290 17 26291
rect 25 26282 27 26291
rect 42 26262 45 26352
rect 71 26321 80 26349
rect 69 26283 80 26321
rect 107 26277 119 26311
rect 129 26283 143 26311
rect 129 26277 141 26283
rect 42 26211 46 26245
rect 72 26211 76 26245
rect 42 26164 76 26168
rect 42 26134 46 26164
rect 72 26134 76 26164
rect 16 26125 38 26131
rect 80 26125 102 26131
rect 144 26125 148 26465
rect 151 26448 156 26482
rect 180 26451 185 26482
rect 400 26465 442 26491
rect 174 26443 246 26451
rect 256 26443 328 26451
rect 332 26449 336 26465
rect 400 26457 438 26465
rect 400 26450 408 26457
rect 434 26450 438 26457
rect 388 26449 454 26450
rect 224 26413 226 26429
rect 196 26405 226 26413
rect 196 26401 230 26405
rect 196 26371 204 26401
rect 216 26371 230 26401
rect 224 26324 226 26371
rect 300 26344 308 26413
rect 332 26411 342 26449
rect 400 26441 404 26449
rect 454 26435 504 26437
rect 494 26431 548 26435
rect 494 26426 514 26431
rect 504 26411 506 26426
rect 336 26399 342 26411
rect 289 26334 308 26344
rect 300 26328 308 26334
rect 332 26365 342 26399
rect 400 26403 404 26411
rect 400 26369 408 26403
rect 434 26369 438 26403
rect 498 26401 506 26411
rect 514 26401 515 26421
rect 504 26385 506 26401
rect 525 26392 528 26426
rect 547 26401 548 26421
rect 557 26401 564 26411
rect 514 26385 530 26391
rect 532 26385 548 26391
rect 332 26337 373 26365
rect 332 26331 351 26337
rect 196 26290 204 26324
rect 216 26290 230 26324
rect 244 26290 257 26324
rect 278 26294 291 26328
rect 300 26312 321 26328
rect 336 26321 351 26331
rect 300 26310 312 26312
rect 300 26294 321 26310
rect 332 26303 351 26321
rect 361 26303 375 26337
rect 400 26331 411 26369
rect 562 26332 612 26334
rect 400 26303 409 26331
rect 466 26323 497 26325
rect 565 26323 596 26325
rect 442 26316 500 26323
rect 466 26315 500 26316
rect 565 26315 599 26323
rect 174 26253 181 26277
rect 224 26243 226 26290
rect 300 26281 308 26294
rect 289 26278 305 26280
rect 332 26253 342 26303
rect 400 26283 404 26303
rect 497 26299 500 26315
rect 596 26299 599 26315
rect 466 26298 500 26299
rect 442 26291 500 26298
rect 565 26291 599 26299
rect 612 26282 614 26332
rect 256 26243 328 26251
rect 336 26245 342 26253
rect 400 26245 404 26253
rect 196 26213 204 26243
rect 216 26213 230 26243
rect 196 26209 230 26213
rect 196 26201 226 26209
rect 224 26185 226 26201
rect 332 26173 336 26241
rect 400 26211 408 26245
rect 434 26211 438 26245
rect 454 26229 504 26231
rect 504 26213 506 26229
rect 514 26223 530 26229
rect 532 26223 548 26229
rect 525 26213 548 26222
rect 400 26203 404 26211
rect 498 26203 506 26213
rect 504 26179 506 26203
rect 514 26193 515 26213
rect 525 26188 528 26213
rect 547 26193 548 26213
rect 557 26203 564 26213
rect 514 26179 548 26183
rect 400 26173 442 26174
rect 174 26163 246 26171
rect 400 26166 404 26173
rect 295 26132 300 26166
rect 324 26132 329 26166
rect 367 26132 438 26166
rect 400 26131 404 26132
rect 378 26125 404 26131
rect 442 26125 464 26131
rect 38 26109 80 26125
rect 400 26109 442 26125
rect -25 26095 25 26097
rect 455 26095 505 26097
rect 557 26095 607 26097
rect 16 26087 102 26095
rect 378 26087 464 26095
rect 8 26053 17 26087
rect 18 26085 51 26087
rect 80 26085 100 26087
rect 18 26053 100 26085
rect 380 26085 404 26087
rect 429 26085 438 26087
rect 442 26085 462 26087
rect 16 26045 102 26053
rect 42 26029 76 26031
rect 16 26009 38 26015
rect 42 26006 76 26010
rect 80 26009 102 26015
rect 42 25976 46 26006
rect 72 25976 76 26006
rect 42 25895 46 25929
rect 72 25895 76 25929
rect -25 25858 25 25860
rect 0 25850 14 25851
rect 0 25849 17 25850
rect 25 25849 27 25858
rect 0 25842 38 25849
rect 0 25841 34 25842
rect 0 25825 8 25841
rect 14 25825 34 25841
rect 0 25824 34 25825
rect 0 25817 38 25824
rect 14 25816 17 25817
rect 25 25808 27 25817
rect 42 25788 45 25878
rect 69 25863 80 25895
rect 107 25863 143 25891
rect 107 25857 119 25863
rect 109 25829 119 25857
rect 129 25829 143 25863
rect 42 25737 46 25771
rect 72 25737 76 25771
rect 38 25699 80 25700
rect 42 25658 76 25692
rect 79 25658 113 25692
rect 42 25579 46 25613
rect 72 25579 76 25613
rect -25 25542 25 25544
rect 0 25534 14 25535
rect 0 25533 17 25534
rect 25 25533 27 25542
rect 0 25526 38 25533
rect 0 25525 34 25526
rect 0 25509 8 25525
rect 14 25509 34 25525
rect 0 25508 34 25509
rect 0 25501 38 25508
rect 14 25500 17 25501
rect 25 25492 27 25501
rect 42 25472 45 25562
rect 71 25531 80 25559
rect 69 25493 80 25531
rect 107 25487 119 25521
rect 129 25493 143 25521
rect 129 25487 141 25493
rect 42 25421 46 25455
rect 72 25421 76 25455
rect 42 25374 76 25378
rect 42 25344 46 25374
rect 72 25344 76 25374
rect 16 25335 38 25341
rect 80 25335 102 25341
rect 144 25335 148 26083
rect 332 26015 336 26083
rect 380 26053 462 26085
rect 463 26053 472 26087
rect 480 26053 497 26087
rect 378 26045 464 26053
rect 505 26045 507 26095
rect 514 26053 548 26087
rect 565 26053 582 26087
rect 607 26045 609 26095
rect 404 26029 438 26031
rect 400 26015 442 26016
rect 378 26009 404 26015
rect 442 26009 464 26015
rect 400 26008 404 26009
rect 174 25969 246 25977
rect 295 25974 300 26008
rect 324 25974 329 26008
rect 224 25939 226 25955
rect 196 25931 226 25939
rect 332 25937 336 26005
rect 367 25974 438 26008
rect 400 25967 404 25974
rect 454 25961 504 25963
rect 494 25957 548 25961
rect 494 25952 514 25957
rect 504 25937 506 25952
rect 196 25927 230 25931
rect 196 25897 204 25927
rect 216 25897 230 25927
rect 400 25929 404 25937
rect 174 25863 181 25889
rect 224 25850 226 25897
rect 256 25889 328 25897
rect 332 25895 336 25925
rect 400 25895 408 25929
rect 434 25895 438 25929
rect 498 25927 506 25937
rect 514 25927 515 25947
rect 504 25911 506 25927
rect 525 25918 528 25952
rect 547 25927 548 25947
rect 557 25927 564 25937
rect 514 25911 530 25917
rect 532 25911 548 25917
rect 289 25860 305 25862
rect 196 25816 204 25850
rect 216 25816 230 25850
rect 244 25816 257 25850
rect 300 25846 308 25859
rect 332 25857 342 25895
rect 400 25887 404 25895
rect 336 25847 342 25857
rect 224 25769 226 25816
rect 278 25812 291 25846
rect 300 25830 321 25846
rect 332 25837 342 25847
rect 400 25847 409 25875
rect 562 25858 612 25860
rect 466 25849 497 25851
rect 565 25849 596 25851
rect 300 25828 312 25830
rect 300 25812 321 25828
rect 300 25806 308 25812
rect 289 25796 308 25806
rect 196 25739 204 25769
rect 216 25739 230 25769
rect 196 25735 230 25739
rect 196 25727 226 25735
rect 300 25727 308 25796
rect 332 25803 351 25837
rect 361 25803 375 25837
rect 400 25803 411 25847
rect 442 25842 500 25849
rect 466 25841 500 25842
rect 565 25841 599 25849
rect 497 25825 500 25841
rect 596 25825 599 25841
rect 466 25824 500 25825
rect 442 25817 500 25824
rect 565 25817 599 25825
rect 612 25808 614 25858
rect 332 25779 342 25803
rect 336 25767 342 25779
rect 224 25711 226 25727
rect 332 25699 342 25767
rect 400 25771 404 25779
rect 400 25737 408 25771
rect 434 25737 438 25771
rect 454 25755 504 25757
rect 504 25739 506 25755
rect 514 25749 530 25755
rect 532 25749 548 25755
rect 525 25739 548 25748
rect 400 25729 404 25737
rect 498 25729 506 25739
rect 504 25705 506 25729
rect 514 25719 515 25739
rect 525 25714 528 25739
rect 547 25719 548 25739
rect 557 25729 564 25739
rect 514 25705 548 25709
rect 151 25658 156 25692
rect 174 25689 246 25697
rect 256 25689 328 25697
rect 336 25691 342 25699
rect 400 25694 404 25699
rect 180 25661 185 25689
rect 174 25653 246 25661
rect 256 25653 328 25661
rect 332 25659 336 25689
rect 400 25660 438 25694
rect 224 25623 226 25639
rect 196 25615 226 25623
rect 196 25611 230 25615
rect 196 25581 204 25611
rect 216 25581 230 25611
rect 224 25534 226 25581
rect 300 25554 308 25623
rect 332 25621 342 25659
rect 400 25651 404 25660
rect 454 25645 504 25647
rect 494 25641 548 25645
rect 494 25636 514 25641
rect 504 25621 506 25636
rect 336 25609 342 25621
rect 289 25544 308 25554
rect 300 25538 308 25544
rect 332 25575 342 25609
rect 400 25613 404 25621
rect 400 25579 408 25613
rect 434 25579 438 25613
rect 498 25611 506 25621
rect 514 25611 515 25631
rect 504 25595 506 25611
rect 525 25602 528 25636
rect 547 25611 548 25631
rect 557 25611 564 25621
rect 514 25595 530 25601
rect 532 25595 548 25601
rect 332 25547 373 25575
rect 332 25541 351 25547
rect 196 25500 204 25534
rect 216 25500 230 25534
rect 244 25500 257 25534
rect 278 25504 291 25538
rect 300 25522 321 25538
rect 336 25531 351 25541
rect 300 25520 312 25522
rect 300 25504 321 25520
rect 332 25513 351 25531
rect 361 25513 375 25547
rect 400 25541 411 25579
rect 562 25542 612 25544
rect 400 25513 409 25541
rect 466 25533 497 25535
rect 565 25533 596 25535
rect 442 25526 500 25533
rect 466 25525 500 25526
rect 565 25525 599 25533
rect 174 25463 181 25487
rect 224 25453 226 25500
rect 300 25491 308 25504
rect 289 25488 305 25490
rect 332 25463 342 25513
rect 400 25493 404 25513
rect 497 25509 500 25525
rect 596 25509 599 25525
rect 466 25508 500 25509
rect 442 25501 500 25508
rect 565 25501 599 25509
rect 612 25492 614 25542
rect 256 25453 328 25461
rect 336 25455 342 25463
rect 400 25455 404 25463
rect 196 25423 204 25453
rect 216 25423 230 25453
rect 196 25419 230 25423
rect 196 25411 226 25419
rect 224 25395 226 25411
rect 332 25383 336 25451
rect 400 25421 408 25455
rect 434 25421 438 25455
rect 454 25439 504 25441
rect 504 25423 506 25439
rect 514 25433 530 25439
rect 532 25433 548 25439
rect 525 25423 548 25432
rect 400 25413 404 25421
rect 498 25413 506 25423
rect 504 25389 506 25413
rect 514 25403 515 25423
rect 525 25398 528 25423
rect 547 25403 548 25423
rect 557 25413 564 25423
rect 514 25389 548 25393
rect 400 25383 442 25384
rect 174 25373 246 25381
rect 400 25376 404 25383
rect 295 25342 300 25376
rect 324 25342 329 25376
rect 367 25342 438 25376
rect 400 25341 404 25342
rect 378 25335 404 25341
rect 442 25335 464 25341
rect 38 25319 80 25335
rect 400 25319 442 25335
rect -25 25305 25 25307
rect 455 25305 505 25307
rect 557 25305 607 25307
rect 16 25297 102 25305
rect 378 25297 464 25305
rect 8 25263 17 25297
rect 18 25295 51 25297
rect 80 25295 100 25297
rect 18 25263 100 25295
rect 380 25295 404 25297
rect 429 25295 438 25297
rect 442 25295 462 25297
rect 16 25255 102 25263
rect 42 25239 76 25241
rect 16 25219 38 25225
rect 42 25216 76 25220
rect 80 25219 102 25225
rect 42 25186 46 25216
rect 72 25186 76 25216
rect 42 25105 46 25139
rect 72 25105 76 25139
rect -25 25068 25 25070
rect 0 25060 14 25061
rect 0 25059 17 25060
rect 25 25059 27 25068
rect 0 25052 38 25059
rect 0 25051 34 25052
rect 0 25035 8 25051
rect 14 25035 34 25051
rect 0 25034 34 25035
rect 0 25027 38 25034
rect 14 25026 17 25027
rect 25 25018 27 25027
rect 42 24998 45 25088
rect 69 25073 80 25105
rect 107 25073 143 25101
rect 107 25067 119 25073
rect 109 25039 119 25067
rect 129 25039 143 25073
rect 42 24947 46 24981
rect 72 24947 76 24981
rect 38 24909 80 24910
rect 42 24868 76 24902
rect 79 24868 113 24902
rect 42 24789 46 24823
rect 72 24789 76 24823
rect -25 24752 25 24754
rect 0 24744 14 24745
rect 0 24743 17 24744
rect 25 24743 27 24752
rect 0 24736 38 24743
rect 0 24735 34 24736
rect 0 24719 8 24735
rect 14 24719 34 24735
rect 0 24718 34 24719
rect 0 24711 38 24718
rect 14 24710 17 24711
rect 25 24702 27 24711
rect 42 24682 45 24772
rect 71 24741 80 24769
rect 69 24703 80 24741
rect 107 24697 119 24731
rect 129 24703 143 24731
rect 129 24697 141 24703
rect 42 24631 46 24665
rect 72 24631 76 24665
rect 42 24584 76 24588
rect 42 24554 46 24584
rect 72 24554 76 24584
rect 16 24545 38 24551
rect 80 24545 102 24551
rect 144 24545 148 25293
rect 332 25225 336 25293
rect 380 25263 462 25295
rect 463 25263 472 25297
rect 480 25263 497 25297
rect 378 25255 464 25263
rect 505 25255 507 25305
rect 514 25263 548 25297
rect 565 25263 582 25297
rect 607 25255 609 25305
rect 404 25239 438 25241
rect 400 25225 442 25226
rect 378 25219 404 25225
rect 442 25219 464 25225
rect 400 25218 404 25219
rect 174 25179 246 25187
rect 295 25184 300 25218
rect 324 25184 329 25218
rect 224 25149 226 25165
rect 196 25141 226 25149
rect 332 25147 336 25215
rect 367 25184 438 25218
rect 400 25177 404 25184
rect 454 25171 504 25173
rect 494 25167 548 25171
rect 494 25162 514 25167
rect 504 25147 506 25162
rect 196 25137 230 25141
rect 196 25107 204 25137
rect 216 25107 230 25137
rect 400 25139 404 25147
rect 174 25073 181 25099
rect 224 25060 226 25107
rect 256 25099 328 25107
rect 332 25105 336 25135
rect 400 25105 408 25139
rect 434 25105 438 25139
rect 498 25137 506 25147
rect 514 25137 515 25157
rect 504 25121 506 25137
rect 525 25128 528 25162
rect 547 25137 548 25157
rect 557 25137 564 25147
rect 514 25121 530 25127
rect 532 25121 548 25127
rect 289 25070 305 25072
rect 196 25026 204 25060
rect 216 25026 230 25060
rect 244 25026 257 25060
rect 300 25056 308 25069
rect 332 25067 342 25105
rect 400 25097 404 25105
rect 336 25057 342 25067
rect 224 24979 226 25026
rect 278 25022 291 25056
rect 300 25040 321 25056
rect 332 25047 342 25057
rect 400 25057 409 25085
rect 562 25068 612 25070
rect 466 25059 497 25061
rect 565 25059 596 25061
rect 300 25038 312 25040
rect 300 25022 321 25038
rect 300 25016 308 25022
rect 289 25006 308 25016
rect 196 24949 204 24979
rect 216 24949 230 24979
rect 196 24945 230 24949
rect 196 24937 226 24945
rect 300 24937 308 25006
rect 332 25013 351 25047
rect 361 25013 375 25047
rect 400 25013 411 25057
rect 442 25052 500 25059
rect 466 25051 500 25052
rect 565 25051 599 25059
rect 497 25035 500 25051
rect 596 25035 599 25051
rect 466 25034 500 25035
rect 442 25027 500 25034
rect 565 25027 599 25035
rect 612 25018 614 25068
rect 332 24989 342 25013
rect 336 24977 342 24989
rect 224 24921 226 24937
rect 332 24909 342 24977
rect 400 24981 404 24989
rect 400 24947 408 24981
rect 434 24947 438 24981
rect 454 24965 504 24967
rect 504 24949 506 24965
rect 514 24959 530 24965
rect 532 24959 548 24965
rect 525 24949 548 24958
rect 400 24939 404 24947
rect 498 24939 506 24949
rect 504 24915 506 24939
rect 514 24929 515 24949
rect 525 24924 528 24949
rect 547 24929 548 24949
rect 557 24939 564 24949
rect 514 24915 548 24919
rect 151 24868 156 24902
rect 174 24899 246 24907
rect 256 24899 328 24907
rect 336 24901 342 24909
rect 400 24904 404 24909
rect 180 24871 185 24899
rect 174 24863 246 24871
rect 256 24863 328 24871
rect 332 24869 336 24899
rect 400 24870 438 24904
rect 224 24833 226 24849
rect 196 24825 226 24833
rect 196 24821 230 24825
rect 196 24791 204 24821
rect 216 24791 230 24821
rect 224 24744 226 24791
rect 300 24764 308 24833
rect 332 24831 342 24869
rect 400 24861 404 24870
rect 454 24855 504 24857
rect 494 24851 548 24855
rect 494 24846 514 24851
rect 504 24831 506 24846
rect 336 24819 342 24831
rect 289 24754 308 24764
rect 300 24748 308 24754
rect 332 24785 342 24819
rect 400 24823 404 24831
rect 400 24789 408 24823
rect 434 24789 438 24823
rect 498 24821 506 24831
rect 514 24821 515 24841
rect 504 24805 506 24821
rect 525 24812 528 24846
rect 547 24821 548 24841
rect 557 24821 564 24831
rect 514 24805 530 24811
rect 532 24805 548 24811
rect 332 24757 373 24785
rect 332 24751 351 24757
rect 196 24710 204 24744
rect 216 24710 230 24744
rect 244 24710 257 24744
rect 278 24714 291 24748
rect 300 24732 321 24748
rect 336 24741 351 24751
rect 300 24730 312 24732
rect 300 24714 321 24730
rect 332 24723 351 24741
rect 361 24723 375 24757
rect 400 24751 411 24789
rect 562 24752 612 24754
rect 400 24723 409 24751
rect 466 24743 497 24745
rect 565 24743 596 24745
rect 442 24736 500 24743
rect 466 24735 500 24736
rect 565 24735 599 24743
rect 174 24673 181 24697
rect 224 24663 226 24710
rect 300 24701 308 24714
rect 289 24698 305 24700
rect 332 24673 342 24723
rect 400 24703 404 24723
rect 497 24719 500 24735
rect 596 24719 599 24735
rect 466 24718 500 24719
rect 442 24711 500 24718
rect 565 24711 599 24719
rect 612 24702 614 24752
rect 256 24663 328 24671
rect 336 24665 342 24673
rect 400 24665 404 24673
rect 196 24633 204 24663
rect 216 24633 230 24663
rect 196 24629 230 24633
rect 196 24621 226 24629
rect 224 24605 226 24621
rect 332 24593 336 24661
rect 400 24631 408 24665
rect 434 24631 438 24665
rect 454 24649 504 24651
rect 504 24633 506 24649
rect 514 24643 530 24649
rect 532 24643 548 24649
rect 525 24633 548 24642
rect 400 24623 404 24631
rect 498 24623 506 24633
rect 504 24599 506 24623
rect 514 24613 515 24633
rect 525 24608 528 24633
rect 547 24613 548 24633
rect 557 24623 564 24633
rect 514 24599 548 24603
rect 400 24593 442 24594
rect 174 24583 246 24591
rect 400 24586 404 24593
rect 295 24552 300 24586
rect 324 24552 329 24586
rect 367 24552 438 24586
rect 400 24551 404 24552
rect 378 24545 404 24551
rect 442 24545 464 24551
rect 38 24529 80 24545
rect 400 24529 442 24545
rect -25 24515 25 24517
rect 455 24515 505 24517
rect 557 24515 607 24517
rect 16 24507 102 24515
rect 378 24507 464 24515
rect 8 24473 17 24507
rect 18 24505 51 24507
rect 80 24505 100 24507
rect 18 24473 100 24505
rect 380 24505 404 24507
rect 429 24505 438 24507
rect 442 24505 462 24507
rect 16 24465 102 24473
rect 42 24449 76 24451
rect 16 24429 38 24435
rect 42 24426 76 24430
rect 80 24429 102 24435
rect 42 24396 46 24426
rect 72 24396 76 24426
rect 42 24315 46 24349
rect 72 24315 76 24349
rect -25 24278 25 24280
rect 0 24270 14 24271
rect 0 24269 17 24270
rect 25 24269 27 24278
rect 0 24262 38 24269
rect 0 24261 34 24262
rect 0 24245 8 24261
rect 14 24245 34 24261
rect 0 24244 34 24245
rect 0 24237 38 24244
rect 14 24236 17 24237
rect 25 24228 27 24237
rect 42 24208 45 24298
rect 69 24283 80 24315
rect 107 24283 143 24311
rect 107 24277 119 24283
rect 109 24249 119 24277
rect 129 24249 143 24283
rect 42 24157 46 24191
rect 72 24157 76 24191
rect 38 24119 80 24120
rect 42 24078 76 24112
rect 79 24078 113 24112
rect 42 23999 46 24033
rect 72 23999 76 24033
rect -25 23962 25 23964
rect 0 23954 14 23955
rect 0 23953 17 23954
rect 25 23953 27 23962
rect 0 23946 38 23953
rect 0 23945 34 23946
rect 0 23929 8 23945
rect 14 23929 34 23945
rect 0 23928 34 23929
rect 0 23921 38 23928
rect 14 23920 17 23921
rect 25 23912 27 23921
rect 42 23892 45 23982
rect 71 23951 80 23979
rect 69 23913 80 23951
rect 107 23907 119 23941
rect 129 23913 143 23941
rect 129 23907 141 23913
rect 42 23841 46 23875
rect 72 23841 76 23875
rect 42 23794 76 23798
rect 42 23764 46 23794
rect 72 23764 76 23794
rect 16 23755 38 23761
rect 80 23755 102 23761
rect 144 23755 148 24503
rect 332 24435 336 24503
rect 380 24473 462 24505
rect 463 24473 472 24507
rect 480 24473 497 24507
rect 378 24465 464 24473
rect 505 24465 507 24515
rect 514 24473 548 24507
rect 565 24473 582 24507
rect 607 24465 609 24515
rect 404 24449 438 24451
rect 400 24435 442 24436
rect 378 24429 404 24435
rect 442 24429 464 24435
rect 400 24428 404 24429
rect 174 24389 246 24397
rect 295 24394 300 24428
rect 324 24394 329 24428
rect 224 24359 226 24375
rect 196 24351 226 24359
rect 332 24357 336 24425
rect 367 24394 438 24428
rect 400 24387 404 24394
rect 454 24381 504 24383
rect 494 24377 548 24381
rect 494 24372 514 24377
rect 504 24357 506 24372
rect 196 24347 230 24351
rect 196 24317 204 24347
rect 216 24317 230 24347
rect 400 24349 404 24357
rect 174 24283 181 24309
rect 224 24270 226 24317
rect 256 24309 328 24317
rect 332 24315 336 24345
rect 400 24315 408 24349
rect 434 24315 438 24349
rect 498 24347 506 24357
rect 514 24347 515 24367
rect 504 24331 506 24347
rect 525 24338 528 24372
rect 547 24347 548 24367
rect 557 24347 564 24357
rect 514 24331 530 24337
rect 532 24331 548 24337
rect 289 24280 305 24282
rect 196 24236 204 24270
rect 216 24236 230 24270
rect 244 24236 257 24270
rect 300 24266 308 24279
rect 332 24277 342 24315
rect 400 24307 404 24315
rect 336 24267 342 24277
rect 224 24189 226 24236
rect 278 24232 291 24266
rect 300 24250 321 24266
rect 332 24257 342 24267
rect 400 24267 409 24295
rect 562 24278 612 24280
rect 466 24269 497 24271
rect 565 24269 596 24271
rect 300 24248 312 24250
rect 300 24232 321 24248
rect 300 24226 308 24232
rect 289 24216 308 24226
rect 196 24159 204 24189
rect 216 24159 230 24189
rect 196 24155 230 24159
rect 196 24147 226 24155
rect 300 24147 308 24216
rect 332 24223 351 24257
rect 361 24223 375 24257
rect 400 24223 411 24267
rect 442 24262 500 24269
rect 466 24261 500 24262
rect 565 24261 599 24269
rect 497 24245 500 24261
rect 596 24245 599 24261
rect 466 24244 500 24245
rect 442 24237 500 24244
rect 565 24237 599 24245
rect 612 24228 614 24278
rect 332 24199 342 24223
rect 336 24187 342 24199
rect 224 24131 226 24147
rect 332 24119 342 24187
rect 400 24191 404 24199
rect 400 24157 408 24191
rect 434 24157 438 24191
rect 454 24175 504 24177
rect 504 24159 506 24175
rect 514 24169 530 24175
rect 532 24169 548 24175
rect 525 24159 548 24168
rect 400 24149 404 24157
rect 498 24149 506 24159
rect 504 24125 506 24149
rect 514 24139 515 24159
rect 525 24134 528 24159
rect 547 24139 548 24159
rect 557 24149 564 24159
rect 514 24125 548 24129
rect 151 24078 156 24112
rect 174 24109 246 24117
rect 256 24109 328 24117
rect 336 24111 342 24119
rect 400 24114 404 24119
rect 180 24081 185 24109
rect 174 24073 246 24081
rect 256 24073 328 24081
rect 332 24079 336 24109
rect 400 24080 438 24114
rect 224 24043 226 24059
rect 196 24035 226 24043
rect 196 24031 230 24035
rect 196 24001 204 24031
rect 216 24001 230 24031
rect 224 23954 226 24001
rect 300 23974 308 24043
rect 332 24041 342 24079
rect 400 24071 404 24080
rect 454 24065 504 24067
rect 494 24061 548 24065
rect 494 24056 514 24061
rect 504 24041 506 24056
rect 336 24029 342 24041
rect 289 23964 308 23974
rect 300 23958 308 23964
rect 332 23995 342 24029
rect 400 24033 404 24041
rect 400 23999 408 24033
rect 434 23999 438 24033
rect 498 24031 506 24041
rect 514 24031 515 24051
rect 504 24015 506 24031
rect 525 24022 528 24056
rect 547 24031 548 24051
rect 557 24031 564 24041
rect 514 24015 530 24021
rect 532 24015 548 24021
rect 332 23967 373 23995
rect 332 23961 351 23967
rect 196 23920 204 23954
rect 216 23920 230 23954
rect 244 23920 257 23954
rect 278 23924 291 23958
rect 300 23942 321 23958
rect 336 23951 351 23961
rect 300 23940 312 23942
rect 300 23924 321 23940
rect 332 23933 351 23951
rect 361 23933 375 23967
rect 400 23961 411 23999
rect 562 23962 612 23964
rect 400 23933 409 23961
rect 466 23953 497 23955
rect 565 23953 596 23955
rect 442 23946 500 23953
rect 466 23945 500 23946
rect 565 23945 599 23953
rect 174 23883 181 23907
rect 224 23873 226 23920
rect 300 23911 308 23924
rect 289 23908 305 23910
rect 332 23883 342 23933
rect 400 23913 404 23933
rect 497 23929 500 23945
rect 596 23929 599 23945
rect 466 23928 500 23929
rect 442 23921 500 23928
rect 565 23921 599 23929
rect 612 23912 614 23962
rect 256 23873 328 23881
rect 336 23875 342 23883
rect 400 23875 404 23883
rect 196 23843 204 23873
rect 216 23843 230 23873
rect 196 23839 230 23843
rect 196 23831 226 23839
rect 224 23815 226 23831
rect 332 23803 336 23871
rect 400 23841 408 23875
rect 434 23841 438 23875
rect 454 23859 504 23861
rect 504 23843 506 23859
rect 514 23853 530 23859
rect 532 23853 548 23859
rect 525 23843 548 23852
rect 400 23833 404 23841
rect 498 23833 506 23843
rect 504 23809 506 23833
rect 514 23823 515 23843
rect 525 23818 528 23843
rect 547 23823 548 23843
rect 557 23833 564 23843
rect 514 23809 548 23813
rect 400 23803 442 23804
rect 174 23793 246 23801
rect 400 23796 404 23803
rect 295 23762 300 23796
rect 324 23762 329 23796
rect 367 23762 438 23796
rect 400 23761 404 23762
rect 378 23755 404 23761
rect 442 23755 464 23761
rect 38 23739 80 23755
rect 400 23739 442 23755
rect -25 23725 25 23727
rect 455 23725 505 23727
rect 557 23725 607 23727
rect 16 23717 102 23725
rect 378 23717 464 23725
rect 8 23683 17 23717
rect 18 23715 51 23717
rect 80 23715 100 23717
rect 18 23683 100 23715
rect 380 23715 404 23717
rect 429 23715 438 23717
rect 442 23715 462 23717
rect 16 23675 102 23683
rect 42 23659 76 23661
rect 16 23639 38 23645
rect 42 23636 76 23640
rect 80 23639 102 23645
rect 42 23606 46 23636
rect 72 23606 76 23636
rect 42 23525 46 23559
rect 72 23525 76 23559
rect -25 23488 25 23490
rect 0 23480 14 23481
rect 0 23479 17 23480
rect 25 23479 27 23488
rect 0 23472 38 23479
rect 0 23471 34 23472
rect 0 23455 8 23471
rect 14 23455 34 23471
rect 0 23454 34 23455
rect 0 23447 38 23454
rect 14 23446 17 23447
rect 25 23438 27 23447
rect 42 23418 45 23508
rect 69 23493 80 23525
rect 107 23493 143 23521
rect 107 23487 119 23493
rect 109 23459 119 23487
rect 129 23459 143 23493
rect 42 23367 46 23401
rect 72 23367 76 23401
rect 38 23329 80 23330
rect 42 23288 76 23322
rect 79 23288 113 23322
rect 42 23209 46 23243
rect 72 23209 76 23243
rect -25 23172 25 23174
rect 0 23164 14 23165
rect 0 23163 17 23164
rect 25 23163 27 23172
rect 0 23156 38 23163
rect 0 23155 34 23156
rect 0 23139 8 23155
rect 14 23139 34 23155
rect 0 23138 34 23139
rect 0 23131 38 23138
rect 14 23130 17 23131
rect 25 23122 27 23131
rect 42 23102 45 23192
rect 71 23161 80 23189
rect 69 23123 80 23161
rect 107 23117 119 23151
rect 129 23123 143 23151
rect 129 23117 141 23123
rect 42 23051 46 23085
rect 72 23051 76 23085
rect 42 23004 76 23008
rect 42 22974 46 23004
rect 72 22974 76 23004
rect 16 22965 38 22971
rect 80 22965 102 22971
rect 144 22965 148 23713
rect 332 23645 336 23713
rect 380 23683 462 23715
rect 463 23683 472 23717
rect 480 23683 497 23717
rect 378 23675 464 23683
rect 505 23675 507 23725
rect 514 23683 548 23717
rect 565 23683 582 23717
rect 607 23675 609 23725
rect 404 23659 438 23661
rect 400 23645 442 23646
rect 378 23639 404 23645
rect 442 23639 464 23645
rect 400 23638 404 23639
rect 174 23599 246 23607
rect 295 23604 300 23638
rect 324 23604 329 23638
rect 224 23569 226 23585
rect 196 23561 226 23569
rect 332 23567 336 23635
rect 367 23604 438 23638
rect 400 23597 404 23604
rect 454 23591 504 23593
rect 494 23587 548 23591
rect 494 23582 514 23587
rect 504 23567 506 23582
rect 196 23557 230 23561
rect 196 23527 204 23557
rect 216 23527 230 23557
rect 400 23559 404 23567
rect 174 23493 181 23519
rect 224 23480 226 23527
rect 256 23519 328 23527
rect 332 23525 336 23555
rect 400 23525 408 23559
rect 434 23525 438 23559
rect 498 23557 506 23567
rect 514 23557 515 23577
rect 504 23541 506 23557
rect 525 23548 528 23582
rect 547 23557 548 23577
rect 557 23557 564 23567
rect 514 23541 530 23547
rect 532 23541 548 23547
rect 289 23490 305 23492
rect 196 23446 204 23480
rect 216 23446 230 23480
rect 244 23446 257 23480
rect 300 23476 308 23489
rect 332 23487 342 23525
rect 400 23517 404 23525
rect 336 23477 342 23487
rect 224 23399 226 23446
rect 278 23442 291 23476
rect 300 23460 321 23476
rect 332 23467 342 23477
rect 400 23477 409 23505
rect 562 23488 612 23490
rect 466 23479 497 23481
rect 565 23479 596 23481
rect 300 23458 312 23460
rect 300 23442 321 23458
rect 300 23436 308 23442
rect 289 23426 308 23436
rect 196 23369 204 23399
rect 216 23369 230 23399
rect 196 23365 230 23369
rect 196 23357 226 23365
rect 300 23357 308 23426
rect 332 23433 351 23467
rect 361 23433 375 23467
rect 400 23433 411 23477
rect 442 23472 500 23479
rect 466 23471 500 23472
rect 565 23471 599 23479
rect 497 23455 500 23471
rect 596 23455 599 23471
rect 466 23454 500 23455
rect 442 23447 500 23454
rect 565 23447 599 23455
rect 612 23438 614 23488
rect 332 23409 342 23433
rect 336 23397 342 23409
rect 224 23341 226 23357
rect 332 23329 342 23397
rect 400 23401 404 23409
rect 400 23367 408 23401
rect 434 23367 438 23401
rect 454 23385 504 23387
rect 504 23369 506 23385
rect 514 23379 530 23385
rect 532 23379 548 23385
rect 525 23369 548 23378
rect 400 23359 404 23367
rect 498 23359 506 23369
rect 504 23335 506 23359
rect 514 23349 515 23369
rect 525 23344 528 23369
rect 547 23349 548 23369
rect 557 23359 564 23369
rect 514 23335 548 23339
rect 151 23288 156 23322
rect 174 23319 246 23327
rect 256 23319 328 23327
rect 336 23321 342 23329
rect 400 23324 404 23329
rect 180 23291 185 23319
rect 174 23283 246 23291
rect 256 23283 328 23291
rect 332 23289 336 23319
rect 400 23290 438 23324
rect 224 23253 226 23269
rect 196 23245 226 23253
rect 196 23241 230 23245
rect 196 23211 204 23241
rect 216 23211 230 23241
rect 224 23164 226 23211
rect 300 23184 308 23253
rect 332 23251 342 23289
rect 400 23281 404 23290
rect 454 23275 504 23277
rect 494 23271 548 23275
rect 494 23266 514 23271
rect 504 23251 506 23266
rect 336 23239 342 23251
rect 289 23174 308 23184
rect 300 23168 308 23174
rect 332 23205 342 23239
rect 400 23243 404 23251
rect 400 23209 408 23243
rect 434 23209 438 23243
rect 498 23241 506 23251
rect 514 23241 515 23261
rect 504 23225 506 23241
rect 525 23232 528 23266
rect 547 23241 548 23261
rect 557 23241 564 23251
rect 514 23225 530 23231
rect 532 23225 548 23231
rect 332 23177 373 23205
rect 332 23171 351 23177
rect 196 23130 204 23164
rect 216 23130 230 23164
rect 244 23130 257 23164
rect 278 23134 291 23168
rect 300 23152 321 23168
rect 336 23161 351 23171
rect 300 23150 312 23152
rect 300 23134 321 23150
rect 332 23143 351 23161
rect 361 23143 375 23177
rect 400 23171 411 23209
rect 562 23172 612 23174
rect 400 23143 409 23171
rect 466 23163 497 23165
rect 565 23163 596 23165
rect 442 23156 500 23163
rect 466 23155 500 23156
rect 565 23155 599 23163
rect 174 23093 181 23117
rect 224 23083 226 23130
rect 300 23121 308 23134
rect 289 23118 305 23120
rect 332 23093 342 23143
rect 400 23123 404 23143
rect 497 23139 500 23155
rect 596 23139 599 23155
rect 466 23138 500 23139
rect 442 23131 500 23138
rect 565 23131 599 23139
rect 612 23122 614 23172
rect 256 23083 328 23091
rect 336 23085 342 23093
rect 400 23085 404 23093
rect 196 23053 204 23083
rect 216 23053 230 23083
rect 196 23049 230 23053
rect 196 23041 226 23049
rect 224 23025 226 23041
rect 332 23013 336 23081
rect 400 23051 408 23085
rect 434 23051 438 23085
rect 454 23069 504 23071
rect 504 23053 506 23069
rect 514 23063 530 23069
rect 532 23063 548 23069
rect 525 23053 548 23062
rect 400 23043 404 23051
rect 498 23043 506 23053
rect 504 23019 506 23043
rect 514 23033 515 23053
rect 525 23028 528 23053
rect 547 23033 548 23053
rect 557 23043 564 23053
rect 514 23019 548 23023
rect 400 23013 442 23014
rect 174 23003 246 23011
rect 400 23006 404 23013
rect 295 22972 300 23006
rect 324 22972 329 23006
rect 367 22972 438 23006
rect 400 22971 404 22972
rect 378 22965 404 22971
rect 442 22965 464 22971
rect 38 22949 80 22965
rect 400 22949 442 22965
rect -25 22935 25 22937
rect 455 22935 505 22937
rect 557 22935 607 22937
rect 16 22927 102 22935
rect 378 22927 464 22935
rect 8 22893 17 22927
rect 18 22925 51 22927
rect 80 22925 100 22927
rect 18 22893 100 22925
rect 380 22925 404 22927
rect 429 22925 438 22927
rect 442 22925 462 22927
rect 16 22885 102 22893
rect 42 22869 76 22871
rect 16 22849 38 22855
rect 42 22846 76 22850
rect 80 22849 102 22855
rect 42 22816 46 22846
rect 72 22816 76 22846
rect 42 22735 46 22769
rect 72 22735 76 22769
rect -25 22698 25 22700
rect 0 22690 14 22691
rect 0 22689 17 22690
rect 25 22689 27 22698
rect 0 22682 38 22689
rect 0 22681 34 22682
rect 0 22665 8 22681
rect 14 22665 34 22681
rect 0 22664 34 22665
rect 0 22657 38 22664
rect 14 22656 17 22657
rect 25 22648 27 22657
rect 42 22628 45 22718
rect 69 22703 80 22735
rect 107 22703 143 22731
rect 107 22697 119 22703
rect 109 22669 119 22697
rect 129 22669 143 22703
rect 42 22577 46 22611
rect 72 22577 76 22611
rect 38 22539 80 22540
rect 42 22498 76 22532
rect 79 22498 113 22532
rect 42 22419 46 22453
rect 72 22419 76 22453
rect -25 22382 25 22384
rect 0 22374 14 22375
rect 0 22373 17 22374
rect 25 22373 27 22382
rect 0 22366 38 22373
rect 0 22365 34 22366
rect 0 22349 8 22365
rect 14 22349 34 22365
rect 0 22348 34 22349
rect 0 22341 38 22348
rect 14 22340 17 22341
rect 25 22332 27 22341
rect 42 22312 45 22402
rect 71 22371 80 22399
rect 69 22333 80 22371
rect 107 22327 119 22361
rect 129 22333 143 22361
rect 129 22327 141 22333
rect 42 22261 46 22295
rect 72 22261 76 22295
rect 42 22214 76 22218
rect 42 22184 46 22214
rect 72 22184 76 22214
rect 16 22175 38 22181
rect 80 22175 102 22181
rect 144 22175 148 22923
rect 332 22855 336 22923
rect 380 22893 462 22925
rect 463 22893 472 22927
rect 480 22893 497 22927
rect 378 22885 464 22893
rect 505 22885 507 22935
rect 514 22893 548 22927
rect 565 22893 582 22927
rect 607 22885 609 22935
rect 404 22869 438 22871
rect 400 22855 442 22856
rect 378 22849 404 22855
rect 442 22849 464 22855
rect 400 22848 404 22849
rect 174 22809 246 22817
rect 295 22814 300 22848
rect 324 22814 329 22848
rect 224 22779 226 22795
rect 196 22771 226 22779
rect 332 22777 336 22845
rect 367 22814 438 22848
rect 400 22807 404 22814
rect 454 22801 504 22803
rect 494 22797 548 22801
rect 494 22792 514 22797
rect 504 22777 506 22792
rect 196 22767 230 22771
rect 196 22737 204 22767
rect 216 22737 230 22767
rect 400 22769 404 22777
rect 174 22703 181 22729
rect 224 22690 226 22737
rect 256 22729 328 22737
rect 332 22735 336 22765
rect 400 22735 408 22769
rect 434 22735 438 22769
rect 498 22767 506 22777
rect 514 22767 515 22787
rect 504 22751 506 22767
rect 525 22758 528 22792
rect 547 22767 548 22787
rect 557 22767 564 22777
rect 514 22751 530 22757
rect 532 22751 548 22757
rect 289 22700 305 22702
rect 196 22656 204 22690
rect 216 22656 230 22690
rect 244 22656 257 22690
rect 300 22686 308 22699
rect 332 22697 342 22735
rect 400 22727 404 22735
rect 336 22687 342 22697
rect 224 22609 226 22656
rect 278 22652 291 22686
rect 300 22670 321 22686
rect 332 22677 342 22687
rect 400 22687 409 22715
rect 562 22698 612 22700
rect 466 22689 497 22691
rect 565 22689 596 22691
rect 300 22668 312 22670
rect 300 22652 321 22668
rect 300 22646 308 22652
rect 289 22636 308 22646
rect 196 22579 204 22609
rect 216 22579 230 22609
rect 196 22575 230 22579
rect 196 22567 226 22575
rect 300 22567 308 22636
rect 332 22643 351 22677
rect 361 22643 375 22677
rect 400 22643 411 22687
rect 442 22682 500 22689
rect 466 22681 500 22682
rect 565 22681 599 22689
rect 497 22665 500 22681
rect 596 22665 599 22681
rect 466 22664 500 22665
rect 442 22657 500 22664
rect 565 22657 599 22665
rect 612 22648 614 22698
rect 332 22619 342 22643
rect 336 22607 342 22619
rect 224 22551 226 22567
rect 332 22539 342 22607
rect 400 22611 404 22619
rect 400 22577 408 22611
rect 434 22577 438 22611
rect 454 22595 504 22597
rect 504 22579 506 22595
rect 514 22589 530 22595
rect 532 22589 548 22595
rect 525 22579 548 22588
rect 400 22569 404 22577
rect 498 22569 506 22579
rect 504 22545 506 22569
rect 514 22559 515 22579
rect 525 22554 528 22579
rect 547 22559 548 22579
rect 557 22569 564 22579
rect 514 22545 548 22549
rect 151 22498 156 22532
rect 174 22529 246 22537
rect 256 22529 328 22537
rect 336 22531 342 22539
rect 400 22534 404 22539
rect 180 22501 185 22529
rect 174 22493 246 22501
rect 256 22493 328 22501
rect 332 22499 336 22529
rect 400 22500 438 22534
rect 224 22463 226 22479
rect 196 22455 226 22463
rect 196 22451 230 22455
rect 196 22421 204 22451
rect 216 22421 230 22451
rect 224 22374 226 22421
rect 300 22394 308 22463
rect 332 22461 342 22499
rect 400 22491 404 22500
rect 454 22485 504 22487
rect 494 22481 548 22485
rect 494 22476 514 22481
rect 504 22461 506 22476
rect 336 22449 342 22461
rect 289 22384 308 22394
rect 300 22378 308 22384
rect 332 22415 342 22449
rect 400 22453 404 22461
rect 400 22419 408 22453
rect 434 22419 438 22453
rect 498 22451 506 22461
rect 514 22451 515 22471
rect 504 22435 506 22451
rect 525 22442 528 22476
rect 547 22451 548 22471
rect 557 22451 564 22461
rect 514 22435 530 22441
rect 532 22435 548 22441
rect 332 22387 373 22415
rect 332 22381 351 22387
rect 196 22340 204 22374
rect 216 22340 230 22374
rect 244 22340 257 22374
rect 278 22344 291 22378
rect 300 22362 321 22378
rect 336 22371 351 22381
rect 300 22360 312 22362
rect 300 22344 321 22360
rect 332 22353 351 22371
rect 361 22353 375 22387
rect 400 22381 411 22419
rect 562 22382 612 22384
rect 400 22353 409 22381
rect 466 22373 497 22375
rect 565 22373 596 22375
rect 442 22366 500 22373
rect 466 22365 500 22366
rect 565 22365 599 22373
rect 174 22303 181 22327
rect 224 22293 226 22340
rect 300 22331 308 22344
rect 289 22328 305 22330
rect 332 22303 342 22353
rect 400 22333 404 22353
rect 497 22349 500 22365
rect 596 22349 599 22365
rect 466 22348 500 22349
rect 442 22341 500 22348
rect 565 22341 599 22349
rect 612 22332 614 22382
rect 256 22293 328 22301
rect 336 22295 342 22303
rect 400 22295 404 22303
rect 196 22263 204 22293
rect 216 22263 230 22293
rect 196 22259 230 22263
rect 196 22251 226 22259
rect 224 22235 226 22251
rect 332 22223 336 22291
rect 400 22261 408 22295
rect 434 22261 438 22295
rect 454 22279 504 22281
rect 504 22263 506 22279
rect 514 22273 530 22279
rect 532 22273 548 22279
rect 525 22263 548 22272
rect 400 22253 404 22261
rect 498 22253 506 22263
rect 504 22229 506 22253
rect 514 22243 515 22263
rect 525 22238 528 22263
rect 547 22243 548 22263
rect 557 22253 564 22263
rect 514 22229 548 22233
rect 400 22223 442 22224
rect 174 22213 246 22221
rect 400 22216 404 22223
rect 295 22182 300 22216
rect 324 22182 329 22216
rect 367 22182 438 22216
rect 400 22181 404 22182
rect 378 22175 404 22181
rect 442 22175 464 22181
rect 38 22159 80 22175
rect 400 22159 442 22175
rect -25 22145 25 22147
rect 455 22145 505 22147
rect 557 22145 607 22147
rect 16 22137 102 22145
rect 378 22137 464 22145
rect 8 22103 17 22137
rect 18 22135 51 22137
rect 80 22135 100 22137
rect 18 22103 100 22135
rect 380 22135 404 22137
rect 429 22135 438 22137
rect 442 22135 462 22137
rect 16 22095 102 22103
rect 42 22079 76 22081
rect 16 22059 38 22065
rect 42 22056 76 22060
rect 80 22059 102 22065
rect 42 22026 46 22056
rect 72 22026 76 22056
rect 42 21945 46 21979
rect 72 21945 76 21979
rect -25 21908 25 21910
rect 0 21900 14 21901
rect 0 21899 17 21900
rect 25 21899 27 21908
rect 0 21892 38 21899
rect 0 21891 34 21892
rect 0 21875 8 21891
rect 14 21875 34 21891
rect 0 21874 34 21875
rect 0 21867 38 21874
rect 14 21866 17 21867
rect 25 21858 27 21867
rect 42 21838 45 21928
rect 69 21913 80 21945
rect 107 21913 143 21941
rect 107 21907 119 21913
rect 109 21879 119 21907
rect 129 21879 143 21913
rect 42 21787 46 21821
rect 72 21787 76 21821
rect 38 21749 80 21750
rect 42 21708 76 21742
rect 79 21708 113 21742
rect 42 21629 46 21663
rect 72 21629 76 21663
rect -25 21592 25 21594
rect 0 21584 14 21585
rect 0 21583 17 21584
rect 25 21583 27 21592
rect 0 21576 38 21583
rect 0 21575 34 21576
rect 0 21559 8 21575
rect 14 21559 34 21575
rect 0 21558 34 21559
rect 0 21551 38 21558
rect 14 21550 17 21551
rect 25 21542 27 21551
rect 42 21522 45 21612
rect 71 21581 80 21609
rect 69 21543 80 21581
rect 107 21537 119 21571
rect 129 21543 143 21571
rect 129 21537 141 21543
rect 42 21471 46 21505
rect 72 21471 76 21505
rect 42 21424 76 21428
rect 42 21394 46 21424
rect 72 21394 76 21424
rect 16 21385 38 21391
rect 80 21385 102 21391
rect 144 21385 148 22133
rect 332 22065 336 22133
rect 380 22103 462 22135
rect 463 22103 472 22137
rect 480 22103 497 22137
rect 378 22095 464 22103
rect 505 22095 507 22145
rect 514 22103 548 22137
rect 565 22103 582 22137
rect 607 22095 609 22145
rect 404 22079 438 22081
rect 400 22065 442 22066
rect 378 22059 404 22065
rect 442 22059 464 22065
rect 400 22058 404 22059
rect 174 22019 246 22027
rect 295 22024 300 22058
rect 324 22024 329 22058
rect 224 21989 226 22005
rect 196 21981 226 21989
rect 332 21987 336 22055
rect 367 22024 438 22058
rect 400 22017 404 22024
rect 454 22011 504 22013
rect 494 22007 548 22011
rect 494 22002 514 22007
rect 504 21987 506 22002
rect 196 21977 230 21981
rect 196 21947 204 21977
rect 216 21947 230 21977
rect 400 21979 404 21987
rect 174 21913 181 21939
rect 224 21900 226 21947
rect 256 21939 328 21947
rect 332 21945 336 21975
rect 400 21945 408 21979
rect 434 21945 438 21979
rect 498 21977 506 21987
rect 514 21977 515 21997
rect 504 21961 506 21977
rect 525 21968 528 22002
rect 547 21977 548 21997
rect 557 21977 564 21987
rect 514 21961 530 21967
rect 532 21961 548 21967
rect 289 21910 305 21912
rect 196 21866 204 21900
rect 216 21866 230 21900
rect 244 21866 257 21900
rect 300 21896 308 21909
rect 332 21907 342 21945
rect 400 21937 404 21945
rect 336 21897 342 21907
rect 224 21819 226 21866
rect 278 21862 291 21896
rect 300 21880 321 21896
rect 332 21887 342 21897
rect 400 21897 409 21925
rect 562 21908 612 21910
rect 466 21899 497 21901
rect 565 21899 596 21901
rect 300 21878 312 21880
rect 300 21862 321 21878
rect 300 21856 308 21862
rect 289 21846 308 21856
rect 196 21789 204 21819
rect 216 21789 230 21819
rect 196 21785 230 21789
rect 196 21777 226 21785
rect 300 21777 308 21846
rect 332 21853 351 21887
rect 361 21853 375 21887
rect 400 21853 411 21897
rect 442 21892 500 21899
rect 466 21891 500 21892
rect 565 21891 599 21899
rect 497 21875 500 21891
rect 596 21875 599 21891
rect 466 21874 500 21875
rect 442 21867 500 21874
rect 565 21867 599 21875
rect 612 21858 614 21908
rect 332 21829 342 21853
rect 336 21817 342 21829
rect 224 21761 226 21777
rect 332 21749 342 21817
rect 400 21821 404 21829
rect 400 21787 408 21821
rect 434 21787 438 21821
rect 454 21805 504 21807
rect 504 21789 506 21805
rect 514 21799 530 21805
rect 532 21799 548 21805
rect 525 21789 548 21798
rect 400 21779 404 21787
rect 498 21779 506 21789
rect 504 21755 506 21779
rect 514 21769 515 21789
rect 525 21764 528 21789
rect 547 21769 548 21789
rect 557 21779 564 21789
rect 514 21755 548 21759
rect 151 21708 156 21742
rect 174 21739 246 21747
rect 256 21739 328 21747
rect 336 21741 342 21749
rect 400 21744 404 21749
rect 180 21711 185 21739
rect 174 21703 246 21711
rect 256 21703 328 21711
rect 332 21709 336 21739
rect 400 21710 438 21744
rect 224 21673 226 21689
rect 196 21665 226 21673
rect 196 21661 230 21665
rect 196 21631 204 21661
rect 216 21631 230 21661
rect 224 21584 226 21631
rect 300 21604 308 21673
rect 332 21671 342 21709
rect 400 21701 404 21710
rect 454 21695 504 21697
rect 494 21691 548 21695
rect 494 21686 514 21691
rect 504 21671 506 21686
rect 336 21659 342 21671
rect 289 21594 308 21604
rect 300 21588 308 21594
rect 332 21625 342 21659
rect 400 21663 404 21671
rect 400 21629 408 21663
rect 434 21629 438 21663
rect 498 21661 506 21671
rect 514 21661 515 21681
rect 504 21645 506 21661
rect 525 21652 528 21686
rect 547 21661 548 21681
rect 557 21661 564 21671
rect 514 21645 530 21651
rect 532 21645 548 21651
rect 332 21597 373 21625
rect 332 21591 351 21597
rect 196 21550 204 21584
rect 216 21550 230 21584
rect 244 21550 257 21584
rect 278 21554 291 21588
rect 300 21572 321 21588
rect 336 21581 351 21591
rect 300 21570 312 21572
rect 300 21554 321 21570
rect 332 21563 351 21581
rect 361 21563 375 21597
rect 400 21591 411 21629
rect 562 21592 612 21594
rect 400 21563 409 21591
rect 466 21583 497 21585
rect 565 21583 596 21585
rect 442 21576 500 21583
rect 466 21575 500 21576
rect 565 21575 599 21583
rect 174 21513 181 21537
rect 224 21503 226 21550
rect 300 21541 308 21554
rect 289 21538 305 21540
rect 332 21513 342 21563
rect 400 21543 404 21563
rect 497 21559 500 21575
rect 596 21559 599 21575
rect 466 21558 500 21559
rect 442 21551 500 21558
rect 565 21551 599 21559
rect 612 21542 614 21592
rect 256 21503 328 21511
rect 336 21505 342 21513
rect 400 21505 404 21513
rect 196 21473 204 21503
rect 216 21473 230 21503
rect 196 21469 230 21473
rect 196 21461 226 21469
rect 224 21445 226 21461
rect 332 21433 336 21501
rect 400 21471 408 21505
rect 434 21471 438 21505
rect 454 21489 504 21491
rect 504 21473 506 21489
rect 514 21483 530 21489
rect 532 21483 548 21489
rect 525 21473 548 21482
rect 400 21463 404 21471
rect 498 21463 506 21473
rect 504 21439 506 21463
rect 514 21453 515 21473
rect 525 21448 528 21473
rect 547 21453 548 21473
rect 557 21463 564 21473
rect 514 21439 548 21443
rect 400 21433 442 21434
rect 174 21423 246 21431
rect 400 21426 404 21433
rect 295 21392 300 21426
rect 324 21392 329 21426
rect 367 21392 438 21426
rect 400 21391 404 21392
rect 378 21385 404 21391
rect 442 21385 464 21391
rect 38 21369 80 21385
rect 400 21369 442 21385
rect -25 21355 25 21357
rect 455 21355 505 21357
rect 557 21355 607 21357
rect 16 21347 102 21355
rect 378 21347 464 21355
rect 8 21313 17 21347
rect 18 21345 51 21347
rect 80 21345 100 21347
rect 18 21313 100 21345
rect 380 21345 404 21347
rect 429 21345 438 21347
rect 442 21345 462 21347
rect 16 21305 102 21313
rect 42 21289 76 21291
rect 16 21269 38 21275
rect 42 21266 76 21270
rect 80 21269 102 21275
rect 42 21236 46 21266
rect 72 21236 76 21266
rect 42 21155 46 21189
rect 72 21155 76 21189
rect -25 21118 25 21120
rect 0 21110 14 21111
rect 0 21109 17 21110
rect 25 21109 27 21118
rect 0 21102 38 21109
rect 0 21101 34 21102
rect 0 21085 8 21101
rect 14 21085 34 21101
rect 0 21084 34 21085
rect 0 21077 38 21084
rect 14 21076 17 21077
rect 25 21068 27 21077
rect 42 21048 45 21138
rect 69 21123 80 21155
rect 107 21123 143 21151
rect 107 21117 119 21123
rect 109 21089 119 21117
rect 129 21089 143 21123
rect 42 20997 46 21031
rect 72 20997 76 21031
rect 38 20959 80 20960
rect 42 20918 76 20952
rect 79 20918 113 20952
rect 42 20839 46 20873
rect 72 20839 76 20873
rect -25 20802 25 20804
rect 0 20794 14 20795
rect 0 20793 17 20794
rect 25 20793 27 20802
rect 0 20786 38 20793
rect 0 20785 34 20786
rect 0 20769 8 20785
rect 14 20769 34 20785
rect 0 20768 34 20769
rect 0 20761 38 20768
rect 14 20760 17 20761
rect 25 20752 27 20761
rect 42 20732 45 20822
rect 71 20791 80 20819
rect 69 20753 80 20791
rect 107 20747 119 20781
rect 129 20753 143 20781
rect 129 20747 141 20753
rect 42 20681 46 20715
rect 72 20681 76 20715
rect 42 20634 76 20638
rect 42 20604 46 20634
rect 72 20604 76 20634
rect 16 20595 38 20601
rect 80 20595 102 20601
rect 144 20595 148 21343
rect 332 21275 336 21343
rect 380 21313 462 21345
rect 463 21313 472 21347
rect 480 21313 497 21347
rect 378 21305 464 21313
rect 505 21305 507 21355
rect 514 21313 548 21347
rect 565 21313 582 21347
rect 607 21305 609 21355
rect 404 21289 438 21291
rect 400 21275 442 21276
rect 378 21269 404 21275
rect 442 21269 464 21275
rect 400 21268 404 21269
rect 174 21229 246 21237
rect 295 21234 300 21268
rect 324 21234 329 21268
rect 224 21199 226 21215
rect 196 21191 226 21199
rect 332 21197 336 21265
rect 367 21234 438 21268
rect 400 21227 404 21234
rect 454 21221 504 21223
rect 494 21217 548 21221
rect 494 21212 514 21217
rect 504 21197 506 21212
rect 196 21187 230 21191
rect 196 21157 204 21187
rect 216 21157 230 21187
rect 400 21189 404 21197
rect 174 21123 181 21149
rect 224 21110 226 21157
rect 256 21149 328 21157
rect 332 21155 336 21185
rect 400 21155 408 21189
rect 434 21155 438 21189
rect 498 21187 506 21197
rect 514 21187 515 21207
rect 504 21171 506 21187
rect 525 21178 528 21212
rect 547 21187 548 21207
rect 557 21187 564 21197
rect 514 21171 530 21177
rect 532 21171 548 21177
rect 289 21120 305 21122
rect 196 21076 204 21110
rect 216 21076 230 21110
rect 244 21076 257 21110
rect 300 21106 308 21119
rect 332 21117 342 21155
rect 400 21147 404 21155
rect 336 21107 342 21117
rect 224 21029 226 21076
rect 278 21072 291 21106
rect 300 21090 321 21106
rect 332 21097 342 21107
rect 400 21107 409 21135
rect 562 21118 612 21120
rect 466 21109 497 21111
rect 565 21109 596 21111
rect 300 21088 312 21090
rect 300 21072 321 21088
rect 300 21066 308 21072
rect 289 21056 308 21066
rect 196 20999 204 21029
rect 216 20999 230 21029
rect 196 20995 230 20999
rect 196 20987 226 20995
rect 300 20987 308 21056
rect 332 21063 351 21097
rect 361 21063 375 21097
rect 400 21063 411 21107
rect 442 21102 500 21109
rect 466 21101 500 21102
rect 565 21101 599 21109
rect 497 21085 500 21101
rect 596 21085 599 21101
rect 466 21084 500 21085
rect 442 21077 500 21084
rect 565 21077 599 21085
rect 612 21068 614 21118
rect 332 21039 342 21063
rect 336 21027 342 21039
rect 224 20971 226 20987
rect 332 20959 342 21027
rect 400 21031 404 21039
rect 400 20997 408 21031
rect 434 20997 438 21031
rect 454 21015 504 21017
rect 504 20999 506 21015
rect 514 21009 530 21015
rect 532 21009 548 21015
rect 525 20999 548 21008
rect 400 20989 404 20997
rect 498 20989 506 20999
rect 504 20965 506 20989
rect 514 20979 515 20999
rect 525 20974 528 20999
rect 547 20979 548 20999
rect 557 20989 564 20999
rect 514 20965 548 20969
rect 151 20918 156 20952
rect 174 20949 246 20957
rect 256 20949 328 20957
rect 336 20951 342 20959
rect 400 20954 404 20959
rect 180 20921 185 20949
rect 174 20913 246 20921
rect 256 20913 328 20921
rect 332 20919 336 20949
rect 400 20920 438 20954
rect 224 20883 226 20899
rect 196 20875 226 20883
rect 196 20871 230 20875
rect 196 20841 204 20871
rect 216 20841 230 20871
rect 224 20794 226 20841
rect 300 20814 308 20883
rect 332 20881 342 20919
rect 400 20911 404 20920
rect 454 20905 504 20907
rect 494 20901 548 20905
rect 494 20896 514 20901
rect 504 20881 506 20896
rect 336 20869 342 20881
rect 289 20804 308 20814
rect 300 20798 308 20804
rect 332 20835 342 20869
rect 400 20873 404 20881
rect 400 20839 408 20873
rect 434 20839 438 20873
rect 498 20871 506 20881
rect 514 20871 515 20891
rect 504 20855 506 20871
rect 525 20862 528 20896
rect 547 20871 548 20891
rect 557 20871 564 20881
rect 514 20855 530 20861
rect 532 20855 548 20861
rect 332 20807 373 20835
rect 332 20801 351 20807
rect 196 20760 204 20794
rect 216 20760 230 20794
rect 244 20760 257 20794
rect 278 20764 291 20798
rect 300 20782 321 20798
rect 336 20791 351 20801
rect 300 20780 312 20782
rect 300 20764 321 20780
rect 332 20773 351 20791
rect 361 20773 375 20807
rect 400 20801 411 20839
rect 562 20802 612 20804
rect 400 20773 409 20801
rect 466 20793 497 20795
rect 565 20793 596 20795
rect 442 20786 500 20793
rect 466 20785 500 20786
rect 565 20785 599 20793
rect 174 20723 181 20747
rect 224 20713 226 20760
rect 300 20751 308 20764
rect 289 20748 305 20750
rect 332 20723 342 20773
rect 400 20753 404 20773
rect 497 20769 500 20785
rect 596 20769 599 20785
rect 466 20768 500 20769
rect 442 20761 500 20768
rect 565 20761 599 20769
rect 612 20752 614 20802
rect 256 20713 328 20721
rect 336 20715 342 20723
rect 400 20715 404 20723
rect 196 20683 204 20713
rect 216 20683 230 20713
rect 196 20679 230 20683
rect 196 20671 226 20679
rect 224 20655 226 20671
rect 332 20643 336 20711
rect 400 20681 408 20715
rect 434 20681 438 20715
rect 454 20699 504 20701
rect 504 20683 506 20699
rect 514 20693 530 20699
rect 532 20693 548 20699
rect 525 20683 548 20692
rect 400 20673 404 20681
rect 498 20673 506 20683
rect 504 20649 506 20673
rect 514 20663 515 20683
rect 525 20658 528 20683
rect 547 20663 548 20683
rect 557 20673 564 20683
rect 514 20649 548 20653
rect 400 20643 442 20644
rect 174 20633 246 20641
rect 400 20636 404 20643
rect 295 20602 300 20636
rect 324 20602 329 20636
rect 367 20602 438 20636
rect 400 20601 404 20602
rect 378 20595 404 20601
rect 442 20595 464 20601
rect 38 20579 80 20595
rect 400 20579 442 20595
rect -25 20565 25 20567
rect 455 20565 505 20567
rect 557 20565 607 20567
rect 16 20557 102 20565
rect 378 20557 464 20565
rect 8 20523 17 20557
rect 18 20555 51 20557
rect 80 20555 100 20557
rect 18 20523 100 20555
rect 380 20555 404 20557
rect 429 20555 438 20557
rect 442 20555 462 20557
rect 16 20515 102 20523
rect 42 20499 76 20501
rect 16 20479 38 20485
rect 42 20476 76 20480
rect 80 20479 102 20485
rect 42 20446 46 20476
rect 72 20446 76 20476
rect 42 20365 46 20399
rect 72 20365 76 20399
rect -25 20328 25 20330
rect 0 20320 14 20321
rect 0 20319 17 20320
rect 25 20319 27 20328
rect 0 20312 38 20319
rect 0 20311 34 20312
rect 0 20295 8 20311
rect 14 20295 34 20311
rect 0 20294 34 20295
rect 0 20287 38 20294
rect 14 20286 17 20287
rect 25 20278 27 20287
rect 42 20258 45 20348
rect 69 20333 80 20365
rect 107 20333 143 20361
rect 107 20327 119 20333
rect 109 20299 119 20327
rect 129 20299 143 20333
rect 42 20207 46 20241
rect 72 20207 76 20241
rect 38 20169 80 20170
rect 42 20128 76 20162
rect 79 20128 113 20162
rect 42 20049 46 20083
rect 72 20049 76 20083
rect -25 20012 25 20014
rect 0 20004 14 20005
rect 0 20003 17 20004
rect 25 20003 27 20012
rect 0 19996 38 20003
rect 0 19995 34 19996
rect 0 19979 8 19995
rect 14 19979 34 19995
rect 0 19978 34 19979
rect 0 19971 38 19978
rect 14 19970 17 19971
rect 25 19962 27 19971
rect 42 19942 45 20032
rect 71 20001 80 20029
rect 69 19963 80 20001
rect 107 19957 119 19991
rect 129 19963 143 19991
rect 129 19957 141 19963
rect 42 19891 46 19925
rect 72 19891 76 19925
rect 42 19844 76 19848
rect 42 19814 46 19844
rect 72 19814 76 19844
rect 16 19805 38 19811
rect 80 19805 102 19811
rect 144 19805 148 20553
rect 332 20485 336 20553
rect 380 20523 462 20555
rect 463 20523 472 20557
rect 480 20523 497 20557
rect 378 20515 464 20523
rect 505 20515 507 20565
rect 514 20523 548 20557
rect 565 20523 582 20557
rect 607 20515 609 20565
rect 404 20499 438 20501
rect 400 20485 442 20486
rect 378 20479 404 20485
rect 442 20479 464 20485
rect 400 20478 404 20479
rect 174 20439 246 20447
rect 295 20444 300 20478
rect 324 20444 329 20478
rect 224 20409 226 20425
rect 196 20401 226 20409
rect 332 20407 336 20475
rect 367 20444 438 20478
rect 400 20437 404 20444
rect 454 20431 504 20433
rect 494 20427 548 20431
rect 494 20422 514 20427
rect 504 20407 506 20422
rect 196 20397 230 20401
rect 196 20367 204 20397
rect 216 20367 230 20397
rect 400 20399 404 20407
rect 174 20333 181 20359
rect 224 20320 226 20367
rect 256 20359 328 20367
rect 332 20365 336 20395
rect 400 20365 408 20399
rect 434 20365 438 20399
rect 498 20397 506 20407
rect 514 20397 515 20417
rect 504 20381 506 20397
rect 525 20388 528 20422
rect 547 20397 548 20417
rect 557 20397 564 20407
rect 514 20381 530 20387
rect 532 20381 548 20387
rect 289 20330 305 20332
rect 196 20286 204 20320
rect 216 20286 230 20320
rect 244 20286 257 20320
rect 300 20316 308 20329
rect 332 20327 342 20365
rect 400 20357 404 20365
rect 336 20317 342 20327
rect 224 20239 226 20286
rect 278 20282 291 20316
rect 300 20300 321 20316
rect 332 20307 342 20317
rect 400 20317 409 20345
rect 562 20328 612 20330
rect 466 20319 497 20321
rect 565 20319 596 20321
rect 300 20298 312 20300
rect 300 20282 321 20298
rect 300 20276 308 20282
rect 289 20266 308 20276
rect 196 20209 204 20239
rect 216 20209 230 20239
rect 196 20205 230 20209
rect 196 20197 226 20205
rect 300 20197 308 20266
rect 332 20273 351 20307
rect 361 20273 375 20307
rect 400 20273 411 20317
rect 442 20312 500 20319
rect 466 20311 500 20312
rect 565 20311 599 20319
rect 497 20295 500 20311
rect 596 20295 599 20311
rect 466 20294 500 20295
rect 442 20287 500 20294
rect 565 20287 599 20295
rect 612 20278 614 20328
rect 332 20249 342 20273
rect 336 20237 342 20249
rect 224 20181 226 20197
rect 332 20169 342 20237
rect 400 20241 404 20249
rect 400 20207 408 20241
rect 434 20207 438 20241
rect 454 20225 504 20227
rect 504 20209 506 20225
rect 514 20219 530 20225
rect 532 20219 548 20225
rect 525 20209 548 20218
rect 400 20199 404 20207
rect 498 20199 506 20209
rect 504 20175 506 20199
rect 514 20189 515 20209
rect 525 20184 528 20209
rect 547 20189 548 20209
rect 557 20199 564 20209
rect 514 20175 548 20179
rect 151 20128 156 20162
rect 174 20159 246 20167
rect 256 20159 328 20167
rect 336 20161 342 20169
rect 400 20164 404 20169
rect 180 20131 185 20159
rect 174 20123 246 20131
rect 256 20123 328 20131
rect 332 20129 336 20159
rect 400 20130 438 20164
rect 224 20093 226 20109
rect 196 20085 226 20093
rect 196 20081 230 20085
rect 196 20051 204 20081
rect 216 20051 230 20081
rect 224 20004 226 20051
rect 300 20024 308 20093
rect 332 20091 342 20129
rect 400 20121 404 20130
rect 454 20115 504 20117
rect 494 20111 548 20115
rect 494 20106 514 20111
rect 504 20091 506 20106
rect 336 20079 342 20091
rect 289 20014 308 20024
rect 300 20008 308 20014
rect 332 20045 342 20079
rect 400 20083 404 20091
rect 400 20049 408 20083
rect 434 20049 438 20083
rect 498 20081 506 20091
rect 514 20081 515 20101
rect 504 20065 506 20081
rect 525 20072 528 20106
rect 547 20081 548 20101
rect 557 20081 564 20091
rect 514 20065 530 20071
rect 532 20065 548 20071
rect 332 20017 373 20045
rect 332 20011 351 20017
rect 196 19970 204 20004
rect 216 19970 230 20004
rect 244 19970 257 20004
rect 278 19974 291 20008
rect 300 19992 321 20008
rect 336 20001 351 20011
rect 300 19990 312 19992
rect 300 19974 321 19990
rect 332 19983 351 20001
rect 361 19983 375 20017
rect 400 20011 411 20049
rect 562 20012 612 20014
rect 400 19983 409 20011
rect 466 20003 497 20005
rect 565 20003 596 20005
rect 442 19996 500 20003
rect 466 19995 500 19996
rect 565 19995 599 20003
rect 174 19933 181 19957
rect 224 19923 226 19970
rect 300 19961 308 19974
rect 289 19958 305 19960
rect 332 19933 342 19983
rect 400 19963 404 19983
rect 497 19979 500 19995
rect 596 19979 599 19995
rect 466 19978 500 19979
rect 442 19971 500 19978
rect 565 19971 599 19979
rect 612 19962 614 20012
rect 256 19923 328 19931
rect 336 19925 342 19933
rect 400 19925 404 19933
rect 196 19893 204 19923
rect 216 19893 230 19923
rect 196 19889 230 19893
rect 196 19881 226 19889
rect 224 19865 226 19881
rect 332 19853 336 19921
rect 400 19891 408 19925
rect 434 19891 438 19925
rect 454 19909 504 19911
rect 504 19893 506 19909
rect 514 19903 530 19909
rect 532 19903 548 19909
rect 525 19893 548 19902
rect 400 19883 404 19891
rect 498 19883 506 19893
rect 504 19859 506 19883
rect 514 19873 515 19893
rect 525 19868 528 19893
rect 547 19873 548 19893
rect 557 19883 564 19893
rect 514 19859 548 19863
rect 400 19853 442 19854
rect 174 19843 246 19851
rect 400 19846 404 19853
rect 295 19812 300 19846
rect 324 19812 329 19846
rect 367 19812 438 19846
rect 400 19811 404 19812
rect 378 19805 404 19811
rect 442 19805 464 19811
rect 38 19789 80 19805
rect 400 19789 442 19805
rect -25 19775 25 19777
rect 455 19775 505 19777
rect 557 19775 607 19777
rect 16 19767 102 19775
rect 378 19767 464 19775
rect 8 19733 17 19767
rect 18 19765 51 19767
rect 80 19765 100 19767
rect 18 19733 100 19765
rect 380 19765 404 19767
rect 429 19765 438 19767
rect 442 19765 462 19767
rect 16 19725 102 19733
rect 42 19709 76 19711
rect 16 19689 38 19695
rect 42 19686 76 19690
rect 80 19689 102 19695
rect 42 19656 46 19686
rect 72 19656 76 19686
rect 42 19575 46 19609
rect 72 19575 76 19609
rect -25 19538 25 19540
rect 0 19530 14 19531
rect 0 19529 17 19530
rect 25 19529 27 19538
rect 0 19522 38 19529
rect 0 19521 34 19522
rect 0 19505 8 19521
rect 14 19505 34 19521
rect 0 19504 34 19505
rect 0 19497 38 19504
rect 14 19496 17 19497
rect 25 19488 27 19497
rect 42 19468 45 19558
rect 69 19543 80 19575
rect 107 19543 143 19571
rect 107 19537 119 19543
rect 109 19509 119 19537
rect 129 19509 143 19543
rect 42 19417 46 19451
rect 72 19417 76 19451
rect 38 19379 80 19380
rect 42 19338 76 19372
rect 79 19338 113 19372
rect 42 19259 46 19293
rect 72 19259 76 19293
rect -25 19222 25 19224
rect 0 19214 14 19215
rect 0 19213 17 19214
rect 25 19213 27 19222
rect 0 19206 38 19213
rect 0 19205 34 19206
rect 0 19189 8 19205
rect 14 19189 34 19205
rect 0 19188 34 19189
rect 0 19181 38 19188
rect 14 19180 17 19181
rect 25 19172 27 19181
rect 42 19152 45 19242
rect 71 19211 80 19239
rect 69 19173 80 19211
rect 107 19167 119 19201
rect 129 19173 143 19201
rect 129 19167 141 19173
rect 42 19101 46 19135
rect 72 19101 76 19135
rect 42 19054 76 19058
rect 42 19024 46 19054
rect 72 19024 76 19054
rect 16 19015 38 19021
rect 80 19015 102 19021
rect 144 19015 148 19763
rect 332 19695 336 19763
rect 380 19733 462 19765
rect 463 19733 472 19767
rect 480 19733 497 19767
rect 378 19725 464 19733
rect 505 19725 507 19775
rect 514 19733 548 19767
rect 565 19733 582 19767
rect 607 19725 609 19775
rect 404 19709 438 19711
rect 400 19695 442 19696
rect 378 19689 404 19695
rect 442 19689 464 19695
rect 400 19688 404 19689
rect 174 19649 246 19657
rect 295 19654 300 19688
rect 324 19654 329 19688
rect 224 19619 226 19635
rect 196 19611 226 19619
rect 332 19617 336 19685
rect 367 19654 438 19688
rect 400 19647 404 19654
rect 454 19641 504 19643
rect 494 19637 548 19641
rect 494 19632 514 19637
rect 504 19617 506 19632
rect 196 19607 230 19611
rect 196 19577 204 19607
rect 216 19577 230 19607
rect 400 19609 404 19617
rect 174 19543 181 19569
rect 224 19530 226 19577
rect 256 19569 328 19577
rect 332 19575 336 19605
rect 400 19575 408 19609
rect 434 19575 438 19609
rect 498 19607 506 19617
rect 514 19607 515 19627
rect 504 19591 506 19607
rect 525 19598 528 19632
rect 547 19607 548 19627
rect 557 19607 564 19617
rect 514 19591 530 19597
rect 532 19591 548 19597
rect 289 19540 305 19542
rect 196 19496 204 19530
rect 216 19496 230 19530
rect 244 19496 257 19530
rect 300 19526 308 19539
rect 332 19537 342 19575
rect 400 19567 404 19575
rect 336 19527 342 19537
rect 224 19449 226 19496
rect 278 19492 291 19526
rect 300 19510 321 19526
rect 332 19517 342 19527
rect 400 19527 409 19555
rect 562 19538 612 19540
rect 466 19529 497 19531
rect 565 19529 596 19531
rect 300 19508 312 19510
rect 300 19492 321 19508
rect 300 19486 308 19492
rect 289 19476 308 19486
rect 196 19419 204 19449
rect 216 19419 230 19449
rect 196 19415 230 19419
rect 196 19407 226 19415
rect 300 19407 308 19476
rect 332 19483 351 19517
rect 361 19483 375 19517
rect 400 19483 411 19527
rect 442 19522 500 19529
rect 466 19521 500 19522
rect 565 19521 599 19529
rect 497 19505 500 19521
rect 596 19505 599 19521
rect 466 19504 500 19505
rect 442 19497 500 19504
rect 565 19497 599 19505
rect 612 19488 614 19538
rect 332 19459 342 19483
rect 336 19447 342 19459
rect 224 19391 226 19407
rect 332 19379 342 19447
rect 400 19451 404 19459
rect 400 19417 408 19451
rect 434 19417 438 19451
rect 454 19435 504 19437
rect 504 19419 506 19435
rect 514 19429 530 19435
rect 532 19429 548 19435
rect 525 19419 548 19428
rect 400 19409 404 19417
rect 498 19409 506 19419
rect 504 19385 506 19409
rect 514 19399 515 19419
rect 525 19394 528 19419
rect 547 19399 548 19419
rect 557 19409 564 19419
rect 514 19385 548 19389
rect 151 19338 156 19372
rect 174 19369 246 19377
rect 256 19369 328 19377
rect 336 19371 342 19379
rect 400 19374 404 19379
rect 180 19341 185 19369
rect 174 19333 246 19341
rect 256 19333 328 19341
rect 332 19339 336 19369
rect 400 19340 438 19374
rect 224 19303 226 19319
rect 196 19295 226 19303
rect 196 19291 230 19295
rect 196 19261 204 19291
rect 216 19261 230 19291
rect 224 19214 226 19261
rect 300 19234 308 19303
rect 332 19301 342 19339
rect 400 19331 404 19340
rect 454 19325 504 19327
rect 494 19321 548 19325
rect 494 19316 514 19321
rect 504 19301 506 19316
rect 336 19289 342 19301
rect 289 19224 308 19234
rect 300 19218 308 19224
rect 332 19255 342 19289
rect 400 19293 404 19301
rect 400 19259 408 19293
rect 434 19259 438 19293
rect 498 19291 506 19301
rect 514 19291 515 19311
rect 504 19275 506 19291
rect 525 19282 528 19316
rect 547 19291 548 19311
rect 557 19291 564 19301
rect 514 19275 530 19281
rect 532 19275 548 19281
rect 332 19227 373 19255
rect 332 19221 351 19227
rect 196 19180 204 19214
rect 216 19180 230 19214
rect 244 19180 257 19214
rect 278 19184 291 19218
rect 300 19202 321 19218
rect 336 19211 351 19221
rect 300 19200 312 19202
rect 300 19184 321 19200
rect 332 19193 351 19211
rect 361 19193 375 19227
rect 400 19221 411 19259
rect 562 19222 612 19224
rect 400 19193 409 19221
rect 466 19213 497 19215
rect 565 19213 596 19215
rect 442 19206 500 19213
rect 466 19205 500 19206
rect 565 19205 599 19213
rect 174 19143 181 19167
rect 224 19133 226 19180
rect 300 19171 308 19184
rect 289 19168 305 19170
rect 332 19143 342 19193
rect 400 19173 404 19193
rect 497 19189 500 19205
rect 596 19189 599 19205
rect 466 19188 500 19189
rect 442 19181 500 19188
rect 565 19181 599 19189
rect 612 19172 614 19222
rect 256 19133 328 19141
rect 336 19135 342 19143
rect 400 19135 404 19143
rect 196 19103 204 19133
rect 216 19103 230 19133
rect 196 19099 230 19103
rect 196 19091 226 19099
rect 224 19075 226 19091
rect 332 19063 336 19131
rect 400 19101 408 19135
rect 434 19101 438 19135
rect 454 19119 504 19121
rect 504 19103 506 19119
rect 514 19113 530 19119
rect 532 19113 548 19119
rect 525 19103 548 19112
rect 400 19093 404 19101
rect 498 19093 506 19103
rect 504 19069 506 19093
rect 514 19083 515 19103
rect 525 19078 528 19103
rect 547 19083 548 19103
rect 557 19093 564 19103
rect 514 19069 548 19073
rect 400 19063 442 19064
rect 174 19053 246 19061
rect 400 19056 404 19063
rect 295 19022 300 19056
rect 324 19022 329 19056
rect 367 19022 438 19056
rect 400 19021 404 19022
rect 378 19015 404 19021
rect 442 19015 464 19021
rect 38 18999 80 19015
rect 400 18999 442 19015
rect -25 18985 25 18987
rect 455 18985 505 18987
rect 557 18985 607 18987
rect 16 18977 102 18985
rect 378 18977 464 18985
rect 8 18943 17 18977
rect 18 18975 51 18977
rect 80 18975 100 18977
rect 18 18943 100 18975
rect 380 18975 404 18977
rect 429 18975 438 18977
rect 442 18975 462 18977
rect 16 18935 102 18943
rect 42 18919 76 18921
rect 16 18899 38 18905
rect 42 18896 76 18900
rect 80 18899 102 18905
rect 42 18866 46 18896
rect 72 18866 76 18896
rect 42 18785 46 18819
rect 72 18785 76 18819
rect -25 18748 25 18750
rect 0 18740 14 18741
rect 0 18739 17 18740
rect 25 18739 27 18748
rect 0 18732 38 18739
rect 0 18731 34 18732
rect 0 18715 8 18731
rect 14 18715 34 18731
rect 0 18714 34 18715
rect 0 18707 38 18714
rect 14 18706 17 18707
rect 25 18698 27 18707
rect 42 18678 45 18768
rect 69 18753 80 18785
rect 107 18753 143 18781
rect 107 18747 119 18753
rect 109 18719 119 18747
rect 129 18719 143 18753
rect 42 18627 46 18661
rect 72 18627 76 18661
rect 38 18589 80 18590
rect 42 18548 76 18582
rect 79 18548 113 18582
rect 42 18469 46 18503
rect 72 18469 76 18503
rect -25 18432 25 18434
rect 0 18424 14 18425
rect 0 18423 17 18424
rect 25 18423 27 18432
rect 0 18416 38 18423
rect 0 18415 34 18416
rect 0 18399 8 18415
rect 14 18399 34 18415
rect 0 18398 34 18399
rect 0 18391 38 18398
rect 14 18390 17 18391
rect 25 18382 27 18391
rect 42 18362 45 18452
rect 71 18421 80 18449
rect 69 18383 80 18421
rect 107 18377 119 18411
rect 129 18383 143 18411
rect 129 18377 141 18383
rect 42 18311 46 18345
rect 72 18311 76 18345
rect 42 18264 76 18268
rect 42 18234 46 18264
rect 72 18234 76 18264
rect 16 18225 38 18231
rect 80 18225 102 18231
rect 144 18225 148 18973
rect 332 18905 336 18973
rect 380 18943 462 18975
rect 463 18943 472 18977
rect 480 18943 497 18977
rect 378 18935 464 18943
rect 505 18935 507 18985
rect 514 18943 548 18977
rect 565 18943 582 18977
rect 607 18935 609 18985
rect 404 18919 438 18921
rect 400 18905 442 18906
rect 378 18899 404 18905
rect 442 18899 464 18905
rect 400 18898 404 18899
rect 174 18859 246 18867
rect 295 18864 300 18898
rect 324 18864 329 18898
rect 224 18829 226 18845
rect 196 18821 226 18829
rect 332 18827 336 18895
rect 367 18864 438 18898
rect 400 18857 404 18864
rect 454 18851 504 18853
rect 494 18847 548 18851
rect 494 18842 514 18847
rect 504 18827 506 18842
rect 196 18817 230 18821
rect 196 18787 204 18817
rect 216 18787 230 18817
rect 400 18819 404 18827
rect 174 18753 181 18779
rect 224 18740 226 18787
rect 256 18779 328 18787
rect 332 18785 336 18815
rect 400 18785 408 18819
rect 434 18785 438 18819
rect 498 18817 506 18827
rect 514 18817 515 18837
rect 504 18801 506 18817
rect 525 18808 528 18842
rect 547 18817 548 18837
rect 557 18817 564 18827
rect 514 18801 530 18807
rect 532 18801 548 18807
rect 289 18750 305 18752
rect 196 18706 204 18740
rect 216 18706 230 18740
rect 244 18706 257 18740
rect 300 18736 308 18749
rect 332 18747 342 18785
rect 400 18777 404 18785
rect 336 18737 342 18747
rect 224 18659 226 18706
rect 278 18702 291 18736
rect 300 18720 321 18736
rect 332 18727 342 18737
rect 400 18737 409 18765
rect 562 18748 612 18750
rect 466 18739 497 18741
rect 565 18739 596 18741
rect 300 18718 312 18720
rect 300 18702 321 18718
rect 300 18696 308 18702
rect 289 18686 308 18696
rect 196 18629 204 18659
rect 216 18629 230 18659
rect 196 18625 230 18629
rect 196 18617 226 18625
rect 300 18617 308 18686
rect 332 18693 351 18727
rect 361 18693 375 18727
rect 400 18693 411 18737
rect 442 18732 500 18739
rect 466 18731 500 18732
rect 565 18731 599 18739
rect 497 18715 500 18731
rect 596 18715 599 18731
rect 466 18714 500 18715
rect 442 18707 500 18714
rect 565 18707 599 18715
rect 612 18698 614 18748
rect 332 18669 342 18693
rect 336 18657 342 18669
rect 224 18601 226 18617
rect 332 18589 342 18657
rect 400 18661 404 18669
rect 400 18627 408 18661
rect 434 18627 438 18661
rect 454 18645 504 18647
rect 504 18629 506 18645
rect 514 18639 530 18645
rect 532 18639 548 18645
rect 525 18629 548 18638
rect 400 18619 404 18627
rect 498 18619 506 18629
rect 504 18595 506 18619
rect 514 18609 515 18629
rect 525 18604 528 18629
rect 547 18609 548 18629
rect 557 18619 564 18629
rect 514 18595 548 18599
rect 151 18548 156 18582
rect 174 18579 246 18587
rect 256 18579 328 18587
rect 336 18581 342 18589
rect 400 18584 404 18589
rect 180 18551 185 18579
rect 174 18543 246 18551
rect 256 18543 328 18551
rect 332 18549 336 18579
rect 400 18550 438 18584
rect 224 18513 226 18529
rect 196 18505 226 18513
rect 196 18501 230 18505
rect 196 18471 204 18501
rect 216 18471 230 18501
rect 224 18424 226 18471
rect 300 18444 308 18513
rect 332 18511 342 18549
rect 400 18541 404 18550
rect 454 18535 504 18537
rect 494 18531 548 18535
rect 494 18526 514 18531
rect 504 18511 506 18526
rect 336 18499 342 18511
rect 289 18434 308 18444
rect 300 18428 308 18434
rect 332 18465 342 18499
rect 400 18503 404 18511
rect 400 18469 408 18503
rect 434 18469 438 18503
rect 498 18501 506 18511
rect 514 18501 515 18521
rect 504 18485 506 18501
rect 525 18492 528 18526
rect 547 18501 548 18521
rect 557 18501 564 18511
rect 514 18485 530 18491
rect 532 18485 548 18491
rect 332 18437 373 18465
rect 332 18431 351 18437
rect 196 18390 204 18424
rect 216 18390 230 18424
rect 244 18390 257 18424
rect 278 18394 291 18428
rect 300 18412 321 18428
rect 336 18421 351 18431
rect 300 18410 312 18412
rect 300 18394 321 18410
rect 332 18403 351 18421
rect 361 18403 375 18437
rect 400 18431 411 18469
rect 562 18432 612 18434
rect 400 18403 409 18431
rect 466 18423 497 18425
rect 565 18423 596 18425
rect 442 18416 500 18423
rect 466 18415 500 18416
rect 565 18415 599 18423
rect 174 18353 181 18377
rect 224 18343 226 18390
rect 300 18381 308 18394
rect 289 18378 305 18380
rect 332 18353 342 18403
rect 400 18383 404 18403
rect 497 18399 500 18415
rect 596 18399 599 18415
rect 466 18398 500 18399
rect 442 18391 500 18398
rect 565 18391 599 18399
rect 612 18382 614 18432
rect 256 18343 328 18351
rect 336 18345 342 18353
rect 400 18345 404 18353
rect 196 18313 204 18343
rect 216 18313 230 18343
rect 196 18309 230 18313
rect 196 18301 226 18309
rect 224 18285 226 18301
rect 332 18273 336 18341
rect 400 18311 408 18345
rect 434 18311 438 18345
rect 454 18329 504 18331
rect 504 18313 506 18329
rect 514 18323 530 18329
rect 532 18323 548 18329
rect 525 18313 548 18322
rect 400 18303 404 18311
rect 498 18303 506 18313
rect 504 18279 506 18303
rect 514 18293 515 18313
rect 525 18288 528 18313
rect 547 18293 548 18313
rect 557 18303 564 18313
rect 514 18279 548 18283
rect 400 18273 442 18274
rect 174 18263 246 18271
rect 400 18266 404 18273
rect 295 18232 300 18266
rect 324 18232 329 18266
rect 367 18232 438 18266
rect 400 18231 404 18232
rect 378 18225 404 18231
rect 442 18225 464 18231
rect 38 18209 80 18225
rect 400 18209 442 18225
rect -25 18195 25 18197
rect 455 18195 505 18197
rect 557 18195 607 18197
rect 16 18187 102 18195
rect 378 18187 464 18195
rect 8 18153 17 18187
rect 18 18185 51 18187
rect 80 18185 100 18187
rect 18 18153 100 18185
rect 380 18185 404 18187
rect 429 18185 438 18187
rect 442 18185 462 18187
rect 16 18145 102 18153
rect 42 18129 76 18131
rect 16 18109 38 18115
rect 42 18106 76 18110
rect 80 18109 102 18115
rect 42 18076 46 18106
rect 72 18076 76 18106
rect 42 17995 46 18029
rect 72 17995 76 18029
rect -25 17958 25 17960
rect 0 17950 14 17951
rect 0 17949 17 17950
rect 25 17949 27 17958
rect 0 17942 38 17949
rect 0 17941 34 17942
rect 0 17925 8 17941
rect 14 17925 34 17941
rect 0 17924 34 17925
rect 0 17917 38 17924
rect 14 17916 17 17917
rect 25 17908 27 17917
rect 42 17888 45 17978
rect 69 17963 80 17995
rect 107 17963 143 17991
rect 107 17957 119 17963
rect 109 17929 119 17957
rect 129 17929 143 17963
rect 42 17837 46 17871
rect 72 17837 76 17871
rect 38 17799 80 17800
rect 42 17758 76 17792
rect 79 17758 113 17792
rect 42 17679 46 17713
rect 72 17679 76 17713
rect -25 17642 25 17644
rect 0 17634 14 17635
rect 0 17633 17 17634
rect 25 17633 27 17642
rect 0 17626 38 17633
rect 0 17625 34 17626
rect 0 17609 8 17625
rect 14 17609 34 17625
rect 0 17608 34 17609
rect 0 17601 38 17608
rect 14 17600 17 17601
rect 25 17592 27 17601
rect 42 17572 45 17662
rect 71 17631 80 17659
rect 69 17593 80 17631
rect 107 17587 119 17621
rect 129 17593 143 17621
rect 129 17587 141 17593
rect 42 17521 46 17555
rect 72 17521 76 17555
rect 42 17474 76 17478
rect 42 17444 46 17474
rect 72 17444 76 17474
rect 16 17435 38 17441
rect 80 17435 102 17441
rect 144 17435 148 18183
rect 332 18115 336 18183
rect 380 18153 462 18185
rect 463 18153 472 18187
rect 480 18153 497 18187
rect 378 18145 464 18153
rect 505 18145 507 18195
rect 514 18153 548 18187
rect 565 18153 582 18187
rect 607 18145 609 18195
rect 404 18129 438 18131
rect 400 18115 442 18116
rect 378 18109 404 18115
rect 442 18109 464 18115
rect 400 18108 404 18109
rect 174 18069 246 18077
rect 295 18074 300 18108
rect 324 18074 329 18108
rect 224 18039 226 18055
rect 196 18031 226 18039
rect 332 18037 336 18105
rect 367 18074 438 18108
rect 400 18067 404 18074
rect 454 18061 504 18063
rect 494 18057 548 18061
rect 494 18052 514 18057
rect 504 18037 506 18052
rect 196 18027 230 18031
rect 196 17997 204 18027
rect 216 17997 230 18027
rect 400 18029 404 18037
rect 174 17963 181 17989
rect 224 17950 226 17997
rect 256 17989 328 17997
rect 332 17995 336 18025
rect 400 17995 408 18029
rect 434 17995 438 18029
rect 498 18027 506 18037
rect 514 18027 515 18047
rect 504 18011 506 18027
rect 525 18018 528 18052
rect 547 18027 548 18047
rect 557 18027 564 18037
rect 514 18011 530 18017
rect 532 18011 548 18017
rect 289 17960 305 17962
rect 196 17916 204 17950
rect 216 17916 230 17950
rect 244 17916 257 17950
rect 300 17946 308 17959
rect 332 17957 342 17995
rect 400 17987 404 17995
rect 336 17947 342 17957
rect 224 17869 226 17916
rect 278 17912 291 17946
rect 300 17930 321 17946
rect 332 17937 342 17947
rect 400 17947 409 17975
rect 562 17958 612 17960
rect 466 17949 497 17951
rect 565 17949 596 17951
rect 300 17928 312 17930
rect 300 17912 321 17928
rect 300 17906 308 17912
rect 289 17896 308 17906
rect 196 17839 204 17869
rect 216 17839 230 17869
rect 196 17835 230 17839
rect 196 17827 226 17835
rect 300 17827 308 17896
rect 332 17903 351 17937
rect 361 17903 375 17937
rect 400 17903 411 17947
rect 442 17942 500 17949
rect 466 17941 500 17942
rect 565 17941 599 17949
rect 497 17925 500 17941
rect 596 17925 599 17941
rect 466 17924 500 17925
rect 442 17917 500 17924
rect 565 17917 599 17925
rect 612 17908 614 17958
rect 332 17879 342 17903
rect 336 17867 342 17879
rect 224 17811 226 17827
rect 332 17799 342 17867
rect 400 17871 404 17879
rect 400 17837 408 17871
rect 434 17837 438 17871
rect 454 17855 504 17857
rect 504 17839 506 17855
rect 514 17849 530 17855
rect 532 17849 548 17855
rect 525 17839 548 17848
rect 400 17829 404 17837
rect 498 17829 506 17839
rect 504 17805 506 17829
rect 514 17819 515 17839
rect 525 17814 528 17839
rect 547 17819 548 17839
rect 557 17829 564 17839
rect 514 17805 548 17809
rect 151 17758 156 17792
rect 174 17789 246 17797
rect 256 17789 328 17797
rect 336 17791 342 17799
rect 400 17794 404 17799
rect 180 17761 185 17789
rect 174 17753 246 17761
rect 256 17753 328 17761
rect 332 17759 336 17789
rect 400 17760 438 17794
rect 224 17723 226 17739
rect 196 17715 226 17723
rect 196 17711 230 17715
rect 196 17681 204 17711
rect 216 17681 230 17711
rect 224 17634 226 17681
rect 300 17654 308 17723
rect 332 17721 342 17759
rect 400 17751 404 17760
rect 454 17745 504 17747
rect 494 17741 548 17745
rect 494 17736 514 17741
rect 504 17721 506 17736
rect 336 17709 342 17721
rect 289 17644 308 17654
rect 300 17638 308 17644
rect 332 17675 342 17709
rect 400 17713 404 17721
rect 400 17679 408 17713
rect 434 17679 438 17713
rect 498 17711 506 17721
rect 514 17711 515 17731
rect 504 17695 506 17711
rect 525 17702 528 17736
rect 547 17711 548 17731
rect 557 17711 564 17721
rect 514 17695 530 17701
rect 532 17695 548 17701
rect 332 17647 373 17675
rect 332 17641 351 17647
rect 196 17600 204 17634
rect 216 17600 230 17634
rect 244 17600 257 17634
rect 278 17604 291 17638
rect 300 17622 321 17638
rect 336 17631 351 17641
rect 300 17620 312 17622
rect 300 17604 321 17620
rect 332 17613 351 17631
rect 361 17613 375 17647
rect 400 17641 411 17679
rect 562 17642 612 17644
rect 400 17613 409 17641
rect 466 17633 497 17635
rect 565 17633 596 17635
rect 442 17626 500 17633
rect 466 17625 500 17626
rect 565 17625 599 17633
rect 174 17563 181 17587
rect 224 17553 226 17600
rect 300 17591 308 17604
rect 289 17588 305 17590
rect 332 17563 342 17613
rect 400 17593 404 17613
rect 497 17609 500 17625
rect 596 17609 599 17625
rect 466 17608 500 17609
rect 442 17601 500 17608
rect 565 17601 599 17609
rect 612 17592 614 17642
rect 256 17553 328 17561
rect 336 17555 342 17563
rect 400 17555 404 17563
rect 196 17523 204 17553
rect 216 17523 230 17553
rect 196 17519 230 17523
rect 196 17511 226 17519
rect 224 17495 226 17511
rect 332 17483 336 17551
rect 400 17521 408 17555
rect 434 17521 438 17555
rect 454 17539 504 17541
rect 504 17523 506 17539
rect 514 17533 530 17539
rect 532 17533 548 17539
rect 525 17523 548 17532
rect 400 17513 404 17521
rect 498 17513 506 17523
rect 504 17489 506 17513
rect 514 17503 515 17523
rect 525 17498 528 17523
rect 547 17503 548 17523
rect 557 17513 564 17523
rect 514 17489 548 17493
rect 400 17483 442 17484
rect 174 17473 246 17481
rect 400 17476 404 17483
rect 295 17442 300 17476
rect 324 17442 329 17476
rect 367 17442 438 17476
rect 400 17441 404 17442
rect 378 17435 404 17441
rect 442 17435 464 17441
rect 38 17419 80 17435
rect 400 17419 442 17435
rect -25 17405 25 17407
rect 455 17405 505 17407
rect 557 17405 607 17407
rect 16 17397 102 17405
rect 378 17397 464 17405
rect 8 17363 17 17397
rect 18 17395 51 17397
rect 80 17395 100 17397
rect 18 17363 100 17395
rect 380 17395 404 17397
rect 429 17395 438 17397
rect 442 17395 462 17397
rect 16 17355 102 17363
rect 42 17339 76 17341
rect 16 17319 38 17325
rect 42 17316 76 17320
rect 80 17319 102 17325
rect 42 17286 46 17316
rect 72 17286 76 17316
rect 42 17205 46 17239
rect 72 17205 76 17239
rect -25 17168 25 17170
rect 0 17160 14 17161
rect 0 17159 17 17160
rect 25 17159 27 17168
rect 0 17152 38 17159
rect 0 17151 34 17152
rect 0 17135 8 17151
rect 14 17135 34 17151
rect 0 17134 34 17135
rect 0 17127 38 17134
rect 14 17126 17 17127
rect 25 17118 27 17127
rect 42 17098 45 17188
rect 69 17173 80 17205
rect 107 17173 143 17201
rect 107 17167 119 17173
rect 109 17139 119 17167
rect 129 17139 143 17173
rect 42 17047 46 17081
rect 72 17047 76 17081
rect 38 17009 80 17010
rect 42 16968 76 17002
rect 79 16968 113 17002
rect 42 16889 46 16923
rect 72 16889 76 16923
rect -25 16852 25 16854
rect 0 16844 14 16845
rect 0 16843 17 16844
rect 25 16843 27 16852
rect 0 16836 38 16843
rect 0 16835 34 16836
rect 0 16819 8 16835
rect 14 16819 34 16835
rect 0 16818 34 16819
rect 0 16811 38 16818
rect 14 16810 17 16811
rect 25 16802 27 16811
rect 42 16782 45 16872
rect 71 16841 80 16869
rect 69 16803 80 16841
rect 107 16797 119 16831
rect 129 16803 143 16831
rect 129 16797 141 16803
rect 42 16731 46 16765
rect 72 16731 76 16765
rect 42 16684 76 16688
rect 42 16654 46 16684
rect 72 16654 76 16684
rect 16 16645 38 16651
rect 80 16645 102 16651
rect 144 16645 148 17393
rect 332 17325 336 17393
rect 380 17363 462 17395
rect 463 17363 472 17397
rect 480 17363 497 17397
rect 378 17355 464 17363
rect 505 17355 507 17405
rect 514 17363 548 17397
rect 565 17363 582 17397
rect 607 17355 609 17405
rect 404 17339 438 17341
rect 400 17325 442 17326
rect 378 17319 404 17325
rect 442 17319 464 17325
rect 400 17318 404 17319
rect 174 17279 246 17287
rect 295 17284 300 17318
rect 324 17284 329 17318
rect 224 17249 226 17265
rect 196 17241 226 17249
rect 332 17247 336 17315
rect 367 17284 438 17318
rect 400 17277 404 17284
rect 454 17271 504 17273
rect 494 17267 548 17271
rect 494 17262 514 17267
rect 504 17247 506 17262
rect 196 17237 230 17241
rect 196 17207 204 17237
rect 216 17207 230 17237
rect 400 17239 404 17247
rect 174 17173 181 17199
rect 224 17160 226 17207
rect 256 17199 328 17207
rect 332 17205 336 17235
rect 400 17205 408 17239
rect 434 17205 438 17239
rect 498 17237 506 17247
rect 514 17237 515 17257
rect 504 17221 506 17237
rect 525 17228 528 17262
rect 547 17237 548 17257
rect 557 17237 564 17247
rect 514 17221 530 17227
rect 532 17221 548 17227
rect 289 17170 305 17172
rect 196 17126 204 17160
rect 216 17126 230 17160
rect 244 17126 257 17160
rect 300 17156 308 17169
rect 332 17167 342 17205
rect 400 17197 404 17205
rect 336 17157 342 17167
rect 224 17079 226 17126
rect 278 17122 291 17156
rect 300 17140 321 17156
rect 332 17147 342 17157
rect 400 17157 409 17185
rect 562 17168 612 17170
rect 466 17159 497 17161
rect 565 17159 596 17161
rect 300 17138 312 17140
rect 300 17122 321 17138
rect 300 17116 308 17122
rect 289 17106 308 17116
rect 196 17049 204 17079
rect 216 17049 230 17079
rect 196 17045 230 17049
rect 196 17037 226 17045
rect 300 17037 308 17106
rect 332 17113 351 17147
rect 361 17113 375 17147
rect 400 17113 411 17157
rect 442 17152 500 17159
rect 466 17151 500 17152
rect 565 17151 599 17159
rect 497 17135 500 17151
rect 596 17135 599 17151
rect 466 17134 500 17135
rect 442 17127 500 17134
rect 565 17127 599 17135
rect 612 17118 614 17168
rect 332 17089 342 17113
rect 336 17077 342 17089
rect 224 17021 226 17037
rect 332 17009 342 17077
rect 400 17081 404 17089
rect 400 17047 408 17081
rect 434 17047 438 17081
rect 454 17065 504 17067
rect 504 17049 506 17065
rect 514 17059 530 17065
rect 532 17059 548 17065
rect 525 17049 548 17058
rect 400 17039 404 17047
rect 498 17039 506 17049
rect 504 17015 506 17039
rect 514 17029 515 17049
rect 525 17024 528 17049
rect 547 17029 548 17049
rect 557 17039 564 17049
rect 514 17015 548 17019
rect 151 16968 156 17002
rect 174 16999 246 17007
rect 256 16999 328 17007
rect 336 17001 342 17009
rect 400 17004 404 17009
rect 180 16971 185 16999
rect 174 16963 246 16971
rect 256 16963 328 16971
rect 332 16969 336 16999
rect 400 16970 438 17004
rect 224 16933 226 16949
rect 196 16925 226 16933
rect 196 16921 230 16925
rect 196 16891 204 16921
rect 216 16891 230 16921
rect 224 16844 226 16891
rect 300 16864 308 16933
rect 332 16931 342 16969
rect 400 16961 404 16970
rect 454 16955 504 16957
rect 494 16951 548 16955
rect 494 16946 514 16951
rect 504 16931 506 16946
rect 336 16919 342 16931
rect 289 16854 308 16864
rect 300 16848 308 16854
rect 332 16885 342 16919
rect 400 16923 404 16931
rect 400 16889 408 16923
rect 434 16889 438 16923
rect 498 16921 506 16931
rect 514 16921 515 16941
rect 504 16905 506 16921
rect 525 16912 528 16946
rect 547 16921 548 16941
rect 557 16921 564 16931
rect 514 16905 530 16911
rect 532 16905 548 16911
rect 332 16857 373 16885
rect 332 16851 351 16857
rect 196 16810 204 16844
rect 216 16810 230 16844
rect 244 16810 257 16844
rect 278 16814 291 16848
rect 300 16832 321 16848
rect 336 16841 351 16851
rect 300 16830 312 16832
rect 300 16814 321 16830
rect 332 16823 351 16841
rect 361 16823 375 16857
rect 400 16851 411 16889
rect 562 16852 612 16854
rect 400 16823 409 16851
rect 466 16843 497 16845
rect 565 16843 596 16845
rect 442 16836 500 16843
rect 466 16835 500 16836
rect 565 16835 599 16843
rect 174 16773 181 16797
rect 224 16763 226 16810
rect 300 16801 308 16814
rect 289 16798 305 16800
rect 332 16773 342 16823
rect 400 16803 404 16823
rect 497 16819 500 16835
rect 596 16819 599 16835
rect 466 16818 500 16819
rect 442 16811 500 16818
rect 565 16811 599 16819
rect 612 16802 614 16852
rect 256 16763 328 16771
rect 336 16765 342 16773
rect 400 16765 404 16773
rect 196 16733 204 16763
rect 216 16733 230 16763
rect 196 16729 230 16733
rect 196 16721 226 16729
rect 224 16705 226 16721
rect 332 16693 336 16761
rect 400 16731 408 16765
rect 434 16731 438 16765
rect 454 16749 504 16751
rect 504 16733 506 16749
rect 514 16743 530 16749
rect 532 16743 548 16749
rect 525 16733 548 16742
rect 400 16723 404 16731
rect 498 16723 506 16733
rect 504 16699 506 16723
rect 514 16713 515 16733
rect 525 16708 528 16733
rect 547 16713 548 16733
rect 557 16723 564 16733
rect 514 16699 548 16703
rect 400 16693 442 16694
rect 174 16683 246 16691
rect 400 16686 404 16693
rect 295 16652 300 16686
rect 324 16652 329 16686
rect 367 16652 438 16686
rect 400 16651 404 16652
rect 378 16645 404 16651
rect 442 16645 464 16651
rect 38 16629 80 16645
rect 400 16629 442 16645
rect -25 16615 25 16617
rect 455 16615 505 16617
rect 557 16615 607 16617
rect 16 16607 102 16615
rect 378 16607 464 16615
rect 8 16573 17 16607
rect 18 16605 51 16607
rect 80 16605 100 16607
rect 18 16573 100 16605
rect 380 16605 404 16607
rect 429 16605 438 16607
rect 442 16605 462 16607
rect 16 16565 102 16573
rect 42 16549 76 16551
rect 16 16529 38 16535
rect 42 16526 76 16530
rect 80 16529 102 16535
rect 42 16496 46 16526
rect 72 16496 76 16526
rect 42 16415 46 16449
rect 72 16415 76 16449
rect -25 16378 25 16380
rect 0 16370 14 16371
rect 0 16369 17 16370
rect 25 16369 27 16378
rect 0 16362 38 16369
rect 0 16361 34 16362
rect 0 16345 8 16361
rect 14 16345 34 16361
rect 0 16344 34 16345
rect 0 16337 38 16344
rect 14 16336 17 16337
rect 25 16328 27 16337
rect 42 16308 45 16398
rect 69 16383 80 16415
rect 107 16383 143 16411
rect 107 16377 119 16383
rect 109 16349 119 16377
rect 129 16349 143 16383
rect 42 16257 46 16291
rect 72 16257 76 16291
rect 38 16219 80 16220
rect 42 16178 76 16212
rect 79 16178 113 16212
rect 42 16099 46 16133
rect 72 16099 76 16133
rect -25 16062 25 16064
rect 0 16054 14 16055
rect 0 16053 17 16054
rect 25 16053 27 16062
rect 0 16046 38 16053
rect 0 16045 34 16046
rect 0 16029 8 16045
rect 14 16029 34 16045
rect 0 16028 34 16029
rect 0 16021 38 16028
rect 14 16020 17 16021
rect 25 16012 27 16021
rect 42 15992 45 16082
rect 71 16051 80 16079
rect 69 16013 80 16051
rect 107 16007 119 16041
rect 129 16013 143 16041
rect 129 16007 141 16013
rect 42 15941 46 15975
rect 72 15941 76 15975
rect 42 15894 76 15898
rect 42 15864 46 15894
rect 72 15864 76 15894
rect 16 15855 38 15861
rect 80 15855 102 15861
rect 144 15855 148 16603
rect 332 16535 336 16603
rect 380 16573 462 16605
rect 463 16573 472 16607
rect 480 16573 497 16607
rect 378 16565 464 16573
rect 505 16565 507 16615
rect 514 16573 548 16607
rect 565 16573 582 16607
rect 607 16565 609 16615
rect 404 16549 438 16551
rect 400 16535 442 16536
rect 378 16529 404 16535
rect 442 16529 464 16535
rect 400 16528 404 16529
rect 174 16489 246 16497
rect 295 16494 300 16528
rect 324 16494 329 16528
rect 224 16459 226 16475
rect 196 16451 226 16459
rect 332 16457 336 16525
rect 367 16494 438 16528
rect 400 16487 404 16494
rect 454 16481 504 16483
rect 494 16477 548 16481
rect 494 16472 514 16477
rect 504 16457 506 16472
rect 196 16447 230 16451
rect 196 16417 204 16447
rect 216 16417 230 16447
rect 400 16449 404 16457
rect 174 16383 181 16409
rect 224 16370 226 16417
rect 256 16409 328 16417
rect 332 16415 336 16445
rect 400 16415 408 16449
rect 434 16415 438 16449
rect 498 16447 506 16457
rect 514 16447 515 16467
rect 504 16431 506 16447
rect 525 16438 528 16472
rect 547 16447 548 16467
rect 557 16447 564 16457
rect 514 16431 530 16437
rect 532 16431 548 16437
rect 289 16380 305 16382
rect 196 16336 204 16370
rect 216 16336 230 16370
rect 244 16336 257 16370
rect 300 16366 308 16379
rect 332 16377 342 16415
rect 400 16407 404 16415
rect 336 16367 342 16377
rect 224 16289 226 16336
rect 278 16332 291 16366
rect 300 16350 321 16366
rect 332 16357 342 16367
rect 400 16367 409 16395
rect 562 16378 612 16380
rect 466 16369 497 16371
rect 565 16369 596 16371
rect 300 16348 312 16350
rect 300 16332 321 16348
rect 300 16326 308 16332
rect 289 16316 308 16326
rect 196 16259 204 16289
rect 216 16259 230 16289
rect 196 16255 230 16259
rect 196 16247 226 16255
rect 300 16247 308 16316
rect 332 16323 351 16357
rect 361 16323 375 16357
rect 400 16323 411 16367
rect 442 16362 500 16369
rect 466 16361 500 16362
rect 565 16361 599 16369
rect 497 16345 500 16361
rect 596 16345 599 16361
rect 466 16344 500 16345
rect 442 16337 500 16344
rect 565 16337 599 16345
rect 612 16328 614 16378
rect 332 16299 342 16323
rect 336 16287 342 16299
rect 224 16231 226 16247
rect 332 16219 342 16287
rect 400 16291 404 16299
rect 400 16257 408 16291
rect 434 16257 438 16291
rect 454 16275 504 16277
rect 504 16259 506 16275
rect 514 16269 530 16275
rect 532 16269 548 16275
rect 525 16259 548 16268
rect 400 16249 404 16257
rect 498 16249 506 16259
rect 504 16225 506 16249
rect 514 16239 515 16259
rect 525 16234 528 16259
rect 547 16239 548 16259
rect 557 16249 564 16259
rect 514 16225 548 16229
rect 151 16178 156 16212
rect 174 16209 246 16217
rect 256 16209 328 16217
rect 336 16211 342 16219
rect 400 16214 404 16219
rect 180 16181 185 16209
rect 174 16173 246 16181
rect 256 16173 328 16181
rect 332 16179 336 16209
rect 400 16180 438 16214
rect 224 16143 226 16159
rect 196 16135 226 16143
rect 196 16131 230 16135
rect 196 16101 204 16131
rect 216 16101 230 16131
rect 224 16054 226 16101
rect 300 16074 308 16143
rect 332 16141 342 16179
rect 400 16171 404 16180
rect 454 16165 504 16167
rect 494 16161 548 16165
rect 494 16156 514 16161
rect 504 16141 506 16156
rect 336 16129 342 16141
rect 289 16064 308 16074
rect 300 16058 308 16064
rect 332 16095 342 16129
rect 400 16133 404 16141
rect 400 16099 408 16133
rect 434 16099 438 16133
rect 498 16131 506 16141
rect 514 16131 515 16151
rect 504 16115 506 16131
rect 525 16122 528 16156
rect 547 16131 548 16151
rect 557 16131 564 16141
rect 514 16115 530 16121
rect 532 16115 548 16121
rect 332 16067 373 16095
rect 332 16061 351 16067
rect 196 16020 204 16054
rect 216 16020 230 16054
rect 244 16020 257 16054
rect 278 16024 291 16058
rect 300 16042 321 16058
rect 336 16051 351 16061
rect 300 16040 312 16042
rect 300 16024 321 16040
rect 332 16033 351 16051
rect 361 16033 375 16067
rect 400 16061 411 16099
rect 562 16062 612 16064
rect 400 16033 409 16061
rect 466 16053 497 16055
rect 565 16053 596 16055
rect 442 16046 500 16053
rect 466 16045 500 16046
rect 565 16045 599 16053
rect 174 15983 181 16007
rect 224 15973 226 16020
rect 300 16011 308 16024
rect 289 16008 305 16010
rect 332 15983 342 16033
rect 400 16013 404 16033
rect 497 16029 500 16045
rect 596 16029 599 16045
rect 466 16028 500 16029
rect 442 16021 500 16028
rect 565 16021 599 16029
rect 612 16012 614 16062
rect 256 15973 328 15981
rect 336 15975 342 15983
rect 400 15975 404 15983
rect 196 15943 204 15973
rect 216 15943 230 15973
rect 196 15939 230 15943
rect 196 15931 226 15939
rect 224 15915 226 15931
rect 332 15903 336 15971
rect 400 15941 408 15975
rect 434 15941 438 15975
rect 454 15959 504 15961
rect 504 15943 506 15959
rect 514 15953 530 15959
rect 532 15953 548 15959
rect 525 15943 548 15952
rect 400 15933 404 15941
rect 498 15933 506 15943
rect 504 15909 506 15933
rect 514 15923 515 15943
rect 525 15918 528 15943
rect 547 15923 548 15943
rect 557 15933 564 15943
rect 514 15909 548 15913
rect 400 15903 442 15904
rect 174 15893 246 15901
rect 400 15896 404 15903
rect 295 15862 300 15896
rect 324 15862 329 15896
rect 367 15862 438 15896
rect 400 15861 404 15862
rect 378 15855 404 15861
rect 442 15855 464 15861
rect 38 15839 80 15855
rect 400 15839 442 15855
rect -25 15825 25 15827
rect 455 15825 505 15827
rect 557 15825 607 15827
rect 16 15817 102 15825
rect 378 15817 464 15825
rect 8 15783 17 15817
rect 18 15815 51 15817
rect 80 15815 100 15817
rect 18 15783 100 15815
rect 380 15815 404 15817
rect 429 15815 438 15817
rect 442 15815 462 15817
rect 16 15775 102 15783
rect 42 15759 76 15761
rect 16 15739 38 15745
rect 42 15736 76 15740
rect 80 15739 102 15745
rect 42 15706 46 15736
rect 72 15706 76 15736
rect 42 15625 46 15659
rect 72 15625 76 15659
rect -25 15588 25 15590
rect 0 15580 14 15581
rect 0 15579 17 15580
rect 25 15579 27 15588
rect 0 15572 38 15579
rect 0 15571 34 15572
rect 0 15555 8 15571
rect 14 15555 34 15571
rect 0 15554 34 15555
rect 0 15547 38 15554
rect 14 15546 17 15547
rect 25 15538 27 15547
rect 42 15518 45 15608
rect 69 15593 80 15625
rect 107 15593 143 15621
rect 107 15587 119 15593
rect 109 15559 119 15587
rect 129 15559 143 15593
rect 42 15467 46 15501
rect 72 15467 76 15501
rect 38 15429 80 15430
rect 42 15388 76 15422
rect 79 15388 113 15422
rect 42 15309 46 15343
rect 72 15309 76 15343
rect -25 15272 25 15274
rect 0 15264 14 15265
rect 0 15263 17 15264
rect 25 15263 27 15272
rect 0 15256 38 15263
rect 0 15255 34 15256
rect 0 15239 8 15255
rect 14 15239 34 15255
rect 0 15238 34 15239
rect 0 15231 38 15238
rect 14 15230 17 15231
rect 25 15222 27 15231
rect 42 15202 45 15292
rect 71 15261 80 15289
rect 69 15223 80 15261
rect 107 15217 119 15251
rect 129 15223 143 15251
rect 129 15217 141 15223
rect 42 15151 46 15185
rect 72 15151 76 15185
rect 42 15104 76 15108
rect 42 15074 46 15104
rect 72 15074 76 15104
rect 16 15065 38 15071
rect 80 15065 102 15071
rect 144 15065 148 15813
rect 332 15745 336 15813
rect 380 15783 462 15815
rect 463 15783 472 15817
rect 480 15783 497 15817
rect 378 15775 464 15783
rect 505 15775 507 15825
rect 514 15783 548 15817
rect 565 15783 582 15817
rect 607 15775 609 15825
rect 404 15759 438 15761
rect 400 15745 442 15746
rect 378 15739 404 15745
rect 442 15739 464 15745
rect 400 15738 404 15739
rect 174 15699 246 15707
rect 295 15704 300 15738
rect 324 15704 329 15738
rect 224 15669 226 15685
rect 196 15661 226 15669
rect 332 15667 336 15735
rect 367 15704 438 15738
rect 400 15697 404 15704
rect 454 15691 504 15693
rect 494 15687 548 15691
rect 494 15682 514 15687
rect 504 15667 506 15682
rect 196 15657 230 15661
rect 196 15627 204 15657
rect 216 15627 230 15657
rect 400 15659 404 15667
rect 174 15593 181 15619
rect 224 15580 226 15627
rect 256 15619 328 15627
rect 332 15625 336 15655
rect 400 15625 408 15659
rect 434 15625 438 15659
rect 498 15657 506 15667
rect 514 15657 515 15677
rect 504 15641 506 15657
rect 525 15648 528 15682
rect 547 15657 548 15677
rect 557 15657 564 15667
rect 514 15641 530 15647
rect 532 15641 548 15647
rect 289 15590 305 15592
rect 196 15546 204 15580
rect 216 15546 230 15580
rect 244 15546 257 15580
rect 300 15576 308 15589
rect 332 15587 342 15625
rect 400 15617 404 15625
rect 336 15577 342 15587
rect 224 15499 226 15546
rect 278 15542 291 15576
rect 300 15560 321 15576
rect 332 15567 342 15577
rect 400 15577 409 15605
rect 562 15588 612 15590
rect 466 15579 497 15581
rect 565 15579 596 15581
rect 300 15558 312 15560
rect 300 15542 321 15558
rect 300 15536 308 15542
rect 289 15526 308 15536
rect 196 15469 204 15499
rect 216 15469 230 15499
rect 196 15465 230 15469
rect 196 15457 226 15465
rect 300 15457 308 15526
rect 332 15533 351 15567
rect 361 15533 375 15567
rect 400 15533 411 15577
rect 442 15572 500 15579
rect 466 15571 500 15572
rect 565 15571 599 15579
rect 497 15555 500 15571
rect 596 15555 599 15571
rect 466 15554 500 15555
rect 442 15547 500 15554
rect 565 15547 599 15555
rect 612 15538 614 15588
rect 332 15509 342 15533
rect 336 15497 342 15509
rect 224 15441 226 15457
rect 332 15429 342 15497
rect 400 15501 404 15509
rect 400 15467 408 15501
rect 434 15467 438 15501
rect 454 15485 504 15487
rect 504 15469 506 15485
rect 514 15479 530 15485
rect 532 15479 548 15485
rect 525 15469 548 15478
rect 400 15459 404 15467
rect 498 15459 506 15469
rect 504 15435 506 15459
rect 514 15449 515 15469
rect 525 15444 528 15469
rect 547 15449 548 15469
rect 557 15459 564 15469
rect 514 15435 548 15439
rect 151 15388 156 15422
rect 174 15419 246 15427
rect 256 15419 328 15427
rect 336 15421 342 15429
rect 400 15424 404 15429
rect 180 15391 185 15419
rect 174 15383 246 15391
rect 256 15383 328 15391
rect 332 15389 336 15419
rect 400 15390 438 15424
rect 224 15353 226 15369
rect 196 15345 226 15353
rect 196 15341 230 15345
rect 196 15311 204 15341
rect 216 15311 230 15341
rect 224 15264 226 15311
rect 300 15284 308 15353
rect 332 15351 342 15389
rect 400 15381 404 15390
rect 454 15375 504 15377
rect 494 15371 548 15375
rect 494 15366 514 15371
rect 504 15351 506 15366
rect 336 15339 342 15351
rect 289 15274 308 15284
rect 300 15268 308 15274
rect 332 15305 342 15339
rect 400 15343 404 15351
rect 400 15309 408 15343
rect 434 15309 438 15343
rect 498 15341 506 15351
rect 514 15341 515 15361
rect 504 15325 506 15341
rect 525 15332 528 15366
rect 547 15341 548 15361
rect 557 15341 564 15351
rect 514 15325 530 15331
rect 532 15325 548 15331
rect 332 15277 373 15305
rect 332 15271 351 15277
rect 196 15230 204 15264
rect 216 15230 230 15264
rect 244 15230 257 15264
rect 278 15234 291 15268
rect 300 15252 321 15268
rect 336 15261 351 15271
rect 300 15250 312 15252
rect 300 15234 321 15250
rect 332 15243 351 15261
rect 361 15243 375 15277
rect 400 15271 411 15309
rect 562 15272 612 15274
rect 400 15243 409 15271
rect 466 15263 497 15265
rect 565 15263 596 15265
rect 442 15256 500 15263
rect 466 15255 500 15256
rect 565 15255 599 15263
rect 174 15193 181 15217
rect 224 15183 226 15230
rect 300 15221 308 15234
rect 289 15218 305 15220
rect 332 15193 342 15243
rect 400 15223 404 15243
rect 497 15239 500 15255
rect 596 15239 599 15255
rect 466 15238 500 15239
rect 442 15231 500 15238
rect 565 15231 599 15239
rect 612 15222 614 15272
rect 256 15183 328 15191
rect 336 15185 342 15193
rect 400 15185 404 15193
rect 196 15153 204 15183
rect 216 15153 230 15183
rect 196 15149 230 15153
rect 196 15141 226 15149
rect 224 15125 226 15141
rect 332 15113 336 15181
rect 400 15151 408 15185
rect 434 15151 438 15185
rect 454 15169 504 15171
rect 504 15153 506 15169
rect 514 15163 530 15169
rect 532 15163 548 15169
rect 525 15153 548 15162
rect 400 15143 404 15151
rect 498 15143 506 15153
rect 504 15119 506 15143
rect 514 15133 515 15153
rect 525 15128 528 15153
rect 547 15133 548 15153
rect 557 15143 564 15153
rect 514 15119 548 15123
rect 400 15113 442 15114
rect 174 15103 246 15111
rect 400 15106 404 15113
rect 295 15072 300 15106
rect 324 15072 329 15106
rect 367 15072 438 15106
rect 400 15071 404 15072
rect 378 15065 404 15071
rect 442 15065 464 15071
rect 38 15049 80 15065
rect 400 15049 442 15065
rect -25 15035 25 15037
rect 455 15035 505 15037
rect 557 15035 607 15037
rect 16 15027 102 15035
rect 378 15027 464 15035
rect 8 14993 17 15027
rect 18 15025 51 15027
rect 80 15025 100 15027
rect 18 14993 100 15025
rect 380 15025 404 15027
rect 429 15025 438 15027
rect 442 15025 462 15027
rect 16 14985 102 14993
rect 42 14969 76 14971
rect 16 14949 38 14955
rect 42 14946 76 14950
rect 80 14949 102 14955
rect 42 14916 46 14946
rect 72 14916 76 14946
rect 42 14835 46 14869
rect 72 14835 76 14869
rect -25 14798 25 14800
rect 0 14790 14 14791
rect 0 14789 17 14790
rect 25 14789 27 14798
rect 0 14782 38 14789
rect 0 14781 34 14782
rect 0 14765 8 14781
rect 14 14765 34 14781
rect 0 14764 34 14765
rect 0 14757 38 14764
rect 14 14756 17 14757
rect 25 14748 27 14757
rect 42 14728 45 14818
rect 69 14803 80 14835
rect 107 14803 143 14831
rect 107 14797 119 14803
rect 109 14769 119 14797
rect 129 14769 143 14803
rect 42 14677 46 14711
rect 72 14677 76 14711
rect 38 14639 80 14640
rect 42 14598 76 14632
rect 79 14598 113 14632
rect 42 14519 46 14553
rect 72 14519 76 14553
rect -25 14482 25 14484
rect 0 14474 14 14475
rect 0 14473 17 14474
rect 25 14473 27 14482
rect 0 14466 38 14473
rect 0 14465 34 14466
rect 0 14449 8 14465
rect 14 14449 34 14465
rect 0 14448 34 14449
rect 0 14441 38 14448
rect 14 14440 17 14441
rect 25 14432 27 14441
rect 42 14412 45 14502
rect 71 14471 80 14499
rect 69 14433 80 14471
rect 107 14427 119 14461
rect 129 14433 143 14461
rect 129 14427 141 14433
rect 42 14361 46 14395
rect 72 14361 76 14395
rect 42 14314 76 14318
rect 42 14284 46 14314
rect 72 14284 76 14314
rect 16 14275 38 14281
rect 80 14275 102 14281
rect 144 14275 148 15023
rect 332 14955 336 15023
rect 380 14993 462 15025
rect 463 14993 472 15027
rect 480 14993 497 15027
rect 378 14985 464 14993
rect 505 14985 507 15035
rect 514 14993 548 15027
rect 565 14993 582 15027
rect 607 14985 609 15035
rect 404 14969 438 14971
rect 400 14955 442 14956
rect 378 14949 404 14955
rect 442 14949 464 14955
rect 400 14948 404 14949
rect 174 14909 246 14917
rect 295 14914 300 14948
rect 324 14914 329 14948
rect 224 14879 226 14895
rect 196 14871 226 14879
rect 332 14877 336 14945
rect 367 14914 438 14948
rect 400 14907 404 14914
rect 454 14901 504 14903
rect 494 14897 548 14901
rect 494 14892 514 14897
rect 504 14877 506 14892
rect 196 14867 230 14871
rect 196 14837 204 14867
rect 216 14837 230 14867
rect 400 14869 404 14877
rect 174 14803 181 14829
rect 224 14790 226 14837
rect 256 14829 328 14837
rect 332 14835 336 14865
rect 400 14835 408 14869
rect 434 14835 438 14869
rect 498 14867 506 14877
rect 514 14867 515 14887
rect 504 14851 506 14867
rect 525 14858 528 14892
rect 547 14867 548 14887
rect 557 14867 564 14877
rect 514 14851 530 14857
rect 532 14851 548 14857
rect 289 14800 305 14802
rect 196 14756 204 14790
rect 216 14756 230 14790
rect 244 14756 257 14790
rect 300 14786 308 14799
rect 332 14797 342 14835
rect 400 14827 404 14835
rect 336 14787 342 14797
rect 224 14709 226 14756
rect 278 14752 291 14786
rect 300 14770 321 14786
rect 332 14777 342 14787
rect 400 14787 409 14815
rect 562 14798 612 14800
rect 466 14789 497 14791
rect 565 14789 596 14791
rect 300 14768 312 14770
rect 300 14752 321 14768
rect 300 14746 308 14752
rect 289 14736 308 14746
rect 196 14679 204 14709
rect 216 14679 230 14709
rect 196 14675 230 14679
rect 196 14667 226 14675
rect 300 14667 308 14736
rect 332 14743 351 14777
rect 361 14743 375 14777
rect 400 14743 411 14787
rect 442 14782 500 14789
rect 466 14781 500 14782
rect 565 14781 599 14789
rect 497 14765 500 14781
rect 596 14765 599 14781
rect 466 14764 500 14765
rect 442 14757 500 14764
rect 565 14757 599 14765
rect 612 14748 614 14798
rect 332 14719 342 14743
rect 336 14707 342 14719
rect 224 14651 226 14667
rect 332 14639 342 14707
rect 400 14711 404 14719
rect 400 14677 408 14711
rect 434 14677 438 14711
rect 454 14695 504 14697
rect 504 14679 506 14695
rect 514 14689 530 14695
rect 532 14689 548 14695
rect 525 14679 548 14688
rect 400 14669 404 14677
rect 498 14669 506 14679
rect 504 14645 506 14669
rect 514 14659 515 14679
rect 525 14654 528 14679
rect 547 14659 548 14679
rect 557 14669 564 14679
rect 514 14645 548 14649
rect 151 14598 156 14632
rect 174 14629 246 14637
rect 256 14629 328 14637
rect 336 14631 342 14639
rect 400 14634 404 14639
rect 180 14601 185 14629
rect 174 14593 246 14601
rect 256 14593 328 14601
rect 332 14599 336 14629
rect 400 14600 438 14634
rect 224 14563 226 14579
rect 196 14555 226 14563
rect 196 14551 230 14555
rect 196 14521 204 14551
rect 216 14521 230 14551
rect 224 14474 226 14521
rect 300 14494 308 14563
rect 332 14561 342 14599
rect 400 14591 404 14600
rect 454 14585 504 14587
rect 494 14581 548 14585
rect 494 14576 514 14581
rect 504 14561 506 14576
rect 336 14549 342 14561
rect 289 14484 308 14494
rect 300 14478 308 14484
rect 332 14515 342 14549
rect 400 14553 404 14561
rect 400 14519 408 14553
rect 434 14519 438 14553
rect 498 14551 506 14561
rect 514 14551 515 14571
rect 504 14535 506 14551
rect 525 14542 528 14576
rect 547 14551 548 14571
rect 557 14551 564 14561
rect 514 14535 530 14541
rect 532 14535 548 14541
rect 332 14487 373 14515
rect 332 14481 351 14487
rect 196 14440 204 14474
rect 216 14440 230 14474
rect 244 14440 257 14474
rect 278 14444 291 14478
rect 300 14462 321 14478
rect 336 14471 351 14481
rect 300 14460 312 14462
rect 300 14444 321 14460
rect 332 14453 351 14471
rect 361 14453 375 14487
rect 400 14481 411 14519
rect 562 14482 612 14484
rect 400 14453 409 14481
rect 466 14473 497 14475
rect 565 14473 596 14475
rect 442 14466 500 14473
rect 466 14465 500 14466
rect 565 14465 599 14473
rect 174 14403 181 14427
rect 224 14393 226 14440
rect 300 14431 308 14444
rect 289 14428 305 14430
rect 332 14403 342 14453
rect 400 14433 404 14453
rect 497 14449 500 14465
rect 596 14449 599 14465
rect 466 14448 500 14449
rect 442 14441 500 14448
rect 565 14441 599 14449
rect 612 14432 614 14482
rect 256 14393 328 14401
rect 336 14395 342 14403
rect 400 14395 404 14403
rect 196 14363 204 14393
rect 216 14363 230 14393
rect 196 14359 230 14363
rect 196 14351 226 14359
rect 224 14335 226 14351
rect 332 14323 336 14391
rect 400 14361 408 14395
rect 434 14361 438 14395
rect 454 14379 504 14381
rect 504 14363 506 14379
rect 514 14373 530 14379
rect 532 14373 548 14379
rect 525 14363 548 14372
rect 400 14353 404 14361
rect 498 14353 506 14363
rect 504 14329 506 14353
rect 514 14343 515 14363
rect 525 14338 528 14363
rect 547 14343 548 14363
rect 557 14353 564 14363
rect 514 14329 548 14333
rect 400 14323 442 14324
rect 174 14313 246 14321
rect 400 14316 404 14323
rect 295 14282 300 14316
rect 324 14282 329 14316
rect 367 14282 438 14316
rect 400 14281 404 14282
rect 378 14275 404 14281
rect 442 14275 464 14281
rect 38 14259 80 14275
rect 400 14259 442 14275
rect -25 14245 25 14247
rect 455 14245 505 14247
rect 557 14245 607 14247
rect 16 14237 102 14245
rect 378 14237 464 14245
rect 8 14203 17 14237
rect 18 14235 51 14237
rect 80 14235 100 14237
rect 18 14203 100 14235
rect 380 14235 404 14237
rect 429 14235 438 14237
rect 442 14235 462 14237
rect 16 14195 102 14203
rect 42 14179 76 14181
rect 16 14159 38 14165
rect 42 14156 76 14160
rect 80 14159 102 14165
rect 42 14126 46 14156
rect 72 14126 76 14156
rect 42 14045 46 14079
rect 72 14045 76 14079
rect -25 14008 25 14010
rect 0 14000 14 14001
rect 0 13999 17 14000
rect 25 13999 27 14008
rect 0 13992 38 13999
rect 0 13991 34 13992
rect 0 13975 8 13991
rect 14 13975 34 13991
rect 0 13974 34 13975
rect 0 13967 38 13974
rect 14 13966 17 13967
rect 25 13958 27 13967
rect 42 13938 45 14028
rect 69 14013 80 14045
rect 107 14013 143 14041
rect 107 14007 119 14013
rect 109 13979 119 14007
rect 129 13979 143 14013
rect 42 13887 46 13921
rect 72 13887 76 13921
rect 38 13849 80 13850
rect 42 13808 76 13842
rect 79 13808 113 13842
rect 42 13729 46 13763
rect 72 13729 76 13763
rect -25 13692 25 13694
rect 0 13684 14 13685
rect 0 13683 17 13684
rect 25 13683 27 13692
rect 0 13676 38 13683
rect 0 13675 34 13676
rect 0 13659 8 13675
rect 14 13659 34 13675
rect 0 13658 34 13659
rect 0 13651 38 13658
rect 14 13650 17 13651
rect 25 13642 27 13651
rect 42 13622 45 13712
rect 71 13681 80 13709
rect 69 13643 80 13681
rect 107 13637 119 13671
rect 129 13643 143 13671
rect 129 13637 141 13643
rect 42 13571 46 13605
rect 72 13571 76 13605
rect 42 13524 76 13528
rect 42 13494 46 13524
rect 72 13494 76 13524
rect 16 13485 38 13491
rect 80 13485 102 13491
rect 144 13485 148 14233
rect 332 14165 336 14233
rect 380 14203 462 14235
rect 463 14203 472 14237
rect 480 14203 497 14237
rect 378 14195 464 14203
rect 505 14195 507 14245
rect 514 14203 548 14237
rect 565 14203 582 14237
rect 607 14195 609 14245
rect 404 14179 438 14181
rect 400 14165 442 14166
rect 378 14159 404 14165
rect 442 14159 464 14165
rect 400 14158 404 14159
rect 174 14119 246 14127
rect 295 14124 300 14158
rect 324 14124 329 14158
rect 224 14089 226 14105
rect 196 14081 226 14089
rect 332 14087 336 14155
rect 367 14124 438 14158
rect 400 14117 404 14124
rect 454 14111 504 14113
rect 494 14107 548 14111
rect 494 14102 514 14107
rect 504 14087 506 14102
rect 196 14077 230 14081
rect 196 14047 204 14077
rect 216 14047 230 14077
rect 400 14079 404 14087
rect 174 14013 181 14039
rect 224 14000 226 14047
rect 256 14039 328 14047
rect 332 14045 336 14075
rect 400 14045 408 14079
rect 434 14045 438 14079
rect 498 14077 506 14087
rect 514 14077 515 14097
rect 504 14061 506 14077
rect 525 14068 528 14102
rect 547 14077 548 14097
rect 557 14077 564 14087
rect 514 14061 530 14067
rect 532 14061 548 14067
rect 289 14010 305 14012
rect 196 13966 204 14000
rect 216 13966 230 14000
rect 244 13966 257 14000
rect 300 13996 308 14009
rect 332 14007 342 14045
rect 400 14037 404 14045
rect 336 13997 342 14007
rect 224 13919 226 13966
rect 278 13962 291 13996
rect 300 13980 321 13996
rect 332 13987 342 13997
rect 400 13997 409 14025
rect 562 14008 612 14010
rect 466 13999 497 14001
rect 565 13999 596 14001
rect 300 13978 312 13980
rect 300 13962 321 13978
rect 300 13956 308 13962
rect 289 13946 308 13956
rect 196 13889 204 13919
rect 216 13889 230 13919
rect 196 13885 230 13889
rect 196 13877 226 13885
rect 300 13877 308 13946
rect 332 13953 351 13987
rect 361 13953 375 13987
rect 400 13953 411 13997
rect 442 13992 500 13999
rect 466 13991 500 13992
rect 565 13991 599 13999
rect 497 13975 500 13991
rect 596 13975 599 13991
rect 466 13974 500 13975
rect 442 13967 500 13974
rect 565 13967 599 13975
rect 612 13958 614 14008
rect 332 13929 342 13953
rect 336 13917 342 13929
rect 224 13861 226 13877
rect 332 13849 342 13917
rect 400 13921 404 13929
rect 400 13887 408 13921
rect 434 13887 438 13921
rect 454 13905 504 13907
rect 504 13889 506 13905
rect 514 13899 530 13905
rect 532 13899 548 13905
rect 525 13889 548 13898
rect 400 13879 404 13887
rect 498 13879 506 13889
rect 504 13855 506 13879
rect 514 13869 515 13889
rect 525 13864 528 13889
rect 547 13869 548 13889
rect 557 13879 564 13889
rect 514 13855 548 13859
rect 151 13808 156 13842
rect 174 13839 246 13847
rect 256 13839 328 13847
rect 336 13841 342 13849
rect 400 13844 404 13849
rect 180 13811 185 13839
rect 174 13803 246 13811
rect 256 13803 328 13811
rect 332 13809 336 13839
rect 400 13810 438 13844
rect 224 13773 226 13789
rect 196 13765 226 13773
rect 196 13761 230 13765
rect 196 13731 204 13761
rect 216 13731 230 13761
rect 224 13684 226 13731
rect 300 13704 308 13773
rect 332 13771 342 13809
rect 400 13801 404 13810
rect 454 13795 504 13797
rect 494 13791 548 13795
rect 494 13786 514 13791
rect 504 13771 506 13786
rect 336 13759 342 13771
rect 289 13694 308 13704
rect 300 13688 308 13694
rect 332 13725 342 13759
rect 400 13763 404 13771
rect 400 13729 408 13763
rect 434 13729 438 13763
rect 498 13761 506 13771
rect 514 13761 515 13781
rect 504 13745 506 13761
rect 525 13752 528 13786
rect 547 13761 548 13781
rect 557 13761 564 13771
rect 514 13745 530 13751
rect 532 13745 548 13751
rect 332 13697 373 13725
rect 332 13691 351 13697
rect 196 13650 204 13684
rect 216 13650 230 13684
rect 244 13650 257 13684
rect 278 13654 291 13688
rect 300 13672 321 13688
rect 336 13681 351 13691
rect 300 13670 312 13672
rect 300 13654 321 13670
rect 332 13663 351 13681
rect 361 13663 375 13697
rect 400 13691 411 13729
rect 562 13692 612 13694
rect 400 13663 409 13691
rect 466 13683 497 13685
rect 565 13683 596 13685
rect 442 13676 500 13683
rect 466 13675 500 13676
rect 565 13675 599 13683
rect 174 13613 181 13637
rect 224 13603 226 13650
rect 300 13641 308 13654
rect 289 13638 305 13640
rect 332 13613 342 13663
rect 400 13643 404 13663
rect 497 13659 500 13675
rect 596 13659 599 13675
rect 466 13658 500 13659
rect 442 13651 500 13658
rect 565 13651 599 13659
rect 612 13642 614 13692
rect 256 13603 328 13611
rect 336 13605 342 13613
rect 400 13605 404 13613
rect 196 13573 204 13603
rect 216 13573 230 13603
rect 196 13569 230 13573
rect 196 13561 226 13569
rect 224 13545 226 13561
rect 332 13533 336 13601
rect 400 13571 408 13605
rect 434 13571 438 13605
rect 454 13589 504 13591
rect 504 13573 506 13589
rect 514 13583 530 13589
rect 532 13583 548 13589
rect 525 13573 548 13582
rect 400 13563 404 13571
rect 498 13563 506 13573
rect 504 13539 506 13563
rect 514 13553 515 13573
rect 525 13548 528 13573
rect 547 13553 548 13573
rect 557 13563 564 13573
rect 514 13539 548 13543
rect 400 13533 442 13534
rect 174 13523 246 13531
rect 400 13526 404 13533
rect 295 13492 300 13526
rect 324 13492 329 13526
rect 367 13492 438 13526
rect 400 13491 404 13492
rect 378 13485 404 13491
rect 442 13485 464 13491
rect 38 13469 80 13485
rect 400 13469 442 13485
rect -25 13455 25 13457
rect 455 13455 505 13457
rect 557 13455 607 13457
rect 16 13447 102 13455
rect 378 13447 464 13455
rect 8 13413 17 13447
rect 18 13445 51 13447
rect 80 13445 100 13447
rect 18 13413 100 13445
rect 380 13445 404 13447
rect 429 13445 438 13447
rect 442 13445 462 13447
rect 16 13405 102 13413
rect 42 13389 76 13391
rect 16 13369 38 13375
rect 42 13366 76 13370
rect 80 13369 102 13375
rect 42 13336 46 13366
rect 72 13336 76 13366
rect 42 13255 46 13289
rect 72 13255 76 13289
rect -25 13218 25 13220
rect 0 13210 14 13211
rect 0 13209 17 13210
rect 25 13209 27 13218
rect 0 13202 38 13209
rect 0 13201 34 13202
rect 0 13185 8 13201
rect 14 13185 34 13201
rect 0 13184 34 13185
rect 0 13177 38 13184
rect 14 13176 17 13177
rect 25 13168 27 13177
rect 42 13148 45 13238
rect 69 13223 80 13255
rect 107 13223 143 13251
rect 107 13217 119 13223
rect 109 13189 119 13217
rect 129 13189 143 13223
rect 42 13097 46 13131
rect 72 13097 76 13131
rect 38 13059 80 13060
rect 42 13018 76 13052
rect 79 13018 113 13052
rect 42 12939 46 12973
rect 72 12939 76 12973
rect -25 12902 25 12904
rect 0 12894 14 12895
rect 0 12893 17 12894
rect 25 12893 27 12902
rect 0 12886 38 12893
rect 0 12885 34 12886
rect 0 12869 8 12885
rect 14 12869 34 12885
rect 0 12868 34 12869
rect 0 12861 38 12868
rect 14 12860 17 12861
rect 25 12852 27 12861
rect 42 12832 45 12922
rect 71 12891 80 12919
rect 69 12853 80 12891
rect 107 12847 119 12881
rect 129 12853 143 12881
rect 129 12847 141 12853
rect 42 12781 46 12815
rect 72 12781 76 12815
rect 42 12734 76 12738
rect 42 12704 46 12734
rect 72 12704 76 12734
rect 16 12695 38 12701
rect 80 12695 102 12701
rect 144 12695 148 13443
rect 332 13375 336 13443
rect 380 13413 462 13445
rect 463 13413 472 13447
rect 480 13413 497 13447
rect 378 13405 464 13413
rect 505 13405 507 13455
rect 514 13413 548 13447
rect 565 13413 582 13447
rect 607 13405 609 13455
rect 404 13389 438 13391
rect 400 13375 442 13376
rect 378 13369 404 13375
rect 442 13369 464 13375
rect 400 13368 404 13369
rect 174 13329 246 13337
rect 295 13334 300 13368
rect 324 13334 329 13368
rect 224 13299 226 13315
rect 196 13291 226 13299
rect 332 13297 336 13365
rect 367 13334 438 13368
rect 400 13327 404 13334
rect 454 13321 504 13323
rect 494 13317 548 13321
rect 494 13312 514 13317
rect 504 13297 506 13312
rect 196 13287 230 13291
rect 196 13257 204 13287
rect 216 13257 230 13287
rect 400 13289 404 13297
rect 174 13223 181 13249
rect 224 13210 226 13257
rect 256 13249 328 13257
rect 332 13255 336 13285
rect 400 13255 408 13289
rect 434 13255 438 13289
rect 498 13287 506 13297
rect 514 13287 515 13307
rect 504 13271 506 13287
rect 525 13278 528 13312
rect 547 13287 548 13307
rect 557 13287 564 13297
rect 514 13271 530 13277
rect 532 13271 548 13277
rect 289 13220 305 13222
rect 196 13176 204 13210
rect 216 13176 230 13210
rect 244 13176 257 13210
rect 300 13206 308 13219
rect 332 13217 342 13255
rect 400 13247 404 13255
rect 336 13207 342 13217
rect 224 13129 226 13176
rect 278 13172 291 13206
rect 300 13190 321 13206
rect 332 13197 342 13207
rect 400 13207 409 13235
rect 562 13218 612 13220
rect 466 13209 497 13211
rect 565 13209 596 13211
rect 300 13188 312 13190
rect 300 13172 321 13188
rect 300 13166 308 13172
rect 289 13156 308 13166
rect 196 13099 204 13129
rect 216 13099 230 13129
rect 196 13095 230 13099
rect 196 13087 226 13095
rect 300 13087 308 13156
rect 332 13163 351 13197
rect 361 13163 375 13197
rect 400 13163 411 13207
rect 442 13202 500 13209
rect 466 13201 500 13202
rect 565 13201 599 13209
rect 497 13185 500 13201
rect 596 13185 599 13201
rect 466 13184 500 13185
rect 442 13177 500 13184
rect 565 13177 599 13185
rect 612 13168 614 13218
rect 332 13139 342 13163
rect 336 13127 342 13139
rect 224 13071 226 13087
rect 332 13059 342 13127
rect 400 13131 404 13139
rect 400 13097 408 13131
rect 434 13097 438 13131
rect 454 13115 504 13117
rect 504 13099 506 13115
rect 514 13109 530 13115
rect 532 13109 548 13115
rect 525 13099 548 13108
rect 400 13089 404 13097
rect 498 13089 506 13099
rect 504 13065 506 13089
rect 514 13079 515 13099
rect 525 13074 528 13099
rect 547 13079 548 13099
rect 557 13089 564 13099
rect 514 13065 548 13069
rect 151 13018 156 13052
rect 174 13049 246 13057
rect 256 13049 328 13057
rect 336 13051 342 13059
rect 400 13054 404 13059
rect 180 13021 185 13049
rect 174 13013 246 13021
rect 256 13013 328 13021
rect 332 13019 336 13049
rect 400 13020 438 13054
rect 224 12983 226 12999
rect 196 12975 226 12983
rect 196 12971 230 12975
rect 196 12941 204 12971
rect 216 12941 230 12971
rect 224 12894 226 12941
rect 300 12914 308 12983
rect 332 12981 342 13019
rect 400 13011 404 13020
rect 454 13005 504 13007
rect 494 13001 548 13005
rect 494 12996 514 13001
rect 504 12981 506 12996
rect 336 12969 342 12981
rect 289 12904 308 12914
rect 300 12898 308 12904
rect 332 12935 342 12969
rect 400 12973 404 12981
rect 400 12939 408 12973
rect 434 12939 438 12973
rect 498 12971 506 12981
rect 514 12971 515 12991
rect 504 12955 506 12971
rect 525 12962 528 12996
rect 547 12971 548 12991
rect 557 12971 564 12981
rect 514 12955 530 12961
rect 532 12955 548 12961
rect 332 12907 373 12935
rect 332 12901 351 12907
rect 196 12860 204 12894
rect 216 12860 230 12894
rect 244 12860 257 12894
rect 278 12864 291 12898
rect 300 12882 321 12898
rect 336 12891 351 12901
rect 300 12880 312 12882
rect 300 12864 321 12880
rect 332 12873 351 12891
rect 361 12873 375 12907
rect 400 12901 411 12939
rect 562 12902 612 12904
rect 400 12873 409 12901
rect 466 12893 497 12895
rect 565 12893 596 12895
rect 442 12886 500 12893
rect 466 12885 500 12886
rect 565 12885 599 12893
rect 174 12823 181 12847
rect 224 12813 226 12860
rect 300 12851 308 12864
rect 289 12848 305 12850
rect 332 12823 342 12873
rect 400 12853 404 12873
rect 497 12869 500 12885
rect 596 12869 599 12885
rect 466 12868 500 12869
rect 442 12861 500 12868
rect 565 12861 599 12869
rect 612 12852 614 12902
rect 256 12813 328 12821
rect 336 12815 342 12823
rect 400 12815 404 12823
rect 196 12783 204 12813
rect 216 12783 230 12813
rect 196 12779 230 12783
rect 196 12771 226 12779
rect 224 12755 226 12771
rect 332 12743 336 12811
rect 400 12781 408 12815
rect 434 12781 438 12815
rect 454 12799 504 12801
rect 504 12783 506 12799
rect 514 12793 530 12799
rect 532 12793 548 12799
rect 525 12783 548 12792
rect 400 12773 404 12781
rect 498 12773 506 12783
rect 504 12749 506 12773
rect 514 12763 515 12783
rect 525 12758 528 12783
rect 547 12763 548 12783
rect 557 12773 564 12783
rect 514 12749 548 12753
rect 400 12743 442 12744
rect 174 12733 246 12741
rect 400 12736 404 12743
rect 295 12702 300 12736
rect 324 12702 329 12736
rect 367 12702 438 12736
rect 400 12701 404 12702
rect 378 12695 404 12701
rect 442 12695 464 12701
rect 38 12679 80 12695
rect 400 12679 442 12695
rect -25 12665 25 12667
rect 455 12665 505 12667
rect 557 12665 607 12667
rect 16 12657 102 12665
rect 378 12657 464 12665
rect 8 12623 17 12657
rect 18 12655 51 12657
rect 80 12655 100 12657
rect 18 12623 100 12655
rect 380 12655 404 12657
rect 429 12655 438 12657
rect 442 12655 462 12657
rect 16 12615 102 12623
rect 42 12599 76 12601
rect 16 12579 38 12585
rect 42 12576 76 12580
rect 80 12579 102 12585
rect 42 12546 46 12576
rect 72 12546 76 12576
rect 42 12465 46 12499
rect 72 12465 76 12499
rect -25 12428 25 12430
rect 0 12420 14 12421
rect 0 12419 17 12420
rect 25 12419 27 12428
rect 0 12412 38 12419
rect 0 12411 34 12412
rect 0 12395 8 12411
rect 14 12395 34 12411
rect 0 12394 34 12395
rect 0 12387 38 12394
rect 14 12386 17 12387
rect 25 12378 27 12387
rect 42 12358 45 12448
rect 69 12433 80 12465
rect 107 12433 143 12461
rect 107 12427 119 12433
rect 109 12399 119 12427
rect 129 12399 143 12433
rect 42 12307 46 12341
rect 72 12307 76 12341
rect 38 12269 80 12270
rect 42 12228 76 12262
rect 79 12228 113 12262
rect 42 12149 46 12183
rect 72 12149 76 12183
rect -25 12112 25 12114
rect 0 12104 14 12105
rect 0 12103 17 12104
rect 25 12103 27 12112
rect 0 12096 38 12103
rect 0 12095 34 12096
rect 0 12079 8 12095
rect 14 12079 34 12095
rect 0 12078 34 12079
rect 0 12071 38 12078
rect 14 12070 17 12071
rect 25 12062 27 12071
rect 42 12042 45 12132
rect 71 12101 80 12129
rect 69 12063 80 12101
rect 107 12057 119 12091
rect 129 12063 143 12091
rect 129 12057 141 12063
rect 42 11991 46 12025
rect 72 11991 76 12025
rect 42 11944 76 11948
rect 42 11914 46 11944
rect 72 11914 76 11944
rect 16 11905 38 11911
rect 80 11905 102 11911
rect 144 11905 148 12653
rect 332 12585 336 12653
rect 380 12623 462 12655
rect 463 12623 472 12657
rect 480 12623 497 12657
rect 378 12615 464 12623
rect 505 12615 507 12665
rect 514 12623 548 12657
rect 565 12623 582 12657
rect 607 12615 609 12665
rect 404 12599 438 12601
rect 400 12585 442 12586
rect 378 12579 404 12585
rect 442 12579 464 12585
rect 400 12578 404 12579
rect 174 12539 246 12547
rect 295 12544 300 12578
rect 324 12544 329 12578
rect 224 12509 226 12525
rect 196 12501 226 12509
rect 332 12507 336 12575
rect 367 12544 438 12578
rect 400 12537 404 12544
rect 454 12531 504 12533
rect 494 12527 548 12531
rect 494 12522 514 12527
rect 504 12507 506 12522
rect 196 12497 230 12501
rect 196 12467 204 12497
rect 216 12467 230 12497
rect 400 12499 404 12507
rect 174 12433 181 12459
rect 224 12420 226 12467
rect 256 12459 328 12467
rect 332 12465 336 12495
rect 400 12465 408 12499
rect 434 12465 438 12499
rect 498 12497 506 12507
rect 514 12497 515 12517
rect 504 12481 506 12497
rect 525 12488 528 12522
rect 547 12497 548 12517
rect 557 12497 564 12507
rect 514 12481 530 12487
rect 532 12481 548 12487
rect 289 12430 305 12432
rect 196 12386 204 12420
rect 216 12386 230 12420
rect 244 12386 257 12420
rect 300 12416 308 12429
rect 332 12427 342 12465
rect 400 12457 404 12465
rect 336 12417 342 12427
rect 224 12339 226 12386
rect 278 12382 291 12416
rect 300 12400 321 12416
rect 332 12407 342 12417
rect 400 12417 409 12445
rect 562 12428 612 12430
rect 466 12419 497 12421
rect 565 12419 596 12421
rect 300 12398 312 12400
rect 300 12382 321 12398
rect 300 12376 308 12382
rect 289 12366 308 12376
rect 196 12309 204 12339
rect 216 12309 230 12339
rect 196 12305 230 12309
rect 196 12297 226 12305
rect 300 12297 308 12366
rect 332 12373 351 12407
rect 361 12373 375 12407
rect 400 12373 411 12417
rect 442 12412 500 12419
rect 466 12411 500 12412
rect 565 12411 599 12419
rect 497 12395 500 12411
rect 596 12395 599 12411
rect 466 12394 500 12395
rect 442 12387 500 12394
rect 565 12387 599 12395
rect 612 12378 614 12428
rect 332 12349 342 12373
rect 336 12337 342 12349
rect 224 12281 226 12297
rect 332 12269 342 12337
rect 400 12341 404 12349
rect 400 12307 408 12341
rect 434 12307 438 12341
rect 454 12325 504 12327
rect 504 12309 506 12325
rect 514 12319 530 12325
rect 532 12319 548 12325
rect 525 12309 548 12318
rect 400 12299 404 12307
rect 498 12299 506 12309
rect 504 12275 506 12299
rect 514 12289 515 12309
rect 525 12284 528 12309
rect 547 12289 548 12309
rect 557 12299 564 12309
rect 514 12275 548 12279
rect 151 12228 156 12262
rect 174 12259 246 12267
rect 256 12259 328 12267
rect 336 12261 342 12269
rect 400 12264 404 12269
rect 180 12231 185 12259
rect 174 12223 246 12231
rect 256 12223 328 12231
rect 332 12229 336 12259
rect 400 12230 438 12264
rect 224 12193 226 12209
rect 196 12185 226 12193
rect 196 12181 230 12185
rect 196 12151 204 12181
rect 216 12151 230 12181
rect 224 12104 226 12151
rect 300 12124 308 12193
rect 332 12191 342 12229
rect 400 12221 404 12230
rect 454 12215 504 12217
rect 494 12211 548 12215
rect 494 12206 514 12211
rect 504 12191 506 12206
rect 336 12179 342 12191
rect 289 12114 308 12124
rect 300 12108 308 12114
rect 332 12145 342 12179
rect 400 12183 404 12191
rect 400 12149 408 12183
rect 434 12149 438 12183
rect 498 12181 506 12191
rect 514 12181 515 12201
rect 504 12165 506 12181
rect 525 12172 528 12206
rect 547 12181 548 12201
rect 557 12181 564 12191
rect 514 12165 530 12171
rect 532 12165 548 12171
rect 332 12117 373 12145
rect 332 12111 351 12117
rect 196 12070 204 12104
rect 216 12070 230 12104
rect 244 12070 257 12104
rect 278 12074 291 12108
rect 300 12092 321 12108
rect 336 12101 351 12111
rect 300 12090 312 12092
rect 300 12074 321 12090
rect 332 12083 351 12101
rect 361 12083 375 12117
rect 400 12111 411 12149
rect 562 12112 612 12114
rect 400 12083 409 12111
rect 466 12103 497 12105
rect 565 12103 596 12105
rect 442 12096 500 12103
rect 466 12095 500 12096
rect 565 12095 599 12103
rect 174 12033 181 12057
rect 224 12023 226 12070
rect 300 12061 308 12074
rect 289 12058 305 12060
rect 332 12033 342 12083
rect 400 12063 404 12083
rect 497 12079 500 12095
rect 596 12079 599 12095
rect 466 12078 500 12079
rect 442 12071 500 12078
rect 565 12071 599 12079
rect 612 12062 614 12112
rect 256 12023 328 12031
rect 336 12025 342 12033
rect 400 12025 404 12033
rect 196 11993 204 12023
rect 216 11993 230 12023
rect 196 11989 230 11993
rect 196 11981 226 11989
rect 224 11965 226 11981
rect 332 11953 336 12021
rect 400 11991 408 12025
rect 434 11991 438 12025
rect 454 12009 504 12011
rect 504 11993 506 12009
rect 514 12003 530 12009
rect 532 12003 548 12009
rect 525 11993 548 12002
rect 400 11983 404 11991
rect 498 11983 506 11993
rect 504 11959 506 11983
rect 514 11973 515 11993
rect 525 11968 528 11993
rect 547 11973 548 11993
rect 557 11983 564 11993
rect 514 11959 548 11963
rect 400 11953 442 11954
rect 174 11943 246 11951
rect 400 11946 404 11953
rect 295 11912 300 11946
rect 324 11912 329 11946
rect 367 11912 438 11946
rect 400 11911 404 11912
rect 378 11905 404 11911
rect 442 11905 464 11911
rect 38 11889 80 11905
rect 400 11889 442 11905
rect -25 11875 25 11877
rect 455 11875 505 11877
rect 557 11875 607 11877
rect 16 11867 102 11875
rect 378 11867 464 11875
rect 8 11833 17 11867
rect 18 11865 51 11867
rect 80 11865 100 11867
rect 18 11833 100 11865
rect 380 11865 404 11867
rect 429 11865 438 11867
rect 442 11865 462 11867
rect 16 11825 102 11833
rect 42 11809 76 11811
rect 16 11789 38 11795
rect 42 11786 76 11790
rect 80 11789 102 11795
rect 42 11756 46 11786
rect 72 11756 76 11786
rect 42 11675 46 11709
rect 72 11675 76 11709
rect -25 11638 25 11640
rect 0 11630 14 11631
rect 0 11629 17 11630
rect 25 11629 27 11638
rect 0 11622 38 11629
rect 0 11621 34 11622
rect 0 11605 8 11621
rect 14 11605 34 11621
rect 0 11604 34 11605
rect 0 11597 38 11604
rect 14 11596 17 11597
rect 25 11588 27 11597
rect 42 11568 45 11658
rect 69 11643 80 11675
rect 107 11643 143 11671
rect 107 11637 119 11643
rect 109 11609 119 11637
rect 129 11609 143 11643
rect 42 11517 46 11551
rect 72 11517 76 11551
rect 38 11479 80 11480
rect 42 11438 76 11472
rect 79 11438 113 11472
rect 42 11359 46 11393
rect 72 11359 76 11393
rect -25 11322 25 11324
rect 0 11314 14 11315
rect 0 11313 17 11314
rect 25 11313 27 11322
rect 0 11306 38 11313
rect 0 11305 34 11306
rect 0 11289 8 11305
rect 14 11289 34 11305
rect 0 11288 34 11289
rect 0 11281 38 11288
rect 14 11280 17 11281
rect 25 11272 27 11281
rect 42 11252 45 11342
rect 71 11311 80 11339
rect 69 11273 80 11311
rect 107 11267 119 11301
rect 129 11273 143 11301
rect 129 11267 141 11273
rect 42 11201 46 11235
rect 72 11201 76 11235
rect 42 11154 76 11158
rect 42 11124 46 11154
rect 72 11124 76 11154
rect 16 11115 38 11121
rect 80 11115 102 11121
rect 144 11115 148 11863
rect 332 11795 336 11863
rect 380 11833 462 11865
rect 463 11833 472 11867
rect 480 11833 497 11867
rect 378 11825 464 11833
rect 505 11825 507 11875
rect 514 11833 548 11867
rect 565 11833 582 11867
rect 607 11825 609 11875
rect 404 11809 438 11811
rect 400 11795 442 11796
rect 378 11789 404 11795
rect 442 11789 464 11795
rect 400 11788 404 11789
rect 174 11749 246 11757
rect 295 11754 300 11788
rect 324 11754 329 11788
rect 224 11719 226 11735
rect 196 11711 226 11719
rect 332 11717 336 11785
rect 367 11754 438 11788
rect 400 11747 404 11754
rect 454 11741 504 11743
rect 494 11737 548 11741
rect 494 11732 514 11737
rect 504 11717 506 11732
rect 196 11707 230 11711
rect 196 11677 204 11707
rect 216 11677 230 11707
rect 400 11709 404 11717
rect 174 11643 181 11669
rect 224 11630 226 11677
rect 256 11669 328 11677
rect 332 11675 336 11705
rect 400 11675 408 11709
rect 434 11675 438 11709
rect 498 11707 506 11717
rect 514 11707 515 11727
rect 504 11691 506 11707
rect 525 11698 528 11732
rect 547 11707 548 11727
rect 557 11707 564 11717
rect 514 11691 530 11697
rect 532 11691 548 11697
rect 289 11640 305 11642
rect 196 11596 204 11630
rect 216 11596 230 11630
rect 244 11596 257 11630
rect 300 11626 308 11639
rect 332 11637 342 11675
rect 400 11667 404 11675
rect 336 11627 342 11637
rect 224 11549 226 11596
rect 278 11592 291 11626
rect 300 11610 321 11626
rect 332 11617 342 11627
rect 400 11627 409 11655
rect 562 11638 612 11640
rect 466 11629 497 11631
rect 565 11629 596 11631
rect 300 11608 312 11610
rect 300 11592 321 11608
rect 300 11586 308 11592
rect 289 11576 308 11586
rect 196 11519 204 11549
rect 216 11519 230 11549
rect 196 11515 230 11519
rect 196 11507 226 11515
rect 300 11507 308 11576
rect 332 11583 351 11617
rect 361 11583 375 11617
rect 400 11583 411 11627
rect 442 11622 500 11629
rect 466 11621 500 11622
rect 565 11621 599 11629
rect 497 11605 500 11621
rect 596 11605 599 11621
rect 466 11604 500 11605
rect 442 11597 500 11604
rect 565 11597 599 11605
rect 612 11588 614 11638
rect 332 11559 342 11583
rect 336 11547 342 11559
rect 224 11491 226 11507
rect 332 11479 342 11547
rect 400 11551 404 11559
rect 400 11517 408 11551
rect 434 11517 438 11551
rect 454 11535 504 11537
rect 504 11519 506 11535
rect 514 11529 530 11535
rect 532 11529 548 11535
rect 525 11519 548 11528
rect 400 11509 404 11517
rect 498 11509 506 11519
rect 504 11485 506 11509
rect 514 11499 515 11519
rect 525 11494 528 11519
rect 547 11499 548 11519
rect 557 11509 564 11519
rect 514 11485 548 11489
rect 151 11438 156 11472
rect 174 11469 246 11477
rect 256 11469 328 11477
rect 336 11471 342 11479
rect 400 11474 404 11479
rect 180 11441 185 11469
rect 174 11433 246 11441
rect 256 11433 328 11441
rect 332 11439 336 11469
rect 400 11440 438 11474
rect 224 11403 226 11419
rect 196 11395 226 11403
rect 196 11391 230 11395
rect 196 11361 204 11391
rect 216 11361 230 11391
rect 224 11314 226 11361
rect 300 11334 308 11403
rect 332 11401 342 11439
rect 400 11431 404 11440
rect 454 11425 504 11427
rect 494 11421 548 11425
rect 494 11416 514 11421
rect 504 11401 506 11416
rect 336 11389 342 11401
rect 289 11324 308 11334
rect 300 11318 308 11324
rect 332 11355 342 11389
rect 400 11393 404 11401
rect 400 11359 408 11393
rect 434 11359 438 11393
rect 498 11391 506 11401
rect 514 11391 515 11411
rect 504 11375 506 11391
rect 525 11382 528 11416
rect 547 11391 548 11411
rect 557 11391 564 11401
rect 514 11375 530 11381
rect 532 11375 548 11381
rect 332 11327 373 11355
rect 332 11321 351 11327
rect 196 11280 204 11314
rect 216 11280 230 11314
rect 244 11280 257 11314
rect 278 11284 291 11318
rect 300 11302 321 11318
rect 336 11311 351 11321
rect 300 11300 312 11302
rect 300 11284 321 11300
rect 332 11293 351 11311
rect 361 11293 375 11327
rect 400 11321 411 11359
rect 562 11322 612 11324
rect 400 11293 409 11321
rect 466 11313 497 11315
rect 565 11313 596 11315
rect 442 11306 500 11313
rect 466 11305 500 11306
rect 565 11305 599 11313
rect 174 11243 181 11267
rect 224 11233 226 11280
rect 300 11271 308 11284
rect 289 11268 305 11270
rect 332 11243 342 11293
rect 400 11273 404 11293
rect 497 11289 500 11305
rect 596 11289 599 11305
rect 466 11288 500 11289
rect 442 11281 500 11288
rect 565 11281 599 11289
rect 612 11272 614 11322
rect 256 11233 328 11241
rect 336 11235 342 11243
rect 400 11235 404 11243
rect 196 11203 204 11233
rect 216 11203 230 11233
rect 196 11199 230 11203
rect 196 11191 226 11199
rect 224 11175 226 11191
rect 332 11163 336 11231
rect 400 11201 408 11235
rect 434 11201 438 11235
rect 454 11219 504 11221
rect 504 11203 506 11219
rect 514 11213 530 11219
rect 532 11213 548 11219
rect 525 11203 548 11212
rect 400 11193 404 11201
rect 498 11193 506 11203
rect 504 11169 506 11193
rect 514 11183 515 11203
rect 525 11178 528 11203
rect 547 11183 548 11203
rect 557 11193 564 11203
rect 514 11169 548 11173
rect 400 11163 442 11164
rect 174 11153 246 11161
rect 400 11156 404 11163
rect 295 11122 300 11156
rect 324 11122 329 11156
rect 367 11122 438 11156
rect 400 11121 404 11122
rect 378 11115 404 11121
rect 442 11115 464 11121
rect 38 11099 80 11115
rect 400 11099 442 11115
rect -25 11085 25 11087
rect 455 11085 505 11087
rect 557 11085 607 11087
rect 16 11077 102 11085
rect 378 11077 464 11085
rect 8 11043 17 11077
rect 18 11075 51 11077
rect 80 11075 100 11077
rect 18 11043 100 11075
rect 380 11075 404 11077
rect 429 11075 438 11077
rect 442 11075 462 11077
rect 16 11035 102 11043
rect 42 11019 76 11021
rect 16 10999 38 11005
rect 42 10996 76 11000
rect 80 10999 102 11005
rect 42 10966 46 10996
rect 72 10966 76 10996
rect 42 10885 46 10919
rect 72 10885 76 10919
rect -25 10848 25 10850
rect 0 10840 14 10841
rect 0 10839 17 10840
rect 25 10839 27 10848
rect 0 10832 38 10839
rect 0 10831 34 10832
rect 0 10815 8 10831
rect 14 10815 34 10831
rect 0 10814 34 10815
rect 0 10807 38 10814
rect 14 10806 17 10807
rect 25 10798 27 10807
rect 42 10778 45 10868
rect 69 10853 80 10885
rect 107 10853 143 10881
rect 107 10847 119 10853
rect 109 10819 119 10847
rect 129 10819 143 10853
rect 42 10727 46 10761
rect 72 10727 76 10761
rect 38 10689 80 10690
rect 42 10648 76 10682
rect 79 10648 113 10682
rect 42 10569 46 10603
rect 72 10569 76 10603
rect -25 10532 25 10534
rect 0 10524 14 10525
rect 0 10523 17 10524
rect 25 10523 27 10532
rect 0 10516 38 10523
rect 0 10515 34 10516
rect 0 10499 8 10515
rect 14 10499 34 10515
rect 0 10498 34 10499
rect 0 10491 38 10498
rect 14 10490 17 10491
rect 25 10482 27 10491
rect 42 10462 45 10552
rect 71 10521 80 10549
rect 69 10483 80 10521
rect 107 10477 119 10511
rect 129 10483 143 10511
rect 129 10477 141 10483
rect 42 10411 46 10445
rect 72 10411 76 10445
rect 42 10364 76 10368
rect 42 10334 46 10364
rect 72 10334 76 10364
rect 16 10325 38 10331
rect 80 10325 102 10331
rect 144 10325 148 11073
rect 332 11005 336 11073
rect 380 11043 462 11075
rect 463 11043 472 11077
rect 480 11043 497 11077
rect 378 11035 464 11043
rect 505 11035 507 11085
rect 514 11043 548 11077
rect 565 11043 582 11077
rect 607 11035 609 11085
rect 404 11019 438 11021
rect 400 11005 442 11006
rect 378 10999 404 11005
rect 442 10999 464 11005
rect 400 10998 404 10999
rect 174 10959 246 10967
rect 295 10964 300 10998
rect 324 10964 329 10998
rect 224 10929 226 10945
rect 196 10921 226 10929
rect 332 10927 336 10995
rect 367 10964 438 10998
rect 400 10957 404 10964
rect 454 10951 504 10953
rect 494 10947 548 10951
rect 494 10942 514 10947
rect 504 10927 506 10942
rect 196 10917 230 10921
rect 196 10887 204 10917
rect 216 10887 230 10917
rect 400 10919 404 10927
rect 174 10853 181 10879
rect 224 10840 226 10887
rect 256 10879 328 10887
rect 332 10885 336 10915
rect 400 10885 408 10919
rect 434 10885 438 10919
rect 498 10917 506 10927
rect 514 10917 515 10937
rect 504 10901 506 10917
rect 525 10908 528 10942
rect 547 10917 548 10937
rect 557 10917 564 10927
rect 514 10901 530 10907
rect 532 10901 548 10907
rect 289 10850 305 10852
rect 196 10806 204 10840
rect 216 10806 230 10840
rect 244 10806 257 10840
rect 300 10836 308 10849
rect 332 10847 342 10885
rect 400 10877 404 10885
rect 336 10837 342 10847
rect 224 10759 226 10806
rect 278 10802 291 10836
rect 300 10820 321 10836
rect 332 10827 342 10837
rect 400 10837 409 10865
rect 562 10848 612 10850
rect 466 10839 497 10841
rect 565 10839 596 10841
rect 300 10818 312 10820
rect 300 10802 321 10818
rect 300 10796 308 10802
rect 289 10786 308 10796
rect 196 10729 204 10759
rect 216 10729 230 10759
rect 196 10725 230 10729
rect 196 10717 226 10725
rect 300 10717 308 10786
rect 332 10793 351 10827
rect 361 10793 375 10827
rect 400 10793 411 10837
rect 442 10832 500 10839
rect 466 10831 500 10832
rect 565 10831 599 10839
rect 497 10815 500 10831
rect 596 10815 599 10831
rect 466 10814 500 10815
rect 442 10807 500 10814
rect 565 10807 599 10815
rect 612 10798 614 10848
rect 332 10769 342 10793
rect 336 10757 342 10769
rect 224 10701 226 10717
rect 332 10689 342 10757
rect 400 10761 404 10769
rect 400 10727 408 10761
rect 434 10727 438 10761
rect 454 10745 504 10747
rect 504 10729 506 10745
rect 514 10739 530 10745
rect 532 10739 548 10745
rect 525 10729 548 10738
rect 400 10719 404 10727
rect 498 10719 506 10729
rect 504 10695 506 10719
rect 514 10709 515 10729
rect 525 10704 528 10729
rect 547 10709 548 10729
rect 557 10719 564 10729
rect 514 10695 548 10699
rect 151 10648 156 10682
rect 174 10679 246 10687
rect 256 10679 328 10687
rect 336 10681 342 10689
rect 400 10684 404 10689
rect 180 10651 185 10679
rect 174 10643 246 10651
rect 256 10643 328 10651
rect 332 10649 336 10679
rect 400 10650 438 10684
rect 224 10613 226 10629
rect 196 10605 226 10613
rect 196 10601 230 10605
rect 196 10571 204 10601
rect 216 10571 230 10601
rect 224 10524 226 10571
rect 300 10544 308 10613
rect 332 10611 342 10649
rect 400 10641 404 10650
rect 454 10635 504 10637
rect 494 10631 548 10635
rect 494 10626 514 10631
rect 504 10611 506 10626
rect 336 10599 342 10611
rect 289 10534 308 10544
rect 300 10528 308 10534
rect 332 10565 342 10599
rect 400 10603 404 10611
rect 400 10569 408 10603
rect 434 10569 438 10603
rect 498 10601 506 10611
rect 514 10601 515 10621
rect 504 10585 506 10601
rect 525 10592 528 10626
rect 547 10601 548 10621
rect 557 10601 564 10611
rect 514 10585 530 10591
rect 532 10585 548 10591
rect 332 10537 373 10565
rect 332 10531 351 10537
rect 196 10490 204 10524
rect 216 10490 230 10524
rect 244 10490 257 10524
rect 278 10494 291 10528
rect 300 10512 321 10528
rect 336 10521 351 10531
rect 300 10510 312 10512
rect 300 10494 321 10510
rect 332 10503 351 10521
rect 361 10503 375 10537
rect 400 10531 411 10569
rect 562 10532 612 10534
rect 400 10503 409 10531
rect 466 10523 497 10525
rect 565 10523 596 10525
rect 442 10516 500 10523
rect 466 10515 500 10516
rect 565 10515 599 10523
rect 174 10453 181 10477
rect 224 10443 226 10490
rect 300 10481 308 10494
rect 289 10478 305 10480
rect 332 10453 342 10503
rect 400 10483 404 10503
rect 497 10499 500 10515
rect 596 10499 599 10515
rect 466 10498 500 10499
rect 442 10491 500 10498
rect 565 10491 599 10499
rect 612 10482 614 10532
rect 256 10443 328 10451
rect 336 10445 342 10453
rect 400 10445 404 10453
rect 196 10413 204 10443
rect 216 10413 230 10443
rect 196 10409 230 10413
rect 196 10401 226 10409
rect 224 10385 226 10401
rect 332 10373 336 10441
rect 400 10411 408 10445
rect 434 10411 438 10445
rect 454 10429 504 10431
rect 504 10413 506 10429
rect 514 10423 530 10429
rect 532 10423 548 10429
rect 525 10413 548 10422
rect 400 10403 404 10411
rect 498 10403 506 10413
rect 504 10379 506 10403
rect 514 10393 515 10413
rect 525 10388 528 10413
rect 547 10393 548 10413
rect 557 10403 564 10413
rect 514 10379 548 10383
rect 400 10373 442 10374
rect 174 10363 246 10371
rect 400 10366 404 10373
rect 295 10332 300 10366
rect 324 10332 329 10366
rect 367 10332 438 10366
rect 400 10331 404 10332
rect 378 10325 404 10331
rect 442 10325 464 10331
rect 38 10309 80 10325
rect 400 10309 442 10325
rect -25 10295 25 10297
rect 455 10295 505 10297
rect 557 10295 607 10297
rect 16 10287 102 10295
rect 378 10287 464 10295
rect 8 10253 17 10287
rect 18 10285 51 10287
rect 80 10285 100 10287
rect 18 10253 100 10285
rect 380 10285 404 10287
rect 429 10285 438 10287
rect 442 10285 462 10287
rect 16 10245 102 10253
rect 42 10229 76 10231
rect 16 10209 38 10215
rect 42 10206 76 10210
rect 80 10209 102 10215
rect 42 10176 46 10206
rect 72 10176 76 10206
rect 42 10095 46 10129
rect 72 10095 76 10129
rect -25 10058 25 10060
rect 0 10050 14 10051
rect 0 10049 17 10050
rect 25 10049 27 10058
rect 0 10042 38 10049
rect 0 10041 34 10042
rect 0 10025 8 10041
rect 14 10025 34 10041
rect 0 10024 34 10025
rect 0 10017 38 10024
rect 14 10016 17 10017
rect 25 10008 27 10017
rect 42 9988 45 10078
rect 69 10063 80 10095
rect 107 10063 143 10091
rect 107 10057 119 10063
rect 109 10029 119 10057
rect 129 10029 143 10063
rect 42 9937 46 9971
rect 72 9937 76 9971
rect 38 9899 80 9900
rect 42 9858 76 9892
rect 79 9858 113 9892
rect 42 9779 46 9813
rect 72 9779 76 9813
rect -25 9742 25 9744
rect 0 9734 14 9735
rect 0 9733 17 9734
rect 25 9733 27 9742
rect 0 9726 38 9733
rect 0 9725 34 9726
rect 0 9709 8 9725
rect 14 9709 34 9725
rect 0 9708 34 9709
rect 0 9701 38 9708
rect 14 9700 17 9701
rect 25 9692 27 9701
rect 42 9672 45 9762
rect 71 9731 80 9759
rect 69 9693 80 9731
rect 107 9687 119 9721
rect 129 9693 143 9721
rect 129 9687 141 9693
rect 42 9621 46 9655
rect 72 9621 76 9655
rect 42 9574 76 9578
rect 42 9544 46 9574
rect 72 9544 76 9574
rect 16 9535 38 9541
rect 80 9535 102 9541
rect 144 9535 148 10283
rect 332 10215 336 10283
rect 380 10253 462 10285
rect 463 10253 472 10287
rect 480 10253 497 10287
rect 378 10245 464 10253
rect 505 10245 507 10295
rect 514 10253 548 10287
rect 565 10253 582 10287
rect 607 10245 609 10295
rect 404 10229 438 10231
rect 400 10215 442 10216
rect 378 10209 404 10215
rect 442 10209 464 10215
rect 400 10208 404 10209
rect 174 10169 246 10177
rect 295 10174 300 10208
rect 324 10174 329 10208
rect 224 10139 226 10155
rect 196 10131 226 10139
rect 332 10137 336 10205
rect 367 10174 438 10208
rect 400 10167 404 10174
rect 454 10161 504 10163
rect 494 10157 548 10161
rect 494 10152 514 10157
rect 504 10137 506 10152
rect 196 10127 230 10131
rect 196 10097 204 10127
rect 216 10097 230 10127
rect 400 10129 404 10137
rect 174 10063 181 10089
rect 224 10050 226 10097
rect 256 10089 328 10097
rect 332 10095 336 10125
rect 400 10095 408 10129
rect 434 10095 438 10129
rect 498 10127 506 10137
rect 514 10127 515 10147
rect 504 10111 506 10127
rect 525 10118 528 10152
rect 547 10127 548 10147
rect 557 10127 564 10137
rect 514 10111 530 10117
rect 532 10111 548 10117
rect 289 10060 305 10062
rect 196 10016 204 10050
rect 216 10016 230 10050
rect 244 10016 257 10050
rect 300 10046 308 10059
rect 332 10057 342 10095
rect 400 10087 404 10095
rect 336 10047 342 10057
rect 224 9969 226 10016
rect 278 10012 291 10046
rect 300 10030 321 10046
rect 332 10037 342 10047
rect 400 10047 409 10075
rect 562 10058 612 10060
rect 466 10049 497 10051
rect 565 10049 596 10051
rect 300 10028 312 10030
rect 300 10012 321 10028
rect 300 10006 308 10012
rect 289 9996 308 10006
rect 196 9939 204 9969
rect 216 9939 230 9969
rect 196 9935 230 9939
rect 196 9927 226 9935
rect 300 9927 308 9996
rect 332 10003 351 10037
rect 361 10003 375 10037
rect 400 10003 411 10047
rect 442 10042 500 10049
rect 466 10041 500 10042
rect 565 10041 599 10049
rect 497 10025 500 10041
rect 596 10025 599 10041
rect 466 10024 500 10025
rect 442 10017 500 10024
rect 565 10017 599 10025
rect 612 10008 614 10058
rect 332 9979 342 10003
rect 336 9967 342 9979
rect 224 9911 226 9927
rect 332 9899 342 9967
rect 400 9971 404 9979
rect 400 9937 408 9971
rect 434 9937 438 9971
rect 454 9955 504 9957
rect 504 9939 506 9955
rect 514 9949 530 9955
rect 532 9949 548 9955
rect 525 9939 548 9948
rect 400 9929 404 9937
rect 498 9929 506 9939
rect 504 9905 506 9929
rect 514 9919 515 9939
rect 525 9914 528 9939
rect 547 9919 548 9939
rect 557 9929 564 9939
rect 514 9905 548 9909
rect 151 9858 156 9892
rect 174 9889 246 9897
rect 256 9889 328 9897
rect 336 9891 342 9899
rect 400 9894 404 9899
rect 180 9861 185 9889
rect 174 9853 246 9861
rect 256 9853 328 9861
rect 332 9859 336 9889
rect 400 9860 438 9894
rect 224 9823 226 9839
rect 196 9815 226 9823
rect 196 9811 230 9815
rect 196 9781 204 9811
rect 216 9781 230 9811
rect 224 9734 226 9781
rect 300 9754 308 9823
rect 332 9821 342 9859
rect 400 9851 404 9860
rect 454 9845 504 9847
rect 494 9841 548 9845
rect 494 9836 514 9841
rect 504 9821 506 9836
rect 336 9809 342 9821
rect 289 9744 308 9754
rect 300 9738 308 9744
rect 332 9775 342 9809
rect 400 9813 404 9821
rect 400 9779 408 9813
rect 434 9779 438 9813
rect 498 9811 506 9821
rect 514 9811 515 9831
rect 504 9795 506 9811
rect 525 9802 528 9836
rect 547 9811 548 9831
rect 557 9811 564 9821
rect 514 9795 530 9801
rect 532 9795 548 9801
rect 332 9747 373 9775
rect 332 9741 351 9747
rect 196 9700 204 9734
rect 216 9700 230 9734
rect 244 9700 257 9734
rect 278 9704 291 9738
rect 300 9722 321 9738
rect 336 9731 351 9741
rect 300 9720 312 9722
rect 300 9704 321 9720
rect 332 9713 351 9731
rect 361 9713 375 9747
rect 400 9741 411 9779
rect 562 9742 612 9744
rect 400 9713 409 9741
rect 466 9733 497 9735
rect 565 9733 596 9735
rect 442 9726 500 9733
rect 466 9725 500 9726
rect 565 9725 599 9733
rect 174 9663 181 9687
rect 224 9653 226 9700
rect 300 9691 308 9704
rect 289 9688 305 9690
rect 332 9663 342 9713
rect 400 9693 404 9713
rect 497 9709 500 9725
rect 596 9709 599 9725
rect 466 9708 500 9709
rect 442 9701 500 9708
rect 565 9701 599 9709
rect 612 9692 614 9742
rect 256 9653 328 9661
rect 336 9655 342 9663
rect 400 9655 404 9663
rect 196 9623 204 9653
rect 216 9623 230 9653
rect 196 9619 230 9623
rect 196 9611 226 9619
rect 224 9595 226 9611
rect 332 9583 336 9651
rect 400 9621 408 9655
rect 434 9621 438 9655
rect 454 9639 504 9641
rect 504 9623 506 9639
rect 514 9633 530 9639
rect 532 9633 548 9639
rect 525 9623 548 9632
rect 400 9613 404 9621
rect 498 9613 506 9623
rect 504 9589 506 9613
rect 514 9603 515 9623
rect 525 9598 528 9623
rect 547 9603 548 9623
rect 557 9613 564 9623
rect 514 9589 548 9593
rect 400 9583 442 9584
rect 174 9573 246 9581
rect 400 9576 404 9583
rect 295 9542 300 9576
rect 324 9542 329 9576
rect 367 9542 438 9576
rect 400 9541 404 9542
rect 378 9535 404 9541
rect 442 9535 464 9541
rect 38 9519 80 9535
rect 400 9519 442 9535
rect -25 9505 25 9507
rect 455 9505 505 9507
rect 557 9505 607 9507
rect 16 9497 102 9505
rect 378 9497 464 9505
rect 8 9463 17 9497
rect 18 9495 51 9497
rect 80 9495 100 9497
rect 18 9463 100 9495
rect 380 9495 404 9497
rect 429 9495 438 9497
rect 442 9495 462 9497
rect 16 9455 102 9463
rect 42 9439 76 9441
rect 16 9419 38 9425
rect 42 9416 76 9420
rect 80 9419 102 9425
rect 42 9386 46 9416
rect 72 9386 76 9416
rect 42 9305 46 9339
rect 72 9305 76 9339
rect -25 9268 25 9270
rect 0 9260 14 9261
rect 0 9259 17 9260
rect 25 9259 27 9268
rect 0 9252 38 9259
rect 0 9251 34 9252
rect 0 9235 8 9251
rect 14 9235 34 9251
rect 0 9234 34 9235
rect 0 9227 38 9234
rect 14 9226 17 9227
rect 25 9218 27 9227
rect 42 9198 45 9288
rect 69 9273 80 9305
rect 107 9273 143 9301
rect 107 9267 119 9273
rect 109 9239 119 9267
rect 129 9239 143 9273
rect 42 9147 46 9181
rect 72 9147 76 9181
rect 38 9109 80 9110
rect 42 9068 76 9102
rect 79 9068 113 9102
rect 42 8989 46 9023
rect 72 8989 76 9023
rect -25 8952 25 8954
rect 0 8944 14 8945
rect 0 8943 17 8944
rect 25 8943 27 8952
rect 0 8936 38 8943
rect 0 8935 34 8936
rect 0 8919 8 8935
rect 14 8919 34 8935
rect 0 8918 34 8919
rect 0 8911 38 8918
rect 14 8910 17 8911
rect 25 8902 27 8911
rect 42 8882 45 8972
rect 71 8941 80 8969
rect 69 8903 80 8941
rect 107 8897 119 8931
rect 129 8903 143 8931
rect 129 8897 141 8903
rect 42 8831 46 8865
rect 72 8831 76 8865
rect 42 8784 76 8788
rect 42 8754 46 8784
rect 72 8754 76 8784
rect 16 8745 38 8751
rect 80 8745 102 8751
rect 144 8745 148 9493
rect 332 9425 336 9493
rect 380 9463 462 9495
rect 463 9463 472 9497
rect 480 9463 497 9497
rect 378 9455 464 9463
rect 505 9455 507 9505
rect 514 9463 548 9497
rect 565 9463 582 9497
rect 607 9455 609 9505
rect 404 9439 438 9441
rect 400 9425 442 9426
rect 378 9419 404 9425
rect 442 9419 464 9425
rect 400 9418 404 9419
rect 174 9379 246 9387
rect 295 9384 300 9418
rect 324 9384 329 9418
rect 224 9349 226 9365
rect 196 9341 226 9349
rect 332 9347 336 9415
rect 367 9384 438 9418
rect 400 9377 404 9384
rect 454 9371 504 9373
rect 494 9367 548 9371
rect 494 9362 514 9367
rect 504 9347 506 9362
rect 196 9337 230 9341
rect 196 9307 204 9337
rect 216 9307 230 9337
rect 400 9339 404 9347
rect 174 9273 181 9299
rect 224 9260 226 9307
rect 256 9299 328 9307
rect 332 9305 336 9335
rect 400 9305 408 9339
rect 434 9305 438 9339
rect 498 9337 506 9347
rect 514 9337 515 9357
rect 504 9321 506 9337
rect 525 9328 528 9362
rect 547 9337 548 9357
rect 557 9337 564 9347
rect 514 9321 530 9327
rect 532 9321 548 9327
rect 289 9270 305 9272
rect 196 9226 204 9260
rect 216 9226 230 9260
rect 244 9226 257 9260
rect 300 9256 308 9269
rect 332 9267 342 9305
rect 400 9297 404 9305
rect 336 9257 342 9267
rect 224 9179 226 9226
rect 278 9222 291 9256
rect 300 9240 321 9256
rect 332 9247 342 9257
rect 400 9257 409 9285
rect 562 9268 612 9270
rect 466 9259 497 9261
rect 565 9259 596 9261
rect 300 9238 312 9240
rect 300 9222 321 9238
rect 300 9216 308 9222
rect 289 9206 308 9216
rect 196 9149 204 9179
rect 216 9149 230 9179
rect 196 9145 230 9149
rect 196 9137 226 9145
rect 300 9137 308 9206
rect 332 9213 351 9247
rect 361 9213 375 9247
rect 400 9213 411 9257
rect 442 9252 500 9259
rect 466 9251 500 9252
rect 565 9251 599 9259
rect 497 9235 500 9251
rect 596 9235 599 9251
rect 466 9234 500 9235
rect 442 9227 500 9234
rect 565 9227 599 9235
rect 612 9218 614 9268
rect 332 9189 342 9213
rect 336 9177 342 9189
rect 224 9121 226 9137
rect 332 9109 342 9177
rect 400 9181 404 9189
rect 400 9147 408 9181
rect 434 9147 438 9181
rect 454 9165 504 9167
rect 504 9149 506 9165
rect 514 9159 530 9165
rect 532 9159 548 9165
rect 525 9149 548 9158
rect 400 9139 404 9147
rect 498 9139 506 9149
rect 504 9115 506 9139
rect 514 9129 515 9149
rect 525 9124 528 9149
rect 547 9129 548 9149
rect 557 9139 564 9149
rect 514 9115 548 9119
rect 151 9068 156 9102
rect 174 9099 246 9107
rect 256 9099 328 9107
rect 336 9101 342 9109
rect 400 9104 404 9109
rect 180 9071 185 9099
rect 174 9063 246 9071
rect 256 9063 328 9071
rect 332 9069 336 9099
rect 400 9070 438 9104
rect 224 9033 226 9049
rect 196 9025 226 9033
rect 196 9021 230 9025
rect 196 8991 204 9021
rect 216 8991 230 9021
rect 224 8944 226 8991
rect 300 8964 308 9033
rect 332 9031 342 9069
rect 400 9061 404 9070
rect 454 9055 504 9057
rect 494 9051 548 9055
rect 494 9046 514 9051
rect 504 9031 506 9046
rect 336 9019 342 9031
rect 289 8954 308 8964
rect 300 8948 308 8954
rect 332 8985 342 9019
rect 400 9023 404 9031
rect 400 8989 408 9023
rect 434 8989 438 9023
rect 498 9021 506 9031
rect 514 9021 515 9041
rect 504 9005 506 9021
rect 525 9012 528 9046
rect 547 9021 548 9041
rect 557 9021 564 9031
rect 514 9005 530 9011
rect 532 9005 548 9011
rect 332 8957 373 8985
rect 332 8951 351 8957
rect 196 8910 204 8944
rect 216 8910 230 8944
rect 244 8910 257 8944
rect 278 8914 291 8948
rect 300 8932 321 8948
rect 336 8941 351 8951
rect 300 8930 312 8932
rect 300 8914 321 8930
rect 332 8923 351 8941
rect 361 8923 375 8957
rect 400 8951 411 8989
rect 562 8952 612 8954
rect 400 8923 409 8951
rect 466 8943 497 8945
rect 565 8943 596 8945
rect 442 8936 500 8943
rect 466 8935 500 8936
rect 565 8935 599 8943
rect 174 8873 181 8897
rect 224 8863 226 8910
rect 300 8901 308 8914
rect 289 8898 305 8900
rect 332 8873 342 8923
rect 400 8903 404 8923
rect 497 8919 500 8935
rect 596 8919 599 8935
rect 466 8918 500 8919
rect 442 8911 500 8918
rect 565 8911 599 8919
rect 612 8902 614 8952
rect 256 8863 328 8871
rect 336 8865 342 8873
rect 400 8865 404 8873
rect 196 8833 204 8863
rect 216 8833 230 8863
rect 196 8829 230 8833
rect 196 8821 226 8829
rect 224 8805 226 8821
rect 332 8793 336 8861
rect 400 8831 408 8865
rect 434 8831 438 8865
rect 454 8849 504 8851
rect 504 8833 506 8849
rect 514 8843 530 8849
rect 532 8843 548 8849
rect 525 8833 548 8842
rect 400 8823 404 8831
rect 498 8823 506 8833
rect 504 8799 506 8823
rect 514 8813 515 8833
rect 525 8808 528 8833
rect 547 8813 548 8833
rect 557 8823 564 8833
rect 514 8799 548 8803
rect 400 8793 442 8794
rect 174 8783 246 8791
rect 400 8786 404 8793
rect 295 8752 300 8786
rect 324 8752 329 8786
rect 367 8752 438 8786
rect 400 8751 404 8752
rect 378 8745 404 8751
rect 442 8745 464 8751
rect 38 8729 80 8745
rect 400 8729 442 8745
rect -25 8715 25 8717
rect 455 8715 505 8717
rect 557 8715 607 8717
rect 16 8707 102 8715
rect 378 8707 464 8715
rect 8 8673 17 8707
rect 18 8705 51 8707
rect 80 8705 100 8707
rect 18 8673 100 8705
rect 380 8705 404 8707
rect 429 8705 438 8707
rect 442 8705 462 8707
rect 16 8665 102 8673
rect 42 8649 76 8651
rect 16 8629 38 8635
rect 42 8626 76 8630
rect 80 8629 102 8635
rect 42 8596 46 8626
rect 72 8596 76 8626
rect 42 8515 46 8549
rect 72 8515 76 8549
rect -25 8478 25 8480
rect 0 8470 14 8471
rect 0 8469 17 8470
rect 25 8469 27 8478
rect 0 8462 38 8469
rect 0 8461 34 8462
rect 0 8445 8 8461
rect 14 8445 34 8461
rect 0 8444 34 8445
rect 0 8437 38 8444
rect 14 8436 17 8437
rect 25 8428 27 8437
rect 42 8408 45 8498
rect 69 8483 80 8515
rect 107 8483 143 8511
rect 107 8477 119 8483
rect 109 8449 119 8477
rect 129 8449 143 8483
rect 42 8357 46 8391
rect 72 8357 76 8391
rect 38 8319 80 8320
rect 42 8278 76 8312
rect 79 8278 113 8312
rect 42 8199 46 8233
rect 72 8199 76 8233
rect -25 8162 25 8164
rect 0 8154 14 8155
rect 0 8153 17 8154
rect 25 8153 27 8162
rect 0 8146 38 8153
rect 0 8145 34 8146
rect 0 8129 8 8145
rect 14 8129 34 8145
rect 0 8128 34 8129
rect 0 8121 38 8128
rect 14 8120 17 8121
rect 25 8112 27 8121
rect 42 8092 45 8182
rect 71 8151 80 8179
rect 69 8113 80 8151
rect 107 8107 119 8141
rect 129 8113 143 8141
rect 129 8107 141 8113
rect 42 8041 46 8075
rect 72 8041 76 8075
rect 42 7994 76 7998
rect 42 7964 46 7994
rect 72 7964 76 7994
rect 16 7955 38 7961
rect 80 7955 102 7961
rect 144 7955 148 8703
rect 332 8635 336 8703
rect 380 8673 462 8705
rect 463 8673 472 8707
rect 480 8673 497 8707
rect 378 8665 464 8673
rect 505 8665 507 8715
rect 514 8673 548 8707
rect 565 8673 582 8707
rect 607 8665 609 8715
rect 404 8649 438 8651
rect 400 8635 442 8636
rect 378 8629 404 8635
rect 442 8629 464 8635
rect 400 8628 404 8629
rect 174 8589 246 8597
rect 295 8594 300 8628
rect 324 8594 329 8628
rect 224 8559 226 8575
rect 196 8551 226 8559
rect 332 8557 336 8625
rect 367 8594 438 8628
rect 400 8587 404 8594
rect 454 8581 504 8583
rect 494 8577 548 8581
rect 494 8572 514 8577
rect 504 8557 506 8572
rect 196 8547 230 8551
rect 196 8517 204 8547
rect 216 8517 230 8547
rect 400 8549 404 8557
rect 174 8483 181 8509
rect 224 8470 226 8517
rect 256 8509 328 8517
rect 332 8515 336 8545
rect 400 8515 408 8549
rect 434 8515 438 8549
rect 498 8547 506 8557
rect 514 8547 515 8567
rect 504 8531 506 8547
rect 525 8538 528 8572
rect 547 8547 548 8567
rect 557 8547 564 8557
rect 514 8531 530 8537
rect 532 8531 548 8537
rect 289 8480 305 8482
rect 196 8436 204 8470
rect 216 8436 230 8470
rect 244 8436 257 8470
rect 300 8466 308 8479
rect 332 8477 342 8515
rect 400 8507 404 8515
rect 336 8467 342 8477
rect 224 8389 226 8436
rect 278 8432 291 8466
rect 300 8450 321 8466
rect 332 8457 342 8467
rect 400 8467 409 8495
rect 562 8478 612 8480
rect 466 8469 497 8471
rect 565 8469 596 8471
rect 300 8448 312 8450
rect 300 8432 321 8448
rect 300 8426 308 8432
rect 289 8416 308 8426
rect 196 8359 204 8389
rect 216 8359 230 8389
rect 196 8355 230 8359
rect 196 8347 226 8355
rect 300 8347 308 8416
rect 332 8423 351 8457
rect 361 8423 375 8457
rect 400 8423 411 8467
rect 442 8462 500 8469
rect 466 8461 500 8462
rect 565 8461 599 8469
rect 497 8445 500 8461
rect 596 8445 599 8461
rect 466 8444 500 8445
rect 442 8437 500 8444
rect 565 8437 599 8445
rect 612 8428 614 8478
rect 332 8399 342 8423
rect 336 8387 342 8399
rect 224 8331 226 8347
rect 332 8319 342 8387
rect 400 8391 404 8399
rect 400 8357 408 8391
rect 434 8357 438 8391
rect 454 8375 504 8377
rect 504 8359 506 8375
rect 514 8369 530 8375
rect 532 8369 548 8375
rect 525 8359 548 8368
rect 400 8349 404 8357
rect 498 8349 506 8359
rect 504 8325 506 8349
rect 514 8339 515 8359
rect 525 8334 528 8359
rect 547 8339 548 8359
rect 557 8349 564 8359
rect 514 8325 548 8329
rect 151 8278 156 8312
rect 174 8309 246 8317
rect 256 8309 328 8317
rect 336 8311 342 8319
rect 400 8314 404 8319
rect 180 8281 185 8309
rect 174 8273 246 8281
rect 256 8273 328 8281
rect 332 8279 336 8309
rect 400 8280 438 8314
rect 224 8243 226 8259
rect 196 8235 226 8243
rect 196 8231 230 8235
rect 196 8201 204 8231
rect 216 8201 230 8231
rect 224 8154 226 8201
rect 300 8174 308 8243
rect 332 8241 342 8279
rect 400 8271 404 8280
rect 454 8265 504 8267
rect 494 8261 548 8265
rect 494 8256 514 8261
rect 504 8241 506 8256
rect 336 8229 342 8241
rect 289 8164 308 8174
rect 300 8158 308 8164
rect 332 8195 342 8229
rect 400 8233 404 8241
rect 400 8199 408 8233
rect 434 8199 438 8233
rect 498 8231 506 8241
rect 514 8231 515 8251
rect 504 8215 506 8231
rect 525 8222 528 8256
rect 547 8231 548 8251
rect 557 8231 564 8241
rect 514 8215 530 8221
rect 532 8215 548 8221
rect 332 8167 373 8195
rect 332 8161 351 8167
rect 196 8120 204 8154
rect 216 8120 230 8154
rect 244 8120 257 8154
rect 278 8124 291 8158
rect 300 8142 321 8158
rect 336 8151 351 8161
rect 300 8140 312 8142
rect 300 8124 321 8140
rect 332 8133 351 8151
rect 361 8133 375 8167
rect 400 8161 411 8199
rect 562 8162 612 8164
rect 400 8133 409 8161
rect 466 8153 497 8155
rect 565 8153 596 8155
rect 442 8146 500 8153
rect 466 8145 500 8146
rect 565 8145 599 8153
rect 174 8083 181 8107
rect 224 8073 226 8120
rect 300 8111 308 8124
rect 289 8108 305 8110
rect 332 8083 342 8133
rect 400 8113 404 8133
rect 497 8129 500 8145
rect 596 8129 599 8145
rect 466 8128 500 8129
rect 442 8121 500 8128
rect 565 8121 599 8129
rect 612 8112 614 8162
rect 256 8073 328 8081
rect 336 8075 342 8083
rect 400 8075 404 8083
rect 196 8043 204 8073
rect 216 8043 230 8073
rect 196 8039 230 8043
rect 196 8031 226 8039
rect 224 8015 226 8031
rect 332 8003 336 8071
rect 400 8041 408 8075
rect 434 8041 438 8075
rect 454 8059 504 8061
rect 504 8043 506 8059
rect 514 8053 530 8059
rect 532 8053 548 8059
rect 525 8043 548 8052
rect 400 8033 404 8041
rect 498 8033 506 8043
rect 504 8009 506 8033
rect 514 8023 515 8043
rect 525 8018 528 8043
rect 547 8023 548 8043
rect 557 8033 564 8043
rect 514 8009 548 8013
rect 400 8003 442 8004
rect 174 7993 246 8001
rect 400 7996 404 8003
rect 295 7962 300 7996
rect 324 7962 329 7996
rect 367 7962 438 7996
rect 400 7961 404 7962
rect 378 7955 404 7961
rect 442 7955 464 7961
rect 38 7939 80 7955
rect 400 7939 442 7955
rect -25 7925 25 7927
rect 455 7925 505 7927
rect 557 7925 607 7927
rect 16 7917 102 7925
rect 378 7917 464 7925
rect 8 7883 17 7917
rect 18 7915 51 7917
rect 80 7915 100 7917
rect 18 7883 100 7915
rect 380 7915 404 7917
rect 429 7915 438 7917
rect 442 7915 462 7917
rect 16 7875 102 7883
rect 42 7859 76 7861
rect 16 7839 38 7845
rect 42 7836 76 7840
rect 80 7839 102 7845
rect 42 7806 46 7836
rect 72 7806 76 7836
rect 42 7725 46 7759
rect 72 7725 76 7759
rect -25 7688 25 7690
rect 0 7680 14 7681
rect 0 7679 17 7680
rect 25 7679 27 7688
rect 0 7672 38 7679
rect 0 7671 34 7672
rect 0 7655 8 7671
rect 14 7655 34 7671
rect 0 7654 34 7655
rect 0 7647 38 7654
rect 14 7646 17 7647
rect 25 7638 27 7647
rect 42 7618 45 7708
rect 69 7693 80 7725
rect 107 7693 143 7721
rect 107 7687 119 7693
rect 109 7659 119 7687
rect 129 7659 143 7693
rect 42 7567 46 7601
rect 72 7567 76 7601
rect 38 7529 80 7530
rect 42 7488 76 7522
rect 79 7488 113 7522
rect 42 7409 46 7443
rect 72 7409 76 7443
rect -25 7372 25 7374
rect 0 7364 14 7365
rect 0 7363 17 7364
rect 25 7363 27 7372
rect 0 7356 38 7363
rect 0 7355 34 7356
rect 0 7339 8 7355
rect 14 7339 34 7355
rect 0 7338 34 7339
rect 0 7331 38 7338
rect 14 7330 17 7331
rect 25 7322 27 7331
rect 42 7302 45 7392
rect 71 7361 80 7389
rect 69 7323 80 7361
rect 107 7317 119 7351
rect 129 7323 143 7351
rect 129 7317 141 7323
rect 42 7251 46 7285
rect 72 7251 76 7285
rect 42 7204 76 7208
rect 42 7174 46 7204
rect 72 7174 76 7204
rect 16 7165 38 7171
rect 80 7165 102 7171
rect 144 7165 148 7913
rect 332 7845 336 7913
rect 380 7883 462 7915
rect 463 7883 472 7917
rect 480 7883 497 7917
rect 378 7875 464 7883
rect 505 7875 507 7925
rect 514 7883 548 7917
rect 565 7883 582 7917
rect 607 7875 609 7925
rect 404 7859 438 7861
rect 400 7845 442 7846
rect 378 7839 404 7845
rect 442 7839 464 7845
rect 400 7838 404 7839
rect 174 7799 246 7807
rect 295 7804 300 7838
rect 324 7804 329 7838
rect 224 7769 226 7785
rect 196 7761 226 7769
rect 332 7767 336 7835
rect 367 7804 438 7838
rect 400 7797 404 7804
rect 454 7791 504 7793
rect 494 7787 548 7791
rect 494 7782 514 7787
rect 504 7767 506 7782
rect 196 7757 230 7761
rect 196 7727 204 7757
rect 216 7727 230 7757
rect 400 7759 404 7767
rect 174 7693 181 7719
rect 224 7680 226 7727
rect 256 7719 328 7727
rect 332 7725 336 7755
rect 400 7725 408 7759
rect 434 7725 438 7759
rect 498 7757 506 7767
rect 514 7757 515 7777
rect 504 7741 506 7757
rect 525 7748 528 7782
rect 547 7757 548 7777
rect 557 7757 564 7767
rect 514 7741 530 7747
rect 532 7741 548 7747
rect 289 7690 305 7692
rect 196 7646 204 7680
rect 216 7646 230 7680
rect 244 7646 257 7680
rect 300 7676 308 7689
rect 332 7687 342 7725
rect 400 7717 404 7725
rect 336 7677 342 7687
rect 224 7599 226 7646
rect 278 7642 291 7676
rect 300 7660 321 7676
rect 332 7667 342 7677
rect 400 7677 409 7705
rect 562 7688 612 7690
rect 466 7679 497 7681
rect 565 7679 596 7681
rect 300 7658 312 7660
rect 300 7642 321 7658
rect 300 7636 308 7642
rect 289 7626 308 7636
rect 196 7569 204 7599
rect 216 7569 230 7599
rect 196 7565 230 7569
rect 196 7557 226 7565
rect 300 7557 308 7626
rect 332 7633 351 7667
rect 361 7633 375 7667
rect 400 7633 411 7677
rect 442 7672 500 7679
rect 466 7671 500 7672
rect 565 7671 599 7679
rect 497 7655 500 7671
rect 596 7655 599 7671
rect 466 7654 500 7655
rect 442 7647 500 7654
rect 565 7647 599 7655
rect 612 7638 614 7688
rect 332 7609 342 7633
rect 336 7597 342 7609
rect 224 7541 226 7557
rect 332 7529 342 7597
rect 400 7601 404 7609
rect 400 7567 408 7601
rect 434 7567 438 7601
rect 454 7585 504 7587
rect 504 7569 506 7585
rect 514 7579 530 7585
rect 532 7579 548 7585
rect 525 7569 548 7578
rect 400 7559 404 7567
rect 498 7559 506 7569
rect 504 7535 506 7559
rect 514 7549 515 7569
rect 525 7544 528 7569
rect 547 7549 548 7569
rect 557 7559 564 7569
rect 514 7535 548 7539
rect 151 7488 156 7522
rect 174 7519 246 7527
rect 256 7519 328 7527
rect 336 7521 342 7529
rect 400 7524 404 7529
rect 180 7491 185 7519
rect 174 7483 246 7491
rect 256 7483 328 7491
rect 332 7489 336 7519
rect 400 7490 438 7524
rect 224 7453 226 7469
rect 196 7445 226 7453
rect 196 7441 230 7445
rect 196 7411 204 7441
rect 216 7411 230 7441
rect 224 7364 226 7411
rect 300 7384 308 7453
rect 332 7451 342 7489
rect 400 7481 404 7490
rect 454 7475 504 7477
rect 494 7471 548 7475
rect 494 7466 514 7471
rect 504 7451 506 7466
rect 336 7439 342 7451
rect 289 7374 308 7384
rect 300 7368 308 7374
rect 332 7405 342 7439
rect 400 7443 404 7451
rect 400 7409 408 7443
rect 434 7409 438 7443
rect 498 7441 506 7451
rect 514 7441 515 7461
rect 504 7425 506 7441
rect 525 7432 528 7466
rect 547 7441 548 7461
rect 557 7441 564 7451
rect 514 7425 530 7431
rect 532 7425 548 7431
rect 332 7377 373 7405
rect 332 7371 351 7377
rect 196 7330 204 7364
rect 216 7330 230 7364
rect 244 7330 257 7364
rect 278 7334 291 7368
rect 300 7352 321 7368
rect 336 7361 351 7371
rect 300 7350 312 7352
rect 300 7334 321 7350
rect 332 7343 351 7361
rect 361 7343 375 7377
rect 400 7371 411 7409
rect 562 7372 612 7374
rect 400 7343 409 7371
rect 466 7363 497 7365
rect 565 7363 596 7365
rect 442 7356 500 7363
rect 466 7355 500 7356
rect 565 7355 599 7363
rect 174 7293 181 7317
rect 224 7283 226 7330
rect 300 7321 308 7334
rect 289 7318 305 7320
rect 332 7293 342 7343
rect 400 7323 404 7343
rect 497 7339 500 7355
rect 596 7339 599 7355
rect 466 7338 500 7339
rect 442 7331 500 7338
rect 565 7331 599 7339
rect 612 7322 614 7372
rect 256 7283 328 7291
rect 336 7285 342 7293
rect 400 7285 404 7293
rect 196 7253 204 7283
rect 216 7253 230 7283
rect 196 7249 230 7253
rect 196 7241 226 7249
rect 224 7225 226 7241
rect 332 7213 336 7281
rect 400 7251 408 7285
rect 434 7251 438 7285
rect 454 7269 504 7271
rect 504 7253 506 7269
rect 514 7263 530 7269
rect 532 7263 548 7269
rect 525 7253 548 7262
rect 400 7243 404 7251
rect 498 7243 506 7253
rect 504 7219 506 7243
rect 514 7233 515 7253
rect 525 7228 528 7253
rect 547 7233 548 7253
rect 557 7243 564 7253
rect 514 7219 548 7223
rect 400 7213 442 7214
rect 174 7203 246 7211
rect 400 7206 404 7213
rect 295 7172 300 7206
rect 324 7172 329 7206
rect 367 7172 438 7206
rect 400 7171 404 7172
rect 378 7165 404 7171
rect 442 7165 464 7171
rect 38 7149 80 7165
rect 400 7149 442 7165
rect -25 7135 25 7137
rect 455 7135 505 7137
rect 557 7135 607 7137
rect 16 7127 102 7135
rect 378 7127 464 7135
rect 8 7093 17 7127
rect 18 7125 51 7127
rect 80 7125 100 7127
rect 18 7093 100 7125
rect 380 7125 404 7127
rect 429 7125 438 7127
rect 442 7125 462 7127
rect 16 7085 102 7093
rect 42 7069 76 7071
rect 16 7049 38 7055
rect 42 7046 76 7050
rect 80 7049 102 7055
rect 42 7016 46 7046
rect 72 7016 76 7046
rect 42 6935 46 6969
rect 72 6935 76 6969
rect -25 6898 25 6900
rect 0 6890 14 6891
rect 0 6889 17 6890
rect 25 6889 27 6898
rect 0 6882 38 6889
rect 0 6881 34 6882
rect 0 6865 8 6881
rect 14 6865 34 6881
rect 0 6864 34 6865
rect 0 6857 38 6864
rect 14 6856 17 6857
rect 25 6848 27 6857
rect 42 6828 45 6918
rect 69 6903 80 6935
rect 107 6903 143 6931
rect 107 6897 119 6903
rect 109 6869 119 6897
rect 129 6869 143 6903
rect 42 6777 46 6811
rect 72 6777 76 6811
rect 38 6739 80 6740
rect 42 6698 76 6732
rect 79 6698 113 6732
rect 42 6619 46 6653
rect 72 6619 76 6653
rect -25 6582 25 6584
rect 0 6574 14 6575
rect 0 6573 17 6574
rect 25 6573 27 6582
rect 0 6566 38 6573
rect 0 6565 34 6566
rect 0 6549 8 6565
rect 14 6549 34 6565
rect 0 6548 34 6549
rect 0 6541 38 6548
rect 14 6540 17 6541
rect 25 6532 27 6541
rect 42 6512 45 6602
rect 71 6571 80 6599
rect 69 6533 80 6571
rect 107 6527 119 6561
rect 129 6533 143 6561
rect 129 6527 141 6533
rect 42 6461 46 6495
rect 72 6461 76 6495
rect 42 6414 76 6418
rect 42 6384 46 6414
rect 72 6384 76 6414
rect 16 6375 38 6381
rect 80 6375 102 6381
rect 144 6375 148 7123
rect 332 7055 336 7123
rect 380 7093 462 7125
rect 463 7093 472 7127
rect 480 7093 497 7127
rect 378 7085 464 7093
rect 505 7085 507 7135
rect 514 7093 548 7127
rect 565 7093 582 7127
rect 607 7085 609 7135
rect 404 7069 438 7071
rect 400 7055 442 7056
rect 378 7049 404 7055
rect 442 7049 464 7055
rect 400 7048 404 7049
rect 174 7009 246 7017
rect 295 7014 300 7048
rect 324 7014 329 7048
rect 224 6979 226 6995
rect 196 6971 226 6979
rect 332 6977 336 7045
rect 367 7014 438 7048
rect 400 7007 404 7014
rect 454 7001 504 7003
rect 494 6997 548 7001
rect 494 6992 514 6997
rect 504 6977 506 6992
rect 196 6967 230 6971
rect 196 6937 204 6967
rect 216 6937 230 6967
rect 400 6969 404 6977
rect 174 6903 181 6929
rect 224 6890 226 6937
rect 256 6929 328 6937
rect 332 6935 336 6965
rect 400 6935 408 6969
rect 434 6935 438 6969
rect 498 6967 506 6977
rect 514 6967 515 6987
rect 504 6951 506 6967
rect 525 6958 528 6992
rect 547 6967 548 6987
rect 557 6967 564 6977
rect 514 6951 530 6957
rect 532 6951 548 6957
rect 289 6900 305 6902
rect 196 6856 204 6890
rect 216 6856 230 6890
rect 244 6856 257 6890
rect 300 6886 308 6899
rect 332 6897 342 6935
rect 400 6927 404 6935
rect 336 6887 342 6897
rect 224 6809 226 6856
rect 278 6852 291 6886
rect 300 6870 321 6886
rect 332 6877 342 6887
rect 400 6887 409 6915
rect 562 6898 612 6900
rect 466 6889 497 6891
rect 565 6889 596 6891
rect 300 6868 312 6870
rect 300 6852 321 6868
rect 300 6846 308 6852
rect 289 6836 308 6846
rect 196 6779 204 6809
rect 216 6779 230 6809
rect 196 6775 230 6779
rect 196 6767 226 6775
rect 300 6767 308 6836
rect 332 6843 351 6877
rect 361 6843 375 6877
rect 400 6843 411 6887
rect 442 6882 500 6889
rect 466 6881 500 6882
rect 565 6881 599 6889
rect 497 6865 500 6881
rect 596 6865 599 6881
rect 466 6864 500 6865
rect 442 6857 500 6864
rect 565 6857 599 6865
rect 612 6848 614 6898
rect 332 6819 342 6843
rect 336 6807 342 6819
rect 224 6751 226 6767
rect 332 6739 342 6807
rect 400 6811 404 6819
rect 400 6777 408 6811
rect 434 6777 438 6811
rect 454 6795 504 6797
rect 504 6779 506 6795
rect 514 6789 530 6795
rect 532 6789 548 6795
rect 525 6779 548 6788
rect 400 6769 404 6777
rect 498 6769 506 6779
rect 504 6745 506 6769
rect 514 6759 515 6779
rect 525 6754 528 6779
rect 547 6759 548 6779
rect 557 6769 564 6779
rect 514 6745 548 6749
rect 151 6698 156 6732
rect 174 6729 246 6737
rect 256 6729 328 6737
rect 336 6731 342 6739
rect 400 6734 404 6739
rect 180 6701 185 6729
rect 174 6693 246 6701
rect 256 6693 328 6701
rect 332 6699 336 6729
rect 400 6700 438 6734
rect 224 6663 226 6679
rect 196 6655 226 6663
rect 196 6651 230 6655
rect 196 6621 204 6651
rect 216 6621 230 6651
rect 224 6574 226 6621
rect 300 6594 308 6663
rect 332 6661 342 6699
rect 400 6691 404 6700
rect 454 6685 504 6687
rect 494 6681 548 6685
rect 494 6676 514 6681
rect 504 6661 506 6676
rect 336 6649 342 6661
rect 289 6584 308 6594
rect 300 6578 308 6584
rect 332 6615 342 6649
rect 400 6653 404 6661
rect 400 6619 408 6653
rect 434 6619 438 6653
rect 498 6651 506 6661
rect 514 6651 515 6671
rect 504 6635 506 6651
rect 525 6642 528 6676
rect 547 6651 548 6671
rect 557 6651 564 6661
rect 514 6635 530 6641
rect 532 6635 548 6641
rect 332 6587 373 6615
rect 332 6581 351 6587
rect 196 6540 204 6574
rect 216 6540 230 6574
rect 244 6540 257 6574
rect 278 6544 291 6578
rect 300 6562 321 6578
rect 336 6571 351 6581
rect 300 6560 312 6562
rect 300 6544 321 6560
rect 332 6553 351 6571
rect 361 6553 375 6587
rect 400 6581 411 6619
rect 562 6582 612 6584
rect 400 6553 409 6581
rect 466 6573 497 6575
rect 565 6573 596 6575
rect 442 6566 500 6573
rect 466 6565 500 6566
rect 565 6565 599 6573
rect 174 6503 181 6527
rect 224 6493 226 6540
rect 300 6531 308 6544
rect 289 6528 305 6530
rect 332 6503 342 6553
rect 400 6533 404 6553
rect 497 6549 500 6565
rect 596 6549 599 6565
rect 466 6548 500 6549
rect 442 6541 500 6548
rect 565 6541 599 6549
rect 612 6532 614 6582
rect 256 6493 328 6501
rect 336 6495 342 6503
rect 400 6495 404 6503
rect 196 6463 204 6493
rect 216 6463 230 6493
rect 196 6459 230 6463
rect 196 6451 226 6459
rect 224 6435 226 6451
rect 332 6423 336 6491
rect 400 6461 408 6495
rect 434 6461 438 6495
rect 454 6479 504 6481
rect 504 6463 506 6479
rect 514 6473 530 6479
rect 532 6473 548 6479
rect 525 6463 548 6472
rect 400 6453 404 6461
rect 498 6453 506 6463
rect 504 6429 506 6453
rect 514 6443 515 6463
rect 525 6438 528 6463
rect 547 6443 548 6463
rect 557 6453 564 6463
rect 514 6429 548 6433
rect 400 6423 442 6424
rect 174 6413 246 6421
rect 400 6416 404 6423
rect 295 6382 300 6416
rect 324 6382 329 6416
rect 367 6382 438 6416
rect 400 6381 404 6382
rect 378 6375 404 6381
rect 442 6375 464 6381
rect 38 6359 80 6375
rect 400 6359 442 6375
rect -25 6345 25 6347
rect 455 6345 505 6347
rect 557 6345 607 6347
rect 16 6337 102 6345
rect 378 6337 464 6345
rect 8 6303 17 6337
rect 18 6335 51 6337
rect 80 6335 100 6337
rect 18 6303 100 6335
rect 380 6335 404 6337
rect 429 6335 438 6337
rect 442 6335 462 6337
rect 16 6295 102 6303
rect 42 6279 76 6281
rect 16 6259 38 6265
rect 42 6256 76 6260
rect 80 6259 102 6265
rect 42 6226 46 6256
rect 72 6226 76 6256
rect 42 6145 46 6179
rect 72 6145 76 6179
rect -25 6108 25 6110
rect 0 6100 14 6101
rect 0 6099 17 6100
rect 25 6099 27 6108
rect 0 6092 38 6099
rect 0 6091 34 6092
rect 0 6075 8 6091
rect 14 6075 34 6091
rect 0 6074 34 6075
rect 0 6067 38 6074
rect 14 6066 17 6067
rect 25 6058 27 6067
rect 42 6038 45 6128
rect 69 6113 80 6145
rect 107 6113 143 6141
rect 107 6107 119 6113
rect 109 6079 119 6107
rect 129 6079 143 6113
rect 42 5987 46 6021
rect 72 5987 76 6021
rect 38 5949 80 5950
rect 42 5908 76 5942
rect 79 5908 113 5942
rect 42 5829 46 5863
rect 72 5829 76 5863
rect -25 5792 25 5794
rect 0 5784 14 5785
rect 0 5783 17 5784
rect 25 5783 27 5792
rect 0 5776 38 5783
rect 0 5775 34 5776
rect 0 5759 8 5775
rect 14 5759 34 5775
rect 0 5758 34 5759
rect 0 5751 38 5758
rect 14 5750 17 5751
rect 25 5742 27 5751
rect 42 5722 45 5812
rect 71 5781 80 5809
rect 69 5743 80 5781
rect 107 5737 119 5771
rect 129 5743 143 5771
rect 129 5737 141 5743
rect 42 5671 46 5705
rect 72 5671 76 5705
rect 42 5624 76 5628
rect 42 5594 46 5624
rect 72 5594 76 5624
rect 16 5585 38 5591
rect 80 5585 102 5591
rect 144 5585 148 6333
rect 332 6265 336 6333
rect 380 6303 462 6335
rect 463 6303 472 6337
rect 480 6303 497 6337
rect 378 6295 464 6303
rect 505 6295 507 6345
rect 514 6303 548 6337
rect 565 6303 582 6337
rect 607 6295 609 6345
rect 404 6279 438 6281
rect 400 6265 442 6266
rect 378 6259 404 6265
rect 442 6259 464 6265
rect 400 6258 404 6259
rect 174 6219 246 6227
rect 295 6224 300 6258
rect 324 6224 329 6258
rect 224 6189 226 6205
rect 196 6181 226 6189
rect 332 6187 336 6255
rect 367 6224 438 6258
rect 400 6217 404 6224
rect 454 6211 504 6213
rect 494 6207 548 6211
rect 494 6202 514 6207
rect 504 6187 506 6202
rect 196 6177 230 6181
rect 196 6147 204 6177
rect 216 6147 230 6177
rect 400 6179 404 6187
rect 174 6113 181 6139
rect 224 6100 226 6147
rect 256 6139 328 6147
rect 332 6145 336 6175
rect 400 6145 408 6179
rect 434 6145 438 6179
rect 498 6177 506 6187
rect 514 6177 515 6197
rect 504 6161 506 6177
rect 525 6168 528 6202
rect 547 6177 548 6197
rect 557 6177 564 6187
rect 514 6161 530 6167
rect 532 6161 548 6167
rect 289 6110 305 6112
rect 196 6066 204 6100
rect 216 6066 230 6100
rect 244 6066 257 6100
rect 300 6096 308 6109
rect 332 6107 342 6145
rect 400 6137 404 6145
rect 336 6097 342 6107
rect 224 6019 226 6066
rect 278 6062 291 6096
rect 300 6080 321 6096
rect 332 6087 342 6097
rect 400 6097 409 6125
rect 562 6108 612 6110
rect 466 6099 497 6101
rect 565 6099 596 6101
rect 300 6078 312 6080
rect 300 6062 321 6078
rect 300 6056 308 6062
rect 289 6046 308 6056
rect 196 5989 204 6019
rect 216 5989 230 6019
rect 196 5985 230 5989
rect 196 5977 226 5985
rect 300 5977 308 6046
rect 332 6053 351 6087
rect 361 6053 375 6087
rect 400 6053 411 6097
rect 442 6092 500 6099
rect 466 6091 500 6092
rect 565 6091 599 6099
rect 497 6075 500 6091
rect 596 6075 599 6091
rect 466 6074 500 6075
rect 442 6067 500 6074
rect 565 6067 599 6075
rect 612 6058 614 6108
rect 332 6029 342 6053
rect 336 6017 342 6029
rect 224 5961 226 5977
rect 332 5949 342 6017
rect 400 6021 404 6029
rect 400 5987 408 6021
rect 434 5987 438 6021
rect 454 6005 504 6007
rect 504 5989 506 6005
rect 514 5999 530 6005
rect 532 5999 548 6005
rect 525 5989 548 5998
rect 400 5979 404 5987
rect 498 5979 506 5989
rect 504 5955 506 5979
rect 514 5969 515 5989
rect 525 5964 528 5989
rect 547 5969 548 5989
rect 557 5979 564 5989
rect 514 5955 548 5959
rect 151 5908 156 5942
rect 174 5939 246 5947
rect 256 5939 328 5947
rect 336 5941 342 5949
rect 400 5944 404 5949
rect 180 5911 185 5939
rect 174 5903 246 5911
rect 256 5903 328 5911
rect 332 5909 336 5939
rect 400 5910 438 5944
rect 224 5873 226 5889
rect 196 5865 226 5873
rect 196 5861 230 5865
rect 196 5831 204 5861
rect 216 5831 230 5861
rect 224 5784 226 5831
rect 300 5804 308 5873
rect 332 5871 342 5909
rect 400 5901 404 5910
rect 454 5895 504 5897
rect 494 5891 548 5895
rect 494 5886 514 5891
rect 504 5871 506 5886
rect 336 5859 342 5871
rect 289 5794 308 5804
rect 300 5788 308 5794
rect 332 5825 342 5859
rect 400 5863 404 5871
rect 400 5829 408 5863
rect 434 5829 438 5863
rect 498 5861 506 5871
rect 514 5861 515 5881
rect 504 5845 506 5861
rect 525 5852 528 5886
rect 547 5861 548 5881
rect 557 5861 564 5871
rect 514 5845 530 5851
rect 532 5845 548 5851
rect 332 5797 373 5825
rect 332 5791 351 5797
rect 196 5750 204 5784
rect 216 5750 230 5784
rect 244 5750 257 5784
rect 278 5754 291 5788
rect 300 5772 321 5788
rect 336 5781 351 5791
rect 300 5770 312 5772
rect 300 5754 321 5770
rect 332 5763 351 5781
rect 361 5763 375 5797
rect 400 5791 411 5829
rect 562 5792 612 5794
rect 400 5763 409 5791
rect 466 5783 497 5785
rect 565 5783 596 5785
rect 442 5776 500 5783
rect 466 5775 500 5776
rect 565 5775 599 5783
rect 174 5713 181 5737
rect 224 5703 226 5750
rect 300 5741 308 5754
rect 289 5738 305 5740
rect 332 5713 342 5763
rect 400 5743 404 5763
rect 497 5759 500 5775
rect 596 5759 599 5775
rect 466 5758 500 5759
rect 442 5751 500 5758
rect 565 5751 599 5759
rect 612 5742 614 5792
rect 256 5703 328 5711
rect 336 5705 342 5713
rect 400 5705 404 5713
rect 196 5673 204 5703
rect 216 5673 230 5703
rect 196 5669 230 5673
rect 196 5661 226 5669
rect 224 5645 226 5661
rect 332 5633 336 5701
rect 400 5671 408 5705
rect 434 5671 438 5705
rect 454 5689 504 5691
rect 504 5673 506 5689
rect 514 5683 530 5689
rect 532 5683 548 5689
rect 525 5673 548 5682
rect 400 5663 404 5671
rect 498 5663 506 5673
rect 504 5639 506 5663
rect 514 5653 515 5673
rect 525 5648 528 5673
rect 547 5653 548 5673
rect 557 5663 564 5673
rect 514 5639 548 5643
rect 400 5633 442 5634
rect 174 5623 246 5631
rect 400 5626 404 5633
rect 295 5592 300 5626
rect 324 5592 329 5626
rect 367 5592 438 5626
rect 400 5591 404 5592
rect 378 5585 404 5591
rect 442 5585 464 5591
rect 38 5569 80 5585
rect 400 5569 442 5585
rect -25 5555 25 5557
rect 455 5555 505 5557
rect 557 5555 607 5557
rect 16 5547 102 5555
rect 378 5547 464 5555
rect 8 5513 17 5547
rect 18 5545 51 5547
rect 80 5545 100 5547
rect 18 5513 100 5545
rect 380 5545 404 5547
rect 429 5545 438 5547
rect 442 5545 462 5547
rect 16 5505 102 5513
rect 42 5489 76 5491
rect 16 5469 38 5475
rect 42 5466 76 5470
rect 80 5469 102 5475
rect 42 5436 46 5466
rect 72 5436 76 5466
rect 42 5355 46 5389
rect 72 5355 76 5389
rect -25 5318 25 5320
rect 0 5310 14 5311
rect 0 5309 17 5310
rect 25 5309 27 5318
rect 0 5302 38 5309
rect 0 5301 34 5302
rect 0 5285 8 5301
rect 14 5285 34 5301
rect 0 5284 34 5285
rect 0 5277 38 5284
rect 14 5276 17 5277
rect 25 5268 27 5277
rect 42 5248 45 5338
rect 69 5323 80 5355
rect 107 5323 143 5351
rect 107 5317 119 5323
rect 109 5289 119 5317
rect 129 5289 143 5323
rect 42 5197 46 5231
rect 72 5197 76 5231
rect 38 5159 80 5160
rect 42 5118 76 5152
rect 79 5118 113 5152
rect 42 5039 46 5073
rect 72 5039 76 5073
rect -25 5002 25 5004
rect 0 4994 14 4995
rect 0 4993 17 4994
rect 25 4993 27 5002
rect 0 4986 38 4993
rect 0 4985 34 4986
rect 0 4969 8 4985
rect 14 4969 34 4985
rect 0 4968 34 4969
rect 0 4961 38 4968
rect 14 4960 17 4961
rect 25 4952 27 4961
rect 42 4932 45 5022
rect 71 4991 80 5019
rect 69 4953 80 4991
rect 107 4947 119 4981
rect 129 4953 143 4981
rect 129 4947 141 4953
rect 42 4881 46 4915
rect 72 4881 76 4915
rect 42 4834 76 4838
rect 42 4804 46 4834
rect 72 4804 76 4834
rect 16 4795 38 4801
rect 80 4795 102 4801
rect 144 4795 148 5543
rect 332 5475 336 5543
rect 380 5513 462 5545
rect 463 5513 472 5547
rect 480 5513 497 5547
rect 378 5505 464 5513
rect 505 5505 507 5555
rect 514 5513 548 5547
rect 565 5513 582 5547
rect 607 5505 609 5555
rect 404 5489 438 5491
rect 400 5475 442 5476
rect 378 5469 404 5475
rect 442 5469 464 5475
rect 400 5468 404 5469
rect 174 5429 246 5437
rect 295 5434 300 5468
rect 324 5434 329 5468
rect 224 5399 226 5415
rect 196 5391 226 5399
rect 332 5397 336 5465
rect 367 5434 438 5468
rect 400 5427 404 5434
rect 454 5421 504 5423
rect 494 5417 548 5421
rect 494 5412 514 5417
rect 504 5397 506 5412
rect 196 5387 230 5391
rect 196 5357 204 5387
rect 216 5357 230 5387
rect 400 5389 404 5397
rect 174 5323 181 5349
rect 224 5310 226 5357
rect 256 5349 328 5357
rect 332 5355 336 5385
rect 400 5355 408 5389
rect 434 5355 438 5389
rect 498 5387 506 5397
rect 514 5387 515 5407
rect 504 5371 506 5387
rect 525 5378 528 5412
rect 547 5387 548 5407
rect 557 5387 564 5397
rect 514 5371 530 5377
rect 532 5371 548 5377
rect 289 5320 305 5322
rect 196 5276 204 5310
rect 216 5276 230 5310
rect 244 5276 257 5310
rect 300 5306 308 5319
rect 332 5317 342 5355
rect 400 5347 404 5355
rect 336 5307 342 5317
rect 224 5229 226 5276
rect 278 5272 291 5306
rect 300 5290 321 5306
rect 332 5297 342 5307
rect 400 5307 409 5335
rect 562 5318 612 5320
rect 466 5309 497 5311
rect 565 5309 596 5311
rect 300 5288 312 5290
rect 300 5272 321 5288
rect 300 5266 308 5272
rect 289 5256 308 5266
rect 196 5199 204 5229
rect 216 5199 230 5229
rect 196 5195 230 5199
rect 196 5187 226 5195
rect 300 5187 308 5256
rect 332 5263 351 5297
rect 361 5263 375 5297
rect 400 5263 411 5307
rect 442 5302 500 5309
rect 466 5301 500 5302
rect 565 5301 599 5309
rect 497 5285 500 5301
rect 596 5285 599 5301
rect 466 5284 500 5285
rect 442 5277 500 5284
rect 565 5277 599 5285
rect 612 5268 614 5318
rect 332 5239 342 5263
rect 336 5227 342 5239
rect 224 5171 226 5187
rect 332 5159 342 5227
rect 400 5231 404 5239
rect 400 5197 408 5231
rect 434 5197 438 5231
rect 454 5215 504 5217
rect 504 5199 506 5215
rect 514 5209 530 5215
rect 532 5209 548 5215
rect 525 5199 548 5208
rect 400 5189 404 5197
rect 498 5189 506 5199
rect 504 5165 506 5189
rect 514 5179 515 5199
rect 525 5174 528 5199
rect 547 5179 548 5199
rect 557 5189 564 5199
rect 514 5165 548 5169
rect 151 5118 156 5152
rect 174 5149 246 5157
rect 256 5149 328 5157
rect 336 5151 342 5159
rect 400 5154 404 5159
rect 180 5121 185 5149
rect 174 5113 246 5121
rect 256 5113 328 5121
rect 332 5119 336 5149
rect 400 5120 438 5154
rect 224 5083 226 5099
rect 196 5075 226 5083
rect 196 5071 230 5075
rect 196 5041 204 5071
rect 216 5041 230 5071
rect 224 4994 226 5041
rect 300 5014 308 5083
rect 332 5081 342 5119
rect 400 5111 404 5120
rect 454 5105 504 5107
rect 494 5101 548 5105
rect 494 5096 514 5101
rect 504 5081 506 5096
rect 336 5069 342 5081
rect 289 5004 308 5014
rect 300 4998 308 5004
rect 332 5035 342 5069
rect 400 5073 404 5081
rect 400 5039 408 5073
rect 434 5039 438 5073
rect 498 5071 506 5081
rect 514 5071 515 5091
rect 504 5055 506 5071
rect 525 5062 528 5096
rect 547 5071 548 5091
rect 557 5071 564 5081
rect 514 5055 530 5061
rect 532 5055 548 5061
rect 332 5007 373 5035
rect 332 5001 351 5007
rect 196 4960 204 4994
rect 216 4960 230 4994
rect 244 4960 257 4994
rect 278 4964 291 4998
rect 300 4982 321 4998
rect 336 4991 351 5001
rect 300 4980 312 4982
rect 300 4964 321 4980
rect 332 4973 351 4991
rect 361 4973 375 5007
rect 400 5001 411 5039
rect 562 5002 612 5004
rect 400 4973 409 5001
rect 466 4993 497 4995
rect 565 4993 596 4995
rect 442 4986 500 4993
rect 466 4985 500 4986
rect 565 4985 599 4993
rect 174 4923 181 4947
rect 224 4913 226 4960
rect 300 4951 308 4964
rect 289 4948 305 4950
rect 332 4923 342 4973
rect 400 4953 404 4973
rect 497 4969 500 4985
rect 596 4969 599 4985
rect 466 4968 500 4969
rect 442 4961 500 4968
rect 565 4961 599 4969
rect 612 4952 614 5002
rect 256 4913 328 4921
rect 336 4915 342 4923
rect 400 4915 404 4923
rect 196 4883 204 4913
rect 216 4883 230 4913
rect 196 4879 230 4883
rect 196 4871 226 4879
rect 224 4855 226 4871
rect 332 4843 336 4911
rect 400 4881 408 4915
rect 434 4881 438 4915
rect 454 4899 504 4901
rect 504 4883 506 4899
rect 514 4893 530 4899
rect 532 4893 548 4899
rect 525 4883 548 4892
rect 400 4873 404 4881
rect 498 4873 506 4883
rect 504 4849 506 4873
rect 514 4863 515 4883
rect 525 4858 528 4883
rect 547 4863 548 4883
rect 557 4873 564 4883
rect 514 4849 548 4853
rect 400 4843 442 4844
rect 174 4833 246 4841
rect 400 4836 404 4843
rect 295 4802 300 4836
rect 324 4802 329 4836
rect 367 4802 438 4836
rect 400 4801 404 4802
rect 378 4795 404 4801
rect 442 4795 464 4801
rect 38 4779 80 4795
rect 400 4779 442 4795
rect -25 4765 25 4767
rect 455 4765 505 4767
rect 557 4765 607 4767
rect 16 4757 102 4765
rect 378 4757 464 4765
rect 8 4723 17 4757
rect 18 4755 51 4757
rect 80 4755 100 4757
rect 18 4723 100 4755
rect 380 4755 404 4757
rect 429 4755 438 4757
rect 442 4755 462 4757
rect 16 4715 102 4723
rect 42 4699 76 4701
rect 16 4679 38 4685
rect 42 4676 76 4680
rect 80 4679 102 4685
rect 42 4646 46 4676
rect 72 4646 76 4676
rect 42 4565 46 4599
rect 72 4565 76 4599
rect -25 4528 25 4530
rect 0 4520 14 4521
rect 0 4519 17 4520
rect 25 4519 27 4528
rect 0 4512 38 4519
rect 0 4511 34 4512
rect 0 4495 8 4511
rect 14 4495 34 4511
rect 0 4494 34 4495
rect 0 4487 38 4494
rect 14 4486 17 4487
rect 25 4478 27 4487
rect 42 4458 45 4548
rect 69 4533 80 4565
rect 107 4533 143 4561
rect 107 4527 119 4533
rect 109 4499 119 4527
rect 129 4499 143 4533
rect 42 4407 46 4441
rect 72 4407 76 4441
rect 38 4369 80 4370
rect 42 4328 76 4362
rect 79 4328 113 4362
rect 42 4249 46 4283
rect 72 4249 76 4283
rect -25 4212 25 4214
rect 0 4204 14 4205
rect 0 4203 17 4204
rect 25 4203 27 4212
rect 0 4196 38 4203
rect 0 4195 34 4196
rect 0 4179 8 4195
rect 14 4179 34 4195
rect 0 4178 34 4179
rect 0 4171 38 4178
rect 14 4170 17 4171
rect 25 4162 27 4171
rect 42 4142 45 4232
rect 71 4201 80 4229
rect 69 4163 80 4201
rect 107 4157 119 4191
rect 129 4163 143 4191
rect 129 4157 141 4163
rect 42 4091 46 4125
rect 72 4091 76 4125
rect 42 4044 76 4048
rect 42 4014 46 4044
rect 72 4014 76 4044
rect 16 4005 38 4011
rect 80 4005 102 4011
rect 144 4005 148 4753
rect 332 4685 336 4753
rect 380 4723 462 4755
rect 463 4723 472 4757
rect 480 4723 497 4757
rect 378 4715 464 4723
rect 505 4715 507 4765
rect 514 4723 548 4757
rect 565 4723 582 4757
rect 607 4715 609 4765
rect 404 4699 438 4701
rect 400 4685 442 4686
rect 378 4679 404 4685
rect 442 4679 464 4685
rect 400 4678 404 4679
rect 174 4639 246 4647
rect 295 4644 300 4678
rect 324 4644 329 4678
rect 224 4609 226 4625
rect 196 4601 226 4609
rect 332 4607 336 4675
rect 367 4644 438 4678
rect 400 4637 404 4644
rect 454 4631 504 4633
rect 494 4627 548 4631
rect 494 4622 514 4627
rect 504 4607 506 4622
rect 196 4597 230 4601
rect 196 4567 204 4597
rect 216 4567 230 4597
rect 400 4599 404 4607
rect 174 4533 181 4559
rect 224 4520 226 4567
rect 256 4559 328 4567
rect 332 4565 336 4595
rect 400 4565 408 4599
rect 434 4565 438 4599
rect 498 4597 506 4607
rect 514 4597 515 4617
rect 504 4581 506 4597
rect 525 4588 528 4622
rect 547 4597 548 4617
rect 557 4597 564 4607
rect 514 4581 530 4587
rect 532 4581 548 4587
rect 289 4530 305 4532
rect 196 4486 204 4520
rect 216 4486 230 4520
rect 244 4486 257 4520
rect 300 4516 308 4529
rect 332 4527 342 4565
rect 400 4557 404 4565
rect 336 4517 342 4527
rect 224 4439 226 4486
rect 278 4482 291 4516
rect 300 4500 321 4516
rect 332 4507 342 4517
rect 400 4517 409 4545
rect 562 4528 612 4530
rect 466 4519 497 4521
rect 565 4519 596 4521
rect 300 4498 312 4500
rect 300 4482 321 4498
rect 300 4476 308 4482
rect 289 4466 308 4476
rect 196 4409 204 4439
rect 216 4409 230 4439
rect 196 4405 230 4409
rect 196 4397 226 4405
rect 300 4397 308 4466
rect 332 4473 351 4507
rect 361 4473 375 4507
rect 400 4473 411 4517
rect 442 4512 500 4519
rect 466 4511 500 4512
rect 565 4511 599 4519
rect 497 4495 500 4511
rect 596 4495 599 4511
rect 466 4494 500 4495
rect 442 4487 500 4494
rect 565 4487 599 4495
rect 612 4478 614 4528
rect 332 4449 342 4473
rect 336 4437 342 4449
rect 224 4381 226 4397
rect 332 4369 342 4437
rect 400 4441 404 4449
rect 400 4407 408 4441
rect 434 4407 438 4441
rect 454 4425 504 4427
rect 504 4409 506 4425
rect 514 4419 530 4425
rect 532 4419 548 4425
rect 525 4409 548 4418
rect 400 4399 404 4407
rect 498 4399 506 4409
rect 504 4375 506 4399
rect 514 4389 515 4409
rect 525 4384 528 4409
rect 547 4389 548 4409
rect 557 4399 564 4409
rect 514 4375 548 4379
rect 151 4328 156 4362
rect 174 4359 246 4367
rect 256 4359 328 4367
rect 336 4361 342 4369
rect 400 4364 404 4369
rect 180 4331 185 4359
rect 174 4323 246 4331
rect 256 4323 328 4331
rect 332 4329 336 4359
rect 400 4330 438 4364
rect 224 4293 226 4309
rect 196 4285 226 4293
rect 196 4281 230 4285
rect 196 4251 204 4281
rect 216 4251 230 4281
rect 224 4204 226 4251
rect 300 4224 308 4293
rect 332 4291 342 4329
rect 400 4321 404 4330
rect 454 4315 504 4317
rect 494 4311 548 4315
rect 494 4306 514 4311
rect 504 4291 506 4306
rect 336 4279 342 4291
rect 289 4214 308 4224
rect 300 4208 308 4214
rect 332 4245 342 4279
rect 400 4283 404 4291
rect 400 4249 408 4283
rect 434 4249 438 4283
rect 498 4281 506 4291
rect 514 4281 515 4301
rect 504 4265 506 4281
rect 525 4272 528 4306
rect 547 4281 548 4301
rect 557 4281 564 4291
rect 514 4265 530 4271
rect 532 4265 548 4271
rect 332 4217 373 4245
rect 332 4211 351 4217
rect 196 4170 204 4204
rect 216 4170 230 4204
rect 244 4170 257 4204
rect 278 4174 291 4208
rect 300 4192 321 4208
rect 336 4201 351 4211
rect 300 4190 312 4192
rect 300 4174 321 4190
rect 332 4183 351 4201
rect 361 4183 375 4217
rect 400 4211 411 4249
rect 562 4212 612 4214
rect 400 4183 409 4211
rect 466 4203 497 4205
rect 565 4203 596 4205
rect 442 4196 500 4203
rect 466 4195 500 4196
rect 565 4195 599 4203
rect 174 4133 181 4157
rect 224 4123 226 4170
rect 300 4161 308 4174
rect 289 4158 305 4160
rect 332 4133 342 4183
rect 400 4163 404 4183
rect 497 4179 500 4195
rect 596 4179 599 4195
rect 466 4178 500 4179
rect 442 4171 500 4178
rect 565 4171 599 4179
rect 612 4162 614 4212
rect 256 4123 328 4131
rect 336 4125 342 4133
rect 400 4125 404 4133
rect 196 4093 204 4123
rect 216 4093 230 4123
rect 196 4089 230 4093
rect 196 4081 226 4089
rect 224 4065 226 4081
rect 332 4053 336 4121
rect 400 4091 408 4125
rect 434 4091 438 4125
rect 454 4109 504 4111
rect 504 4093 506 4109
rect 514 4103 530 4109
rect 532 4103 548 4109
rect 525 4093 548 4102
rect 400 4083 404 4091
rect 498 4083 506 4093
rect 504 4059 506 4083
rect 514 4073 515 4093
rect 525 4068 528 4093
rect 547 4073 548 4093
rect 557 4083 564 4093
rect 514 4059 548 4063
rect 400 4053 442 4054
rect 174 4043 246 4051
rect 400 4046 404 4053
rect 295 4012 300 4046
rect 324 4012 329 4046
rect 367 4012 438 4046
rect 400 4011 404 4012
rect 378 4005 404 4011
rect 442 4005 464 4011
rect 38 3989 80 4005
rect 400 3989 442 4005
rect -25 3975 25 3977
rect 455 3975 505 3977
rect 557 3975 607 3977
rect 16 3967 102 3975
rect 378 3967 464 3975
rect 8 3933 17 3967
rect 18 3965 51 3967
rect 80 3965 100 3967
rect 18 3933 100 3965
rect 380 3965 404 3967
rect 429 3965 438 3967
rect 442 3965 462 3967
rect 16 3925 102 3933
rect 42 3909 76 3911
rect 16 3889 38 3895
rect 42 3886 76 3890
rect 80 3889 102 3895
rect 42 3856 46 3886
rect 72 3856 76 3886
rect 42 3775 46 3809
rect 72 3775 76 3809
rect -25 3738 25 3740
rect 0 3730 14 3731
rect 0 3729 17 3730
rect 25 3729 27 3738
rect 0 3722 38 3729
rect 0 3721 34 3722
rect 0 3705 8 3721
rect 14 3705 34 3721
rect 0 3704 34 3705
rect 0 3697 38 3704
rect 14 3696 17 3697
rect 25 3688 27 3697
rect 42 3668 45 3758
rect 69 3743 80 3775
rect 107 3743 143 3771
rect 107 3737 119 3743
rect 109 3709 119 3737
rect 129 3709 143 3743
rect 42 3617 46 3651
rect 72 3617 76 3651
rect 38 3579 80 3580
rect 42 3538 76 3572
rect 79 3538 113 3572
rect 42 3459 46 3493
rect 72 3459 76 3493
rect -25 3422 25 3424
rect 0 3414 14 3415
rect 0 3413 17 3414
rect 25 3413 27 3422
rect 0 3406 38 3413
rect 0 3405 34 3406
rect 0 3389 8 3405
rect 14 3389 34 3405
rect 0 3388 34 3389
rect 0 3381 38 3388
rect 14 3380 17 3381
rect 25 3372 27 3381
rect 42 3352 45 3442
rect 71 3411 80 3439
rect 69 3373 80 3411
rect 107 3367 119 3401
rect 129 3373 143 3401
rect 129 3367 141 3373
rect 42 3301 46 3335
rect 72 3301 76 3335
rect 42 3254 76 3258
rect 42 3224 46 3254
rect 72 3224 76 3254
rect 16 3215 38 3221
rect 80 3215 102 3221
rect 144 3215 148 3963
rect 332 3895 336 3963
rect 380 3933 462 3965
rect 463 3933 472 3967
rect 480 3933 497 3967
rect 378 3925 464 3933
rect 505 3925 507 3975
rect 514 3933 548 3967
rect 565 3933 582 3967
rect 607 3925 609 3975
rect 404 3909 438 3911
rect 400 3895 442 3896
rect 378 3889 404 3895
rect 442 3889 464 3895
rect 400 3888 404 3889
rect 174 3849 246 3857
rect 295 3854 300 3888
rect 324 3854 329 3888
rect 224 3819 226 3835
rect 196 3811 226 3819
rect 332 3817 336 3885
rect 367 3854 438 3888
rect 400 3847 404 3854
rect 454 3841 504 3843
rect 494 3837 548 3841
rect 494 3832 514 3837
rect 504 3817 506 3832
rect 196 3807 230 3811
rect 196 3777 204 3807
rect 216 3777 230 3807
rect 400 3809 404 3817
rect 174 3743 181 3769
rect 224 3730 226 3777
rect 256 3769 328 3777
rect 332 3775 336 3805
rect 400 3775 408 3809
rect 434 3775 438 3809
rect 498 3807 506 3817
rect 514 3807 515 3827
rect 504 3791 506 3807
rect 525 3798 528 3832
rect 547 3807 548 3827
rect 557 3807 564 3817
rect 514 3791 530 3797
rect 532 3791 548 3797
rect 289 3740 305 3742
rect 196 3696 204 3730
rect 216 3696 230 3730
rect 244 3696 257 3730
rect 300 3726 308 3739
rect 332 3737 342 3775
rect 400 3767 404 3775
rect 336 3727 342 3737
rect 224 3649 226 3696
rect 278 3692 291 3726
rect 300 3710 321 3726
rect 332 3717 342 3727
rect 400 3727 409 3755
rect 562 3738 612 3740
rect 466 3729 497 3731
rect 565 3729 596 3731
rect 300 3708 312 3710
rect 300 3692 321 3708
rect 300 3686 308 3692
rect 289 3676 308 3686
rect 196 3619 204 3649
rect 216 3619 230 3649
rect 196 3615 230 3619
rect 196 3607 226 3615
rect 300 3607 308 3676
rect 332 3683 351 3717
rect 361 3683 375 3717
rect 400 3683 411 3727
rect 442 3722 500 3729
rect 466 3721 500 3722
rect 565 3721 599 3729
rect 497 3705 500 3721
rect 596 3705 599 3721
rect 466 3704 500 3705
rect 442 3697 500 3704
rect 565 3697 599 3705
rect 612 3688 614 3738
rect 332 3659 342 3683
rect 336 3647 342 3659
rect 224 3591 226 3607
rect 332 3579 342 3647
rect 400 3651 404 3659
rect 400 3617 408 3651
rect 434 3617 438 3651
rect 454 3635 504 3637
rect 504 3619 506 3635
rect 514 3629 530 3635
rect 532 3629 548 3635
rect 525 3619 548 3628
rect 400 3609 404 3617
rect 498 3609 506 3619
rect 504 3585 506 3609
rect 514 3599 515 3619
rect 525 3594 528 3619
rect 547 3599 548 3619
rect 557 3609 564 3619
rect 514 3585 548 3589
rect 151 3538 156 3572
rect 174 3569 246 3577
rect 256 3569 328 3577
rect 336 3571 342 3579
rect 400 3574 404 3579
rect 180 3541 185 3569
rect 174 3533 246 3541
rect 256 3533 328 3541
rect 332 3539 336 3569
rect 400 3540 438 3574
rect 224 3503 226 3519
rect 196 3495 226 3503
rect 196 3491 230 3495
rect 196 3461 204 3491
rect 216 3461 230 3491
rect 224 3414 226 3461
rect 300 3434 308 3503
rect 332 3501 342 3539
rect 400 3531 404 3540
rect 454 3525 504 3527
rect 494 3521 548 3525
rect 494 3516 514 3521
rect 504 3501 506 3516
rect 336 3489 342 3501
rect 289 3424 308 3434
rect 300 3418 308 3424
rect 332 3455 342 3489
rect 400 3493 404 3501
rect 400 3459 408 3493
rect 434 3459 438 3493
rect 498 3491 506 3501
rect 514 3491 515 3511
rect 504 3475 506 3491
rect 525 3482 528 3516
rect 547 3491 548 3511
rect 557 3491 564 3501
rect 514 3475 530 3481
rect 532 3475 548 3481
rect 332 3427 373 3455
rect 332 3421 351 3427
rect 196 3380 204 3414
rect 216 3380 230 3414
rect 244 3380 257 3414
rect 278 3384 291 3418
rect 300 3402 321 3418
rect 336 3411 351 3421
rect 300 3400 312 3402
rect 300 3384 321 3400
rect 332 3393 351 3411
rect 361 3393 375 3427
rect 400 3421 411 3459
rect 562 3422 612 3424
rect 400 3393 409 3421
rect 466 3413 497 3415
rect 565 3413 596 3415
rect 442 3406 500 3413
rect 466 3405 500 3406
rect 565 3405 599 3413
rect 174 3343 181 3367
rect 224 3333 226 3380
rect 300 3371 308 3384
rect 289 3368 305 3370
rect 332 3343 342 3393
rect 400 3373 404 3393
rect 497 3389 500 3405
rect 596 3389 599 3405
rect 466 3388 500 3389
rect 442 3381 500 3388
rect 565 3381 599 3389
rect 612 3372 614 3422
rect 256 3333 328 3341
rect 336 3335 342 3343
rect 400 3335 404 3343
rect 196 3303 204 3333
rect 216 3303 230 3333
rect 196 3299 230 3303
rect 196 3291 226 3299
rect 224 3275 226 3291
rect 332 3263 336 3331
rect 400 3301 408 3335
rect 434 3301 438 3335
rect 454 3319 504 3321
rect 504 3303 506 3319
rect 514 3313 530 3319
rect 532 3313 548 3319
rect 525 3303 548 3312
rect 400 3293 404 3301
rect 498 3293 506 3303
rect 504 3269 506 3293
rect 514 3283 515 3303
rect 525 3278 528 3303
rect 547 3283 548 3303
rect 557 3293 564 3303
rect 514 3269 548 3273
rect 400 3263 442 3264
rect 174 3253 246 3261
rect 400 3256 404 3263
rect 295 3222 300 3256
rect 324 3222 329 3256
rect 367 3222 438 3256
rect 400 3221 404 3222
rect 378 3215 404 3221
rect 442 3215 464 3221
rect 38 3199 80 3215
rect 400 3199 442 3215
rect -25 3185 25 3187
rect 455 3185 505 3187
rect 557 3185 607 3187
rect 16 3177 102 3185
rect 378 3177 464 3185
rect 8 3143 17 3177
rect 18 3175 51 3177
rect 80 3175 100 3177
rect 18 3143 100 3175
rect 380 3175 404 3177
rect 429 3175 438 3177
rect 442 3175 462 3177
rect 16 3135 102 3143
rect 42 3119 76 3121
rect 16 3099 38 3105
rect 42 3096 76 3100
rect 80 3099 102 3105
rect 42 3066 46 3096
rect 72 3066 76 3096
rect 42 2985 46 3019
rect 72 2985 76 3019
rect -25 2948 25 2950
rect 0 2940 14 2941
rect 0 2939 17 2940
rect 25 2939 27 2948
rect 0 2932 38 2939
rect 0 2931 34 2932
rect 0 2915 8 2931
rect 14 2915 34 2931
rect 0 2914 34 2915
rect 0 2907 38 2914
rect 14 2906 17 2907
rect 25 2898 27 2907
rect 42 2878 45 2968
rect 69 2953 80 2985
rect 107 2953 143 2981
rect 107 2947 119 2953
rect 109 2919 119 2947
rect 129 2919 143 2953
rect 42 2827 46 2861
rect 72 2827 76 2861
rect 38 2789 80 2790
rect 42 2748 76 2782
rect 79 2748 113 2782
rect 42 2669 46 2703
rect 72 2669 76 2703
rect -25 2632 25 2634
rect 0 2624 14 2625
rect 0 2623 17 2624
rect 25 2623 27 2632
rect 0 2616 38 2623
rect 0 2615 34 2616
rect 0 2599 8 2615
rect 14 2599 34 2615
rect 0 2598 34 2599
rect 0 2591 38 2598
rect 14 2590 17 2591
rect 25 2582 27 2591
rect 42 2562 45 2652
rect 71 2621 80 2649
rect 69 2583 80 2621
rect 107 2577 119 2611
rect 129 2583 143 2611
rect 129 2577 141 2583
rect 42 2511 46 2545
rect 72 2511 76 2545
rect 42 2464 76 2468
rect 42 2434 46 2464
rect 72 2434 76 2464
rect 16 2425 38 2431
rect 80 2425 102 2431
rect 144 2425 148 3173
rect 332 3105 336 3173
rect 380 3143 462 3175
rect 463 3143 472 3177
rect 480 3143 497 3177
rect 378 3135 464 3143
rect 505 3135 507 3185
rect 514 3143 548 3177
rect 565 3143 582 3177
rect 607 3135 609 3185
rect 404 3119 438 3121
rect 400 3105 442 3106
rect 378 3099 404 3105
rect 442 3099 464 3105
rect 400 3098 404 3099
rect 174 3059 246 3067
rect 295 3064 300 3098
rect 324 3064 329 3098
rect 224 3029 226 3045
rect 196 3021 226 3029
rect 332 3027 336 3095
rect 367 3064 438 3098
rect 400 3057 404 3064
rect 454 3051 504 3053
rect 494 3047 548 3051
rect 494 3042 514 3047
rect 504 3027 506 3042
rect 196 3017 230 3021
rect 196 2987 204 3017
rect 216 2987 230 3017
rect 400 3019 404 3027
rect 174 2953 181 2979
rect 224 2940 226 2987
rect 256 2979 328 2987
rect 332 2985 336 3015
rect 400 2985 408 3019
rect 434 2985 438 3019
rect 498 3017 506 3027
rect 514 3017 515 3037
rect 504 3001 506 3017
rect 525 3008 528 3042
rect 547 3017 548 3037
rect 557 3017 564 3027
rect 514 3001 530 3007
rect 532 3001 548 3007
rect 289 2950 305 2952
rect 196 2906 204 2940
rect 216 2906 230 2940
rect 244 2906 257 2940
rect 300 2936 308 2949
rect 332 2947 342 2985
rect 400 2977 404 2985
rect 336 2937 342 2947
rect 224 2859 226 2906
rect 278 2902 291 2936
rect 300 2920 321 2936
rect 332 2927 342 2937
rect 400 2937 409 2965
rect 562 2948 612 2950
rect 466 2939 497 2941
rect 565 2939 596 2941
rect 300 2918 312 2920
rect 300 2902 321 2918
rect 300 2896 308 2902
rect 289 2886 308 2896
rect 196 2829 204 2859
rect 216 2829 230 2859
rect 196 2825 230 2829
rect 196 2817 226 2825
rect 300 2817 308 2886
rect 332 2893 351 2927
rect 361 2893 375 2927
rect 400 2893 411 2937
rect 442 2932 500 2939
rect 466 2931 500 2932
rect 565 2931 599 2939
rect 497 2915 500 2931
rect 596 2915 599 2931
rect 466 2914 500 2915
rect 442 2907 500 2914
rect 565 2907 599 2915
rect 612 2898 614 2948
rect 332 2869 342 2893
rect 336 2857 342 2869
rect 224 2801 226 2817
rect 332 2789 342 2857
rect 400 2861 404 2869
rect 400 2827 408 2861
rect 434 2827 438 2861
rect 454 2845 504 2847
rect 504 2829 506 2845
rect 514 2839 530 2845
rect 532 2839 548 2845
rect 525 2829 548 2838
rect 400 2819 404 2827
rect 498 2819 506 2829
rect 504 2795 506 2819
rect 514 2809 515 2829
rect 525 2804 528 2829
rect 547 2809 548 2829
rect 557 2819 564 2829
rect 514 2795 548 2799
rect 151 2748 156 2782
rect 174 2779 246 2787
rect 256 2779 328 2787
rect 336 2781 342 2789
rect 400 2784 404 2789
rect 180 2751 185 2779
rect 174 2743 246 2751
rect 256 2743 328 2751
rect 332 2749 336 2779
rect 400 2750 438 2784
rect 224 2713 226 2729
rect 196 2705 226 2713
rect 196 2701 230 2705
rect 196 2671 204 2701
rect 216 2671 230 2701
rect 224 2624 226 2671
rect 300 2644 308 2713
rect 332 2711 342 2749
rect 400 2741 404 2750
rect 454 2735 504 2737
rect 494 2731 548 2735
rect 494 2726 514 2731
rect 504 2711 506 2726
rect 336 2699 342 2711
rect 289 2634 308 2644
rect 300 2628 308 2634
rect 332 2665 342 2699
rect 400 2703 404 2711
rect 400 2669 408 2703
rect 434 2669 438 2703
rect 498 2701 506 2711
rect 514 2701 515 2721
rect 504 2685 506 2701
rect 525 2692 528 2726
rect 547 2701 548 2721
rect 557 2701 564 2711
rect 514 2685 530 2691
rect 532 2685 548 2691
rect 332 2637 373 2665
rect 332 2631 351 2637
rect 196 2590 204 2624
rect 216 2590 230 2624
rect 244 2590 257 2624
rect 278 2594 291 2628
rect 300 2612 321 2628
rect 336 2621 351 2631
rect 300 2610 312 2612
rect 300 2594 321 2610
rect 332 2603 351 2621
rect 361 2603 375 2637
rect 400 2631 411 2669
rect 562 2632 612 2634
rect 400 2603 409 2631
rect 466 2623 497 2625
rect 565 2623 596 2625
rect 442 2616 500 2623
rect 466 2615 500 2616
rect 565 2615 599 2623
rect 174 2553 181 2577
rect 224 2543 226 2590
rect 300 2581 308 2594
rect 289 2578 305 2580
rect 332 2553 342 2603
rect 400 2583 404 2603
rect 497 2599 500 2615
rect 596 2599 599 2615
rect 466 2598 500 2599
rect 442 2591 500 2598
rect 565 2591 599 2599
rect 612 2582 614 2632
rect 256 2543 328 2551
rect 336 2545 342 2553
rect 400 2545 404 2553
rect 196 2513 204 2543
rect 216 2513 230 2543
rect 196 2509 230 2513
rect 196 2501 226 2509
rect 224 2485 226 2501
rect 332 2473 336 2541
rect 400 2511 408 2545
rect 434 2511 438 2545
rect 454 2529 504 2531
rect 504 2513 506 2529
rect 514 2523 530 2529
rect 532 2523 548 2529
rect 525 2513 548 2522
rect 400 2503 404 2511
rect 498 2503 506 2513
rect 504 2479 506 2503
rect 514 2493 515 2513
rect 525 2488 528 2513
rect 547 2493 548 2513
rect 557 2503 564 2513
rect 514 2479 548 2483
rect 400 2473 442 2474
rect 174 2463 246 2471
rect 400 2466 404 2473
rect 295 2432 300 2466
rect 324 2432 329 2466
rect 367 2432 438 2466
rect 400 2431 404 2432
rect 378 2425 404 2431
rect 442 2425 464 2431
rect 38 2409 80 2425
rect 400 2409 442 2425
rect -25 2395 25 2397
rect 455 2395 505 2397
rect 557 2395 607 2397
rect 16 2387 102 2395
rect 378 2387 464 2395
rect 8 2353 17 2387
rect 18 2385 51 2387
rect 80 2385 100 2387
rect 18 2353 100 2385
rect 380 2385 404 2387
rect 429 2385 438 2387
rect 442 2385 462 2387
rect 16 2345 102 2353
rect 42 2329 76 2331
rect 16 2309 38 2315
rect 42 2306 76 2310
rect 80 2309 102 2315
rect 42 2276 46 2306
rect 72 2276 76 2306
rect 42 2195 46 2229
rect 72 2195 76 2229
rect -25 2158 25 2160
rect 0 2150 14 2151
rect 0 2149 17 2150
rect 25 2149 27 2158
rect 0 2142 38 2149
rect 0 2141 34 2142
rect 0 2125 8 2141
rect 14 2125 34 2141
rect 0 2124 34 2125
rect 0 2117 38 2124
rect 14 2116 17 2117
rect 25 2108 27 2117
rect 42 2088 45 2178
rect 69 2163 80 2195
rect 107 2163 143 2191
rect 107 2157 119 2163
rect 109 2129 119 2157
rect 129 2129 143 2163
rect 42 2037 46 2071
rect 72 2037 76 2071
rect 38 1999 80 2000
rect 42 1958 76 1992
rect 79 1958 113 1992
rect 42 1879 46 1913
rect 72 1879 76 1913
rect -25 1842 25 1844
rect 0 1834 14 1835
rect 0 1833 17 1834
rect 25 1833 27 1842
rect 0 1826 38 1833
rect 0 1825 34 1826
rect 0 1809 8 1825
rect 14 1809 34 1825
rect 0 1808 34 1809
rect 0 1801 38 1808
rect 14 1800 17 1801
rect 25 1792 27 1801
rect 42 1772 45 1862
rect 71 1831 80 1859
rect 69 1793 80 1831
rect 107 1787 119 1821
rect 129 1793 143 1821
rect 129 1787 141 1793
rect 42 1721 46 1755
rect 72 1721 76 1755
rect 42 1674 76 1678
rect 42 1644 46 1674
rect 72 1644 76 1674
rect 16 1635 38 1641
rect 80 1635 102 1641
rect 144 1635 148 2383
rect 332 2315 336 2383
rect 380 2353 462 2385
rect 463 2353 472 2387
rect 480 2353 497 2387
rect 378 2345 464 2353
rect 505 2345 507 2395
rect 514 2353 548 2387
rect 565 2353 582 2387
rect 607 2345 609 2395
rect 404 2329 438 2331
rect 400 2315 442 2316
rect 378 2309 404 2315
rect 442 2309 464 2315
rect 400 2308 404 2309
rect 174 2269 246 2277
rect 295 2274 300 2308
rect 324 2274 329 2308
rect 224 2239 226 2255
rect 196 2231 226 2239
rect 332 2237 336 2305
rect 367 2274 438 2308
rect 400 2267 404 2274
rect 454 2261 504 2263
rect 494 2257 548 2261
rect 494 2252 514 2257
rect 504 2237 506 2252
rect 196 2227 230 2231
rect 196 2197 204 2227
rect 216 2197 230 2227
rect 400 2229 404 2237
rect 174 2163 181 2189
rect 224 2150 226 2197
rect 256 2189 328 2197
rect 332 2195 336 2225
rect 400 2195 408 2229
rect 434 2195 438 2229
rect 498 2227 506 2237
rect 514 2227 515 2247
rect 504 2211 506 2227
rect 525 2218 528 2252
rect 547 2227 548 2247
rect 557 2227 564 2237
rect 514 2211 530 2217
rect 532 2211 548 2217
rect 289 2160 305 2162
rect 196 2116 204 2150
rect 216 2116 230 2150
rect 244 2116 257 2150
rect 300 2146 308 2159
rect 332 2157 342 2195
rect 400 2187 404 2195
rect 336 2147 342 2157
rect 224 2069 226 2116
rect 278 2112 291 2146
rect 300 2130 321 2146
rect 332 2137 342 2147
rect 400 2147 409 2175
rect 562 2158 612 2160
rect 466 2149 497 2151
rect 565 2149 596 2151
rect 300 2128 312 2130
rect 300 2112 321 2128
rect 300 2106 308 2112
rect 289 2096 308 2106
rect 196 2039 204 2069
rect 216 2039 230 2069
rect 196 2035 230 2039
rect 196 2027 226 2035
rect 300 2027 308 2096
rect 332 2103 351 2137
rect 361 2103 375 2137
rect 400 2103 411 2147
rect 442 2142 500 2149
rect 466 2141 500 2142
rect 565 2141 599 2149
rect 497 2125 500 2141
rect 596 2125 599 2141
rect 466 2124 500 2125
rect 442 2117 500 2124
rect 565 2117 599 2125
rect 612 2108 614 2158
rect 332 2079 342 2103
rect 336 2067 342 2079
rect 224 2011 226 2027
rect 332 1999 342 2067
rect 400 2071 404 2079
rect 400 2037 408 2071
rect 434 2037 438 2071
rect 454 2055 504 2057
rect 504 2039 506 2055
rect 514 2049 530 2055
rect 532 2049 548 2055
rect 525 2039 548 2048
rect 400 2029 404 2037
rect 498 2029 506 2039
rect 504 2005 506 2029
rect 514 2019 515 2039
rect 525 2014 528 2039
rect 547 2019 548 2039
rect 557 2029 564 2039
rect 514 2005 548 2009
rect 151 1958 156 1992
rect 174 1989 246 1997
rect 256 1989 328 1997
rect 336 1991 342 1999
rect 400 1994 404 1999
rect 180 1961 185 1989
rect 174 1953 246 1961
rect 256 1953 328 1961
rect 332 1959 336 1989
rect 400 1960 438 1994
rect 224 1923 226 1939
rect 196 1915 226 1923
rect 196 1911 230 1915
rect 196 1881 204 1911
rect 216 1881 230 1911
rect 224 1834 226 1881
rect 300 1854 308 1923
rect 332 1921 342 1959
rect 400 1951 404 1960
rect 454 1945 504 1947
rect 494 1941 548 1945
rect 494 1936 514 1941
rect 504 1921 506 1936
rect 336 1909 342 1921
rect 289 1844 308 1854
rect 300 1838 308 1844
rect 332 1875 342 1909
rect 400 1913 404 1921
rect 400 1879 408 1913
rect 434 1879 438 1913
rect 498 1911 506 1921
rect 514 1911 515 1931
rect 504 1895 506 1911
rect 525 1902 528 1936
rect 547 1911 548 1931
rect 557 1911 564 1921
rect 514 1895 530 1901
rect 532 1895 548 1901
rect 332 1847 373 1875
rect 332 1841 351 1847
rect 196 1800 204 1834
rect 216 1800 230 1834
rect 244 1800 257 1834
rect 278 1804 291 1838
rect 300 1822 321 1838
rect 336 1831 351 1841
rect 300 1820 312 1822
rect 300 1804 321 1820
rect 332 1813 351 1831
rect 361 1813 375 1847
rect 400 1841 411 1879
rect 562 1842 612 1844
rect 400 1813 409 1841
rect 466 1833 497 1835
rect 565 1833 596 1835
rect 442 1826 500 1833
rect 466 1825 500 1826
rect 565 1825 599 1833
rect 174 1763 181 1787
rect 224 1753 226 1800
rect 300 1791 308 1804
rect 289 1788 305 1790
rect 332 1763 342 1813
rect 400 1793 404 1813
rect 497 1809 500 1825
rect 596 1809 599 1825
rect 466 1808 500 1809
rect 442 1801 500 1808
rect 565 1801 599 1809
rect 612 1792 614 1842
rect 256 1753 328 1761
rect 336 1755 342 1763
rect 400 1755 404 1763
rect 196 1723 204 1753
rect 216 1723 230 1753
rect 196 1719 230 1723
rect 196 1711 226 1719
rect 224 1695 226 1711
rect 332 1683 336 1751
rect 400 1721 408 1755
rect 434 1721 438 1755
rect 454 1739 504 1741
rect 504 1723 506 1739
rect 514 1733 530 1739
rect 532 1733 548 1739
rect 525 1723 548 1732
rect 400 1713 404 1721
rect 498 1713 506 1723
rect 504 1689 506 1713
rect 514 1703 515 1723
rect 525 1698 528 1723
rect 547 1703 548 1723
rect 557 1713 564 1723
rect 514 1689 548 1693
rect 400 1683 442 1684
rect 174 1673 246 1681
rect 400 1676 404 1683
rect 295 1642 300 1676
rect 324 1642 329 1676
rect 367 1642 438 1676
rect 400 1641 404 1642
rect 378 1635 404 1641
rect 442 1635 464 1641
rect 38 1619 80 1635
rect 400 1619 442 1635
rect -25 1605 25 1607
rect 455 1605 505 1607
rect 557 1605 607 1607
rect 16 1597 102 1605
rect 378 1597 464 1605
rect 8 1563 17 1597
rect 18 1595 51 1597
rect 80 1595 100 1597
rect 18 1563 100 1595
rect 380 1595 404 1597
rect 429 1595 438 1597
rect 442 1595 462 1597
rect 16 1555 102 1563
rect 42 1539 76 1541
rect 16 1519 38 1525
rect 42 1516 76 1520
rect 80 1519 102 1525
rect 42 1486 46 1516
rect 72 1486 76 1516
rect 42 1405 46 1439
rect 72 1405 76 1439
rect -25 1368 25 1370
rect 0 1360 14 1361
rect 0 1359 17 1360
rect 25 1359 27 1368
rect 0 1352 38 1359
rect 0 1351 34 1352
rect 0 1335 8 1351
rect 14 1335 34 1351
rect 0 1334 34 1335
rect 0 1327 38 1334
rect 14 1326 17 1327
rect 25 1318 27 1327
rect 42 1298 45 1388
rect 69 1373 80 1405
rect 107 1373 143 1401
rect 107 1367 119 1373
rect 109 1339 119 1367
rect 129 1339 143 1373
rect 42 1247 46 1281
rect 72 1247 76 1281
rect 38 1209 80 1210
rect 42 1168 76 1202
rect 79 1168 113 1202
rect 42 1089 46 1123
rect 72 1089 76 1123
rect -25 1052 25 1054
rect 0 1044 14 1045
rect 0 1043 17 1044
rect 25 1043 27 1052
rect 0 1036 38 1043
rect 0 1035 34 1036
rect 0 1019 8 1035
rect 14 1019 34 1035
rect 0 1018 34 1019
rect 0 1011 38 1018
rect 14 1010 17 1011
rect 25 1002 27 1011
rect 42 982 45 1072
rect 71 1041 80 1069
rect 69 1003 80 1041
rect 107 997 119 1031
rect 129 1003 143 1031
rect 129 997 141 1003
rect 42 931 46 965
rect 72 931 76 965
rect 42 884 76 888
rect 42 854 46 884
rect 72 854 76 884
rect 16 845 38 851
rect 80 845 102 851
rect 144 845 148 1593
rect 332 1525 336 1593
rect 380 1563 462 1595
rect 463 1563 472 1597
rect 480 1563 497 1597
rect 378 1555 464 1563
rect 505 1555 507 1605
rect 514 1563 548 1597
rect 565 1563 582 1597
rect 607 1555 609 1605
rect 404 1539 438 1541
rect 400 1525 442 1526
rect 378 1519 404 1525
rect 442 1519 464 1525
rect 400 1518 404 1519
rect 174 1479 246 1487
rect 295 1484 300 1518
rect 324 1484 329 1518
rect 224 1449 226 1465
rect 196 1441 226 1449
rect 332 1447 336 1515
rect 367 1484 438 1518
rect 400 1477 404 1484
rect 454 1471 504 1473
rect 494 1467 548 1471
rect 494 1462 514 1467
rect 504 1447 506 1462
rect 196 1437 230 1441
rect 196 1407 204 1437
rect 216 1407 230 1437
rect 400 1439 404 1447
rect 174 1373 181 1399
rect 224 1360 226 1407
rect 256 1399 328 1407
rect 332 1405 336 1435
rect 400 1405 408 1439
rect 434 1405 438 1439
rect 498 1437 506 1447
rect 514 1437 515 1457
rect 504 1421 506 1437
rect 525 1428 528 1462
rect 547 1437 548 1457
rect 557 1437 564 1447
rect 514 1421 530 1427
rect 532 1421 548 1427
rect 289 1370 305 1372
rect 196 1326 204 1360
rect 216 1326 230 1360
rect 244 1326 257 1360
rect 300 1356 308 1369
rect 332 1367 342 1405
rect 400 1397 404 1405
rect 336 1357 342 1367
rect 224 1279 226 1326
rect 278 1322 291 1356
rect 300 1340 321 1356
rect 332 1347 342 1357
rect 400 1357 409 1385
rect 562 1368 612 1370
rect 466 1359 497 1361
rect 565 1359 596 1361
rect 300 1338 312 1340
rect 300 1322 321 1338
rect 300 1316 308 1322
rect 289 1306 308 1316
rect 196 1249 204 1279
rect 216 1249 230 1279
rect 196 1245 230 1249
rect 196 1237 226 1245
rect 300 1237 308 1306
rect 332 1313 351 1347
rect 361 1313 375 1347
rect 400 1313 411 1357
rect 442 1352 500 1359
rect 466 1351 500 1352
rect 565 1351 599 1359
rect 497 1335 500 1351
rect 596 1335 599 1351
rect 466 1334 500 1335
rect 442 1327 500 1334
rect 565 1327 599 1335
rect 612 1318 614 1368
rect 332 1289 342 1313
rect 336 1277 342 1289
rect 224 1221 226 1237
rect 332 1209 342 1277
rect 400 1281 404 1289
rect 400 1247 408 1281
rect 434 1247 438 1281
rect 454 1265 504 1267
rect 504 1249 506 1265
rect 514 1259 530 1265
rect 532 1259 548 1265
rect 525 1249 548 1258
rect 400 1239 404 1247
rect 498 1239 506 1249
rect 504 1215 506 1239
rect 514 1229 515 1249
rect 525 1224 528 1249
rect 547 1229 548 1249
rect 557 1239 564 1249
rect 514 1215 548 1219
rect 151 1168 156 1202
rect 174 1199 246 1207
rect 256 1199 328 1207
rect 336 1201 342 1209
rect 400 1204 404 1209
rect 180 1171 185 1199
rect 174 1163 246 1171
rect 256 1163 328 1171
rect 332 1169 336 1199
rect 400 1170 438 1204
rect 224 1133 226 1149
rect 196 1125 226 1133
rect 196 1121 230 1125
rect 196 1091 204 1121
rect 216 1091 230 1121
rect 224 1044 226 1091
rect 300 1064 308 1133
rect 332 1131 342 1169
rect 400 1161 404 1170
rect 454 1155 504 1157
rect 494 1151 548 1155
rect 494 1146 514 1151
rect 504 1131 506 1146
rect 336 1119 342 1131
rect 289 1054 308 1064
rect 300 1048 308 1054
rect 332 1085 342 1119
rect 400 1123 404 1131
rect 400 1089 408 1123
rect 434 1089 438 1123
rect 498 1121 506 1131
rect 514 1121 515 1141
rect 504 1105 506 1121
rect 525 1112 528 1146
rect 547 1121 548 1141
rect 557 1121 564 1131
rect 514 1105 530 1111
rect 532 1105 548 1111
rect 332 1057 373 1085
rect 332 1051 351 1057
rect 196 1010 204 1044
rect 216 1010 230 1044
rect 244 1010 257 1044
rect 278 1014 291 1048
rect 300 1032 321 1048
rect 336 1041 351 1051
rect 300 1030 312 1032
rect 300 1014 321 1030
rect 332 1023 351 1041
rect 361 1023 375 1057
rect 400 1051 411 1089
rect 562 1052 612 1054
rect 400 1023 409 1051
rect 466 1043 497 1045
rect 565 1043 596 1045
rect 442 1036 500 1043
rect 466 1035 500 1036
rect 565 1035 599 1043
rect 174 973 181 997
rect 224 963 226 1010
rect 300 1001 308 1014
rect 289 998 305 1000
rect 332 973 342 1023
rect 400 1003 404 1023
rect 497 1019 500 1035
rect 596 1019 599 1035
rect 466 1018 500 1019
rect 442 1011 500 1018
rect 565 1011 599 1019
rect 612 1002 614 1052
rect 256 963 328 971
rect 336 965 342 973
rect 400 965 404 973
rect 196 933 204 963
rect 216 933 230 963
rect 196 929 230 933
rect 196 921 226 929
rect 224 905 226 921
rect 332 893 336 961
rect 400 931 408 965
rect 434 931 438 965
rect 454 949 504 951
rect 504 933 506 949
rect 514 943 530 949
rect 532 943 548 949
rect 525 933 548 942
rect 400 923 404 931
rect 498 923 506 933
rect 504 899 506 923
rect 514 913 515 933
rect 525 908 528 933
rect 547 913 548 933
rect 557 923 564 933
rect 514 899 548 903
rect 400 893 442 894
rect 174 883 246 891
rect 400 886 404 893
rect 295 852 300 886
rect 324 852 329 886
rect 367 852 438 886
rect 400 851 404 852
rect 378 845 404 851
rect 442 845 464 851
rect 38 829 80 845
rect 400 829 442 845
rect -25 815 25 817
rect 455 815 505 817
rect 557 815 607 817
rect 16 807 102 815
rect 378 807 464 815
rect 8 773 17 807
rect 18 805 51 807
rect 80 805 100 807
rect 18 773 100 805
rect 380 805 404 807
rect 429 805 438 807
rect 442 805 462 807
rect 16 765 102 773
rect 42 749 76 751
rect 16 729 38 735
rect 42 726 76 730
rect 80 729 102 735
rect 42 696 46 726
rect 72 696 76 726
rect 69 583 80 621
rect 107 583 143 611
rect -25 578 25 580
rect 0 569 17 571
rect 25 569 27 578
rect 107 577 119 583
rect 0 562 38 569
rect 0 561 34 562
rect 0 545 8 561
rect 17 545 34 561
rect 109 549 119 577
rect 129 549 143 583
rect 0 544 34 545
rect 0 537 38 544
rect 25 528 27 537
rect 42 420 76 429
rect 38 419 80 420
rect 42 395 76 419
rect 79 395 113 412
rect 144 395 148 803
rect 332 735 336 803
rect 380 773 462 805
rect 463 773 472 807
rect 480 773 497 807
rect 378 765 464 773
rect 505 765 507 815
rect 514 773 548 807
rect 565 773 582 807
rect 607 765 609 815
rect 404 749 438 751
rect 400 735 442 736
rect 378 729 404 735
rect 442 729 464 735
rect 400 728 404 729
rect 295 694 300 728
rect 324 694 329 728
rect 332 657 336 725
rect 367 694 438 728
rect 400 687 404 694
rect 454 681 504 683
rect 494 677 548 681
rect 494 672 514 677
rect 504 657 506 672
rect 174 583 181 609
rect 332 577 336 645
rect 400 607 404 657
rect 498 647 506 657
rect 514 647 515 667
rect 504 631 506 647
rect 525 638 528 672
rect 547 647 548 667
rect 557 647 564 657
rect 514 631 530 637
rect 532 631 548 637
rect 400 567 409 595
rect 562 578 612 580
rect 463 569 497 571
rect 332 499 336 567
rect 341 523 351 557
rect 361 523 375 557
rect 400 523 411 567
rect 442 562 497 569
rect 463 561 497 562
rect 565 569 596 571
rect 565 561 599 569
rect 596 545 599 561
rect 463 544 497 545
rect 442 537 497 544
rect 565 537 599 545
rect 612 528 614 578
rect 332 419 336 487
rect 400 449 404 499
rect 454 475 504 477
rect 504 459 506 475
rect 514 469 530 475
rect 532 469 548 475
rect 525 459 548 468
rect 498 449 506 459
rect 404 419 438 429
rect 504 425 506 449
rect 514 439 515 459
rect 525 434 528 459
rect 547 439 548 459
rect 557 449 564 459
rect 514 425 548 429
rect 38 378 113 395
rect 151 378 156 412
rect 180 378 185 412
rect 400 411 438 419
rect 388 410 454 411
rect 400 403 408 410
rect 434 403 438 410
rect 400 395 438 403
rect 38 369 80 378
rect 400 369 442 395
<< metal1 >>
rect 78 0 114 26860
rect 150 0 186 26860
rect 222 26149 258 26490
rect 222 25359 258 25991
rect 222 24569 258 25201
rect 222 23779 258 24411
rect 222 22989 258 23621
rect 222 22199 258 22831
rect 222 21409 258 22041
rect 222 20619 258 21251
rect 222 19829 258 20461
rect 222 19039 258 19671
rect 222 18249 258 18881
rect 222 17459 258 18091
rect 222 16669 258 17301
rect 222 15879 258 16511
rect 222 15089 258 15721
rect 222 14299 258 14931
rect 222 13509 258 14141
rect 222 12719 258 13351
rect 222 11929 258 12561
rect 222 11139 258 11771
rect 222 10349 258 10981
rect 222 9559 258 10191
rect 222 8769 258 9401
rect 222 7979 258 8611
rect 222 7189 258 7821
rect 222 6399 258 7031
rect 222 5609 258 6241
rect 222 4819 258 5451
rect 222 4029 258 4661
rect 222 3239 258 3871
rect 222 2449 258 3081
rect 222 1659 258 2291
rect 222 869 258 1501
rect 222 370 258 711
rect 294 0 330 26860
rect 366 0 402 26860
<< metal2 >>
rect 0 26576 624 26686
rect 0 26393 624 26441
rect 186 26269 294 26345
rect 0 26173 624 26221
rect 186 26015 294 26125
rect 0 25919 624 25967
rect 186 25795 294 25871
rect 0 25699 624 25747
rect 0 25603 624 25651
rect 186 25479 294 25555
rect 0 25383 624 25431
rect 186 25225 294 25335
rect 0 25129 624 25177
rect 186 25005 294 25081
rect 0 24909 624 24957
rect 0 24813 624 24861
rect 186 24689 294 24765
rect 0 24593 624 24641
rect 186 24435 294 24545
rect 0 24339 624 24387
rect 186 24215 294 24291
rect 0 24119 624 24167
rect 0 24023 624 24071
rect 186 23899 294 23975
rect 0 23803 624 23851
rect 186 23645 294 23755
rect 0 23549 624 23597
rect 186 23425 294 23501
rect 0 23329 624 23377
rect 0 23233 624 23281
rect 186 23109 294 23185
rect 0 23013 624 23061
rect 186 22855 294 22965
rect 0 22759 624 22807
rect 186 22635 294 22711
rect 0 22539 624 22587
rect 0 22443 624 22491
rect 186 22319 294 22395
rect 0 22223 624 22271
rect 186 22065 294 22175
rect 0 21969 624 22017
rect 186 21845 294 21921
rect 0 21749 624 21797
rect 0 21653 624 21701
rect 186 21529 294 21605
rect 0 21433 624 21481
rect 186 21275 294 21385
rect 0 21179 624 21227
rect 186 21055 294 21131
rect 0 20959 624 21007
rect 0 20863 624 20911
rect 186 20739 294 20815
rect 0 20643 624 20691
rect 186 20485 294 20595
rect 0 20389 624 20437
rect 186 20265 294 20341
rect 0 20169 624 20217
rect 0 20073 624 20121
rect 186 19949 294 20025
rect 0 19853 624 19901
rect 186 19695 294 19805
rect 0 19599 624 19647
rect 186 19475 294 19551
rect 0 19379 624 19427
rect 0 19283 624 19331
rect 186 19159 294 19235
rect 0 19063 624 19111
rect 186 18905 294 19015
rect 0 18809 624 18857
rect 186 18685 294 18761
rect 0 18589 624 18637
rect 0 18493 624 18541
rect 186 18369 294 18445
rect 0 18273 624 18321
rect 186 18115 294 18225
rect 0 18019 624 18067
rect 186 17895 294 17971
rect 0 17799 624 17847
rect 0 17703 624 17751
rect 186 17579 294 17655
rect 0 17483 624 17531
rect 186 17325 294 17435
rect 0 17229 624 17277
rect 186 17105 294 17181
rect 0 17009 624 17057
rect 0 16913 624 16961
rect 186 16789 294 16865
rect 0 16693 624 16741
rect 186 16535 294 16645
rect 0 16439 624 16487
rect 186 16315 294 16391
rect 0 16219 624 16267
rect 0 16123 624 16171
rect 186 15999 294 16075
rect 0 15903 624 15951
rect 186 15745 294 15855
rect 0 15649 624 15697
rect 186 15525 294 15601
rect 0 15429 624 15477
rect 0 15333 624 15381
rect 186 15209 294 15285
rect 0 15113 624 15161
rect 186 14955 294 15065
rect 0 14859 624 14907
rect 186 14735 294 14811
rect 0 14639 624 14687
rect 0 14543 624 14591
rect 186 14419 294 14495
rect 0 14323 624 14371
rect 186 14165 294 14275
rect 0 14069 624 14117
rect 186 13945 294 14021
rect 0 13849 624 13897
rect 0 13753 624 13801
rect 186 13629 294 13705
rect 0 13533 624 13581
rect 186 13375 294 13485
rect 0 13279 624 13327
rect 186 13155 294 13231
rect 0 13059 624 13107
rect 0 12963 624 13011
rect 186 12839 294 12915
rect 0 12743 624 12791
rect 186 12585 294 12695
rect 0 12489 624 12537
rect 186 12365 294 12441
rect 0 12269 624 12317
rect 0 12173 624 12221
rect 186 12049 294 12125
rect 0 11953 624 12001
rect 186 11795 294 11905
rect 0 11699 624 11747
rect 186 11575 294 11651
rect 0 11479 624 11527
rect 0 11383 624 11431
rect 186 11259 294 11335
rect 0 11163 624 11211
rect 186 11005 294 11115
rect 0 10909 624 10957
rect 186 10785 294 10861
rect 0 10689 624 10737
rect 0 10593 624 10641
rect 186 10469 294 10545
rect 0 10373 624 10421
rect 186 10215 294 10325
rect 0 10119 624 10167
rect 186 9995 294 10071
rect 0 9899 624 9947
rect 0 9803 624 9851
rect 186 9679 294 9755
rect 0 9583 624 9631
rect 186 9425 294 9535
rect 0 9329 624 9377
rect 186 9205 294 9281
rect 0 9109 624 9157
rect 0 9013 624 9061
rect 186 8889 294 8965
rect 0 8793 624 8841
rect 186 8635 294 8745
rect 0 8539 624 8587
rect 186 8415 294 8491
rect 0 8319 624 8367
rect 0 8223 624 8271
rect 186 8099 294 8175
rect 0 8003 624 8051
rect 186 7845 294 7955
rect 0 7749 624 7797
rect 186 7625 294 7701
rect 0 7529 624 7577
rect 0 7433 624 7481
rect 186 7309 294 7385
rect 0 7213 624 7261
rect 186 7055 294 7165
rect 0 6959 624 7007
rect 186 6835 294 6911
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 186 6519 294 6595
rect 0 6423 624 6471
rect 186 6265 294 6375
rect 0 6169 624 6217
rect 186 6045 294 6121
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 186 5729 294 5805
rect 0 5633 624 5681
rect 186 5475 294 5585
rect 0 5379 624 5427
rect 186 5255 294 5331
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 186 4939 294 5015
rect 0 4843 624 4891
rect 186 4685 294 4795
rect 0 4589 624 4637
rect 186 4465 294 4541
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 186 4149 294 4225
rect 0 4053 624 4101
rect 186 3895 294 4005
rect 0 3799 624 3847
rect 186 3675 294 3751
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 186 3359 294 3435
rect 0 3263 624 3311
rect 186 3105 294 3215
rect 0 3009 624 3057
rect 186 2885 294 2961
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 186 2569 294 2645
rect 0 2473 624 2521
rect 186 2315 294 2425
rect 0 2219 624 2267
rect 186 2095 294 2171
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 186 1779 294 1855
rect 0 1683 624 1731
rect 186 1525 294 1635
rect 0 1429 624 1477
rect 186 1305 294 1381
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 186 989 294 1065
rect 0 893 624 941
rect 186 735 294 845
rect 0 639 624 687
rect 186 515 294 591
rect 0 419 624 467
rect 0 174 624 284
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_0
timestamp 1661296025
transform 1 0 0 0 -1 26860
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_1
timestamp 1661296025
transform 1 0 0 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1661296025
transform 1 0 0 0 -1 790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_0
timestamp 1661296025
transform 1 0 0 0 1 26070
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_1
timestamp 1661296025
transform 1 0 0 0 -1 26070
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_2
timestamp 1661296025
transform 1 0 0 0 1 25280
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_3
timestamp 1661296025
transform 1 0 0 0 -1 25280
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_4
timestamp 1661296025
transform 1 0 0 0 1 24490
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_5
timestamp 1661296025
transform 1 0 0 0 -1 24490
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_6
timestamp 1661296025
transform 1 0 0 0 1 23700
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_7
timestamp 1661296025
transform 1 0 0 0 -1 23700
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_8
timestamp 1661296025
transform 1 0 0 0 1 22910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_9
timestamp 1661296025
transform 1 0 0 0 -1 22910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_10
timestamp 1661296025
transform 1 0 0 0 1 22120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_11
timestamp 1661296025
transform 1 0 0 0 -1 22120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_12
timestamp 1661296025
transform 1 0 0 0 1 21330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_13
timestamp 1661296025
transform 1 0 0 0 -1 21330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_14
timestamp 1661296025
transform 1 0 0 0 1 20540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_15
timestamp 1661296025
transform 1 0 0 0 -1 20540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_16
timestamp 1661296025
transform 1 0 0 0 1 19750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_17
timestamp 1661296025
transform 1 0 0 0 -1 19750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_18
timestamp 1661296025
transform 1 0 0 0 1 18960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_19
timestamp 1661296025
transform 1 0 0 0 -1 18960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_20
timestamp 1661296025
transform 1 0 0 0 1 18170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_21
timestamp 1661296025
transform 1 0 0 0 -1 18170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_22
timestamp 1661296025
transform 1 0 0 0 1 17380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_23
timestamp 1661296025
transform 1 0 0 0 -1 17380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_24
timestamp 1661296025
transform 1 0 0 0 1 16590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_25
timestamp 1661296025
transform 1 0 0 0 -1 16590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_26
timestamp 1661296025
transform 1 0 0 0 1 15800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_27
timestamp 1661296025
transform 1 0 0 0 -1 15800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_28
timestamp 1661296025
transform 1 0 0 0 1 15010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_29
timestamp 1661296025
transform 1 0 0 0 -1 15010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_30
timestamp 1661296025
transform 1 0 0 0 1 14220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_31
timestamp 1661296025
transform 1 0 0 0 -1 14220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_32
timestamp 1661296025
transform 1 0 0 0 1 13430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_33
timestamp 1661296025
transform 1 0 0 0 -1 13430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_34
timestamp 1661296025
transform 1 0 0 0 1 12640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_35
timestamp 1661296025
transform 1 0 0 0 -1 12640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_36
timestamp 1661296025
transform 1 0 0 0 1 11850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_37
timestamp 1661296025
transform 1 0 0 0 -1 11850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_38
timestamp 1661296025
transform 1 0 0 0 1 11060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_39
timestamp 1661296025
transform 1 0 0 0 -1 11060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_40
timestamp 1661296025
transform 1 0 0 0 1 10270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_41
timestamp 1661296025
transform 1 0 0 0 -1 10270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_42
timestamp 1661296025
transform 1 0 0 0 1 9480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_43
timestamp 1661296025
transform 1 0 0 0 -1 9480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_44
timestamp 1661296025
transform 1 0 0 0 1 8690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_45
timestamp 1661296025
transform 1 0 0 0 -1 8690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_46
timestamp 1661296025
transform 1 0 0 0 1 7900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_47
timestamp 1661296025
transform 1 0 0 0 -1 7900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_48
timestamp 1661296025
transform 1 0 0 0 1 7110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_49
timestamp 1661296025
transform 1 0 0 0 -1 7110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_50
timestamp 1661296025
transform 1 0 0 0 1 6320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_51
timestamp 1661296025
transform 1 0 0 0 -1 6320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_52
timestamp 1661296025
transform 1 0 0 0 1 5530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_53
timestamp 1661296025
transform 1 0 0 0 -1 5530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_54
timestamp 1661296025
transform 1 0 0 0 1 4740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_55
timestamp 1661296025
transform 1 0 0 0 -1 4740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_56
timestamp 1661296025
transform 1 0 0 0 1 3950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_57
timestamp 1661296025
transform 1 0 0 0 -1 3950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_58
timestamp 1661296025
transform 1 0 0 0 1 3160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_59
timestamp 1661296025
transform 1 0 0 0 -1 3160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_60
timestamp 1661296025
transform 1 0 0 0 1 2370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_61
timestamp 1661296025
transform 1 0 0 0 -1 2370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_62
timestamp 1661296025
transform 1 0 0 0 1 1580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_63
timestamp 1661296025
transform 1 0 0 0 -1 1580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_64
timestamp 1661296025
transform 1 0 0 0 1 790
box -42 -105 650 424
<< labels >>
rlabel metal1 s 78 0 114 26860 4 bl_0_0
port 1 nsew
rlabel metal1 s 150 0 186 26860 4 br_0_0
port 2 nsew
rlabel metal1 s 294 0 330 26860 4 bl_1_0
port 3 nsew
rlabel metal1 s 366 0 402 26860 4 br_1_0
port 4 nsew
rlabel metal2 s 0 419 624 467 4 wl_0_0
port 5 nsew
rlabel metal2 s 0 1113 624 1161 4 wl_0_1
port 6 nsew
rlabel metal2 s 0 1209 624 1257 4 wl_0_2
port 7 nsew
rlabel metal2 s 0 1903 624 1951 4 wl_0_3
port 8 nsew
rlabel metal2 s 0 1999 624 2047 4 wl_0_4
port 9 nsew
rlabel metal2 s 0 2693 624 2741 4 wl_0_5
port 10 nsew
rlabel metal2 s 0 2789 624 2837 4 wl_0_6
port 11 nsew
rlabel metal2 s 0 3483 624 3531 4 wl_0_7
port 12 nsew
rlabel metal2 s 0 3579 624 3627 4 wl_0_8
port 13 nsew
rlabel metal2 s 0 4273 624 4321 4 wl_0_9
port 14 nsew
rlabel metal2 s 0 4369 624 4417 4 wl_0_10
port 15 nsew
rlabel metal2 s 0 5063 624 5111 4 wl_0_11
port 16 nsew
rlabel metal2 s 0 5159 624 5207 4 wl_0_12
port 17 nsew
rlabel metal2 s 0 5853 624 5901 4 wl_0_13
port 18 nsew
rlabel metal2 s 0 5949 624 5997 4 wl_0_14
port 19 nsew
rlabel metal2 s 0 6643 624 6691 4 wl_0_15
port 20 nsew
rlabel metal2 s 0 6739 624 6787 4 wl_0_16
port 21 nsew
rlabel metal2 s 0 7433 624 7481 4 wl_0_17
port 22 nsew
rlabel metal2 s 0 7529 624 7577 4 wl_0_18
port 23 nsew
rlabel metal2 s 0 8223 624 8271 4 wl_0_19
port 24 nsew
rlabel metal2 s 0 8319 624 8367 4 wl_0_20
port 25 nsew
rlabel metal2 s 0 9013 624 9061 4 wl_0_21
port 26 nsew
rlabel metal2 s 0 9109 624 9157 4 wl_0_22
port 27 nsew
rlabel metal2 s 0 9803 624 9851 4 wl_0_23
port 28 nsew
rlabel metal2 s 0 9899 624 9947 4 wl_0_24
port 29 nsew
rlabel metal2 s 0 10593 624 10641 4 wl_0_25
port 30 nsew
rlabel metal2 s 0 10689 624 10737 4 wl_0_26
port 31 nsew
rlabel metal2 s 0 11383 624 11431 4 wl_0_27
port 32 nsew
rlabel metal2 s 0 11479 624 11527 4 wl_0_28
port 33 nsew
rlabel metal2 s 0 12173 624 12221 4 wl_0_29
port 34 nsew
rlabel metal2 s 0 12269 624 12317 4 wl_0_30
port 35 nsew
rlabel metal2 s 0 12963 624 13011 4 wl_0_31
port 36 nsew
rlabel metal2 s 0 13059 624 13107 4 wl_0_32
port 37 nsew
rlabel metal2 s 0 13753 624 13801 4 wl_0_33
port 38 nsew
rlabel metal2 s 0 13849 624 13897 4 wl_0_34
port 39 nsew
rlabel metal2 s 0 14543 624 14591 4 wl_0_35
port 40 nsew
rlabel metal2 s 0 14639 624 14687 4 wl_0_36
port 41 nsew
rlabel metal2 s 0 15333 624 15381 4 wl_0_37
port 42 nsew
rlabel metal2 s 0 15429 624 15477 4 wl_0_38
port 43 nsew
rlabel metal2 s 0 16123 624 16171 4 wl_0_39
port 44 nsew
rlabel metal2 s 0 16219 624 16267 4 wl_0_40
port 45 nsew
rlabel metal2 s 0 16913 624 16961 4 wl_0_41
port 46 nsew
rlabel metal2 s 0 17009 624 17057 4 wl_0_42
port 47 nsew
rlabel metal2 s 0 17703 624 17751 4 wl_0_43
port 48 nsew
rlabel metal2 s 0 17799 624 17847 4 wl_0_44
port 49 nsew
rlabel metal2 s 0 18493 624 18541 4 wl_0_45
port 50 nsew
rlabel metal2 s 0 18589 624 18637 4 wl_0_46
port 51 nsew
rlabel metal2 s 0 19283 624 19331 4 wl_0_47
port 52 nsew
rlabel metal2 s 0 19379 624 19427 4 wl_0_48
port 53 nsew
rlabel metal2 s 0 20073 624 20121 4 wl_0_49
port 54 nsew
rlabel metal2 s 0 20169 624 20217 4 wl_0_50
port 55 nsew
rlabel metal2 s 0 20863 624 20911 4 wl_0_51
port 56 nsew
rlabel metal2 s 0 20959 624 21007 4 wl_0_52
port 57 nsew
rlabel metal2 s 0 21653 624 21701 4 wl_0_53
port 58 nsew
rlabel metal2 s 0 21749 624 21797 4 wl_0_54
port 59 nsew
rlabel metal2 s 0 22443 624 22491 4 wl_0_55
port 60 nsew
rlabel metal2 s 0 22539 624 22587 4 wl_0_56
port 61 nsew
rlabel metal2 s 0 23233 624 23281 4 wl_0_57
port 62 nsew
rlabel metal2 s 0 23329 624 23377 4 wl_0_58
port 63 nsew
rlabel metal2 s 0 24023 624 24071 4 wl_0_59
port 64 nsew
rlabel metal2 s 0 24119 624 24167 4 wl_0_60
port 65 nsew
rlabel metal2 s 0 24813 624 24861 4 wl_0_61
port 66 nsew
rlabel metal2 s 0 24909 624 24957 4 wl_0_62
port 67 nsew
rlabel metal2 s 0 25603 624 25651 4 wl_0_63
port 68 nsew
rlabel metal2 s 0 25699 624 25747 4 wl_0_64
port 69 nsew
rlabel metal2 s 0 26393 624 26441 4 wl_0_65
port 70 nsew
rlabel metal2 s 0 639 624 687 4 wl_1_0
port 71 nsew
rlabel metal2 s 0 893 624 941 4 wl_1_1
port 72 nsew
rlabel metal2 s 0 1429 624 1477 4 wl_1_2
port 73 nsew
rlabel metal2 s 0 1683 624 1731 4 wl_1_3
port 74 nsew
rlabel metal2 s 0 2219 624 2267 4 wl_1_4
port 75 nsew
rlabel metal2 s 0 2473 624 2521 4 wl_1_5
port 76 nsew
rlabel metal2 s 0 3009 624 3057 4 wl_1_6
port 77 nsew
rlabel metal2 s 0 3263 624 3311 4 wl_1_7
port 78 nsew
rlabel metal2 s 0 3799 624 3847 4 wl_1_8
port 79 nsew
rlabel metal2 s 0 4053 624 4101 4 wl_1_9
port 80 nsew
rlabel metal2 s 0 4589 624 4637 4 wl_1_10
port 81 nsew
rlabel metal2 s 0 4843 624 4891 4 wl_1_11
port 82 nsew
rlabel metal2 s 0 5379 624 5427 4 wl_1_12
port 83 nsew
rlabel metal2 s 0 5633 624 5681 4 wl_1_13
port 84 nsew
rlabel metal2 s 0 6169 624 6217 4 wl_1_14
port 85 nsew
rlabel metal2 s 0 6423 624 6471 4 wl_1_15
port 86 nsew
rlabel metal2 s 0 6959 624 7007 4 wl_1_16
port 87 nsew
rlabel metal2 s 0 7213 624 7261 4 wl_1_17
port 88 nsew
rlabel metal2 s 0 7749 624 7797 4 wl_1_18
port 89 nsew
rlabel metal2 s 0 8003 624 8051 4 wl_1_19
port 90 nsew
rlabel metal2 s 0 8539 624 8587 4 wl_1_20
port 91 nsew
rlabel metal2 s 0 8793 624 8841 4 wl_1_21
port 92 nsew
rlabel metal2 s 0 9329 624 9377 4 wl_1_22
port 93 nsew
rlabel metal2 s 0 9583 624 9631 4 wl_1_23
port 94 nsew
rlabel metal2 s 0 10119 624 10167 4 wl_1_24
port 95 nsew
rlabel metal2 s 0 10373 624 10421 4 wl_1_25
port 96 nsew
rlabel metal2 s 0 10909 624 10957 4 wl_1_26
port 97 nsew
rlabel metal2 s 0 11163 624 11211 4 wl_1_27
port 98 nsew
rlabel metal2 s 0 11699 624 11747 4 wl_1_28
port 99 nsew
rlabel metal2 s 0 11953 624 12001 4 wl_1_29
port 100 nsew
rlabel metal2 s 0 12489 624 12537 4 wl_1_30
port 101 nsew
rlabel metal2 s 0 12743 624 12791 4 wl_1_31
port 102 nsew
rlabel metal2 s 0 13279 624 13327 4 wl_1_32
port 103 nsew
rlabel metal2 s 0 13533 624 13581 4 wl_1_33
port 104 nsew
rlabel metal2 s 0 14069 624 14117 4 wl_1_34
port 105 nsew
rlabel metal2 s 0 14323 624 14371 4 wl_1_35
port 106 nsew
rlabel metal2 s 0 14859 624 14907 4 wl_1_36
port 107 nsew
rlabel metal2 s 0 15113 624 15161 4 wl_1_37
port 108 nsew
rlabel metal2 s 0 15649 624 15697 4 wl_1_38
port 109 nsew
rlabel metal2 s 0 15903 624 15951 4 wl_1_39
port 110 nsew
rlabel metal2 s 0 16439 624 16487 4 wl_1_40
port 111 nsew
rlabel metal2 s 0 16693 624 16741 4 wl_1_41
port 112 nsew
rlabel metal2 s 0 17229 624 17277 4 wl_1_42
port 113 nsew
rlabel metal2 s 0 17483 624 17531 4 wl_1_43
port 114 nsew
rlabel metal2 s 0 18019 624 18067 4 wl_1_44
port 115 nsew
rlabel metal2 s 0 18273 624 18321 4 wl_1_45
port 116 nsew
rlabel metal2 s 0 18809 624 18857 4 wl_1_46
port 117 nsew
rlabel metal2 s 0 19063 624 19111 4 wl_1_47
port 118 nsew
rlabel metal2 s 0 19599 624 19647 4 wl_1_48
port 119 nsew
rlabel metal2 s 0 19853 624 19901 4 wl_1_49
port 120 nsew
rlabel metal2 s 0 20389 624 20437 4 wl_1_50
port 121 nsew
rlabel metal2 s 0 20643 624 20691 4 wl_1_51
port 122 nsew
rlabel metal2 s 0 21179 624 21227 4 wl_1_52
port 123 nsew
rlabel metal2 s 0 21433 624 21481 4 wl_1_53
port 124 nsew
rlabel metal2 s 0 21969 624 22017 4 wl_1_54
port 125 nsew
rlabel metal2 s 0 22223 624 22271 4 wl_1_55
port 126 nsew
rlabel metal2 s 0 22759 624 22807 4 wl_1_56
port 127 nsew
rlabel metal2 s 0 23013 624 23061 4 wl_1_57
port 128 nsew
rlabel metal2 s 0 23549 624 23597 4 wl_1_58
port 129 nsew
rlabel metal2 s 0 23803 624 23851 4 wl_1_59
port 130 nsew
rlabel metal2 s 0 24339 624 24387 4 wl_1_60
port 131 nsew
rlabel metal2 s 0 24593 624 24641 4 wl_1_61
port 132 nsew
rlabel metal2 s 0 25129 624 25177 4 wl_1_62
port 133 nsew
rlabel metal2 s 0 25383 624 25431 4 wl_1_63
port 134 nsew
rlabel metal2 s 0 25919 624 25967 4 wl_1_64
port 135 nsew
rlabel metal2 s 0 26173 624 26221 4 wl_1_65
port 136 nsew
rlabel metal1 s 222 14590 258 14931 4 vdd
port 137 nsew
rlabel metal1 s 222 10640 258 10981 4 vdd
port 137 nsew
rlabel metal1 s 222 22490 258 22831 4 vdd
port 137 nsew
rlabel metal2 s 0 174 624 284 4 vdd
port 137 nsew
rlabel metal1 s 222 18249 258 18590 4 vdd
port 137 nsew
rlabel metal1 s 222 20120 258 20461 4 vdd
port 137 nsew
rlabel metal1 s 222 6399 258 6740 4 vdd
port 137 nsew
rlabel metal1 s 222 9060 258 9401 4 vdd
port 137 nsew
rlabel metal1 s 222 12220 258 12561 4 vdd
port 137 nsew
rlabel metal1 s 222 3530 258 3871 4 vdd
port 137 nsew
rlabel metal1 s 222 24569 258 24910 4 vdd
port 137 nsew
rlabel metal1 s 222 8769 258 9110 4 vdd
port 137 nsew
rlabel metal1 s 222 13509 258 13850 4 vdd
port 137 nsew
rlabel metal1 s 222 15089 258 15430 4 vdd
port 137 nsew
rlabel metal1 s 222 22199 258 22540 4 vdd
port 137 nsew
rlabel metal1 s 222 21409 258 21750 4 vdd
port 137 nsew
rlabel metal1 s 222 16669 258 17010 4 vdd
port 137 nsew
rlabel metal1 s 222 1659 258 2000 4 vdd
port 137 nsew
rlabel metal1 s 222 2449 258 2790 4 vdd
port 137 nsew
rlabel metal1 s 222 11430 258 11771 4 vdd
port 137 nsew
rlabel metal1 s 222 16170 258 16511 4 vdd
port 137 nsew
rlabel metal1 s 222 11139 258 11480 4 vdd
port 137 nsew
rlabel metal1 s 222 17459 258 17800 4 vdd
port 137 nsew
rlabel metal1 s 222 7189 258 7530 4 vdd
port 137 nsew
rlabel metal1 s 222 9850 258 10191 4 vdd
port 137 nsew
rlabel metal1 s 222 6690 258 7031 4 vdd
port 137 nsew
rlabel metal1 s 222 18540 258 18881 4 vdd
port 137 nsew
rlabel metal1 s 222 24070 258 24411 4 vdd
port 137 nsew
rlabel metal1 s 222 25650 258 25991 4 vdd
port 137 nsew
rlabel metal1 s 222 7480 258 7821 4 vdd
port 137 nsew
rlabel metal1 s 222 19039 258 19380 4 vdd
port 137 nsew
rlabel metal1 s 222 7979 258 8320 4 vdd
port 137 nsew
rlabel metal1 s 222 12719 258 13060 4 vdd
port 137 nsew
rlabel metal1 s 222 22989 258 23330 4 vdd
port 137 nsew
rlabel metal1 s 222 23779 258 24120 4 vdd
port 137 nsew
rlabel metal1 s 222 5609 258 5950 4 vdd
port 137 nsew
rlabel metal1 s 222 5900 258 6241 4 vdd
port 137 nsew
rlabel metal1 s 222 8270 258 8611 4 vdd
port 137 nsew
rlabel metal1 s 222 4320 258 4661 4 vdd
port 137 nsew
rlabel metal1 s 222 4819 258 5160 4 vdd
port 137 nsew
rlabel metal1 s 222 10349 258 10690 4 vdd
port 137 nsew
rlabel metal1 s 222 13800 258 14141 4 vdd
port 137 nsew
rlabel metal1 s 222 15380 258 15721 4 vdd
port 137 nsew
rlabel metal1 s 222 15879 258 16220 4 vdd
port 137 nsew
rlabel metal1 s 222 25359 258 25700 4 vdd
port 137 nsew
rlabel metal1 s 222 24860 258 25201 4 vdd
port 137 nsew
rlabel metal2 s 0 26576 624 26686 4 vdd
port 137 nsew
rlabel metal1 s 222 4029 258 4370 4 vdd
port 137 nsew
rlabel metal1 s 222 21700 258 22041 4 vdd
port 137 nsew
rlabel metal1 s 222 26149 258 26490 4 vdd
port 137 nsew
rlabel metal1 s 222 2740 258 3081 4 vdd
port 137 nsew
rlabel metal1 s 222 11929 258 12270 4 vdd
port 137 nsew
rlabel metal1 s 222 19829 258 20170 4 vdd
port 137 nsew
rlabel metal1 s 222 9559 258 9900 4 vdd
port 137 nsew
rlabel metal1 s 222 370 258 711 4 vdd
port 137 nsew
rlabel metal1 s 222 13010 258 13351 4 vdd
port 137 nsew
rlabel metal1 s 222 16960 258 17301 4 vdd
port 137 nsew
rlabel metal1 s 222 19330 258 19671 4 vdd
port 137 nsew
rlabel metal1 s 222 17750 258 18091 4 vdd
port 137 nsew
rlabel metal1 s 222 20619 258 20960 4 vdd
port 137 nsew
rlabel metal1 s 222 20910 258 21251 4 vdd
port 137 nsew
rlabel metal1 s 222 23280 258 23621 4 vdd
port 137 nsew
rlabel metal1 s 222 14299 258 14640 4 vdd
port 137 nsew
rlabel metal1 s 222 1950 258 2291 4 vdd
port 137 nsew
rlabel metal1 s 222 1160 258 1501 4 vdd
port 137 nsew
rlabel metal1 s 222 869 258 1210 4 vdd
port 137 nsew
rlabel metal1 s 222 5110 258 5451 4 vdd
port 137 nsew
rlabel metal1 s 222 3239 258 3580 4 vdd
port 137 nsew
rlabel metal2 s 186 9995 294 10071 4 gnd
port 138 nsew
rlabel metal2 s 186 1305 294 1381 4 gnd
port 138 nsew
rlabel metal2 s 186 23425 294 23501 4 gnd
port 138 nsew
rlabel metal2 s 186 15209 294 15285 4 gnd
port 138 nsew
rlabel metal2 s 186 20739 294 20815 4 gnd
port 138 nsew
rlabel metal2 s 186 14735 294 14811 4 gnd
port 138 nsew
rlabel metal2 s 186 5475 294 5585 4 gnd
port 138 nsew
rlabel metal2 s 186 22065 294 22175 4 gnd
port 138 nsew
rlabel metal2 s 186 10785 294 10861 4 gnd
port 138 nsew
rlabel metal2 s 186 12365 294 12441 4 gnd
port 138 nsew
rlabel metal2 s 186 2569 294 2645 4 gnd
port 138 nsew
rlabel metal2 s 186 5255 294 5331 4 gnd
port 138 nsew
rlabel metal2 s 186 26015 294 26125 4 gnd
port 138 nsew
rlabel metal2 s 186 11575 294 11651 4 gnd
port 138 nsew
rlabel metal2 s 186 26269 294 26345 4 gnd
port 138 nsew
rlabel metal2 s 186 18685 294 18761 4 gnd
port 138 nsew
rlabel metal2 s 186 25005 294 25081 4 gnd
port 138 nsew
rlabel metal2 s 186 12585 294 12695 4 gnd
port 138 nsew
rlabel metal2 s 186 13375 294 13485 4 gnd
port 138 nsew
rlabel metal2 s 186 18905 294 19015 4 gnd
port 138 nsew
rlabel metal2 s 186 735 294 845 4 gnd
port 138 nsew
rlabel metal2 s 186 17895 294 17971 4 gnd
port 138 nsew
rlabel metal2 s 186 22635 294 22711 4 gnd
port 138 nsew
rlabel metal2 s 186 10215 294 10325 4 gnd
port 138 nsew
rlabel metal2 s 186 7845 294 7955 4 gnd
port 138 nsew
rlabel metal2 s 186 8415 294 8491 4 gnd
port 138 nsew
rlabel metal2 s 186 9425 294 9535 4 gnd
port 138 nsew
rlabel metal2 s 186 6519 294 6595 4 gnd
port 138 nsew
rlabel metal2 s 186 8099 294 8175 4 gnd
port 138 nsew
rlabel metal2 s 186 8635 294 8745 4 gnd
port 138 nsew
rlabel metal2 s 186 24215 294 24291 4 gnd
port 138 nsew
rlabel metal2 s 186 22855 294 22965 4 gnd
port 138 nsew
rlabel metal2 s 186 25479 294 25555 4 gnd
port 138 nsew
rlabel metal2 s 186 21529 294 21605 4 gnd
port 138 nsew
rlabel metal2 s 186 19159 294 19235 4 gnd
port 138 nsew
rlabel metal2 s 186 11259 294 11335 4 gnd
port 138 nsew
rlabel metal2 s 186 23899 294 23975 4 gnd
port 138 nsew
rlabel metal2 s 186 25225 294 25335 4 gnd
port 138 nsew
rlabel metal2 s 186 16789 294 16865 4 gnd
port 138 nsew
rlabel metal2 s 186 4465 294 4541 4 gnd
port 138 nsew
rlabel metal2 s 186 8889 294 8965 4 gnd
port 138 nsew
rlabel metal2 s 186 4939 294 5015 4 gnd
port 138 nsew
rlabel metal2 s 186 24435 294 24545 4 gnd
port 138 nsew
rlabel metal2 s 186 6265 294 6375 4 gnd
port 138 nsew
rlabel metal2 s 186 17325 294 17435 4 gnd
port 138 nsew
rlabel metal2 s 186 23645 294 23755 4 gnd
port 138 nsew
rlabel metal2 s 186 15745 294 15855 4 gnd
port 138 nsew
rlabel metal2 s 186 11795 294 11905 4 gnd
port 138 nsew
rlabel metal2 s 186 515 294 591 4 gnd
port 138 nsew
rlabel metal2 s 186 7625 294 7701 4 gnd
port 138 nsew
rlabel metal2 s 186 21275 294 21385 4 gnd
port 138 nsew
rlabel metal2 s 186 9205 294 9281 4 gnd
port 138 nsew
rlabel metal2 s 186 2095 294 2171 4 gnd
port 138 nsew
rlabel metal2 s 186 12049 294 12125 4 gnd
port 138 nsew
rlabel metal2 s 186 3105 294 3215 4 gnd
port 138 nsew
rlabel metal2 s 186 4685 294 4795 4 gnd
port 138 nsew
rlabel metal2 s 186 18115 294 18225 4 gnd
port 138 nsew
rlabel metal2 s 186 10469 294 10545 4 gnd
port 138 nsew
rlabel metal2 s 186 18369 294 18445 4 gnd
port 138 nsew
rlabel metal2 s 186 1779 294 1855 4 gnd
port 138 nsew
rlabel metal2 s 186 17105 294 17181 4 gnd
port 138 nsew
rlabel metal2 s 186 13629 294 13705 4 gnd
port 138 nsew
rlabel metal2 s 186 24689 294 24765 4 gnd
port 138 nsew
rlabel metal2 s 186 3359 294 3435 4 gnd
port 138 nsew
rlabel metal2 s 186 21845 294 21921 4 gnd
port 138 nsew
rlabel metal2 s 186 1525 294 1635 4 gnd
port 138 nsew
rlabel metal2 s 186 19949 294 20025 4 gnd
port 138 nsew
rlabel metal2 s 186 22319 294 22395 4 gnd
port 138 nsew
rlabel metal2 s 186 20485 294 20595 4 gnd
port 138 nsew
rlabel metal2 s 186 4149 294 4225 4 gnd
port 138 nsew
rlabel metal2 s 186 6835 294 6911 4 gnd
port 138 nsew
rlabel metal2 s 186 9679 294 9755 4 gnd
port 138 nsew
rlabel metal2 s 186 13155 294 13231 4 gnd
port 138 nsew
rlabel metal2 s 186 14419 294 14495 4 gnd
port 138 nsew
rlabel metal2 s 186 5729 294 5805 4 gnd
port 138 nsew
rlabel metal2 s 186 13945 294 14021 4 gnd
port 138 nsew
rlabel metal2 s 186 14165 294 14275 4 gnd
port 138 nsew
rlabel metal2 s 186 21055 294 21131 4 gnd
port 138 nsew
rlabel metal2 s 186 25795 294 25871 4 gnd
port 138 nsew
rlabel metal2 s 186 23109 294 23185 4 gnd
port 138 nsew
rlabel metal2 s 186 14955 294 15065 4 gnd
port 138 nsew
rlabel metal2 s 186 19695 294 19805 4 gnd
port 138 nsew
rlabel metal2 s 186 15999 294 16075 4 gnd
port 138 nsew
rlabel metal2 s 186 7309 294 7385 4 gnd
port 138 nsew
rlabel metal2 s 186 11005 294 11115 4 gnd
port 138 nsew
rlabel metal2 s 186 7055 294 7165 4 gnd
port 138 nsew
rlabel metal2 s 186 19475 294 19551 4 gnd
port 138 nsew
rlabel metal2 s 186 3895 294 4005 4 gnd
port 138 nsew
rlabel metal2 s 186 6045 294 6121 4 gnd
port 138 nsew
rlabel metal2 s 186 16535 294 16645 4 gnd
port 138 nsew
rlabel metal2 s 186 17579 294 17655 4 gnd
port 138 nsew
rlabel metal2 s 186 989 294 1065 4 gnd
port 138 nsew
rlabel metal2 s 186 2885 294 2961 4 gnd
port 138 nsew
rlabel metal2 s 186 15525 294 15601 4 gnd
port 138 nsew
rlabel metal2 s 186 3675 294 3751 4 gnd
port 138 nsew
rlabel metal2 s 186 20265 294 20341 4 gnd
port 138 nsew
rlabel metal2 s 186 12839 294 12915 4 gnd
port 138 nsew
rlabel metal2 s 186 16315 294 16391 4 gnd
port 138 nsew
rlabel metal2 s 186 2315 294 2425 4 gnd
port 138 nsew
<< properties >>
string FIXED_BBOX 0 0 624 26860
<< end >>
