magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< nwell >>
rect -54 -54 204 278
<< scpmos >>
rect 60 0 90 224
<< pdiff >>
rect 0 0 60 224
rect 90 0 150 224
<< poly >>
rect 60 224 90 250
rect 60 -26 90 0
<< locali >>
rect 8 79 42 145
rect 108 79 142 145
use sky130_sram_1r1w_24x128_8_contact_11  sky130_sram_1r1w_24x128_8_contact_11_0
timestamp 1661296025
transform 1 0 100 0 1 79
box -59 -51 109 117
use sky130_sram_1r1w_24x128_8_contact_11  sky130_sram_1r1w_24x128_8_contact_11_1
timestamp 1661296025
transform 1 0 0 0 1 79
box -59 -51 109 117
<< labels >>
rlabel poly s 75 112 75 112 4 G
port 1 nsew
rlabel locali s 25 112 25 112 4 S
port 2 nsew
rlabel locali s 125 112 125 112 4 D
port 3 nsew
<< properties >>
string FIXED_BBOX -54 -54 204 278
<< end >>
