magic
tech sky130B
magscale 1 2
timestamp 1662225218
<< metal4 >>
rect -17000 400 -10000 500
rect -17000 -1900 -12000 400
rect -10100 -1900 -10000 400
rect -17000 -2000 -10000 -1900
<< via4 >>
rect -12000 -1900 -10100 400
<< metal5 >>
tri -13852 6000 -11852 8000 se
rect -11852 6000 9252 8000
tri 9252 6000 11252 8000 sw
tri -15300 4552 -13852 6000 se
rect -13852 5400 -11624 6000
tri -11624 5400 -11024 6000 nw
tri 8424 5400 9024 6000 ne
rect 9024 5400 11252 6000
rect -13852 4552 -12473 5400
tri -15528 4324 -15300 4552 se
rect -15300 4551 -12473 4552
tri -12473 4551 -11624 5400 nw
tri -11624 4551 -10775 5400 se
rect -10775 4551 8175 5400
tri 8175 4551 9024 5400 sw
tri 9024 4551 9873 5400 ne
rect 9873 4551 11252 5400
rect -15300 4324 -12700 4551
tri -12700 4324 -12473 4551 nw
tri -11851 4324 -11624 4551 se
rect -11624 4324 9024 4551
tri -17300 2552 -15528 4324 se
rect -15528 3475 -13549 4324
tri -13549 3475 -12700 4324 nw
tri -12700 3475 -11851 4324 se
rect -11851 4249 9024 4324
tri 9024 4249 9326 4551 sw
tri 9873 4249 10175 4551 ne
rect 10175 4249 11252 4551
rect -11851 3475 9326 4249
rect -15528 3247 -13777 3475
tri -13777 3247 -13549 3475 nw
tri -12928 3247 -12700 3475 se
rect -12700 3400 9326 3475
tri 9326 3400 10175 4249 sw
tri 10175 3400 11024 4249 ne
rect 11024 3400 11252 4249
tri 11252 3400 13852 6000 sw
rect -15528 2552 -14626 3247
rect -17300 2398 -14626 2552
tri -14626 2398 -13777 3247 nw
tri -13777 2398 -12928 3247 se
rect -12928 2398 -12700 3247
rect -17300 1500 -15300 2398
tri -15300 1724 -14626 2398 nw
tri -14451 1724 -13777 2398 se
rect -13777 1724 -12700 2398
tri -14700 1475 -14451 1724 se
rect -14451 1475 -12700 1724
rect -14700 -3085 -12700 1475
tri -12700 647 -9947 3400 nw
tri 7347 647 10100 3400 ne
rect 10100 2551 10175 3400
tri 10175 2551 11024 3400 sw
tri 11024 2551 11873 3400 ne
rect 11873 2552 13852 3400
tri 13852 2552 14700 3400 sw
rect 11873 2551 14700 2552
rect 10100 1724 11024 2551
tri 11024 1724 11851 2551 sw
tri 11873 1724 12700 2551 ne
rect 10100 1475 11851 1724
tri 11851 1475 12100 1724 sw
tri -12100 398 -12000 498 se
rect -12000 400 -10000 500
rect -12100 -1900 -12000 398
rect -10100 -1900 -10000 400
rect -12100 -2237 -10000 -1900
tri -12700 -3085 -12100 -2485 sw
tri -12100 -3085 -11252 -2237 ne
rect -11252 -3085 -10000 -2237
rect -14700 -3314 -12100 -3085
tri -14700 -3400 -14614 -3314 ne
rect -14614 -3400 -12100 -3314
tri -12100 -3400 -11785 -3085 sw
tri -11252 -3400 -10937 -3085 ne
rect -10937 -3400 -10000 -3085
tri -10000 -3400 -8108 -1508 sw
tri 8108 -3400 10100 -1408 se
rect 10100 -2237 12100 1475
rect 10100 -3085 11252 -2237
tri 11252 -3085 12100 -2237 nw
tri 12100 -3085 12700 -2485 se
rect 12700 -3085 14700 2551
rect 10100 -3400 10937 -3085
tri 10937 -3400 11252 -3085 nw
tri 11785 -3400 12100 -3085 se
rect 12100 -3314 14700 -3085
rect 12100 -3400 12700 -3314
tri -14614 -6000 -12014 -3400 ne
rect -12014 -4248 -11785 -3400
tri -11785 -4248 -10937 -3400 sw
tri -10937 -4248 -10089 -3400 ne
rect -10089 -4237 10100 -3400
tri 10100 -4237 10937 -3400 nw
tri 10948 -4237 11785 -3400 se
rect 11785 -4237 12700 -3400
rect -10089 -4248 9252 -4237
rect -12014 -4552 -10937 -4248
tri -10937 -4552 -10633 -4248 sw
tri -10089 -4552 -9785 -4248 ne
rect -9785 -4552 9252 -4248
rect -12014 -5400 -10633 -4552
tri -10633 -5400 -9785 -4552 sw
tri -9785 -5400 -8937 -4552 ne
rect -8937 -5085 9252 -4552
tri 9252 -5085 10100 -4237 nw
tri 10100 -5085 10948 -4237 se
rect 10948 -5085 12700 -4237
rect -8937 -5400 8937 -5085
tri 8937 -5400 9252 -5085 nw
tri 9785 -5400 10100 -5085 se
rect 10100 -5314 12700 -5085
tri 12700 -5314 14700 -3314 nw
rect -12014 -6000 -9785 -5400
tri -9785 -6000 -9185 -5400 sw
tri 9185 -6000 9785 -5400 se
rect 9785 -6000 10100 -5400
tri -12014 -8000 -10014 -6000 ne
rect -10014 -7914 10100 -6000
tri 10100 -7914 12700 -5314 nw
rect -10014 -8000 10014 -7914
tri 10014 -8000 10100 -7914 nw
<< end >>
