magic
tech sky130B
magscale 1 2
timestamp 1660789662
<< pwell >>
rect 2400 100 3014 1146
<< locali >>
rect 2880 980 2960 990
rect 2880 920 2890 980
rect 2950 920 2960 980
rect 2880 910 2960 920
rect 2660 330 2740 340
rect 2660 270 2670 330
rect 2730 270 2740 330
rect 2660 260 2740 270
<< viali >>
rect 2540 1080 3080 1120
rect 2890 920 2950 980
rect 2670 270 2730 330
<< metal1 >>
rect -100 1400 3100 1500
rect 2500 1120 3100 1400
rect 2500 1080 2540 1120
rect 3080 1080 3100 1120
rect 2500 1060 3100 1080
rect 2870 990 2970 1000
rect 2870 910 2880 990
rect 2960 910 2970 990
rect 2870 900 2970 910
rect 2650 340 2750 350
rect 2650 260 2660 340
rect 2740 260 2750 340
rect 2650 250 2750 260
<< via1 >>
rect 2880 980 2960 990
rect 2880 920 2890 980
rect 2890 920 2950 980
rect 2950 920 2960 980
rect 2880 910 2960 920
rect 2660 330 2740 340
rect 2660 270 2670 330
rect 2670 270 2730 330
rect 2730 270 2740 330
rect 2660 260 2740 270
<< metal2 >>
rect -100 1400 2600 1500
rect -100 700 100 1400
rect 2400 700 2600 1400
rect 2770 990 2970 1000
rect 2770 910 2780 990
rect 2960 910 2970 990
rect 2770 900 2970 910
rect 2650 340 2850 350
rect 2650 260 2660 340
rect 2840 260 2850 340
rect 2650 250 2850 260
<< via2 >>
rect 2780 910 2880 990
rect 2880 910 2960 990
rect 980 220 1460 500
rect 2660 260 2740 340
rect 2740 260 2840 340
<< metal3 >>
rect 2420 990 2970 1100
rect 2420 910 2780 990
rect 2960 910 2970 990
rect 2420 900 2970 910
rect -650 530 500 790
rect 2420 760 2570 900
rect 2050 540 2570 760
rect 960 500 1520 540
rect 960 220 980 500
rect 1460 220 1520 500
rect 960 180 1520 220
rect 2650 340 2850 350
rect 2650 160 2660 340
rect 2840 160 2850 340
rect 2650 150 2850 160
<< via3 >>
rect 980 220 1460 500
rect 2660 260 2840 340
rect 2660 160 2840 260
<< metal4 >>
rect 960 500 2000 551
rect 960 220 980 500
rect 1460 220 2000 500
rect 960 30 2000 220
rect 600 -80 2000 30
rect 2650 340 2850 350
rect 2650 160 2660 340
rect 2840 160 2850 340
rect 2650 -80 2850 160
rect 600 -610 3840 -80
rect 600 -800 2000 -610
use RF_nfet_6xaM02W5p0L0p15  RF_nfet_6xaM02W5p0L0p15_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660736647
transform 1 0 0 0 1 0
box 0 0 2474 1440
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660275339
transform 1 0 -200 0 1 2600
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_1
timestamp 1660275339
transform 1 0 300 0 1 2600
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_2
timestamp 1660275339
transform 1 0 800 0 1 2600
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_3
timestamp 1660275339
transform 1 0 1300 0 1 2600
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_4
timestamp 1660275339
transform 1 0 1800 0 1 2600
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_5
timestamp 1660275339
transform 1 0 2300 0 1 2600
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_6
timestamp 1660275339
transform 1 0 -700 0 1 2600
box 100 -1100 600 -600
use sky130_fd_pr__res_generic_po_JFYRVD  sky130_fd_pr__res_generic_po_JFYRVD_0
timestamp 1659754026
transform 1 0 2807 0 1 623
box -307 -523 307 523
<< labels >>
rlabel metal4 600 -800 2000 -10 1 NDRAIN
rlabel metal3 -650 530 -300 790 1 NGATE
rlabel space -100 1390 2610 1500 1 NSOURCE
<< end >>
