magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< locali >>
rect 2583 1443 3160 1477
rect 174 1372 1662 1406
rect 94 1264 1662 1298
rect 1156 1072 1662 1106
rect 1396 964 1662 998
rect 2583 893 3160 927
rect 2583 653 3160 687
rect 174 603 414 637
rect 1236 582 1662 616
rect 1316 474 1662 508
rect 1156 282 1662 316
rect 94 153 414 187
rect 1236 174 1662 208
rect 2583 103 3160 137
<< metal1 >>
rect 80 199 108 1580
rect 160 649 188 1580
rect 151 591 197 649
rect 71 141 117 199
rect 80 80 108 141
rect 160 80 188 591
rect 504 421 532 790
rect 900 421 928 790
rect 1030 644 1094 696
rect 486 369 550 421
rect 882 369 946 421
rect 504 80 532 369
rect 900 80 928 369
rect 1030 94 1094 146
rect 1142 80 1170 1580
rect 1222 80 1250 1580
rect 1302 80 1330 1580
rect 1382 80 1410 1580
rect 1788 1218 1836 1610
rect 2212 1218 2262 1612
rect 1780 1166 1844 1218
rect 2205 1166 2269 1218
rect 2602 1211 2630 1580
rect 2998 1211 3026 1580
rect 1788 428 1836 1166
rect 2212 428 2262 1166
rect 2584 1159 2648 1211
rect 2980 1159 3044 1211
rect 1780 376 1844 428
rect 2205 376 2269 428
rect 2602 421 2630 1159
rect 2998 421 3026 1159
rect 1788 80 1836 376
rect 2212 80 2262 376
rect 2584 369 2648 421
rect 2980 369 3044 421
rect 2602 80 2630 369
rect 2998 80 3026 369
<< metal2 >>
rect 1784 1168 1840 1216
rect 2209 1168 2265 1216
rect 2588 1161 2644 1209
rect 2984 1161 3040 1209
rect 1048 692 1236 720
rect 1048 670 1076 692
rect 490 371 546 419
rect 886 371 942 419
rect 1784 378 1840 426
rect 2209 378 2265 426
rect 2588 371 2644 419
rect 2984 371 3040 419
rect 1048 297 1156 325
rect 1048 120 1076 297
<< metal3 >>
rect 1763 1143 1861 1241
rect 2188 1143 2286 1241
rect 2567 1136 2665 1234
rect 2963 1136 3061 1234
rect 469 346 567 444
rect 865 346 963 444
rect 1763 353 1861 451
rect 2188 353 2286 451
rect 2567 346 2665 444
rect 2963 346 3061 444
use sky130_sram_1r1w_24x128_8_and2_dec  sky130_sram_1r1w_24x128_8_and2_dec_0
timestamp 1661296025
transform 1 0 1542 0 -1 1580
box 70 -56 1636 490
use sky130_sram_1r1w_24x128_8_and2_dec  sky130_sram_1r1w_24x128_8_and2_dec_1
timestamp 1661296025
transform 1 0 1542 0 1 790
box 70 -56 1636 490
use sky130_sram_1r1w_24x128_8_and2_dec  sky130_sram_1r1w_24x128_8_and2_dec_2
timestamp 1661296025
transform 1 0 1542 0 -1 790
box 70 -56 1636 490
use sky130_sram_1r1w_24x128_8_and2_dec  sky130_sram_1r1w_24x128_8_and2_dec_3
timestamp 1661296025
transform 1 0 1542 0 1 0
box 70 -56 1636 490
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 1033 0 1 637
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 1033 0 1 87
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_0
timestamp 1661296025
transform 1 0 1363 0 1 1360
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_1
timestamp 1661296025
transform 1 0 1283 0 1 1252
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_2
timestamp 1661296025
transform 1 0 1363 0 1 952
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_3
timestamp 1661296025
transform 1 0 1123 0 1 1060
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_4
timestamp 1661296025
transform 1 0 1203 0 1 570
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_5
timestamp 1661296025
transform 1 0 1283 0 1 462
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_6
timestamp 1661296025
transform 1 0 1203 0 1 162
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_7
timestamp 1661296025
transform 1 0 1123 0 1 270
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_8
timestamp 1661296025
transform 1 0 141 0 1 591
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_16  sky130_sram_1r1w_24x128_8_contact_16_9
timestamp 1661296025
transform 1 0 61 0 1 141
box 0 0 66 58
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_0
timestamp 1661296025
transform 1 0 2584 0 1 1153
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_1
timestamp 1661296025
transform 1 0 1780 0 1 1160
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_2
timestamp 1661296025
transform 1 0 2584 0 1 363
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_3
timestamp 1661296025
transform 1 0 1780 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_4
timestamp 1661296025
transform 1 0 486 0 1 363
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_5
timestamp 1661296025
transform 1 0 486 0 1 363
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_6
timestamp 1661296025
transform 1 0 2205 0 1 1160
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_7
timestamp 1661296025
transform 1 0 2980 0 1 1153
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_8
timestamp 1661296025
transform 1 0 2205 0 1 370
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_9
timestamp 1661296025
transform 1 0 2980 0 1 363
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_10
timestamp 1661296025
transform 1 0 882 0 1 363
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_11
timestamp 1661296025
transform 1 0 882 0 1 363
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_12
timestamp 1661296025
transform 1 0 1030 0 1 638
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_13
timestamp 1661296025
transform 1 0 1030 0 1 88
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_0
timestamp 1661296025
transform 1 0 1204 0 1 674
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_19  sky130_sram_1r1w_24x128_8_contact_19_1
timestamp 1661296025
transform 1 0 1124 0 1 279
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_20  sky130_sram_1r1w_24x128_8_contact_20_0
timestamp 1661296025
transform 1 0 1363 0 1 1366
box 0 0 66 46
use sky130_sram_1r1w_24x128_8_contact_20  sky130_sram_1r1w_24x128_8_contact_20_1
timestamp 1661296025
transform 1 0 141 0 1 1366
box 0 0 66 46
use sky130_sram_1r1w_24x128_8_contact_20  sky130_sram_1r1w_24x128_8_contact_20_2
timestamp 1661296025
transform 1 0 1283 0 1 1258
box 0 0 66 46
use sky130_sram_1r1w_24x128_8_contact_20  sky130_sram_1r1w_24x128_8_contact_20_3
timestamp 1661296025
transform 1 0 61 0 1 1258
box 0 0 66 46
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_0
timestamp 1661296025
transform 1 0 2583 0 1 1148
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_1
timestamp 1661296025
transform 1 0 1779 0 1 1155
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_2
timestamp 1661296025
transform 1 0 2583 0 1 358
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_3
timestamp 1661296025
transform 1 0 1779 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_4
timestamp 1661296025
transform 1 0 485 0 1 358
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_5
timestamp 1661296025
transform 1 0 485 0 1 358
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_6
timestamp 1661296025
transform 1 0 2204 0 1 1155
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_7
timestamp 1661296025
transform 1 0 2979 0 1 1148
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_8
timestamp 1661296025
transform 1 0 2204 0 1 365
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_9
timestamp 1661296025
transform 1 0 2979 0 1 358
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_10
timestamp 1661296025
transform 1 0 881 0 1 358
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_11
timestamp 1661296025
transform 1 0 881 0 1 358
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_pinv_dec  sky130_sram_1r1w_24x128_8_pinv_dec_0
timestamp 1661296025
transform 1 0 320 0 -1 790
box 44 0 760 490
use sky130_sram_1r1w_24x128_8_pinv_dec  sky130_sram_1r1w_24x128_8_pinv_dec_1
timestamp 1661296025
transform 1 0 320 0 1 0
box 44 0 760 490
<< labels >>
rlabel metal1 s 71 141 117 199 4 in_0
port 1 nsew
rlabel metal1 s 151 591 197 649 4 in_1
port 2 nsew
rlabel locali s 2871 120 2871 120 4 out_0
port 3 nsew
rlabel locali s 2871 670 2871 670 4 out_1
port 4 nsew
rlabel locali s 2871 910 2871 910 4 out_2
port 5 nsew
rlabel locali s 2871 1460 2871 1460 4 out_3
port 6 nsew
rlabel metal3 s 2188 353 2286 451 4 vdd
port 7 nsew
rlabel metal3 s 2963 346 3061 444 4 vdd
port 7 nsew
rlabel metal3 s 2963 1136 3061 1234 4 vdd
port 7 nsew
rlabel metal3 s 865 346 963 444 4 vdd
port 7 nsew
rlabel metal3 s 2188 1143 2286 1241 4 vdd
port 7 nsew
rlabel metal3 s 2567 346 2665 444 4 gnd
port 8 nsew
rlabel metal3 s 469 346 567 444 4 gnd
port 8 nsew
rlabel metal3 s 2567 1136 2665 1234 4 gnd
port 8 nsew
rlabel metal3 s 1763 1143 1861 1241 4 gnd
port 8 nsew
rlabel metal3 s 1763 353 1861 451 4 gnd
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 3160 1580
<< end >>
