* NGSPICE file created from NMOS_30_0p5_30_diff4x_1_flat.ext - technology: sky130B

X0 SD2L.t119 GL SD1L.t79 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X1 SD1R.t119 GL SD2R.t94 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X2 SD1R.t59 GR SD2R.t26 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X3 SD2L.t118 GL SD1L.t99 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X4 SD1R.t118 GL SD2R.t101 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X5 SD2L.t117 GL SD1L.t70 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X6 SD1R.t58 GR SD2R.t41 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X7 SD1L.t24 GR SD2L.t59 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X8 SD1L.t118 GL SD2L.t116 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X9 SD1L.t103 GL SD2L.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X10 SD2R.t75 GL SD1R.t117 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X11 SD1L.t71 GL SD2L.t114 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X12 SD1R.t116 GL SD2R.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X13 SD1L.t84 GL SD2L.t113 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X14 SD2R.t69 GL SD1R.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X15 SD2R.t0 GR SD1R.t57 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X16 SD2R.t23 GR SD1R.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X17 SD2L.t58 GR SD1L.t52 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X18 SD2R.t105 GL SD1R.t114 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X19 SD2L.t57 GR SD1L.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X20 SD2R.t33 GR SD1R.t55 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X21 SD1L.t94 GL SD2L.t112 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X22 SD1R.t54 GR SD2R.t59 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X23 SD2R.t107 GL SD1R.t113 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X24 SD2L.t111 GL SD1L.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X25 SD1L.t20 GR SD2L.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X26 SD1R.t53 GR SD2R.t54 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X27 SD2L.t110 GL SD1L.t60 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X28 SD2L.t109 GL SD1L.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X29 SD1R.t52 GR SD2R.t19 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X30 SD2L.t108 GL SD1L.t85 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X31 SD1L.t34 GR SD2L.t55 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X32 SD1R.t51 GR SD2R.t1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X33 SD1R.t112 GL SD2R.t85 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X34 SD2R.t37 GR SD1R.t50 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X35 SD1R.t111 GL SD2R.t82 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X36 SD1R.t110 GL SD2R.t114 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X37 SD1L.t100 GL SD2L.t107 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X38 SD1R.t109 GL SD2R.t88 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X39 SD1R.t108 GL SD2R.t63 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X40 SD1L.t80 GL SD2L.t106 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X41 SD1L.t40 GR SD2L.t54 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X42 SD2L.t53 GR SD1L.t6 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X43 SD1L.t105 GL SD2L.t105 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X44 SD2L.t52 GR SD1L.t46 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X45 SD1R.t107 GL SD2R.t70 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X46 SD2R.t71 GL SD1R.t106 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X47 SD2L.t51 GR SD1L.t25 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X48 SD2R.t5 GR SD1R.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X49 SD1R.t48 GR SD2R.t48 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X50 SD1R.t47 GR SD2R.t38 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X51 SD2L.t50 GR SD1L.t53 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X52 SD2R.t49 GR SD1R.t46 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X53 SD1L.t66 GL SD2L.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X54 SD2L.t49 GR SD1L.t17 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X55 SD2L.t103 GL SD1L.t95 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X56 SD1R.t105 GL SD2R.t95 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X57 SD2R.t76 GL SD1R.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X58 SD2L.t48 GR SD1L.t26 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X59 SD1R.t45 GR SD2R.t34 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X60 SD2R.t89 GL SD1R.t103 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X61 SD2R.t79 GL SD1R.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X62 SD1L.t13 GR SD2L.t47 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X63 SD2L.t102 GL SD1L.t106 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X64 SD1L.t38 GR SD2L.t46 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X65 SD1R.t44 GR SD2R.t36 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X66 SD1L.t7 GR SD2L.t45 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X67 SD1R.t101 GL SD2R.t92 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X68 SD1L.t61 GL SD2L.t101 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X69 SD2L.t44 GR SD1L.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X70 SD1L.t41 GR SD2L.t43 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X71 SD2R.t12 GR SD1R.t43 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X72 SD2L.t42 GR SD1L.t8 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X73 SD1L.t21 GR SD2L.t41 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X74 SD2R.t6 GR SD1R.t42 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X75 SD1R.t100 GL SD2R.t64 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X76 SD1R.t99 GL SD2R.t61 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X77 SD2R.t3 GR SD1R.t41 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X78 SD1R.t98 GL SD2R.t106 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X79 SD1R.t40 GR SD2R.t51 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X80 SD2R.t108 GL SD1R.t97 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X81 SD2L.t40 GR SD1L.t35 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X82 SD1R.t39 GR SD2R.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X83 SD2L.t39 GR SD1L.t42 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X84 SD1R.t38 GR SD2R.t24 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X85 SD2R.t118 GL SD1R.t96 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X86 SD2L.t38 GR SD1L.t0 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X87 SD1L.t9 GR SD2L.t37 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X88 SD2L.t36 GR SD1L.t22 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X89 SD2R.t115 GL SD1R.t95 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X90 SD1L.t39 GR SD2L.t35 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X91 SD2R.t21 GR SD1R.t37 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X92 SD2L.t100 GL SD1L.t92 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X93 SD2R.t111 GL SD1R.t94 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X94 SD1L.t73 GL SD2L.t99 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X95 SD2R.t56 GR SD1R.t36 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X96 SD1L.t14 GR SD2L.t34 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X97 SD1L.t43 GR SD2L.t33 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X98 SD2L.t32 GR SD1L.t4 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X99 SD1L.t67 GL SD2L.t98 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X100 SD1L.t36 GR SD2L.t31 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X101 SD2R.t55 GR SD1R.t35 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X102 SD1R.t93 GL SD2R.t100 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X103 SD2R.t30 GR SD1R.t34 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X104 SD2L.t30 GR SD1L.t44 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X105 SD1R.t92 GL SD2R.t96 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X106 SD2R.t39 GR SD1R.t33 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X107 SD2R.t90 GL SD1R.t91 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X108 SD2L.t97 GL SD1L.t64 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X109 SD1R.t32 GR SD2R.t50 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X110 SD2L.t96 GL SD1L.t112 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X111 SD2L.t95 GL SD1L.t89 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X112 SD2R.t119 GL SD1R.t90 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X113 SD1L.t1 GR SD2L.t29 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X114 SD1R.t89 GL SD2R.t112 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X115 SD1L.t30 GR SD2L.t28 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X116 SD2L.t94 GL SD1L.t116 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X117 SD1R.t88 GL SD2R.t81 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X118 SD1L.t10 GR SD2L.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X119 SD2R.t17 GR SD1R.t31 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X120 SD1L.t115 GL SD2L.t93 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X121 SD1L.t86 GL SD2L.t92 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X122 SD1L.t96 GL SD2L.t91 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X123 SD2R.t18 GR SD1R.t30 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X124 SD1L.t107 GL SD2L.t90 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X125 SD2R.t13 GR SD1R.t29 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X126 SD1L.t74 GL SD2L.t89 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X127 SD2L.t88 GL SD1L.t113 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X128 SD1L.t90 GL SD2L.t87 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X129 SD1L.t5 GR SD2L.t26 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X130 SD2R.t52 GR SD1R.t28 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X131 SD2L.t86 GL SD1L.t117 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X132 SD2R.t60 GL SD1R.t87 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X133 SD2R.t97 GL SD1R.t86 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X134 SD2R.t65 GL SD1R.t85 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X135 SD2L.t85 GL SD1L.t83 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X136 SD2L.t25 GR SD1L.t3 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X137 SD2L.t84 GL SD1L.t91 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X138 SD2R.t68 GL SD1R.t84 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X139 SD2L.t83 GL SD1L.t81 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X140 SD1L.t47 GR SD2L.t24 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X141 SD2L.t82 GL SD1L.t101 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X142 SD1R.t83 GL SD2R.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X143 SD1L.t75 GL SD2L.t81 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X144 SD2R.t28 GR SD1R.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X145 SD2L.t80 GL SD1L.t119 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X146 SD2R.t25 GR SD1R.t26 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X147 SD1L.t108 GL SD2L.t79 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X148 SD1L.t76 GL SD2L.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X149 SD2R.t98 GL SD1R.t82 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X150 SD1R.t81 GL SD2R.t103 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X151 SD1L.t87 GL SD2L.t77 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X152 SD1L.t97 GL SD2L.t76 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X153 SD2R.t91 GL SD1R.t80 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X154 SD1L.t109 GL SD2L.t75 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X155 SD2L.t23 GR SD1L.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X156 SD2R.t22 GR SD1R.t25 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X157 SD2L.t22 GR SD1L.t54 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X158 SD2L.t74 GL SD1L.t62 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X159 SD2L.t21 GR SD1L.t50 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X160 SD1L.t23 GR SD2L.t20 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X161 SD2R.t93 GL SD1R.t79 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X162 SD1R.t24 GR SD2R.t57 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X163 SD2L.t73 GL SD1L.t77 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X164 SD2L.t72 GL SD1L.t88 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X165 SD1R.t23 GR SD2R.t31 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X166 SD2R.t72 GL SD1R.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X167 SD2L.t71 GL SD1L.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X168 SD2L.t70 GL SD1L.t82 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X169 SD1L.t37 GR SD2L.t19 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X170 SD1R.t22 GR SD2R.t7 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X171 SD1R.t77 GL SD2R.t66 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X172 SD2R.t14 GR SD1R.t21 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X173 SD1L.t45 GR SD2L.t18 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X174 SD1R.t76 GL SD2R.t62 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X175 SD2L.t17 GR SD1L.t11 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X176 SD2R.t20 GR SD1R.t20 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X177 SD1L.t110 GL SD2L.t69 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X178 SD2L.t16 GR SD1L.t48 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X179 SD1L.t68 GL SD2L.t68 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X180 SD1R.t19 GR SD2R.t32 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X181 SD2R.t109 GL SD1R.t75 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X182 SD1L.t98 GL SD2L.t67 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X183 SD1L.t28 GR SD2L.t15 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X184 SD1R.t18 GR SD2R.t42 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X185 SD2R.t86 GL SD1R.t74 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X186 SD2R.t83 GL SD1R.t73 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X187 SD2L.t14 GR SD1L.t55 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X188 SD1L.t18 GR SD2L.t13 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X189 SD1L.t29 GR SD2L.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X190 SD2L.t11 GR SD1L.t15 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X191 SD1R.t17 GR SD2R.t43 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X192 SD2R.t44 GR SD1R.t16 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X193 SD2R.t116 GL SD1R.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X194 SD2R.t113 GL SD1R.t71 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X195 SD1L.t12 GR SD2L.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X196 SD1R.t15 GR SD2R.t45 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X197 SD2R.t16 GR SD1R.t14 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X198 SD1R.t13 GR SD2R.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X199 SD2R.t15 GR SD1R.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X200 SD1L.t57 GR SD2L.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X201 SD1L.t111 GL SD2L.t66 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X202 SD1R.t70 GL SD2R.t99 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X203 SD1R.t69 GL SD2R.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X204 SD2L.t8 GR SD1L.t32 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X205 SD1L.t2 GR SD2L.t7 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X206 SD2L.t6 GR SD1L.t59 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X207 SD1R.t68 GL SD2R.t77 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X208 SD1R.t67 GL SD2R.t80 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X209 SD1L.t31 GR SD2L.t5 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X210 SD2L.t4 GR SD1L.t58 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X211 SD2R.t73 GL SD1R.t66 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X212 SD1R.t11 GR SD2R.t46 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X213 SD2R.t110 GL SD1R.t65 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X214 SD2R.t87 GL SD1R.t64 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X215 SD1R.t10 GR SD2R.t2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X216 SD2L.t3 GR SD1L.t51 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X217 SD2L.t65 GL SD1L.t63 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X218 SD1R.t9 GR SD2R.t8 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X219 SD1R.t8 GR SD2R.t40 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X220 SD2R.t47 GR SD1R.t7 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X221 SD1L.t19 GR SD2L.t2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X222 SD2R.t35 GR SD1R.t6 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X223 SD1R.t63 GL SD2R.t84 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X224 SD2L.t1 GR SD1L.t16 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X225 SD2L.t64 GL SD1L.t93 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X226 SD1L.t78 GL SD2L.t63 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X227 SD1R.t5 GR SD2R.t11 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X228 SD1R.t62 GL SD2R.t117 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X229 SD2R.t9 GR SD1R.t4 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X230 SD1R.t61 GL SD2R.t67 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X231 SD1R.t3 GR SD2R.t4 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X232 SD1L.t69 GL SD2L.t62 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X233 SD1R.t60 GL SD2R.t74 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X234 SD2L.t61 GL SD1L.t65 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X235 SD2L.t0 GR SD1L.t33 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X236 SD2R.t53 GR SD1R.t2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X237 SD2L.t60 GL SD1L.t114 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X238 SD1R.t1 GR SD2R.t29 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X239 SD1R.t0 GR SD2R.t58 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
C0 SD1R GR 57.73fF
C1 SD1L GL 46.26fF
C2 SD1R SD1L 45.81fF
C3 SD2R SD2L 60.85fF
C4 SD2L GL 65.11fF
C5 SD1R SD2L 60.66fF
C6 GR SD1L 44.48fF
C7 SD2R GL 47.75fF
C8 SD2R SD1R 847.92fF
C9 GR SD2L 59.66fF
C10 SD1R GL 57.84fF
C11 SD2R GR 53.53fF
C12 GR GL 28.28fF
C13 SD1L SD2L 789.80fF
R0 SD1L.n6 SD1L.n40 1.435
R1 SD1L.n4 SD1L.n55 1.435
R2 SD1L.n2 SD1L.n25 1.435
R3 SD1L.n0 SD1L.n74 1.435
R4 SD1L.n14 SD1L.n30 1.428
R5 SD1L.n14 SD1L.n31 1.428
R6 SD1L.n13 SD1L.n32 1.428
R7 SD1L.n13 SD1L.n33 1.428
R8 SD1L.n7 SD1L.n34 1.428
R9 SD1L.n7 SD1L.n35 1.428
R10 SD1L.n7 SD1L.n36 1.428
R11 SD1L.n7 SD1L.n37 1.428
R12 SD1L.n6 SD1L.n38 1.428
R13 SD1L.n6 SD1L.n39 1.428
R14 SD1L.n12 SD1L.n45 1.428
R15 SD1L.n12 SD1L.n46 1.428
R16 SD1L.n11 SD1L.n47 1.428
R17 SD1L.n11 SD1L.n48 1.428
R18 SD1L.n5 SD1L.n49 1.428
R19 SD1L.n5 SD1L.n50 1.428
R20 SD1L.n5 SD1L.n51 1.428
R21 SD1L.n5 SD1L.n52 1.428
R22 SD1L.n4 SD1L.n53 1.428
R23 SD1L.n4 SD1L.n54 1.428
R24 SD1L.n8 SD1L.n15 1.428
R25 SD1L.n8 SD1L.n16 1.428
R26 SD1L.n8 SD1L.n17 1.428
R27 SD1L.n3 SD1L.n18 1.428
R28 SD1L.n3 SD1L.n19 1.428
R29 SD1L.n3 SD1L.n20 1.428
R30 SD1L.n3 SD1L.n21 1.428
R31 SD1L.n2 SD1L.n22 1.428
R32 SD1L.n2 SD1L.n23 1.428
R33 SD1L.n2 SD1L.n24 1.428
R34 SD1L.n10 SD1L.n65 1.428
R35 SD1L.n10 SD1L.n66 1.428
R36 SD1L.n9 SD1L.n67 1.428
R37 SD1L.n9 SD1L.n68 1.428
R38 SD1L.n1 SD1L.n69 1.428
R39 SD1L.n1 SD1L.n70 1.428
R40 SD1L.n1 SD1L.n71 1.428
R41 SD1L.n0 SD1L.n72 1.428
R42 SD1L.n0 SD1L.n73 1.428
R43 SD1L.n1 SD1L.n75 1.427
R44 SD1L.n14 SD1L.n41 0.895
R45 SD1L.n12 SD1L.n56 0.895
R46 SD1L.n10 SD1L.n64 0.895
R47 SD1L.n14 SD1L.n42 0.894
R48 SD1L.n14 SD1L.n43 0.894
R49 SD1L.n12 SD1L.n57 0.894
R50 SD1L.n12 SD1L.n58 0.894
R51 SD1L.n8 SD1L.n29 0.894
R52 SD1L.n8 SD1L.n28 0.894
R53 SD1L.n8 SD1L.n27 0.894
R54 SD1L.n10 SD1L.n62 0.894
R55 SD1L.n10 SD1L.n61 0.894
R56 SD1L.n14 SD1L.n44 0.893
R57 SD1L.n12 SD1L.n59 0.893
R58 SD1L.n10 SD1L.n63 0.893
R59 SD1L.n8 SD1L.n26 0.892
R60 SD1L.n30 SD1L.t79 0.551
R61 SD1L.n30 SD1L.t78 0.551
R62 SD1L.n31 SD1L.t93 0.551
R63 SD1L.n31 SD1L.t94 0.551
R64 SD1L.n32 SD1L.t117 0.551
R65 SD1L.n32 SD1L.t68 0.551
R66 SD1L.n33 SD1L.t116 0.551
R67 SD1L.n33 SD1L.t76 0.551
R68 SD1L.n34 SD1L.t119 0.551
R69 SD1L.n34 SD1L.t74 0.551
R70 SD1L.n35 SD1L.t95 0.551
R71 SD1L.n35 SD1L.t100 0.551
R72 SD1L.n36 SD1L.t85 0.551
R73 SD1L.n36 SD1L.t84 0.551
R74 SD1L.n37 SD1L.t99 0.551
R75 SD1L.n37 SD1L.t66 0.551
R76 SD1L.n38 SD1L.t102 0.551
R77 SD1L.n38 SD1L.t111 0.551
R78 SD1L.n39 SD1L.t91 0.551
R79 SD1L.n39 SD1L.t98 0.551
R80 SD1L.n40 SD1L.t82 0.551
R81 SD1L.n40 SD1L.t97 0.551
R82 SD1L.n41 SD1L.t72 0.551
R83 SD1L.n41 SD1L.t103 0.551
R84 SD1L.n42 SD1L.t106 0.551
R85 SD1L.n42 SD1L.t67 0.551
R86 SD1L.n43 SD1L.t101 0.551
R87 SD1L.n43 SD1L.t107 0.551
R88 SD1L.n44 SD1L.t89 0.551
R89 SD1L.n44 SD1L.t87 0.551
R90 SD1L.n45 SD1L.t27 0.551
R91 SD1L.n45 SD1L.t47 0.551
R92 SD1L.n46 SD1L.t3 0.551
R93 SD1L.n46 SD1L.t28 0.551
R94 SD1L.n47 SD1L.t46 0.551
R95 SD1L.n47 SD1L.t43 0.551
R96 SD1L.n48 SD1L.t49 0.551
R97 SD1L.n48 SD1L.t38 0.551
R98 SD1L.n49 SD1L.t26 0.551
R99 SD1L.n49 SD1L.t40 0.551
R100 SD1L.n50 SD1L.t58 0.551
R101 SD1L.n50 SD1L.t12 0.551
R102 SD1L.n51 SD1L.t15 0.551
R103 SD1L.n51 SD1L.t45 0.551
R104 SD1L.n52 SD1L.t50 0.551
R105 SD1L.n52 SD1L.t2 0.551
R106 SD1L.n53 SD1L.t42 0.551
R107 SD1L.n53 SD1L.t10 0.551
R108 SD1L.n54 SD1L.t53 0.551
R109 SD1L.n54 SD1L.t36 0.551
R110 SD1L.n55 SD1L.t22 0.551
R111 SD1L.n55 SD1L.t41 0.551
R112 SD1L.n56 SD1L.t55 0.551
R113 SD1L.n56 SD1L.t37 0.551
R114 SD1L.n57 SD1L.t51 0.551
R115 SD1L.n57 SD1L.t24 0.551
R116 SD1L.n58 SD1L.t17 0.551
R117 SD1L.n58 SD1L.t34 0.551
R118 SD1L.n59 SD1L.t52 0.551
R119 SD1L.n59 SD1L.t21 0.551
R120 SD1L.n15 SD1L.t64 0.551
R121 SD1L.n15 SD1L.t73 0.551
R122 SD1L.n16 SD1L.t92 0.551
R123 SD1L.n16 SD1L.t90 0.551
R124 SD1L.n17 SD1L.t65 0.551
R125 SD1L.n17 SD1L.t80 0.551
R126 SD1L.n18 SD1L.t63 0.551
R127 SD1L.n18 SD1L.t118 0.551
R128 SD1L.n19 SD1L.t70 0.551
R129 SD1L.n19 SD1L.t69 0.551
R130 SD1L.n20 SD1L.t62 0.551
R131 SD1L.n20 SD1L.t75 0.551
R132 SD1L.n21 SD1L.t81 0.551
R133 SD1L.n21 SD1L.t96 0.551
R134 SD1L.n22 SD1L.t112 0.551
R135 SD1L.n22 SD1L.t109 0.551
R136 SD1L.n23 SD1L.t104 0.551
R137 SD1L.n23 SD1L.t61 0.551
R138 SD1L.n24 SD1L.t114 0.551
R139 SD1L.n24 SD1L.t105 0.551
R140 SD1L.n25 SD1L.t60 0.551
R141 SD1L.n25 SD1L.t71 0.551
R142 SD1L.n29 SD1L.t83 0.551
R143 SD1L.n29 SD1L.t86 0.551
R144 SD1L.n28 SD1L.t88 0.551
R145 SD1L.n28 SD1L.t115 0.551
R146 SD1L.n27 SD1L.t77 0.551
R147 SD1L.n27 SD1L.t108 0.551
R148 SD1L.n26 SD1L.t113 0.551
R149 SD1L.n26 SD1L.t110 0.551
R150 SD1L.n65 SD1L.t48 0.551
R151 SD1L.n65 SD1L.t23 0.551
R152 SD1L.n66 SD1L.t54 0.551
R153 SD1L.n66 SD1L.t57 0.551
R154 SD1L.n67 SD1L.t8 0.551
R155 SD1L.n67 SD1L.t30 0.551
R156 SD1L.n68 SD1L.t25 0.551
R157 SD1L.n68 SD1L.t39 0.551
R158 SD1L.n69 SD1L.t16 0.551
R159 SD1L.n69 SD1L.t31 0.551
R160 SD1L.n70 SD1L.t32 0.551
R161 SD1L.n70 SD1L.t18 0.551
R162 SD1L.n71 SD1L.t11 0.551
R163 SD1L.n71 SD1L.t19 0.551
R164 SD1L.n72 SD1L.t4 0.551
R165 SD1L.n72 SD1L.t5 0.551
R166 SD1L.n73 SD1L.t56 0.551
R167 SD1L.n73 SD1L.t1 0.551
R168 SD1L.n74 SD1L.t44 0.551
R169 SD1L.n74 SD1L.t9 0.551
R170 SD1L.n64 SD1L.t59 0.551
R171 SD1L.n64 SD1L.t29 0.551
R172 SD1L.n63 SD1L.t33 0.551
R173 SD1L.n63 SD1L.t20 0.551
R174 SD1L.n62 SD1L.t35 0.551
R175 SD1L.n62 SD1L.t13 0.551
R176 SD1L.n61 SD1L.t6 0.551
R177 SD1L.n61 SD1L.t14 0.551
R178 SD1L.n75 SD1L.t0 0.551
R179 SD1L.n75 SD1L.t7 0.551
R180 SD1L.n60 SD1L.n12 0.185
R181 SD1L.n76 SD1L.n60 0.112
R182 SD1L.n77 SD1L.n76 0.08
R183 SD1L.n60 SD1L.n14 0.073
R184 SD1L.n77 SD1L.n8 0.073
R185 SD1L.n76 SD1L.n10 0.073
R186 SD1L.n8 SD1L.n3 0.041
R187 SD1L SD1L.n77 0.04
R188 SD1L.n13 SD1L.n7 0.028
R189 SD1L.n11 SD1L.n5 0.028
R190 SD1L.n3 SD1L.n2 0.028
R191 SD1L.n9 SD1L.n1 0.028
R192 SD1L.n14 SD1L.n13 0.022
R193 SD1L.n12 SD1L.n11 0.022
R194 SD1L.n10 SD1L.n9 0.022
R195 SD1L.n1 SD1L.n0 0.021
R196 SD1L.n5 SD1L.n4 0.021
R197 SD1L.n7 SD1L.n6 0.021
R198 SD2L.n37 SD2L.t30 1.972
R199 SD2L.n63 SD2L.t70 1.972
R200 SD2L.n14 SD2L.t110 1.972
R201 SD2L.n90 SD2L.t36 1.972
R202 SD2L.n25 SD2L.t69 1.826
R203 SD2L.n51 SD2L.t34 1.824
R204 SD2L.n77 SD2L.t77 1.824
R205 SD2L.n103 SD2L.t41 1.824
R206 SD2L.n47 SD2L.n26 1.414
R207 SD2L.n46 SD2L.n27 1.414
R208 SD2L.n45 SD2L.n28 1.414
R209 SD2L.n44 SD2L.n29 1.414
R210 SD2L.n43 SD2L.n30 1.414
R211 SD2L.n42 SD2L.n31 1.414
R212 SD2L.n41 SD2L.n32 1.414
R213 SD2L.n40 SD2L.n33 1.414
R214 SD2L.n39 SD2L.n34 1.414
R215 SD2L.n38 SD2L.n35 1.414
R216 SD2L.n37 SD2L.n36 1.414
R217 SD2L.n73 SD2L.n52 1.414
R218 SD2L.n72 SD2L.n53 1.414
R219 SD2L.n71 SD2L.n54 1.414
R220 SD2L.n70 SD2L.n55 1.414
R221 SD2L.n69 SD2L.n56 1.414
R222 SD2L.n68 SD2L.n57 1.414
R223 SD2L.n67 SD2L.n58 1.414
R224 SD2L.n66 SD2L.n59 1.414
R225 SD2L.n65 SD2L.n60 1.414
R226 SD2L.n64 SD2L.n61 1.414
R227 SD2L.n63 SD2L.n62 1.414
R228 SD2L.n24 SD2L.n3 1.414
R229 SD2L.n23 SD2L.n4 1.414
R230 SD2L.n22 SD2L.n5 1.414
R231 SD2L.n21 SD2L.n6 1.414
R232 SD2L.n20 SD2L.n7 1.414
R233 SD2L.n19 SD2L.n8 1.414
R234 SD2L.n18 SD2L.n9 1.414
R235 SD2L.n17 SD2L.n10 1.414
R236 SD2L.n16 SD2L.n11 1.414
R237 SD2L.n15 SD2L.n12 1.414
R238 SD2L.n14 SD2L.n13 1.414
R239 SD2L.n100 SD2L.n79 1.414
R240 SD2L.n99 SD2L.n80 1.414
R241 SD2L.n98 SD2L.n81 1.414
R242 SD2L.n97 SD2L.n82 1.414
R243 SD2L.n96 SD2L.n83 1.414
R244 SD2L.n95 SD2L.n84 1.414
R245 SD2L.n94 SD2L.n85 1.414
R246 SD2L.n93 SD2L.n86 1.414
R247 SD2L.n92 SD2L.n87 1.414
R248 SD2L.n91 SD2L.n88 1.414
R249 SD2L.n90 SD2L.n89 1.414
R250 SD2L.n51 SD2L.n49 1.261
R251 SD2L.n51 SD2L.n48 1.261
R252 SD2L.n77 SD2L.n75 1.261
R253 SD2L.n77 SD2L.n74 1.261
R254 SD2L.n25 SD2L.n0 1.261
R255 SD2L.n25 SD2L.n1 1.261
R256 SD2L.n103 SD2L.n102 1.261
R257 SD2L.n103 SD2L.n101 1.261
R258 SD2L.n51 SD2L.n50 1.261
R259 SD2L.n77 SD2L.n76 1.261
R260 SD2L.n25 SD2L.n2 1.261
R261 SD2L.n103 SD2L.n78 1.26
R262 SD2L.n26 SD2L.t20 0.551
R263 SD2L.n26 SD2L.t6 0.551
R264 SD2L.n27 SD2L.t9 0.551
R265 SD2L.n27 SD2L.t16 0.551
R266 SD2L.n28 SD2L.t28 0.551
R267 SD2L.n28 SD2L.t22 0.551
R268 SD2L.n29 SD2L.t35 0.551
R269 SD2L.n29 SD2L.t42 0.551
R270 SD2L.n30 SD2L.t45 0.551
R271 SD2L.n30 SD2L.t51 0.551
R272 SD2L.n31 SD2L.t5 0.551
R273 SD2L.n31 SD2L.t38 0.551
R274 SD2L.n32 SD2L.t13 0.551
R275 SD2L.n32 SD2L.t1 0.551
R276 SD2L.n33 SD2L.t2 0.551
R277 SD2L.n33 SD2L.t8 0.551
R278 SD2L.n34 SD2L.t26 0.551
R279 SD2L.n34 SD2L.t17 0.551
R280 SD2L.n35 SD2L.t29 0.551
R281 SD2L.n35 SD2L.t32 0.551
R282 SD2L.n36 SD2L.t37 0.551
R283 SD2L.n36 SD2L.t44 0.551
R284 SD2L.n48 SD2L.t12 0.551
R285 SD2L.n48 SD2L.t0 0.551
R286 SD2L.n50 SD2L.t56 0.551
R287 SD2L.n50 SD2L.t40 0.551
R288 SD2L.n49 SD2L.t47 0.551
R289 SD2L.n49 SD2L.t53 0.551
R290 SD2L.n52 SD2L.t63 0.551
R291 SD2L.n52 SD2L.t109 0.551
R292 SD2L.n53 SD2L.t112 0.551
R293 SD2L.n53 SD2L.t119 0.551
R294 SD2L.n54 SD2L.t68 0.551
R295 SD2L.n54 SD2L.t64 0.551
R296 SD2L.n55 SD2L.t78 0.551
R297 SD2L.n55 SD2L.t86 0.551
R298 SD2L.n56 SD2L.t89 0.551
R299 SD2L.n56 SD2L.t94 0.551
R300 SD2L.n57 SD2L.t107 0.551
R301 SD2L.n57 SD2L.t80 0.551
R302 SD2L.n58 SD2L.t113 0.551
R303 SD2L.n58 SD2L.t103 0.551
R304 SD2L.n59 SD2L.t104 0.551
R305 SD2L.n59 SD2L.t108 0.551
R306 SD2L.n60 SD2L.t66 0.551
R307 SD2L.n60 SD2L.t118 0.551
R308 SD2L.n61 SD2L.t67 0.551
R309 SD2L.n61 SD2L.t71 0.551
R310 SD2L.n62 SD2L.t76 0.551
R311 SD2L.n62 SD2L.t84 0.551
R312 SD2L.n74 SD2L.t115 0.551
R313 SD2L.n74 SD2L.t102 0.551
R314 SD2L.n76 SD2L.t98 0.551
R315 SD2L.n76 SD2L.t82 0.551
R316 SD2L.n75 SD2L.t90 0.551
R317 SD2L.n75 SD2L.t95 0.551
R318 SD2L.n3 SD2L.t99 0.551
R319 SD2L.n3 SD2L.t85 0.551
R320 SD2L.n4 SD2L.t87 0.551
R321 SD2L.n4 SD2L.t97 0.551
R322 SD2L.n5 SD2L.t106 0.551
R323 SD2L.n5 SD2L.t100 0.551
R324 SD2L.n6 SD2L.t116 0.551
R325 SD2L.n6 SD2L.t61 0.551
R326 SD2L.n7 SD2L.t62 0.551
R327 SD2L.n7 SD2L.t65 0.551
R328 SD2L.n8 SD2L.t81 0.551
R329 SD2L.n8 SD2L.t117 0.551
R330 SD2L.n9 SD2L.t91 0.551
R331 SD2L.n9 SD2L.t74 0.551
R332 SD2L.n10 SD2L.t75 0.551
R333 SD2L.n10 SD2L.t83 0.551
R334 SD2L.n11 SD2L.t101 0.551
R335 SD2L.n11 SD2L.t96 0.551
R336 SD2L.n12 SD2L.t105 0.551
R337 SD2L.n12 SD2L.t111 0.551
R338 SD2L.n13 SD2L.t114 0.551
R339 SD2L.n13 SD2L.t60 0.551
R340 SD2L.n1 SD2L.t92 0.551
R341 SD2L.n1 SD2L.t72 0.551
R342 SD2L.n2 SD2L.t93 0.551
R343 SD2L.n2 SD2L.t73 0.551
R344 SD2L.n0 SD2L.t79 0.551
R345 SD2L.n0 SD2L.t88 0.551
R346 SD2L.n79 SD2L.t24 0.551
R347 SD2L.n79 SD2L.t14 0.551
R348 SD2L.n80 SD2L.t15 0.551
R349 SD2L.n80 SD2L.t23 0.551
R350 SD2L.n81 SD2L.t33 0.551
R351 SD2L.n81 SD2L.t25 0.551
R352 SD2L.n82 SD2L.t46 0.551
R353 SD2L.n82 SD2L.t52 0.551
R354 SD2L.n83 SD2L.t54 0.551
R355 SD2L.n83 SD2L.t57 0.551
R356 SD2L.n84 SD2L.t10 0.551
R357 SD2L.n84 SD2L.t48 0.551
R358 SD2L.n85 SD2L.t18 0.551
R359 SD2L.n85 SD2L.t4 0.551
R360 SD2L.n86 SD2L.t7 0.551
R361 SD2L.n86 SD2L.t11 0.551
R362 SD2L.n87 SD2L.t27 0.551
R363 SD2L.n87 SD2L.t21 0.551
R364 SD2L.n88 SD2L.t31 0.551
R365 SD2L.n88 SD2L.t39 0.551
R366 SD2L.n89 SD2L.t43 0.551
R367 SD2L.n89 SD2L.t50 0.551
R368 SD2L.n101 SD2L.t19 0.551
R369 SD2L.n101 SD2L.t3 0.551
R370 SD2L.n102 SD2L.t55 0.551
R371 SD2L.n102 SD2L.t58 0.551
R372 SD2L.n78 SD2L.t59 0.551
R373 SD2L.n78 SD2L.t49 0.551
R374 SD2L.n104 SD2L.n103 0.479
R375 SD2L.n105 SD2L.n51 0.367
R376 SD2L.n104 SD2L.n77 0.367
R377 SD2L.n106 SD2L.n25 0.367
R378 SD2L.n105 SD2L.n104 0.112
R379 SD2L.n106 SD2L.n105 0.109
R380 SD2L SD2L.n106 0.011
R381 SD2L.n38 SD2L.n37 0.007
R382 SD2L.n39 SD2L.n38 0.007
R383 SD2L.n40 SD2L.n39 0.007
R384 SD2L.n41 SD2L.n40 0.007
R385 SD2L.n42 SD2L.n41 0.007
R386 SD2L.n43 SD2L.n42 0.007
R387 SD2L.n44 SD2L.n43 0.007
R388 SD2L.n45 SD2L.n44 0.007
R389 SD2L.n46 SD2L.n45 0.007
R390 SD2L.n47 SD2L.n46 0.007
R391 SD2L.n64 SD2L.n63 0.007
R392 SD2L.n65 SD2L.n64 0.007
R393 SD2L.n66 SD2L.n65 0.007
R394 SD2L.n67 SD2L.n66 0.007
R395 SD2L.n68 SD2L.n67 0.007
R396 SD2L.n69 SD2L.n68 0.007
R397 SD2L.n70 SD2L.n69 0.007
R398 SD2L.n71 SD2L.n70 0.007
R399 SD2L.n72 SD2L.n71 0.007
R400 SD2L.n73 SD2L.n72 0.007
R401 SD2L.n15 SD2L.n14 0.007
R402 SD2L.n16 SD2L.n15 0.007
R403 SD2L.n17 SD2L.n16 0.007
R404 SD2L.n18 SD2L.n17 0.007
R405 SD2L.n19 SD2L.n18 0.007
R406 SD2L.n20 SD2L.n19 0.007
R407 SD2L.n21 SD2L.n20 0.007
R408 SD2L.n22 SD2L.n21 0.007
R409 SD2L.n23 SD2L.n22 0.007
R410 SD2L.n24 SD2L.n23 0.007
R411 SD2L.n91 SD2L.n90 0.007
R412 SD2L.n92 SD2L.n91 0.007
R413 SD2L.n93 SD2L.n92 0.007
R414 SD2L.n94 SD2L.n93 0.007
R415 SD2L.n95 SD2L.n94 0.007
R416 SD2L.n96 SD2L.n95 0.007
R417 SD2L.n97 SD2L.n96 0.007
R418 SD2L.n98 SD2L.n97 0.007
R419 SD2L.n99 SD2L.n98 0.007
R420 SD2L.n100 SD2L.n99 0.007
R421 SD2L.n51 SD2L.n47 0.004
R422 SD2L.n77 SD2L.n73 0.004
R423 SD2L.n25 SD2L.n24 0.004
R424 SD2L.n103 SD2L.n100 0.004
R425 SD2R.n11 SD2R.n56 1.435
R426 SD2R.n8 SD2R.n30 1.435
R427 SD2R.n6 SD2R.n41 1.435
R428 SD2R.n5 SD2R.n15 1.435
R429 SD2R.n3 SD2R.n26 1.435
R430 SD2R.n2 SD2R.n71 1.435
R431 SD2R.n0 SD2R.n64 1.435
R432 SD2R.n9 SD2R.n52 1.434
R433 SD2R.n9 SD2R.n51 1.428
R434 SD2R.n9 SD2R.n50 1.428
R435 SD2R.n10 SD2R.n49 1.428
R436 SD2R.n10 SD2R.n48 1.428
R437 SD2R.n10 SD2R.n47 1.428
R438 SD2R.n10 SD2R.n46 1.428
R439 SD2R.n11 SD2R.n53 1.428
R440 SD2R.n11 SD2R.n54 1.428
R441 SD2R.n11 SD2R.n55 1.428
R442 SD2R.n8 SD2R.n27 1.428
R443 SD2R.n8 SD2R.n28 1.428
R444 SD2R.n8 SD2R.n29 1.428
R445 SD2R.n6 SD2R.n40 1.428
R446 SD2R.n6 SD2R.n39 1.428
R447 SD2R.n7 SD2R.n38 1.428
R448 SD2R.n7 SD2R.n37 1.428
R449 SD2R.n7 SD2R.n36 1.428
R450 SD2R.n8 SD2R.n35 1.428
R451 SD2R.n5 SD2R.n12 1.428
R452 SD2R.n5 SD2R.n13 1.428
R453 SD2R.n5 SD2R.n14 1.428
R454 SD2R.n3 SD2R.n25 1.428
R455 SD2R.n3 SD2R.n24 1.428
R456 SD2R.n4 SD2R.n23 1.428
R457 SD2R.n4 SD2R.n22 1.428
R458 SD2R.n4 SD2R.n21 1.428
R459 SD2R.n5 SD2R.n20 1.428
R460 SD2R.n2 SD2R.n69 1.428
R461 SD2R.n2 SD2R.n70 1.428
R462 SD2R.n0 SD2R.n63 1.428
R463 SD2R.n0 SD2R.n62 1.428
R464 SD2R.n1 SD2R.n61 1.428
R465 SD2R.n1 SD2R.n60 1.428
R466 SD2R.n1 SD2R.n59 1.428
R467 SD2R.n2 SD2R.n58 1.428
R468 SD2R.n2 SD2R.n72 1.427
R469 SD2R.n8 SD2R.n31 0.895
R470 SD2R.n5 SD2R.n16 0.895
R471 SD2R.n2 SD2R.n68 0.895
R472 SD2R.n8 SD2R.n32 0.894
R473 SD2R.n8 SD2R.n33 0.894
R474 SD2R.n5 SD2R.n17 0.894
R475 SD2R.n5 SD2R.n18 0.894
R476 SD2R.n2 SD2R.n66 0.894
R477 SD2R.n2 SD2R.n65 0.894
R478 SD2R.n10 SD2R.n42 0.893
R479 SD2R.n10 SD2R.n43 0.893
R480 SD2R.n10 SD2R.n44 0.893
R481 SD2R.n10 SD2R.n45 0.893
R482 SD2R.n8 SD2R.n34 0.893
R483 SD2R.n5 SD2R.n19 0.893
R484 SD2R.n2 SD2R.n67 0.893
R485 SD2R.n52 SD2R.t1 0.551
R486 SD2R.n52 SD2R.t33 0.551
R487 SD2R.n51 SD2R.t11 0.551
R488 SD2R.n51 SD2R.t52 0.551
R489 SD2R.n50 SD2R.t50 0.551
R490 SD2R.n50 SD2R.t53 0.551
R491 SD2R.n49 SD2R.t46 0.551
R492 SD2R.n49 SD2R.t17 0.551
R493 SD2R.n48 SD2R.t51 0.551
R494 SD2R.n48 SD2R.t35 0.551
R495 SD2R.n47 SD2R.t29 0.551
R496 SD2R.n47 SD2R.t9 0.551
R497 SD2R.n46 SD2R.t24 0.551
R498 SD2R.n46 SD2R.t12 0.551
R499 SD2R.n53 SD2R.t34 0.551
R500 SD2R.n53 SD2R.t5 0.551
R501 SD2R.n54 SD2R.t10 0.551
R502 SD2R.n54 SD2R.t18 0.551
R503 SD2R.n55 SD2R.t36 0.551
R504 SD2R.n55 SD2R.t49 0.551
R505 SD2R.n56 SD2R.t41 0.551
R506 SD2R.n56 SD2R.t22 0.551
R507 SD2R.n42 SD2R.t45 0.551
R508 SD2R.n42 SD2R.t39 0.551
R509 SD2R.n43 SD2R.t59 0.551
R510 SD2R.n43 SD2R.t20 0.551
R511 SD2R.n44 SD2R.t43 0.551
R512 SD2R.n44 SD2R.t55 0.551
R513 SD2R.n45 SD2R.t26 0.551
R514 SD2R.n45 SD2R.t14 0.551
R515 SD2R.n27 SD2R.t64 0.551
R516 SD2R.n27 SD2R.t76 0.551
R517 SD2R.n28 SD2R.t77 0.551
R518 SD2R.n28 SD2R.t97 0.551
R519 SD2R.n29 SD2R.t106 0.551
R520 SD2R.n29 SD2R.t89 0.551
R521 SD2R.n30 SD2R.t78 0.551
R522 SD2R.n30 SD2R.t72 0.551
R523 SD2R.n41 SD2R.t84 0.551
R524 SD2R.n41 SD2R.t110 0.551
R525 SD2R.n40 SD2R.t66 0.551
R526 SD2R.n40 SD2R.t108 0.551
R527 SD2R.n39 SD2R.t61 0.551
R528 SD2R.n39 SD2R.t109 0.551
R529 SD2R.n38 SD2R.t62 0.551
R530 SD2R.n38 SD2R.t118 0.551
R531 SD2R.n37 SD2R.t114 0.551
R532 SD2R.n37 SD2R.t83 0.551
R533 SD2R.n36 SD2R.t104 0.551
R534 SD2R.n36 SD2R.t113 0.551
R535 SD2R.n35 SD2R.t63 0.551
R536 SD2R.n35 SD2R.t107 0.551
R537 SD2R.n31 SD2R.t99 0.551
R538 SD2R.n31 SD2R.t119 0.551
R539 SD2R.n32 SD2R.t82 0.551
R540 SD2R.n32 SD2R.t86 0.551
R541 SD2R.n33 SD2R.t103 0.551
R542 SD2R.n33 SD2R.t79 0.551
R543 SD2R.n34 SD2R.t80 0.551
R544 SD2R.n34 SD2R.t65 0.551
R545 SD2R.n12 SD2R.t100 0.551
R546 SD2R.n12 SD2R.t115 0.551
R547 SD2R.n13 SD2R.t74 0.551
R548 SD2R.n13 SD2R.t93 0.551
R549 SD2R.n14 SD2R.t96 0.551
R550 SD2R.n14 SD2R.t111 0.551
R551 SD2R.n15 SD2R.t70 0.551
R552 SD2R.n15 SD2R.t116 0.551
R553 SD2R.n26 SD2R.t95 0.551
R554 SD2R.n26 SD2R.t71 0.551
R555 SD2R.n25 SD2R.t94 0.551
R556 SD2R.n25 SD2R.t98 0.551
R557 SD2R.n24 SD2R.t102 0.551
R558 SD2R.n24 SD2R.t75 0.551
R559 SD2R.n23 SD2R.t101 0.551
R560 SD2R.n23 SD2R.t91 0.551
R561 SD2R.n22 SD2R.t112 0.551
R562 SD2R.n22 SD2R.t69 0.551
R563 SD2R.n21 SD2R.t85 0.551
R564 SD2R.n21 SD2R.t105 0.551
R565 SD2R.n20 SD2R.t81 0.551
R566 SD2R.n20 SD2R.t90 0.551
R567 SD2R.n16 SD2R.t67 0.551
R568 SD2R.n16 SD2R.t68 0.551
R569 SD2R.n17 SD2R.t92 0.551
R570 SD2R.n17 SD2R.t87 0.551
R571 SD2R.n18 SD2R.t117 0.551
R572 SD2R.n18 SD2R.t60 0.551
R573 SD2R.n19 SD2R.t88 0.551
R574 SD2R.n19 SD2R.t73 0.551
R575 SD2R.n69 SD2R.t7 0.551
R576 SD2R.n69 SD2R.t30 0.551
R577 SD2R.n70 SD2R.t19 0.551
R578 SD2R.n70 SD2R.t23 0.551
R579 SD2R.n71 SD2R.t40 0.551
R580 SD2R.n71 SD2R.t13 0.551
R581 SD2R.n64 SD2R.t4 0.551
R582 SD2R.n64 SD2R.t47 0.551
R583 SD2R.n63 SD2R.t32 0.551
R584 SD2R.n63 SD2R.t21 0.551
R585 SD2R.n62 SD2R.t27 0.551
R586 SD2R.n62 SD2R.t44 0.551
R587 SD2R.n61 SD2R.t42 0.551
R588 SD2R.n61 SD2R.t56 0.551
R589 SD2R.n60 SD2R.t48 0.551
R590 SD2R.n60 SD2R.t16 0.551
R591 SD2R.n59 SD2R.t2 0.551
R592 SD2R.n59 SD2R.t15 0.551
R593 SD2R.n58 SD2R.t38 0.551
R594 SD2R.n58 SD2R.t37 0.551
R595 SD2R.n68 SD2R.t31 0.551
R596 SD2R.n68 SD2R.t3 0.551
R597 SD2R.n67 SD2R.t58 0.551
R598 SD2R.n67 SD2R.t25 0.551
R599 SD2R.n66 SD2R.t57 0.551
R600 SD2R.n66 SD2R.t6 0.551
R601 SD2R.n65 SD2R.t8 0.551
R602 SD2R.n65 SD2R.t28 0.551
R603 SD2R.n72 SD2R.t54 0.551
R604 SD2R.n72 SD2R.t0 0.551
R605 SD2R.n57 SD2R.n10 0.273
R606 SD2R.n57 SD2R.n8 0.161
R607 SD2R.n74 SD2R.n5 0.161
R608 SD2R.n73 SD2R.n2 0.161
R609 SD2R.n74 SD2R.n73 0.112
R610 SD2R.n73 SD2R.n57 0.112
R611 SD2R SD2R.n74 0.045
R612 SD2R.n8 SD2R.n7 0.035
R613 SD2R.n5 SD2R.n4 0.035
R614 SD2R.n2 SD2R.n1 0.035
R615 SD2R.n10 SD2R.n11 0.033
R616 SD2R.n10 SD2R.n9 0.028
R617 SD2R.n7 SD2R.n6 0.028
R618 SD2R.n4 SD2R.n3 0.028
R619 SD2R.n1 SD2R.n0 0.028
R620 SD1R.n72 SD1R.t65 1.972
R621 SD1R.n43 SD1R.t7 1.972
R622 SD1R.n14 SD1R.t106 1.972
R623 SD1R.n99 SD1R.t55 1.972
R624 SD1R.n86 SD1R.t116 1.812
R625 SD1R.n57 SD1R.t8 1.812
R626 SD1R.n28 SD1R.t107 1.812
R627 SD1R.n115 SD1R.t58 1.812
R628 SD1R.n99 SD1R.n98 1.414
R629 SD1R.n100 SD1R.n97 1.414
R630 SD1R.n101 SD1R.n96 1.414
R631 SD1R.n102 SD1R.n95 1.414
R632 SD1R.n103 SD1R.n94 1.414
R633 SD1R.n104 SD1R.n93 1.414
R634 SD1R.n105 SD1R.n92 1.414
R635 SD1R.n108 SD1R.n91 1.414
R636 SD1R.n109 SD1R.n90 1.414
R637 SD1R.n110 SD1R.n89 1.414
R638 SD1R.n111 SD1R.n88 1.414
R639 SD1R.n112 SD1R.n87 1.414
R640 SD1R.n72 SD1R.n71 1.414
R641 SD1R.n73 SD1R.n70 1.414
R642 SD1R.n74 SD1R.n69 1.414
R643 SD1R.n75 SD1R.n68 1.414
R644 SD1R.n76 SD1R.n67 1.414
R645 SD1R.n77 SD1R.n66 1.414
R646 SD1R.n78 SD1R.n65 1.414
R647 SD1R.n79 SD1R.n64 1.414
R648 SD1R.n80 SD1R.n63 1.414
R649 SD1R.n81 SD1R.n62 1.414
R650 SD1R.n82 SD1R.n61 1.414
R651 SD1R.n83 SD1R.n60 1.414
R652 SD1R.n84 SD1R.n59 1.414
R653 SD1R.n43 SD1R.n42 1.414
R654 SD1R.n44 SD1R.n41 1.414
R655 SD1R.n45 SD1R.n40 1.414
R656 SD1R.n46 SD1R.n39 1.414
R657 SD1R.n47 SD1R.n38 1.414
R658 SD1R.n48 SD1R.n37 1.414
R659 SD1R.n49 SD1R.n36 1.414
R660 SD1R.n50 SD1R.n35 1.414
R661 SD1R.n51 SD1R.n34 1.414
R662 SD1R.n52 SD1R.n33 1.414
R663 SD1R.n53 SD1R.n32 1.414
R664 SD1R.n54 SD1R.n31 1.414
R665 SD1R.n55 SD1R.n30 1.414
R666 SD1R.n14 SD1R.n13 1.414
R667 SD1R.n15 SD1R.n12 1.414
R668 SD1R.n16 SD1R.n11 1.414
R669 SD1R.n17 SD1R.n10 1.414
R670 SD1R.n18 SD1R.n9 1.414
R671 SD1R.n19 SD1R.n8 1.414
R672 SD1R.n20 SD1R.n7 1.414
R673 SD1R.n21 SD1R.n6 1.414
R674 SD1R.n22 SD1R.n5 1.414
R675 SD1R.n23 SD1R.n4 1.414
R676 SD1R.n24 SD1R.n3 1.414
R677 SD1R.n25 SD1R.n2 1.414
R678 SD1R.n26 SD1R.n1 1.414
R679 SD1R.n107 SD1R.n106 1.413
R680 SD1R.n114 SD1R.n113 1.271
R681 SD1R.n85 SD1R.n58 1.27
R682 SD1R.n56 SD1R.n29 1.27
R683 SD1R.n27 SD1R.n0 1.27
R684 SD1R.n116 SD1R.n115 0.567
R685 SD1R.n98 SD1R.t28 0.551
R686 SD1R.n98 SD1R.t51 0.551
R687 SD1R.n97 SD1R.t2 0.551
R688 SD1R.n97 SD1R.t5 0.551
R689 SD1R.n96 SD1R.t31 0.551
R690 SD1R.n96 SD1R.t32 0.551
R691 SD1R.n95 SD1R.t6 0.551
R692 SD1R.n95 SD1R.t11 0.551
R693 SD1R.n94 SD1R.t4 0.551
R694 SD1R.n94 SD1R.t40 0.551
R695 SD1R.n93 SD1R.t43 0.551
R696 SD1R.n93 SD1R.t1 0.551
R697 SD1R.n92 SD1R.t21 0.551
R698 SD1R.n92 SD1R.t38 0.551
R699 SD1R.n91 SD1R.t20 0.551
R700 SD1R.n91 SD1R.t17 0.551
R701 SD1R.n90 SD1R.t33 0.551
R702 SD1R.n90 SD1R.t54 0.551
R703 SD1R.n89 SD1R.t49 0.551
R704 SD1R.n89 SD1R.t15 0.551
R705 SD1R.n88 SD1R.t30 0.551
R706 SD1R.n88 SD1R.t45 0.551
R707 SD1R.n87 SD1R.t46 0.551
R708 SD1R.n87 SD1R.t13 0.551
R709 SD1R.n71 SD1R.t97 0.551
R710 SD1R.n71 SD1R.t63 0.551
R711 SD1R.n70 SD1R.t75 0.551
R712 SD1R.n70 SD1R.t77 0.551
R713 SD1R.n69 SD1R.t96 0.551
R714 SD1R.n69 SD1R.t99 0.551
R715 SD1R.n68 SD1R.t73 0.551
R716 SD1R.n68 SD1R.t76 0.551
R717 SD1R.n67 SD1R.t71 0.551
R718 SD1R.n67 SD1R.t110 0.551
R719 SD1R.n66 SD1R.t113 0.551
R720 SD1R.n66 SD1R.t69 0.551
R721 SD1R.n65 SD1R.t85 0.551
R722 SD1R.n65 SD1R.t108 0.551
R723 SD1R.n64 SD1R.t102 0.551
R724 SD1R.n64 SD1R.t67 0.551
R725 SD1R.n63 SD1R.t74 0.551
R726 SD1R.n63 SD1R.t81 0.551
R727 SD1R.n62 SD1R.t90 0.551
R728 SD1R.n62 SD1R.t111 0.551
R729 SD1R.n61 SD1R.t104 0.551
R730 SD1R.n61 SD1R.t70 0.551
R731 SD1R.n60 SD1R.t86 0.551
R732 SD1R.n60 SD1R.t100 0.551
R733 SD1R.n59 SD1R.t103 0.551
R734 SD1R.n59 SD1R.t68 0.551
R735 SD1R.n58 SD1R.t78 0.551
R736 SD1R.n58 SD1R.t98 0.551
R737 SD1R.n42 SD1R.t37 0.551
R738 SD1R.n42 SD1R.t3 0.551
R739 SD1R.n41 SD1R.t16 0.551
R740 SD1R.n41 SD1R.t19 0.551
R741 SD1R.n40 SD1R.t36 0.551
R742 SD1R.n40 SD1R.t39 0.551
R743 SD1R.n39 SD1R.t14 0.551
R744 SD1R.n39 SD1R.t18 0.551
R745 SD1R.n38 SD1R.t12 0.551
R746 SD1R.n38 SD1R.t48 0.551
R747 SD1R.n37 SD1R.t50 0.551
R748 SD1R.n37 SD1R.t10 0.551
R749 SD1R.n36 SD1R.t27 0.551
R750 SD1R.n36 SD1R.t47 0.551
R751 SD1R.n35 SD1R.t42 0.551
R752 SD1R.n35 SD1R.t9 0.551
R753 SD1R.n34 SD1R.t26 0.551
R754 SD1R.n34 SD1R.t24 0.551
R755 SD1R.n33 SD1R.t41 0.551
R756 SD1R.n33 SD1R.t0 0.551
R757 SD1R.n32 SD1R.t57 0.551
R758 SD1R.n32 SD1R.t23 0.551
R759 SD1R.n31 SD1R.t34 0.551
R760 SD1R.n31 SD1R.t53 0.551
R761 SD1R.n30 SD1R.t56 0.551
R762 SD1R.n30 SD1R.t22 0.551
R763 SD1R.n29 SD1R.t29 0.551
R764 SD1R.n29 SD1R.t52 0.551
R765 SD1R.n13 SD1R.t82 0.551
R766 SD1R.n13 SD1R.t105 0.551
R767 SD1R.n12 SD1R.t117 0.551
R768 SD1R.n12 SD1R.t119 0.551
R769 SD1R.n11 SD1R.t80 0.551
R770 SD1R.n11 SD1R.t83 0.551
R771 SD1R.n10 SD1R.t115 0.551
R772 SD1R.n10 SD1R.t118 0.551
R773 SD1R.n9 SD1R.t114 0.551
R774 SD1R.n9 SD1R.t89 0.551
R775 SD1R.n8 SD1R.t91 0.551
R776 SD1R.n8 SD1R.t112 0.551
R777 SD1R.n7 SD1R.t66 0.551
R778 SD1R.n7 SD1R.t88 0.551
R779 SD1R.n6 SD1R.t87 0.551
R780 SD1R.n6 SD1R.t109 0.551
R781 SD1R.n5 SD1R.t64 0.551
R782 SD1R.n5 SD1R.t62 0.551
R783 SD1R.n4 SD1R.t84 0.551
R784 SD1R.n4 SD1R.t101 0.551
R785 SD1R.n3 SD1R.t95 0.551
R786 SD1R.n3 SD1R.t61 0.551
R787 SD1R.n2 SD1R.t79 0.551
R788 SD1R.n2 SD1R.t93 0.551
R789 SD1R.n1 SD1R.t94 0.551
R790 SD1R.n1 SD1R.t60 0.551
R791 SD1R.n0 SD1R.t72 0.551
R792 SD1R.n0 SD1R.t92 0.551
R793 SD1R.n113 SD1R.t25 0.551
R794 SD1R.n113 SD1R.t44 0.551
R795 SD1R.n106 SD1R.t35 0.551
R796 SD1R.n106 SD1R.t59 0.551
R797 SD1R SD1R.n28 0.484
R798 SD1R.n116 SD1R.n86 0.455
R799 SD1R.n117 SD1R.n57 0.455
R800 SD1R.n117 SD1R.n116 0.112
R801 SD1R SD1R.n117 0.08
R802 SD1R.n84 SD1R.n83 0.007
R803 SD1R.n83 SD1R.n82 0.007
R804 SD1R.n82 SD1R.n81 0.007
R805 SD1R.n81 SD1R.n80 0.007
R806 SD1R.n80 SD1R.n79 0.007
R807 SD1R.n79 SD1R.n78 0.007
R808 SD1R.n78 SD1R.n77 0.007
R809 SD1R.n77 SD1R.n76 0.007
R810 SD1R.n76 SD1R.n75 0.007
R811 SD1R.n75 SD1R.n74 0.007
R812 SD1R.n74 SD1R.n73 0.007
R813 SD1R.n73 SD1R.n72 0.007
R814 SD1R.n55 SD1R.n54 0.007
R815 SD1R.n54 SD1R.n53 0.007
R816 SD1R.n53 SD1R.n52 0.007
R817 SD1R.n52 SD1R.n51 0.007
R818 SD1R.n51 SD1R.n50 0.007
R819 SD1R.n50 SD1R.n49 0.007
R820 SD1R.n49 SD1R.n48 0.007
R821 SD1R.n48 SD1R.n47 0.007
R822 SD1R.n47 SD1R.n46 0.007
R823 SD1R.n46 SD1R.n45 0.007
R824 SD1R.n45 SD1R.n44 0.007
R825 SD1R.n44 SD1R.n43 0.007
R826 SD1R.n26 SD1R.n25 0.007
R827 SD1R.n25 SD1R.n24 0.007
R828 SD1R.n24 SD1R.n23 0.007
R829 SD1R.n23 SD1R.n22 0.007
R830 SD1R.n22 SD1R.n21 0.007
R831 SD1R.n21 SD1R.n20 0.007
R832 SD1R.n20 SD1R.n19 0.007
R833 SD1R.n19 SD1R.n18 0.007
R834 SD1R.n18 SD1R.n17 0.007
R835 SD1R.n17 SD1R.n16 0.007
R836 SD1R.n16 SD1R.n15 0.007
R837 SD1R.n15 SD1R.n14 0.007
R838 SD1R.n112 SD1R.n111 0.007
R839 SD1R.n111 SD1R.n110 0.007
R840 SD1R.n110 SD1R.n109 0.007
R841 SD1R.n109 SD1R.n108 0.007
R842 SD1R.n108 SD1R.n107 0.007
R843 SD1R.n107 SD1R.n105 0.007
R844 SD1R.n105 SD1R.n104 0.007
R845 SD1R.n104 SD1R.n103 0.007
R846 SD1R.n103 SD1R.n102 0.007
R847 SD1R.n102 SD1R.n101 0.007
R848 SD1R.n101 SD1R.n100 0.007
R849 SD1R.n100 SD1R.n99 0.007
R850 SD1R.n85 SD1R.n84 0.006
R851 SD1R.n56 SD1R.n55 0.006
R852 SD1R.n27 SD1R.n26 0.006
R853 SD1R.n114 SD1R.n112 0.006
R854 SD1R.n86 SD1R.n85 0.003
R855 SD1R.n57 SD1R.n56 0.003
R856 SD1R.n28 SD1R.n27 0.003
R857 SD1R.n115 SD1R.n114 0.003
C14 SD2R SUB 47.32fF
C15 SD1R SUB 209.24fF
C16 GR SUB 98.13fF $ **FLOATING
C17 SD1L SUB 52.73fF
C18 SD2L SUB 93.29fF
C19 GL SUB 98.70fF $ **FLOATING
C20 SD1R.n0 SUB 3.36fF
C21 SD1R.n1 SUB 3.38fF
C22 SD1R.n2 SUB 3.38fF
C23 SD1R.n3 SUB 3.38fF
C24 SD1R.n4 SUB 3.38fF
C25 SD1R.n5 SUB 3.38fF
C26 SD1R.n6 SUB 3.38fF
C27 SD1R.n7 SUB 3.38fF
C28 SD1R.n8 SUB 3.38fF
C29 SD1R.n9 SUB 3.38fF
C30 SD1R.n10 SUB 3.38fF
C31 SD1R.n11 SUB 3.38fF
C32 SD1R.n12 SUB 3.38fF
C33 SD1R.n13 SUB 3.38fF
C34 SD1R.t106 SUB 3.07fF $ **FLOATING
C35 SD1R.n14 SUB 9.18fF
C36 SD1R.n15 SUB 4.03fF
C37 SD1R.n16 SUB 4.03fF
C38 SD1R.n17 SUB 4.03fF
C39 SD1R.n18 SUB 4.03fF
C40 SD1R.n19 SUB 4.03fF
C41 SD1R.n20 SUB 4.03fF
C42 SD1R.n21 SUB 4.03fF
C43 SD1R.n22 SUB 4.03fF
C44 SD1R.n23 SUB 4.03fF
C45 SD1R.n24 SUB 4.03fF
C46 SD1R.n25 SUB 4.03fF
C47 SD1R.n26 SUB 3.92fF
C48 SD1R.n27 SUB 3.54fF
C49 SD1R.t107 SUB 2.94fF $ **FLOATING
C50 SD1R.n28 SUB 76.81fF
C51 SD1R.n29 SUB 3.36fF
C52 SD1R.n30 SUB 3.38fF
C53 SD1R.n31 SUB 3.38fF
C54 SD1R.n32 SUB 3.38fF
C55 SD1R.n33 SUB 3.38fF
C56 SD1R.n34 SUB 3.38fF
C57 SD1R.n35 SUB 3.38fF
C58 SD1R.n36 SUB 3.38fF
C59 SD1R.n37 SUB 3.38fF
C60 SD1R.n38 SUB 3.38fF
C61 SD1R.n39 SUB 3.38fF
C62 SD1R.n40 SUB 3.38fF
C63 SD1R.n41 SUB 3.38fF
C64 SD1R.n42 SUB 3.38fF
C65 SD1R.t7 SUB 3.07fF $ **FLOATING
C66 SD1R.n43 SUB 9.18fF
C67 SD1R.n44 SUB 4.03fF
C68 SD1R.n45 SUB 4.03fF
C69 SD1R.n46 SUB 4.03fF
C70 SD1R.n47 SUB 4.03fF
C71 SD1R.n48 SUB 4.03fF
C72 SD1R.n49 SUB 4.03fF
C73 SD1R.n50 SUB 4.03fF
C74 SD1R.n51 SUB 4.03fF
C75 SD1R.n52 SUB 4.03fF
C76 SD1R.n53 SUB 4.03fF
C77 SD1R.n54 SUB 4.03fF
C78 SD1R.n55 SUB 3.92fF
C79 SD1R.n56 SUB 3.54fF
C80 SD1R.t8 SUB 2.94fF $ **FLOATING
C81 SD1R.n57 SUB 72.51fF
C82 SD1R.n58 SUB 3.36fF
C83 SD1R.n59 SUB 3.38fF
C84 SD1R.n60 SUB 3.38fF
C85 SD1R.n61 SUB 3.38fF
C86 SD1R.n62 SUB 3.38fF
C87 SD1R.n63 SUB 3.38fF
C88 SD1R.n64 SUB 3.38fF
C89 SD1R.n65 SUB 3.38fF
C90 SD1R.n66 SUB 3.38fF
C91 SD1R.n67 SUB 3.38fF
C92 SD1R.n68 SUB 3.38fF
C93 SD1R.n69 SUB 3.38fF
C94 SD1R.n70 SUB 3.38fF
C95 SD1R.n71 SUB 3.38fF
C96 SD1R.t65 SUB 3.07fF $ **FLOATING
C97 SD1R.n72 SUB 9.18fF
C98 SD1R.n73 SUB 4.03fF
C99 SD1R.n74 SUB 4.03fF
C100 SD1R.n75 SUB 4.03fF
C101 SD1R.n76 SUB 4.03fF
C102 SD1R.n77 SUB 4.03fF
C103 SD1R.n78 SUB 4.03fF
C104 SD1R.n79 SUB 4.03fF
C105 SD1R.n80 SUB 4.03fF
C106 SD1R.n81 SUB 4.03fF
C107 SD1R.n82 SUB 4.03fF
C108 SD1R.n83 SUB 4.03fF
C109 SD1R.n84 SUB 3.92fF
C110 SD1R.n85 SUB 3.54fF
C111 SD1R.t116 SUB 2.94fF $ **FLOATING
C112 SD1R.n86 SUB 72.51fF
C113 SD1R.t58 SUB 2.94fF $ **FLOATING
C114 SD1R.n87 SUB 3.38fF
C115 SD1R.n88 SUB 3.38fF
C116 SD1R.n89 SUB 3.38fF
C117 SD1R.n90 SUB 3.38fF
C118 SD1R.n91 SUB 3.38fF
C119 SD1R.n92 SUB 3.38fF
C120 SD1R.n93 SUB 3.38fF
C121 SD1R.n94 SUB 3.38fF
C122 SD1R.n95 SUB 3.38fF
C123 SD1R.n96 SUB 3.38fF
C124 SD1R.n97 SUB 3.38fF
C125 SD1R.n98 SUB 3.38fF
C126 SD1R.t55 SUB 3.07fF $ **FLOATING
C127 SD1R.n99 SUB 9.18fF
C128 SD1R.n100 SUB 4.03fF
C129 SD1R.n101 SUB 4.03fF
C130 SD1R.n102 SUB 4.03fF
C131 SD1R.n103 SUB 4.03fF
C132 SD1R.n104 SUB 4.03fF
C133 SD1R.n105 SUB 4.03fF
C134 SD1R.n106 SUB 3.38fF
C135 SD1R.n107 SUB 4.03fF
C136 SD1R.n108 SUB 4.03fF
C137 SD1R.n109 SUB 4.03fF
C138 SD1R.n110 SUB 4.03fF
C139 SD1R.n111 SUB 4.03fF
C140 SD1R.n112 SUB 3.92fF
C141 SD1R.n113 SUB 3.36fF
C142 SD1R.n114 SUB 3.54fF
C143 SD1R.n115 SUB 90.05fF
C144 SD1R.n116 SUB 180.05fF
C145 SD1R.n117 SUB 101.39fF
C146 SD2R.n0 SUB 15.12fF
C147 SD2R.n1 SUB 13.60fF
C148 SD2R.n2 SUB 70.61fF
C149 SD2R.n3 SUB 15.12fF
C150 SD2R.n4 SUB 13.60fF
C151 SD2R.n5 SUB 70.61fF
C152 SD2R.n6 SUB 15.12fF
C153 SD2R.n7 SUB 13.60fF
C154 SD2R.n8 SUB 70.61fF
C155 SD2R.n9 SUB 15.12fF
C156 SD2R.n10 SUB 90.36fF
C157 SD2R.n11 SUB 19.63fF
C158 SD2R.n12 SUB 3.81fF
C159 SD2R.n13 SUB 3.81fF
C160 SD2R.n14 SUB 3.81fF
C161 SD2R.n15 SUB 3.84fF
C162 SD2R.n16 SUB 3.68fF
C163 SD2R.n17 SUB 3.68fF
C164 SD2R.n18 SUB 3.68fF
C165 SD2R.n19 SUB 3.68fF
C166 SD2R.n20 SUB 3.81fF
C167 SD2R.n21 SUB 3.81fF
C168 SD2R.n22 SUB 3.81fF
C169 SD2R.n23 SUB 3.81fF
C170 SD2R.n24 SUB 3.81fF
C171 SD2R.n25 SUB 3.81fF
C172 SD2R.n26 SUB 3.84fF
C173 SD2R.n27 SUB 3.81fF
C174 SD2R.n28 SUB 3.81fF
C175 SD2R.n29 SUB 3.81fF
C176 SD2R.n30 SUB 3.84fF
C177 SD2R.n31 SUB 3.68fF
C178 SD2R.n32 SUB 3.68fF
C179 SD2R.n33 SUB 3.68fF
C180 SD2R.n34 SUB 3.68fF
C181 SD2R.n35 SUB 3.81fF
C182 SD2R.n36 SUB 3.81fF
C183 SD2R.n37 SUB 3.81fF
C184 SD2R.n38 SUB 3.81fF
C185 SD2R.n39 SUB 3.81fF
C186 SD2R.n40 SUB 3.81fF
C187 SD2R.n41 SUB 3.84fF
C188 SD2R.n42 SUB 3.68fF
C189 SD2R.n43 SUB 3.68fF
C190 SD2R.n44 SUB 3.68fF
C191 SD2R.n45 SUB 3.68fF
C192 SD2R.n46 SUB 3.81fF
C193 SD2R.n47 SUB 3.81fF
C194 SD2R.n48 SUB 3.81fF
C195 SD2R.n49 SUB 3.81fF
C196 SD2R.n50 SUB 3.81fF
C197 SD2R.n51 SUB 3.81fF
C198 SD2R.n52 SUB 3.84fF
C199 SD2R.n53 SUB 3.81fF
C200 SD2R.n54 SUB 3.81fF
C201 SD2R.n55 SUB 3.81fF
C202 SD2R.n56 SUB 3.84fF
C203 SD2R.n57 SUB 122.36fF
C204 SD2R.n58 SUB 3.81fF
C205 SD2R.n59 SUB 3.81fF
C206 SD2R.n60 SUB 3.81fF
C207 SD2R.n61 SUB 3.81fF
C208 SD2R.n62 SUB 3.81fF
C209 SD2R.n63 SUB 3.81fF
C210 SD2R.n64 SUB 3.84fF
C211 SD2R.n65 SUB 3.68fF
C212 SD2R.n66 SUB 3.68fF
C213 SD2R.n67 SUB 3.68fF
C214 SD2R.n68 SUB 3.68fF
C215 SD2R.n69 SUB 3.81fF
C216 SD2R.n70 SUB 3.81fF
C217 SD2R.n71 SUB 3.84fF
C218 SD2R.n72 SUB 3.81fF
C219 SD2R.n73 SUB 85.31fF
C220 SD2R.n74 SUB 93.44fF
C221 SD2L.n0 SUB 3.53fF
C222 SD2L.t69 SUB 3.12fF $ **FLOATING
C223 SD2L.n1 SUB 3.53fF
C224 SD2L.n2 SUB 3.53fF
C225 SD2L.n3 SUB 3.56fF
C226 SD2L.n4 SUB 3.56fF
C227 SD2L.n5 SUB 3.56fF
C228 SD2L.n6 SUB 3.56fF
C229 SD2L.n7 SUB 3.56fF
C230 SD2L.n8 SUB 3.56fF
C231 SD2L.n9 SUB 3.56fF
C232 SD2L.n10 SUB 3.56fF
C233 SD2L.n11 SUB 3.56fF
C234 SD2L.n12 SUB 3.56fF
C235 SD2L.n13 SUB 3.56fF
C236 SD2L.t110 SUB 3.23fF $ **FLOATING
C237 SD2L.n14 SUB 9.69fF
C238 SD2L.n15 SUB 4.24fF
C239 SD2L.n16 SUB 4.24fF
C240 SD2L.n17 SUB 4.24fF
C241 SD2L.n18 SUB 4.24fF
C242 SD2L.n19 SUB 4.24fF
C243 SD2L.n20 SUB 4.24fF
C244 SD2L.n21 SUB 4.24fF
C245 SD2L.n22 SUB 4.24fF
C246 SD2L.n23 SUB 4.24fF
C247 SD2L.n24 SUB 3.62fF
C248 SD2L.n25 SUB 69.17fF
C249 SD2L.t34 SUB 3.11fF $ **FLOATING
C250 SD2L.n26 SUB 3.56fF
C251 SD2L.n27 SUB 3.56fF
C252 SD2L.n28 SUB 3.56fF
C253 SD2L.n29 SUB 3.56fF
C254 SD2L.n30 SUB 3.56fF
C255 SD2L.n31 SUB 3.56fF
C256 SD2L.n32 SUB 3.56fF
C257 SD2L.n33 SUB 3.56fF
C258 SD2L.n34 SUB 3.56fF
C259 SD2L.n35 SUB 3.56fF
C260 SD2L.n36 SUB 3.56fF
C261 SD2L.t30 SUB 3.23fF $ **FLOATING
C262 SD2L.n37 SUB 9.69fF
C263 SD2L.n38 SUB 4.24fF
C264 SD2L.n39 SUB 4.24fF
C265 SD2L.n40 SUB 4.24fF
C266 SD2L.n41 SUB 4.24fF
C267 SD2L.n42 SUB 4.24fF
C268 SD2L.n43 SUB 4.24fF
C269 SD2L.n44 SUB 4.24fF
C270 SD2L.n45 SUB 4.24fF
C271 SD2L.n46 SUB 4.24fF
C272 SD2L.n47 SUB 3.62fF
C273 SD2L.n48 SUB 3.53fF
C274 SD2L.n49 SUB 3.53fF
C275 SD2L.n50 SUB 3.53fF
C276 SD2L.n51 SUB 69.18fF
C277 SD2L.t77 SUB 3.11fF $ **FLOATING
C278 SD2L.n52 SUB 3.56fF
C279 SD2L.n53 SUB 3.56fF
C280 SD2L.n54 SUB 3.56fF
C281 SD2L.n55 SUB 3.56fF
C282 SD2L.n56 SUB 3.56fF
C283 SD2L.n57 SUB 3.56fF
C284 SD2L.n58 SUB 3.56fF
C285 SD2L.n59 SUB 3.56fF
C286 SD2L.n60 SUB 3.56fF
C287 SD2L.n61 SUB 3.56fF
C288 SD2L.n62 SUB 3.56fF
C289 SD2L.t70 SUB 3.23fF $ **FLOATING
C290 SD2L.n63 SUB 9.69fF
C291 SD2L.n64 SUB 4.24fF
C292 SD2L.n65 SUB 4.24fF
C293 SD2L.n66 SUB 4.24fF
C294 SD2L.n67 SUB 4.24fF
C295 SD2L.n68 SUB 4.24fF
C296 SD2L.n69 SUB 4.24fF
C297 SD2L.n70 SUB 4.24fF
C298 SD2L.n71 SUB 4.24fF
C299 SD2L.n72 SUB 4.24fF
C300 SD2L.n73 SUB 3.62fF
C301 SD2L.n74 SUB 3.53fF
C302 SD2L.n75 SUB 3.53fF
C303 SD2L.n76 SUB 3.53fF
C304 SD2L.n77 SUB 69.18fF
C305 SD2L.n78 SUB 3.53fF
C306 SD2L.t41 SUB 3.11fF $ **FLOATING
C307 SD2L.n79 SUB 3.56fF
C308 SD2L.n80 SUB 3.56fF
C309 SD2L.n81 SUB 3.56fF
C310 SD2L.n82 SUB 3.56fF
C311 SD2L.n83 SUB 3.56fF
C312 SD2L.n84 SUB 3.56fF
C313 SD2L.n85 SUB 3.56fF
C314 SD2L.n86 SUB 3.56fF
C315 SD2L.n87 SUB 3.56fF
C316 SD2L.n88 SUB 3.56fF
C317 SD2L.n89 SUB 3.56fF
C318 SD2L.t36 SUB 3.23fF $ **FLOATING
C319 SD2L.n90 SUB 9.69fF
C320 SD2L.n91 SUB 4.24fF
C321 SD2L.n92 SUB 4.24fF
C322 SD2L.n93 SUB 4.24fF
C323 SD2L.n94 SUB 4.24fF
C324 SD2L.n95 SUB 4.24fF
C325 SD2L.n96 SUB 4.24fF
C326 SD2L.n97 SUB 4.24fF
C327 SD2L.n98 SUB 4.24fF
C328 SD2L.n99 SUB 4.24fF
C329 SD2L.n100 SUB 3.62fF
C330 SD2L.n101 SUB 3.53fF
C331 SD2L.n102 SUB 3.53fF
C332 SD2L.n103 SUB 88.59fF
C333 SD2L.n104 SUB 167.69fF
C334 SD2L.n105 SUB 103.77fF
C335 SD2L.n106 SUB 82.30fF
C336 SD1L.n0 SUB 15.64fF
C337 SD1L.n1 SUB 18.70fF
C338 SD1L.n2 SUB 20.32fF
C339 SD1L.n3 SUB 18.70fF
C340 SD1L.n4 SUB 15.64fF
C341 SD1L.n5 SUB 18.70fF
C342 SD1L.n6 SUB 15.64fF
C343 SD1L.n7 SUB 18.70fF
C344 SD1L.n8 SUB 52.04fF
C345 SD1L.n9 SUB 9.35fF
C346 SD1L.n10 SUB 47.37fF
C347 SD1L.n11 SUB 9.35fF
C348 SD1L.n12 SUB 79.67fF
C349 SD1L.n13 SUB 9.35fF
C350 SD1L.n14 SUB 47.37fF
C351 SD1L.n15 SUB 3.93fF
C352 SD1L.n16 SUB 3.93fF
C353 SD1L.n17 SUB 3.93fF
C354 SD1L.n18 SUB 3.93fF
C355 SD1L.n19 SUB 3.93fF
C356 SD1L.n20 SUB 3.93fF
C357 SD1L.n21 SUB 3.93fF
C358 SD1L.n22 SUB 3.93fF
C359 SD1L.n23 SUB 3.93fF
C360 SD1L.n24 SUB 3.93fF
C361 SD1L.n25 SUB 3.96fF
C362 SD1L.n26 SUB 3.80fF
C363 SD1L.n27 SUB 3.80fF
C364 SD1L.n28 SUB 3.80fF
C365 SD1L.n29 SUB 3.80fF
C366 SD1L.n30 SUB 3.93fF
C367 SD1L.n31 SUB 3.93fF
C368 SD1L.n32 SUB 3.93fF
C369 SD1L.n33 SUB 3.93fF
C370 SD1L.n34 SUB 3.93fF
C371 SD1L.n35 SUB 3.93fF
C372 SD1L.n36 SUB 3.93fF
C373 SD1L.n37 SUB 3.93fF
C374 SD1L.n38 SUB 3.93fF
C375 SD1L.n39 SUB 3.93fF
C376 SD1L.n40 SUB 3.96fF
C377 SD1L.n41 SUB 3.80fF
C378 SD1L.n42 SUB 3.80fF
C379 SD1L.n43 SUB 3.80fF
C380 SD1L.n44 SUB 3.79fF
C381 SD1L.n45 SUB 3.93fF
C382 SD1L.n46 SUB 3.93fF
C383 SD1L.n47 SUB 3.93fF
C384 SD1L.n48 SUB 3.93fF
C385 SD1L.n49 SUB 3.93fF
C386 SD1L.n50 SUB 3.93fF
C387 SD1L.n51 SUB 3.93fF
C388 SD1L.n52 SUB 3.93fF
C389 SD1L.n53 SUB 3.93fF
C390 SD1L.n54 SUB 3.93fF
C391 SD1L.n55 SUB 3.96fF
C392 SD1L.n56 SUB 3.80fF
C393 SD1L.n57 SUB 3.80fF
C394 SD1L.n58 SUB 3.80fF
C395 SD1L.n59 SUB 3.79fF
C396 SD1L.n60 SUB 97.62fF
C397 SD1L.n61 SUB 3.80fF
C398 SD1L.n62 SUB 3.80fF
C399 SD1L.n63 SUB 3.79fF
C400 SD1L.n64 SUB 3.80fF
C401 SD1L.n65 SUB 3.93fF
C402 SD1L.n66 SUB 3.93fF
C403 SD1L.n67 SUB 3.93fF
C404 SD1L.n68 SUB 3.93fF
C405 SD1L.n69 SUB 3.93fF
C406 SD1L.n70 SUB 3.93fF
C407 SD1L.n71 SUB 3.93fF
C408 SD1L.n72 SUB 3.93fF
C409 SD1L.n73 SUB 3.93fF
C410 SD1L.n74 SUB 3.96fF
C411 SD1L.n75 SUB 3.93fF
C412 SD1L.n76 SUB 67.97fF
C413 SD1L.n77 SUB 75.99fF
