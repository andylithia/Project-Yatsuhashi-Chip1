* NGSPICE file created from cascode_flat.ext - technology: sky130A

X0 SD4R.t119 G34R SD3R.t75 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X1 SD1L.t119 G12L SD2L.t224 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X2 SD1R.t119 G12R SD2R.t155 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X3 SD3L.t239 G23L SD2L.t59 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X4 SD3L.t238 G23L SD2L.t58 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X5 SD1L.t118 G12L SD2L.t223 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X6 SD3R.t123 G23R SD2R.t119 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X7 SD4L.t119 G34L SD3L.t19 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X8 SD4L.t118 G34L SD3L.t86 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X9 SD4L.t117 G34L SD3L.t27 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X10 SD4R.t118 G34R SD3R.t74 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X11 SD2L.t81 G23L SD3L.t237 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X12 SD3R.t47 G34R SD4R.t117 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X13 SD3R.t122 G23R SD2R.t118 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X14 SD3L.t236 G23L SD2L.t80 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X15 SD1L.t117 G12L SD2L.t131 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X16 SD3L.t107 G34L SD4L.t116 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X17 SD1L.t116 G12L SD2L.t130 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X18 SD3R.t175 G23R SD2R.t117 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X19 SD3R.t46 G34R SD4R.t116 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X20 SD2R.t138 G12R SD1R.t118 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X21 SD3R.t174 G23R SD2R.t116 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X22 SD1L.t115 G12L SD2L.t149 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X23 SD3R.t63 G34R SD4R.t115 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X24 SD3R.t62 G34R SD4R.t114 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X25 SD3R.t157 G23R SD2R.t115 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X26 SD1L.t114 G12L SD2L.t148 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X27 SD4L.t115 G34L SD3L.t49 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X28 SD2R.t114 G23R SD3R.t156 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X29 SD3R.t57 G34R SD4R.t113 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X30 SD2R.t182 G12R SD1R.t117 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X31 SD2R.t219 G12R SD1R.t116 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X32 SD2R.t236 G12R SD1R.t115 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X33 SD3R.t159 G23R SD2R.t113 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X34 SD1R.t114 G12R SD2R.t160 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X35 SD3L.t235 G23L SD2L.t103 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X36 SD4L.t114 G34L SD3L.t0 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X37 SD3R.t56 G34R SD4R.t112 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X38 SD2R.t112 G23R SD3R.t158 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X39 SD2R.t161 G12R SD1R.t113 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X40 SD2L.t188 G12L SD1L.t113 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X41 SD3R.t59 G34R SD4R.t111 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X42 SD2L.t187 G12L SD1L.t112 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X43 SD3R.t207 G23R SD2R.t111 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X44 SD3R.t206 G23R SD2R.t110 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X45 SD4L.t113 G34L SD3L.t69 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X46 SD4L.t112 G34L SD3L.t61 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X47 SD3L.t234 G23L SD2L.t102 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X48 SD2L.t99 G23L SD3L.t233 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X49 SD2R.t109 G23R SD3R.t139 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X50 SD4R.t110 G34R SD3R.t58 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X51 SD2L.t182 G12L SD1L.t111 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X52 SD2L.t98 G23L SD3L.t232 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X53 SD2L.t119 G23L SD3L.t231 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X54 SD3L.t63 G34L SD4L.t111 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X55 SD2R.t108 G23R SD3R.t138 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X56 SD2L.t181 G12L SD1L.t110 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X57 SD4R.t109 G34R SD3R.t115 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X58 SD3L.t73 G34L SD4L.t110 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X59 SD1L.t109 G12L SD2L.t212 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X60 SD4L.t109 G34L SD3L.t79 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X61 SD4R.t108 G34R SD3R.t114 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X62 SD2L.t118 G23L SD3L.t230 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X63 SD2L.t211 G12L SD1L.t108 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X64 SD2L.t91 G23L SD3L.t229 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X65 SD2L.t202 G12L SD1L.t107 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X66 SD3R.t179 G23R SD2R.t107 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X67 SD4L.t108 G34L SD3L.t103 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X68 SD4R.t107 G34R SD3R.t41 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X69 SD2L.t90 G23L SD3L.t228 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X70 SD4R.t106 G34R SD3R.t40 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X71 SD2L.t13 G23L SD3L.t227 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X72 SD4L.t107 G34L SD3L.t115 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X73 SD3R.t23 G34R SD4R.t105 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X74 SD4R.t104 G34R SD3R.t22 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X75 SD3R.t51 G34R SD4R.t103 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X76 SD2R.t163 G12R SD1R.t112 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X77 SD2L.t201 G12L SD1L.t106 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X78 SD3R.t178 G23R SD2R.t106 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X79 SD1L.t105 G12L SD2L.t129 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X80 SD3L.t226 G23L SD2L.t12 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X81 SD3R.t221 G23R SD2R.t105 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X82 SD1L.t104 G12L SD2L.t128 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X83 SD1L.t103 G12L SD2L.t200 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X84 SD4L.t106 G34L SD3L.t98 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X85 SD2R.t232 G12R SD1R.t111 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X86 SD3R.t220 G23R SD2R.t104 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X87 SD4L.t105 G34L SD3L.t38 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X88 SD3R.t50 G34R SD4R.t102 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X89 SD1R.t110 G12R SD2R.t213 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X90 SD3L.t106 G34L SD4L.t104 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X91 SD3R.t93 G34R SD4R.t101 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X92 SD3R.t121 G23R SD2R.t103 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X93 SD3R.t120 G23R SD2R.t102 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X94 SD3L.t225 G23L SD2L.t101 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X95 SD1L.t102 G12L SD2L.t199 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X96 SD1R.t109 G12R SD2R.t168 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X97 SD2R.t180 G12R SD1R.t108 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X98 SD2L.t100 G23L SD3L.t224 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X99 SD3R.t92 G34R SD4R.t100 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X100 SD3R.t53 G34R SD4R.t99 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X101 SD3L.t50 G34L SD4L.t103 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X102 SD3L.t117 G34L SD4L.t102 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X103 SD3L.t44 G34L SD4L.t101 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X104 SD3R.t52 G34R SD4R.t98 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X105 SD3L.t223 G23L SD2L.t71 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X106 SD3L.t222 G23L SD2L.t70 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X107 SD1R.t107 G12R SD2R.t197 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X108 SD1R.t106 G12R SD2R.t169 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X109 SD1L.t101 G12L SD2L.t123 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X110 SD3R.t129 G23R SD2R.t101 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X111 SD2R.t167 G12R SD1R.t105 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X112 SD2L.t69 G23L SD3L.t221 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X113 SD2L.t68 G23L SD3L.t220 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X114 SD2L.t122 G12L SD1L.t100 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X115 SD3L.t14 G34L SD4L.t100 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X116 SD3L.t60 G34L SD4L.t99 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X117 SD3L.t219 G23L SD2L.t67 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X118 SD1R.t104 G12R SD2R.t202 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X119 SD4R.t97 G34R SD3R.t49 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X120 SD2L.t198 G12L SD1L.t99 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X121 SD1L.t98 G12L SD2L.t197 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X122 SD1L.t97 G12L SD2L.t222 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X123 SD1R.t103 G12R SD2R.t235 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X124 SD2R.t100 G23R SD3R.t128 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X125 SD2R.t129 G12R SD1R.t102 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X126 SD2R.t233 G12R SD1R.t101 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X127 SD4R.t96 G34R SD3R.t48 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X128 SD2R.t99 G23R SD3R.t183 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X129 SD3L.t218 G23L SD2L.t66 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X130 SD4R.t95 G34R SD3R.t73 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X131 SD4R.t94 G34R SD3R.t72 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X132 SD4L.t98 G34L SD3L.t76 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X133 SD4L.t97 G34L SD3L.t15 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X134 SD2L.t79 G23L SD3L.t217 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X135 SD1R.t100 G12R SD2R.t191 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X136 SD4R.t93 G34R SD3R.t65 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X137 SD2R.t231 G12R SD1R.t99 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X138 SD1R.t98 G12R SD2R.t205 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X139 SD2R.t226 G12R SD1R.t97 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X140 SD1L.t96 G12L SD2L.t221 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X141 SD2R.t98 G23R SD3R.t182 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X142 SD1L.t95 G12L SD2L.t147 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X143 SD1R.t96 G12R SD2R.t149 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X144 SD1L.t94 G12L SD2L.t146 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X145 SD4L.t96 G34L SD3L.t97 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X146 SD4R.t92 G34R SD3R.t64 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X147 SD2R.t97 G23R SD3R.t143 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X148 SD2L.t78 G23L SD3L.t216 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X149 SD2L.t19 G23L SD3L.t215 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X150 SD3L.t2 G34L SD4L.t95 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X151 SD1R.t95 G12R SD2R.t225 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X152 SD3R.t142 G23R SD2R.t96 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X153 SD1R.t94 G12R SD2R.t178 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X154 SD1R.t93 G12R SD2R.t217 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X155 SD4R.t91 G34R SD3R.t99 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X156 SD2R.t176 G12R SD1R.t92 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X157 SD4L.t94 G34L SD3L.t51 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X158 SD2R.t95 G23R SD3R.t181 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X159 SD2R.t94 G23R SD3R.t180 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X160 SD2L.t18 G23L SD3L.t214 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X161 SD3L.t57 G34L SD4L.t93 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X162 SD4R.t90 G34R SD3R.t98 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X163 SD3L.t3 G34L SD4L.t92 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X164 SD3L.t213 G23L SD2L.t15 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X165 SD3L.t212 G23L SD2L.t14 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X166 SD1L.t93 G12L SD2L.t186 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X167 SD4R.t89 G34R SD3R.t61 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X168 SD4R.t88 G34R SD3R.t60 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X169 SD1R.t91 G12R SD2R.t207 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X170 SD3L.t211 G23L SD2L.t93 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X171 SD4L.t91 G34L SD3L.t62 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X172 SD3R.t21 G34R SD4R.t87 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X173 SD2R.t93 G23R SD3R.t131 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X174 SD3R.t130 G23R SD2R.t92 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X175 SD3L.t90 G34L SD4L.t90 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X176 SD1L.t92 G12L SD2L.t185 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X177 SD1L.t91 G12L SD2L.t239 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X178 SD2L.t238 G12L SD1L.t90 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X179 SD2R.t200 G12R SD1R.t90 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X180 SD2L.t210 G12L SD1L.t89 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X181 SD1L.t88 G12L SD2L.t209 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X182 SD2R.t91 G23R SD3R.t133 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X183 SD3R.t20 G34R SD4R.t86 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X184 SD3R.t132 G23R SD2R.t90 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X185 SD3R.t227 G23R SD2R.t89 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X186 SD2L.t232 G12L SD1L.t87 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X187 SD1R.t89 G12R SD2R.t185 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X188 SD3R.t39 G34R SD4R.t85 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X189 SD2R.t221 G12R SD1R.t88 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X190 SD1L.t86 G12L SD2L.t231 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X191 SD2R.t165 G12R SD1R.t87 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X192 SD1R.t86 G12R SD2R.t135 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X193 SD1L.t85 G12L SD2L.t237 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X194 SD3R.t38 G34R SD4R.t84 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X195 SD3R.t43 G34R SD4R.t83 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X196 SD3R.t42 G34R SD4R.t82 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X197 SD2L.t92 G23L SD3L.t210 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X198 SD3R.t226 G23R SD2R.t88 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X199 SD3R.t141 G23R SD2R.t87 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X200 SD4L.t89 G34L SD3L.t20 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X201 SD3R.t101 G34R SD4R.t81 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X202 SD2R.t86 G23R SD3R.t140 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X203 SD2L.t95 G23L SD3L.t209 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X204 SD2L.t236 G12L SD1L.t84 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X205 SD2L.t94 G23L SD3L.t208 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X206 SD3R.t100 G34R SD4R.t80 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X207 SD3R.t67 G34R SD4R.t79 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X208 SD3L.t25 G34L SD4L.t88 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X209 SD3L.t17 G34L SD4L.t87 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X210 SD4L.t86 G34L SD3L.t65 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X211 SD1L.t83 G12L SD2L.t180 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X212 SD1R.t85 G12R SD2R.t216 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X213 SD4R.t78 G34R SD3R.t66 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X214 SD2R.t85 G23R SD3R.t197 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X215 SD2R.t84 G23R SD3R.t196 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X216 SD2L.t179 G12L SD1L.t82 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X217 SD1R.t84 G12R SD2R.t209 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X218 SD2L.t89 G23L SD3L.t207 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X219 SD4R.t77 G34R SD3R.t111 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X220 SD4L.t85 G34L SD3L.t47 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X221 SD4L.t84 G34L SD3L.t88 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X222 SD2L.t196 G12L SD1L.t81 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X223 SD2L.t88 G23L SD3L.t206 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X224 SD2R.t158 G12R SD1R.t83 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X225 SD4L.t83 G34L SD3L.t46 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X226 SD4R.t76 G34R SD3R.t110 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X227 SD2L.t83 G23L SD3L.t205 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X228 SD2L.t82 G23L SD3L.t204 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X229 SD2R.t83 G23R SD3R.t161 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X230 SD2L.t195 G12L SD1L.t80 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X231 SD3R.t160 G23R SD2R.t82 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X232 SD2L.t33 G23L SD3L.t203 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X233 SD3R.t117 G34R SD4R.t75 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X234 SD3R.t171 G23R SD2R.t81 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X235 SD3R.t116 G34R SD4R.t74 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X236 SD3R.t170 G23R SD2R.t80 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X237 SD2L.t145 G12L SD1L.t79 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X238 SD3R.t113 G34R SD4R.t73 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X239 SD3R.t135 G23R SD2R.t79 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X240 SD2L.t32 G23L SD3L.t202 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X241 SD3R.t134 G23R SD2R.t78 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X242 SD1L.t78 G12L SD2L.t144 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X243 SD2L.t17 G23L SD3L.t201 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X244 SD3R.t185 G23R SD2R.t77 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X245 SD2L.t166 G12L SD1L.t77 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X246 SD1R.t82 G12R SD2R.t120 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X247 SD1R.t81 G12R SD2R.t208 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X248 SD1R.t80 G12R SD2R.t139 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X249 SD3R.t184 G23R SD2R.t76 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X250 SD3R.t112 G34R SD4R.t72 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X251 SD3R.t103 G34R SD4R.t71 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X252 SD1R.t79 G12R SD2R.t187 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X253 SD3L.t101 G34L SD4L.t82 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X254 SD3L.t13 G34L SD4L.t81 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X255 SD3L.t200 G23L SD2L.t16 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X256 SD1R.t78 G12R SD2R.t134 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X257 SD4R.t70 G34R SD3R.t102 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X258 SD2R.t75 G23R SD3R.t199 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X259 SD3L.t28 G34L SD4L.t80 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X260 SD2L.t73 G23L SD3L.t199 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X261 SD3L.t198 G23L SD2L.t72 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X262 SD1R.t77 G12R SD2R.t203 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X263 SD3L.t1 G34L SD4L.t79 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X264 SD1R.t76 G12R SD2R.t199 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X265 SD3L.t30 G34L SD4L.t78 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X266 SD3L.t92 G34L SD4L.t77 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X267 SD3L.t197 G23L SD2L.t111 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X268 SD1R.t75 G12R SD2R.t237 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X269 SD2L.t110 G23L SD3L.t196 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X270 SD2R.t74 G23R SD3R.t198 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X271 SD3R.t127 G23R SD2R.t73 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X272 SD3L.t99 G34L SD4L.t76 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X273 SD3L.t102 G34L SD4L.t75 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X274 SD1L.t76 G12L SD2L.t165 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X275 SD1L.t75 G12L SD2L.t230 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X276 SD3R.t95 G34R SD4R.t69 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X277 SD3L.t195 G23L SD2L.t105 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X278 SD4R.t68 G34R SD3R.t94 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X279 SD2R.t210 G12R SD1R.t74 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X280 SD2R.t72 G23R SD3R.t126 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X281 SD2L.t229 G12L SD1L.t74 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X282 SD2R.t71 G23R SD3R.t125 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X283 SD4L.t74 G34L SD3L.t18 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X284 SD4R.t67 G34R SD3R.t97 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X285 SD2L.t235 G12L SD1L.t73 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X286 SD2R.t70 G23R SD3R.t124 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X287 SD3R.t96 G34R SD4R.t66 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X288 SD4L.t73 G34L SD3L.t4 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X289 SD4R.t65 G34R SD3R.t45 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X290 SD2R.t69 G23R SD3R.t187 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X291 SD2R.t174 G12R SD1R.t73 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X292 SD2R.t68 G23R SD3R.t186 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X293 SD2L.t234 G12L SD1L.t72 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X294 SD2L.t164 G12L SD1L.t71 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X295 SD4R.t64 G34R SD3R.t44 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X296 SD2R.t177 G12R SD1R.t72 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X297 SD1R.t71 G12R SD2R.t229 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X298 SD1L.t70 G12L SD2L.t163 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X299 SD1L.t69 G12L SD2L.t220 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X300 SD1R.t70 G12R SD2R.t190 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X301 SD2R.t136 G12R SD1R.t69 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X302 SD4L.t72 G34L SD3L.t6 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X303 SD2L.t219 G12L SD1L.t68 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X304 SD4R.t63 G34R SD3R.t119 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X305 SD4R.t62 G34R SD3R.t118 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X306 SD4L.t71 G34L SD3L.t32 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X307 SD2R.t67 G23R SD3R.t215 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X308 SD2L.t127 G12L SD1L.t67 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X309 SD2R.t66 G23R SD3R.t214 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X310 SD3L.t59 G34L SD4L.t70 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X311 SD1R.t68 G12R SD2R.t215 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X312 SD2R.t201 G12R SD1R.t67 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X313 SD4R.t61 G34R SD3R.t55 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X314 SD3R.t229 G23R SD2R.t65 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X315 SD1R.t66 G12R SD2R.t122 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X316 SD2R.t64 G23R SD3R.t228 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X317 SD1L.t66 G12L SD2L.t126 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X318 SD3L.t26 G34L SD4L.t69 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X319 SD2R.t63 G23R SD3R.t211 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X320 SD3L.t43 G34L SD4L.t68 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X321 SD3R.t54 G34R SD4R.t60 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X322 SD2R.t198 G12R SD1R.t65 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X323 SD1R.t64 G12R SD2R.t123 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X324 SD3R.t210 G23R SD2R.t62 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X325 SD3L.t194 G23L SD2L.t104 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X326 SD1L.t65 G12L SD2L.t143 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X327 SD2L.t61 G23L SD3L.t193 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X328 SD2L.t142 G12L SD1L.t64 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X329 SD3R.t167 G23R SD2R.t61 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X330 SD3R.t71 G34R SD4R.t59 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X331 SD3L.t192 G23L SD2L.t60 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X332 SD1L.t63 G12L SD2L.t184 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X333 SD3R.t70 G34R SD4R.t58 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X334 SD3L.t191 G23L SD2L.t41 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X335 SD3L.t190 G23L SD2L.t40 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X336 SD1L.t62 G12L SD2L.t183 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X337 SD3R.t166 G23R SD2R.t60 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X338 SD1L.t61 G12L SD2L.t178 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X339 SD2R.t59 G23R SD3R.t165 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X340 SD3L.t24 G34L SD4L.t67 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X341 SD3R.t69 G34R SD4R.t57 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X342 SD3L.t189 G23L SD2L.t51 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X343 SD3L.t52 G34L SD4L.t66 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X344 SD3R.t68 G34R SD4R.t56 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X345 SD3L.t188 G23L SD2L.t50 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X346 SD3L.t78 G34L SD4L.t65 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X347 SD3L.t187 G23L SD2L.t21 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X348 SD4R.t55 G34R SD3R.t105 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X349 SD2R.t58 G23R SD3R.t164 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X350 SD3R.t163 G23R SD2R.t57 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X351 SD2R.t173 G12R SD1R.t63 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X352 SD2L.t20 G23L SD3L.t186 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X353 SD2L.t35 G23L SD3L.t185 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X354 SD1L.t60 G12L SD2L.t177 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X355 SD2R.t206 G12R SD1R.t62 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X356 SD4R.t54 G34R SD3R.t104 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X357 SD3L.t83 G34L SD4L.t64 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X358 SD4R.t53 G34R SD3R.t25 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X359 SD2L.t208 G12L SD1L.t59 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X360 SD3R.t24 G34R SD4R.t52 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X361 SD3L.t184 G23L SD2L.t34 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X362 SD4R.t51 G34R SD3R.t77 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X363 SD2R.t56 G23R SD3R.t162 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X364 SD2R.t133 G12R SD1R.t61 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X365 SD2L.t63 G23L SD3L.t183 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X366 SD2L.t62 G23L SD3L.t182 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X367 SD2R.t128 G12R SD1R.t60 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X368 SD2L.t207 G12L SD1L.t58 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X369 SD2L.t85 G23L SD3L.t181 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X370 SD3R.t209 G23R SD2R.t55 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X371 SD2R.t140 G12R SD1R.t59 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X372 SD3R.t208 G23R SD2R.t54 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X373 SD3L.t180 G23L SD2L.t84 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X374 SD4L.t63 G34L SD3L.t100 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X375 SD4R.t50 G34R SD3R.t76 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X376 SD2R.t53 G23R SD3R.t233 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X377 SD2L.t107 G23L SD3L.t179 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X378 SD2R.t172 G12R SD1R.t58 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X379 SD2L.t194 G12L SD1L.t57 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X380 SD2R.t148 G12R SD1R.t57 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X381 SD3L.t178 G23L SD2L.t106 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X382 SD3L.t177 G23L SD2L.t5 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X383 SD4L.t62 G34L SD3L.t110 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X384 SD4L.t61 G34L SD3L.t114 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X385 SD4L.t60 G34L SD3L.t109 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X386 SD4L.t59 G34L SD3L.t23 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X387 SD4R.t49 G34R SD3R.t107 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X388 SD2L.t4 G23L SD3L.t176 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X389 SD2R.t137 G12R SD1R.t56 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X390 SD2R.t211 G12R SD1R.t55 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X391 SD3R.t106 G34R SD4R.t48 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X392 SD1R.t54 G12R SD2R.t192 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X393 SD2L.t193 G12L SD1L.t56 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X394 SD1L.t55 G12L SD2L.t141 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X395 SD1L.t54 G12L SD2L.t140 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X396 SD1L.t53 G12L SD2L.t156 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X397 SD3R.t232 G23R SD2R.t52 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X398 SD1L.t52 G12L SD2L.t155 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X399 SD4L.t58 G34L SD3L.t9 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X400 SD4L.t57 G34L SD3L.t54 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X401 SD4R.t47 G34R SD3R.t109 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X402 SD3R.t219 G23R SD2R.t51 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X403 SD2R.t152 G12R SD1R.t53 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X404 SD3L.t36 G34L SD4L.t56 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X405 SD2L.t75 G23L SD3L.t175 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X406 SD3R.t218 G23R SD2R.t50 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X407 SD3L.t33 G34L SD4L.t55 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X408 SD3L.t89 G34L SD4L.t54 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X409 SD3R.t239 G23R SD2R.t49 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X410 SD3L.t174 G23L SD2L.t74 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X411 SD1R.t52 G12R SD2R.t193 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X412 SD1R.t51 G12R SD2R.t223 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X413 SD1R.t50 G12R SD2R.t220 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X414 SD3R.t108 G34R SD4R.t46 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X415 SD2L.t23 G23L SD3L.t173 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X416 SD3R.t238 G23R SD2R.t48 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X417 SD2L.t22 G23L SD3L.t172 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X418 SD3R.t237 G23R SD2R.t47 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X419 SD2L.t154 G12L SD1L.t51 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X420 SD3R.t79 G34R SD4R.t45 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X421 SD3L.t41 G34L SD4L.t53 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X422 SD3L.t70 G34L SD4L.t52 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X423 SD4R.t44 G34R SD3R.t78 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X424 SD3L.t48 G34L SD4L.t51 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X425 SD3L.t171 G23L SD2L.t43 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X426 SD1R.t49 G12R SD2R.t222 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X427 SD1R.t48 G12R SD2R.t212 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X428 SD4L.t50 G34L SD3L.t37 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X429 SD4R.t43 G34R SD3R.t19 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X430 SD2R.t238 G12R SD1R.t47 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X431 SD1L.t50 G12L SD2L.t153 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X432 SD2R.t46 G23R SD3R.t236 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X433 SD2L.t158 G12L SD1L.t49 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X434 SD2R.t214 G12R SD1R.t46 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X435 SD3R.t235 G23R SD2R.t45 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X436 SD3L.t170 G23L SD2L.t42 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X437 SD3L.t169 G23L SD2L.t53 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X438 SD4L.t49 G34L SD3L.t22 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X439 SD4L.t48 G34L SD3L.t58 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X440 SD4L.t47 G34L SD3L.t111 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X441 SD2R.t44 G23R SD3R.t234 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X442 SD2R.t228 G12R SD1R.t45 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X443 SD2L.t157 G12L SD1L.t48 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X444 SD3R.t217 G23R SD2R.t43 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X445 SD3R.t216 G23R SD2R.t42 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X446 SD2R.t41 G23R SD3R.t231 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X447 SD3L.t168 G23L SD2L.t52 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X448 SD2R.t40 G23R SD3R.t230 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X449 SD4R.t42 G34R SD3R.t18 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X450 SD2L.t7 G23L SD3L.t167 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X451 SD2L.t6 G23L SD3L.t166 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X452 SD2L.t228 G12L SD1L.t47 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X453 SD4R.t41 G34R SD3R.t17 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X454 SD1L.t46 G12L SD2L.t227 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X455 SD1R.t44 G12R SD2R.t204 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X456 SD2R.t39 G23R SD3R.t213 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X457 SD1L.t45 G12L SD2L.t226 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X458 SD2L.t225 G12L SD1L.t44 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X459 SD4R.t40 G34R SD3R.t16 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X460 SD3L.t113 G34L SD4L.t46 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X461 SD1L.t43 G12L SD2L.t135 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X462 SD1R.t43 G12R SD2R.t224 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X463 SD1R.t42 G12R SD2R.t124 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X464 SD2R.t218 G12R SD1R.t41 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X465 SD4R.t39 G34R SD3R.t91 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X466 SD2R.t38 G23R SD3R.t212 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X467 SD2R.t37 G23R SD3R.t155 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X468 SD2R.t36 G23R SD3R.t154 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X469 SD3L.t82 G34L SD4L.t45 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X470 SD4R.t38 G34R SD3R.t90 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X471 SD3L.t29 G34L SD4L.t44 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X472 SD4R.t37 G34R SD3R.t89 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X473 SD3L.t165 G23L SD2L.t113 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X474 SD1R.t40 G12R SD2R.t186 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X475 SD1R.t39 G12R SD2R.t162 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X476 SD3L.t164 G23L SD2L.t112 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X477 SD3L.t163 G23L SD2L.t29 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X478 SD1L.t42 G12L SD2L.t134 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X479 SD4R.t36 G34R SD3R.t88 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X480 SD4R.t35 G34R SD3R.t35 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X481 SD4L.t43 G34L SD3L.t84 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X482 SD2R.t35 G23R SD3R.t203 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X483 SD2R.t34 G23R SD3R.t202 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X484 SD3L.t67 G34L SD4L.t42 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X485 SD2L.t28 G23L SD3L.t162 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X486 SD2R.t157 G12R SD1R.t38 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X487 SD3R.t34 G34R SD4R.t34 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X488 SD3L.t161 G23L SD2L.t77 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X489 SD3L.t160 G23L SD2L.t76 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X490 SD1L.t41 G12L SD2L.t125 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X491 SD4L.t41 G34L SD3L.t11 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X492 SD2R.t151 G12R SD1R.t37 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X493 SD3L.t116 G34L SD4L.t40 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X494 SD1R.t36 G12R SD2R.t125 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X495 SD3R.t15 G34R SD4R.t33 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X496 SD3R.t201 G23R SD2R.t33 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X497 SD1L.t40 G12L SD2L.t124 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X498 SD3L.t159 G23L SD2L.t115 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X499 SD3L.t158 G23L SD2L.t114 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X500 SD1L.t39 G12L SD2L.t139 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X501 SD3L.t105 G34L SD4L.t39 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X502 SD3L.t157 G23L SD2L.t1 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X503 SD3R.t14 G34R SD4R.t32 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X504 SD3L.t34 G34L SD4L.t38 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X505 SD3L.t55 G34L SD4L.t37 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X506 SD3R.t200 G23R SD2R.t32 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X507 SD3R.t13 G34R SD4R.t31 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X508 SD2R.t31 G23R SD3R.t223 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X509 SD2L.t138 G12L SD1L.t38 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X510 SD2L.t0 G23L SD3L.t156 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X511 SD2L.t176 G12L SD1L.t37 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X512 SD2R.t30 G23R SD3R.t222 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X513 SD2R.t188 G12R SD1R.t35 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X514 SD4R.t30 G34R SD3R.t12 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X515 SD1R.t34 G12R SD2R.t175 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X516 SD2R.t29 G23R SD3R.t225 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X517 SD2R.t28 G23R SD3R.t224 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X518 SD2L.t175 G12L SD1L.t36 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X519 SD2L.t206 G12L SD1L.t35 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X520 SD1L.t34 G12L SD2L.t205 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X521 SD4R.t29 G34R SD3R.t1 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X522 SD2R.t159 G12R SD1R.t33 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X523 SD4L.t36 G34L SD3L.t5 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X524 SD4L.t35 G34L SD3L.t119 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X525 SD4L.t34 G34L SD3L.t104 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X526 SD2R.t27 G23R SD3R.t177 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X527 SD2L.t192 G12L SD1L.t33 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X528 SD2R.t26 G23R SD3R.t176 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X529 SD2R.t25 G23R SD3R.t149 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X530 SD2L.t45 G23L SD3L.t155 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X531 SD1R.t32 G12R SD2R.t126 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X532 SD2R.t171 G12R SD1R.t31 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X533 SD2R.t181 G12R SD1R.t30 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X534 SD2L.t191 G12L SD1L.t32 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X535 SD3L.t154 G23L SD2L.t44 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X536 SD2L.t55 G23L SD3L.t153 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X537 SD3R.t148 G23R SD2R.t24 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X538 SD4L.t33 G34L SD3L.t71 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X539 SD4L.t32 G34L SD3L.t81 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X540 SD4L.t31 G34L SD3L.t12 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X541 SD2L.t54 G23L SD3L.t152 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X542 SD2R.t234 G12R SD1R.t29 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X543 SD2R.t23 G23R SD3R.t145 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X544 SD1R.t28 G12R SD2R.t196 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X545 SD1L.t31 G12L SD2L.t204 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X546 SD4L.t30 G34L SD3L.t16 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X547 SD4L.t29 G34L SD3L.t74 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X548 SD2L.t117 G23L SD3L.t151 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X549 SD2L.t203 G12L SD1L.t30 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X550 SD3L.t150 G23L SD2L.t116 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X551 SD2L.t9 G23L SD3L.t149 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X552 SD3R.t144 G23R SD2R.t22 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X553 SD4L.t28 G34L SD3L.t95 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X554 SD1L.t29 G12L SD2L.t190 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X555 SD2L.t189 G12L SD1L.t28 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X556 SD2L.t137 G12L SD1L.t27 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X557 SD3L.t148 G23L SD2L.t8 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X558 SD3R.t205 G23R SD2R.t21 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X559 SD4R.t28 G34R SD3R.t0 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X560 SD3L.t108 G34L SD4L.t27 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X561 SD3L.t147 G23L SD2L.t25 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X562 SD3R.t33 G34R SD4R.t27 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X563 SD1R.t27 G12R SD2R.t143 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X564 SD1R.t26 G12R SD2R.t141 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X565 SD1L.t26 G12L SD2L.t136 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X566 SD1R.t25 G12R SD2R.t127 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X567 SD4L.t26 G34L SD3L.t96 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X568 SD2R.t144 G12R SD1R.t24 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X569 SD1L.t25 G12L SD2L.t133 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X570 SD3R.t204 G23R SD2R.t20 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X571 SD2R.t19 G23R SD3R.t169 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X572 SD3L.t91 G34L SD4L.t25 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X573 SD3R.t32 G34R SD4R.t26 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X574 SD3L.t146 G23L SD2L.t24 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X575 SD1L.t24 G12L SD2L.t132 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X576 SD2L.t172 G12L SD1L.t23 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X577 SD2L.t171 G12L SD1L.t22 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X578 SD2R.t239 G12R SD1R.t23 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X579 SD2L.t121 G12L SD1L.t21 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X580 SD3R.t87 G34R SD4R.t25 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X581 SD3L.t77 G34L SD4L.t24 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X582 SD3R.t86 G34R SD4R.t24 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X583 SD3L.t145 G23L SD2L.t31 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X584 SD3R.t168 G23R SD2R.t18 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X585 SD3R.t173 G23R SD2R.t17 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X586 SD3L.t144 G23L SD2L.t30 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X587 SD2R.t230 G12R SD1R.t22 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X588 SD4L.t23 G34L SD3L.t31 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X589 SD1R.t21 G12R SD2R.t142 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X590 SD3L.t64 G34L SD4L.t22 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X591 SD1L.t20 G12L SD2L.t120 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X592 SD2L.t47 G23L SD3L.t143 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X593 SD2R.t131 G12R SD1R.t20 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X594 SD2R.t183 G12R SD1R.t19 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X595 SD1R.t18 G12R SD2R.t150 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X596 SD3R.t31 G34R SD4R.t23 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X597 SD3R.t30 G34R SD4R.t22 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X598 SD2L.t46 G23L SD3L.t142 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X599 SD3L.t118 G34L SD4L.t21 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X600 SD3R.t172 G23R SD2R.t16 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X601 SD2R.t15 G23R SD3R.t137 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X602 SD4L.t20 G34L SD3L.t94 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X603 SD3R.t11 G34R SD4R.t21 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X604 SD1L.t19 G12L SD2L.t218 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X605 SD2L.t57 G23L SD3L.t141 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X606 SD4L.t19 G34L SD3L.t45 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X607 SD3R.t10 G34R SD4R.t20 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X608 SD4R.t19 G34R SD3R.t85 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X609 SD2R.t14 G23R SD3R.t136 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X610 SD4L.t18 G34L SD3L.t39 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X611 SD1L.t18 G12L SD2L.t217 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X612 SD2L.t170 G12L SD1L.t17 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X613 SD4R.t18 G34R SD3R.t84 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X614 SD2L.t169 G12L SD1L.t16 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X615 SD2L.t152 G12L SD1L.t15 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X616 SD2L.t56 G23L SD3L.t140 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X617 SD2L.t151 G12L SD1L.t14 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X618 SD2R.t13 G23R SD3R.t189 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X619 SD2L.t160 G12L SD1L.t13 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X620 SD2L.t159 G12L SD1L.t12 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X621 SD4R.t17 G34R SD3R.t5 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X622 SD4R.t16 G34R SD3R.t4 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X623 SD2L.t49 G23L SD3L.t139 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X624 SD2R.t12 G23R SD3R.t188 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X625 SD2L.t48 G23L SD3L.t138 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X626 SD4R.t15 G34R SD3R.t9 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X627 SD2L.t3 G23L SD3L.t137 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X628 SD2L.t2 G23L SD3L.t136 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X629 SD2L.t162 G12L SD1L.t11 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X630 SD3L.t135 G23L SD2L.t87 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X631 SD2R.t11 G23R SD3R.t153 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X632 SD1R.t17 G12R SD2R.t184 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X633 SD3R.t152 G23R SD2R.t10 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X634 SD4R.t14 G34R SD3R.t8 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X635 SD3L.t112 G34L SD4L.t17 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X636 SD4R.t13 G34R SD3R.t83 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X637 SD2L.t86 G23L SD3L.t134 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X638 SD3R.t82 G34R SD4R.t12 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X639 SD3L.t53 G34L SD4L.t16 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X640 SD2R.t156 G12R SD1R.t16 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X641 SD3R.t151 G23R SD2R.t9 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X642 SD1R.t15 G12R SD2R.t194 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X643 SD1L.t10 G12L SD2L.t161 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X644 SD1R.t14 G12R SD2R.t146 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X645 SD3R.t81 G34R SD4R.t11 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X646 SD3R.t80 G34R SD4R.t10 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X647 SD2L.t168 G12L SD1L.t9 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X648 SD3L.t7 G34L SD4L.t15 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X649 SD3R.t150 G23R SD2R.t8 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X650 SD2L.t11 G23L SD3L.t133 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X651 SD3R.t147 G23R SD2R.t7 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X652 SD2R.t227 G12R SD1R.t13 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X653 SD1R.t12 G12R SD2R.t195 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X654 SD3L.t35 G34L SD4L.t14 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X655 SD2R.t145 G12R SD1R.t11 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X656 SD3R.t29 G34R SD4R.t9 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X657 SD3L.t132 G23L SD2L.t10 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X658 SD3L.t131 G23L SD2L.t109 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X659 SD3L.t130 G23L SD2L.t108 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X660 SD1R.t10 G12R SD2R.t166 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X661 SD1R.t9 G12R SD2R.t189 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X662 SD1L.t8 G12L SD2L.t167 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X663 SD3L.t42 G34L SD4L.t13 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X664 SD2R.t6 G23R SD3R.t146 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X665 SD3R.t28 G34R SD4R.t8 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X666 SD3L.t129 G23L SD2L.t27 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X667 SD3L.t128 G23L SD2L.t26 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X668 SD3R.t191 G23R SD2R.t5 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X669 SD1R.t8 G12R SD2R.t164 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X670 SD2R.t4 G23R SD3R.t190 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X671 SD3L.t80 G34L SD4L.t12 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X672 SD2L.t214 G12L SD1L.t7 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X673 SD3L.t127 G23L SD2L.t97 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X674 SD4R.t7 G34R SD3R.t7 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X675 SD3L.t85 G34L SD4L.t11 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X676 SD3R.t6 G34R SD4R.t6 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X677 SD3L.t126 G23L SD2L.t96 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X678 SD1L.t6 G12L SD2L.t213 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X679 SD2L.t37 G23L SD3L.t125 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X680 SD2L.t216 G12L SD1L.t5 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X681 SD2R.t3 G23R SD3R.t195 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X682 SD1L.t4 G12L SD2L.t215 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X683 SD4R.t5 G34R SD3R.t27 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X684 SD3L.t66 G34L SD4L.t10 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X685 SD4R.t4 G34R SD3R.t26 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X686 SD3L.t87 G34L SD4L.t9 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X687 SD3L.t75 G34L SD4L.t8 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X688 SD2L.t174 G12L SD1L.t3 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X689 SD3L.t10 G34L SD4L.t7 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X690 SD3R.t3 G34R SD4R.t3 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X691 SD4L.t6 G34L SD3L.t8 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X692 SD3L.t124 G23L SD2L.t36 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X693 SD4R.t2 G34R SD3R.t2 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X694 SD2L.t173 G12L SD1L.t2 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X695 SD2R.t130 G12R SD1R.t7 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X696 SD2R.t154 G12R SD1R.t6 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X697 SD3R.t194 G23R SD2R.t2 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X698 SD1R.t5 G12R SD2R.t147 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X699 SD4L.t5 G34L SD3L.t72 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X700 SD3L.t123 G23L SD2L.t65 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X701 SD2L.t64 G23L SD3L.t122 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X702 SD3R.t37 G34R SD4R.t1 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X703 SD2R.t170 G12R SD1R.t4 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X704 SD4L.t4 G34L SD3L.t93 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X705 SD3L.t121 G23L SD2L.t39 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X706 SD2R.t1 G23R SD3R.t193 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X707 SD4L.t3 G34L SD3L.t56 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X708 SD4L.t2 G34L SD3L.t68 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X709 SD2R.t121 G12R SD1R.t3 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X710 SD2L.t233 G12L SD1L.t1 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X711 SD4L.t1 G34L SD3L.t40 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X712 SD2R.t0 G23R SD3R.t192 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X713 SD2L.t38 G23L SD3L.t120 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X714 SD2R.t179 G12R SD1R.t2 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X715 SD2R.t153 G12R SD1R.t1 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X716 SD4L.t0 G34L SD3L.t21 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X717 SD3R.t36 G34R SD4R.t0 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X718 SD2R.t132 G12R SD1R.t0 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X719 SD2L.t150 G12L SD1L.t0 a_n13364_5836# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
C0 SD3R SD4R 830.88fF
C1 G34L SD4R 14.35fF
C2 SD3L SD3R 126.14fF
C3 SD4L G34R 16.27fF
C4 SD2L SD2R 126.14fF
C5 G34L SD3L 101.57fF
C6 G23L SD3R 17.37fF
C7 SD4L SD3R 37.66fF
C8 SD3L SD4R 38.12fF
C9 SD2L G12L 95.72fF
C10 G23R SD2R 97.56fF
C11 G34L SD4L 96.22fF
C12 SD2L SD3R 38.67fF
C13 G23L SD3L 95.38fF
C14 SD4L SD4R 62.36fF
C15 SD2L SD1L 837.17fF
C16 SD2R G12R 96.55fF
C17 SD3L SD4L 836.09fF
C18 G23R SD3R 96.55fF
C19 SD2L SD3L 835.89fF
C20 G23L SD2L 101.57fF
C21 SD2R SD1R 831.76fF
C22 G12L G12R 28.25fF
C23 G23R SD3L 16.02fF
C24 G23L G23R 28.25fF
C25 SD1L G12R 16.11fF
C26 G12L SD1R 16.25fF
C27 SD2L G23R 18.09fF
C28 SD1L SD1R 55.20fF
C29 SD2L G12R 16.02fF
C30 SD2L SD1R 38.04fF
C31 SD2R G12L 17.37fF
C32 SD2R SD3R 831.34fF
C33 G34R SD3R 97.56fF
C34 SD2R SD1L 44.36fF
C35 G34L G34R 28.25fF
C36 G12R SD1R 98.95fF
C37 SD3L SD2R 37.51fF
C38 G34R SD4R 94.65fF
C39 G12L SD1L 97.03fF
C40 SD3L G34R 18.09fF
C41 G34L SD3R 14.33fF
C42 G23L SD2R 14.33fF
R0 SD3R.n12 SD3R.t139 1.972
R1 SD3R.n7 SD3R.t48 1.972
R2 SD3R.n3 SD3R.t213 1.972
R3 SD3R.n15 SD3R.t22 1.972
R4 SD3R.n27 SD3R.t220 1.963
R5 SD3R.n28 SD3R.t42 1.963
R6 SD3R.n29 SD3R.t185 1.963
R7 SD3R.n26 SD3R.t23 1.96
R8 SD3R.n22 SD3R.n140 1.435
R9 SD3R.n0 SD3R.n145 1.435
R10 SD3R.n10 SD3R.n112 1.435
R11 SD3R.n24 SD3R.n40 1.435
R12 SD3R.n6 SD3R.n35 1.435
R13 SD3R.n1 SD3R.n69 1.435
R14 SD3R.n23 SD3R.n136 1.428
R15 SD3R.n23 SD3R.n137 1.428
R16 SD3R.n22 SD3R.n138 1.428
R17 SD3R.n22 SD3R.n139 1.428
R18 SD3R.n0 SD3R.n144 1.428
R19 SD3R.n0 SD3R.n143 1.428
R20 SD3R.n0 SD3R.n142 1.428
R21 SD3R.n23 SD3R.n141 1.428
R22 SD3R.n21 SD3R.n102 1.428
R23 SD3R.n21 SD3R.n103 1.428
R24 SD3R.n20 SD3R.n104 1.428
R25 SD3R.n20 SD3R.n105 1.428
R26 SD3R.n11 SD3R.n106 1.428
R27 SD3R.n11 SD3R.n107 1.428
R28 SD3R.n11 SD3R.n108 1.428
R29 SD3R.n11 SD3R.n109 1.428
R30 SD3R.n10 SD3R.n110 1.428
R31 SD3R.n10 SD3R.n111 1.428
R32 SD3R.n25 SD3R.n36 1.428
R33 SD3R.n25 SD3R.n37 1.428
R34 SD3R.n24 SD3R.n38 1.428
R35 SD3R.n24 SD3R.n39 1.428
R36 SD3R.n6 SD3R.n34 1.428
R37 SD3R.n6 SD3R.n33 1.428
R38 SD3R.n6 SD3R.n32 1.428
R39 SD3R.n6 SD3R.n31 1.428
R40 SD3R.n25 SD3R.n30 1.428
R41 SD3R.n19 SD3R.n59 1.428
R42 SD3R.n19 SD3R.n60 1.428
R43 SD3R.n18 SD3R.n61 1.428
R44 SD3R.n18 SD3R.n62 1.428
R45 SD3R.n2 SD3R.n63 1.428
R46 SD3R.n2 SD3R.n64 1.428
R47 SD3R.n2 SD3R.n65 1.428
R48 SD3R.n2 SD3R.n66 1.428
R49 SD3R.n1 SD3R.n67 1.428
R50 SD3R.n1 SD3R.n68 1.428
R51 SD3R.n0 SD3R.n146 1.427
R52 SD3R.n15 SD3R.n84 1.414
R53 SD3R.n15 SD3R.n83 1.414
R54 SD3R.n16 SD3R.n82 1.414
R55 SD3R.n16 SD3R.n81 1.414
R56 SD3R.n16 SD3R.n80 1.414
R57 SD3R.n16 SD3R.n79 1.414
R58 SD3R.n17 SD3R.n78 1.414
R59 SD3R.n17 SD3R.n77 1.414
R60 SD3R.n17 SD3R.n76 1.414
R61 SD3R.n17 SD3R.n75 1.414
R62 SD3R.n26 SD3R.n74 1.414
R63 SD3R.n27 SD3R.n88 1.414
R64 SD3R.n14 SD3R.n89 1.414
R65 SD3R.n14 SD3R.n90 1.414
R66 SD3R.n14 SD3R.n91 1.414
R67 SD3R.n14 SD3R.n92 1.414
R68 SD3R.n13 SD3R.n93 1.414
R69 SD3R.n13 SD3R.n94 1.414
R70 SD3R.n13 SD3R.n95 1.414
R71 SD3R.n13 SD3R.n96 1.414
R72 SD3R.n12 SD3R.n97 1.414
R73 SD3R.n12 SD3R.n98 1.414
R74 SD3R.n28 SD3R.n117 1.414
R75 SD3R.n9 SD3R.n118 1.414
R76 SD3R.n9 SD3R.n119 1.414
R77 SD3R.n9 SD3R.n120 1.414
R78 SD3R.n9 SD3R.n121 1.414
R79 SD3R.n8 SD3R.n122 1.414
R80 SD3R.n8 SD3R.n123 1.414
R81 SD3R.n8 SD3R.n124 1.414
R82 SD3R.n8 SD3R.n125 1.414
R83 SD3R.n7 SD3R.n126 1.414
R84 SD3R.n7 SD3R.n127 1.414
R85 SD3R.n29 SD3R.n45 1.414
R86 SD3R.n5 SD3R.n46 1.414
R87 SD3R.n5 SD3R.n47 1.414
R88 SD3R.n5 SD3R.n48 1.414
R89 SD3R.n5 SD3R.n49 1.414
R90 SD3R.n4 SD3R.n50 1.414
R91 SD3R.n4 SD3R.n51 1.414
R92 SD3R.n4 SD3R.n52 1.414
R93 SD3R.n4 SD3R.n53 1.414
R94 SD3R.n3 SD3R.n54 1.414
R95 SD3R.n3 SD3R.n55 1.414
R96 SD3R.n27 SD3R.n101 1.412
R97 SD3R.n27 SD3R.n100 1.412
R98 SD3R.n27 SD3R.n99 1.412
R99 SD3R.n28 SD3R.n130 1.412
R100 SD3R.n28 SD3R.n129 1.412
R101 SD3R.n28 SD3R.n128 1.412
R102 SD3R.n29 SD3R.n58 1.412
R103 SD3R.n29 SD3R.n57 1.412
R104 SD3R.n29 SD3R.n56 1.412
R105 SD3R.n26 SD3R.n85 1.41
R106 SD3R.n26 SD3R.n86 1.409
R107 SD3R.n26 SD3R.n87 1.409
R108 SD3R.n21 SD3R.n113 1.282
R109 SD3R.n19 SD3R.n70 1.282
R110 SD3R.n21 SD3R.n114 1.28
R111 SD3R.n21 SD3R.n116 1.28
R112 SD3R.n21 SD3R.n115 1.28
R113 SD3R.n25 SD3R.n41 1.28
R114 SD3R.n25 SD3R.n42 1.28
R115 SD3R.n25 SD3R.n43 1.28
R116 SD3R.n25 SD3R.n44 1.28
R117 SD3R.n19 SD3R.n71 1.28
R118 SD3R.n19 SD3R.n73 1.28
R119 SD3R.n19 SD3R.n72 1.28
R120 SD3R.n23 SD3R.n135 1.28
R121 SD3R.n23 SD3R.n134 1.28
R122 SD3R.n23 SD3R.n133 1.28
R123 SD3R.n23 SD3R.n132 1.28
R124 SD3R.n136 SD3R.t114 0.551
R125 SD3R.n136 SD3R.t15 0.551
R126 SD3R.n137 SD3R.t97 0.551
R127 SD3R.n137 SD3R.t71 0.551
R128 SD3R.n138 SD3R.t40 0.551
R129 SD3R.n138 SD3R.t33 0.551
R130 SD3R.n139 SD3R.t76 0.551
R131 SD3R.n139 SD3R.t68 0.551
R132 SD3R.n140 SD3R.t65 0.551
R133 SD3R.n140 SD3R.t28 0.551
R134 SD3R.n145 SD3R.t41 0.551
R135 SD3R.n145 SD3R.t53 0.551
R136 SD3R.n144 SD3R.t78 0.551
R137 SD3R.n144 SD3R.t14 0.551
R138 SD3R.n143 SD3R.t98 0.551
R139 SD3R.n143 SD3R.t11 0.551
R140 SD3R.n142 SD3R.t90 0.551
R141 SD3R.n142 SD3R.t101 0.551
R142 SD3R.n141 SD3R.t49 0.551
R143 SD3R.n141 SD3R.t51 0.551
R144 SD3R.n135 SD3R.t94 0.551
R145 SD3R.n135 SD3R.t47 0.551
R146 SD3R.n134 SD3R.t2 0.551
R147 SD3R.n134 SD3R.t34 0.551
R148 SD3R.n133 SD3R.t66 0.551
R149 SD3R.n133 SD3R.t36 0.551
R150 SD3R.n132 SD3R.t19 0.551
R151 SD3R.n132 SD3R.t106 0.551
R152 SD3R.n84 SD3R.t88 0.551
R153 SD3R.n84 SD3R.t59 0.551
R154 SD3R.n83 SD3R.t61 0.551
R155 SD3R.n83 SD3R.t100 0.551
R156 SD3R.n82 SD3R.t91 0.551
R157 SD3R.n82 SD3R.t79 0.551
R158 SD3R.n81 SD3R.t99 0.551
R159 SD3R.n81 SD3R.t38 0.551
R160 SD3R.n80 SD3R.t73 0.551
R161 SD3R.n80 SD3R.t31 0.551
R162 SD3R.n79 SD3R.t5 0.551
R163 SD3R.n79 SD3R.t92 0.551
R164 SD3R.n78 SD3R.t119 0.551
R165 SD3R.n78 SD3R.t87 0.551
R166 SD3R.n77 SD3R.t1 0.551
R167 SD3R.n77 SD3R.t50 0.551
R168 SD3R.n76 SD3R.t111 0.551
R169 SD3R.n76 SD3R.t112 0.551
R170 SD3R.n75 SD3R.t12 0.551
R171 SD3R.n75 SD3R.t63 0.551
R172 SD3R.n74 SD3R.t27 0.551
R173 SD3R.n74 SD3R.t113 0.551
R174 SD3R.n85 SD3R.t104 0.551
R175 SD3R.n85 SD3R.t81 0.551
R176 SD3R.n86 SD3R.t7 0.551
R177 SD3R.n86 SD3R.t117 0.551
R178 SD3R.n87 SD3R.t105 0.551
R179 SD3R.n87 SD3R.t82 0.551
R180 SD3R.n88 SD3R.t126 0.551
R181 SD3R.n88 SD3R.t122 0.551
R182 SD3R.n89 SD3R.t234 0.551
R183 SD3R.n89 SD3R.t160 0.551
R184 SD3R.n90 SD3R.t190 0.551
R185 SD3R.n90 SD3R.t152 0.551
R186 SD3R.n91 SD3R.t236 0.551
R187 SD3R.n91 SD3R.t142 0.551
R188 SD3R.n92 SD3R.t146 0.551
R189 SD3R.n92 SD3R.t208 0.551
R190 SD3R.n93 SD3R.t165 0.551
R191 SD3R.n93 SD3R.t179 0.551
R192 SD3R.n94 SD3R.t156 0.551
R193 SD3R.n94 SD3R.t238 0.551
R194 SD3R.n95 SD3R.t182 0.551
R195 SD3R.n95 SD3R.t129 0.551
R196 SD3R.n96 SD3R.t145 0.551
R197 SD3R.n96 SD3R.t200 0.551
R198 SD3R.n97 SD3R.t214 0.551
R199 SD3R.n97 SD3R.t209 0.551
R200 SD3R.n98 SD3R.t230 0.551
R201 SD3R.n98 SD3R.t175 0.551
R202 SD3R.n99 SD3R.t136 0.551
R203 SD3R.n99 SD3R.t210 0.551
R204 SD3R.n100 SD3R.t124 0.551
R205 SD3R.n100 SD3R.t174 0.551
R206 SD3R.n101 SD3R.t222 0.551
R207 SD3R.n101 SD3R.t170 0.551
R208 SD3R.n102 SD3R.t149 0.551
R209 SD3R.n102 SD3R.t167 0.551
R210 SD3R.n103 SD3R.t215 0.551
R211 SD3R.n103 SD3R.t127 0.551
R212 SD3R.n104 SD3R.t188 0.551
R213 SD3R.n104 SD3R.t173 0.551
R214 SD3R.n105 SD3R.t228 0.551
R215 SD3R.n105 SD3R.t227 0.551
R216 SD3R.n106 SD3R.t180 0.551
R217 SD3R.n106 SD3R.t172 0.551
R218 SD3R.n107 SD3R.t155 0.551
R219 SD3R.n107 SD3R.t141 0.551
R220 SD3R.n108 SD3R.t131 0.551
R221 SD3R.n108 SD3R.t194 0.551
R222 SD3R.n109 SD3R.t202 0.551
R223 SD3R.n109 SD3R.t216 0.551
R224 SD3R.n110 SD3R.t199 0.551
R225 SD3R.n110 SD3R.t206 0.551
R226 SD3R.n111 SD3R.t169 0.551
R227 SD3R.n111 SD3R.t148 0.551
R228 SD3R.n112 SD3R.t154 0.551
R229 SD3R.n112 SD3R.t226 0.551
R230 SD3R.n113 SD3R.t186 0.551
R231 SD3R.n113 SD3R.t157 0.551
R232 SD3R.n114 SD3R.t193 0.551
R233 SD3R.n114 SD3R.t134 0.551
R234 SD3R.n116 SD3R.t196 0.551
R235 SD3R.n116 SD3R.t147 0.551
R236 SD3R.n115 SD3R.t231 0.551
R237 SD3R.n115 SD3R.t218 0.551
R238 SD3R.n117 SD3R.t60 0.551
R239 SD3R.n117 SD3R.t10 0.551
R240 SD3R.n118 SD3R.t109 0.551
R241 SD3R.n118 SD3R.t43 0.551
R242 SD3R.n119 SD3R.t8 0.551
R243 SD3R.n119 SD3R.t30 0.551
R244 SD3R.n120 SD3R.t55 0.551
R245 SD3R.n120 SD3R.t56 0.551
R246 SD3R.n121 SD3R.t4 0.551
R247 SD3R.n121 SD3R.t69 0.551
R248 SD3R.n122 SD3R.t118 0.551
R249 SD3R.n122 SD3R.t57 0.551
R250 SD3R.n123 SD3R.t75 0.551
R251 SD3R.n123 SD3R.t103 0.551
R252 SD3R.n124 SD3R.t115 0.551
R253 SD3R.n124 SD3R.t62 0.551
R254 SD3R.n125 SD3R.t17 0.551
R255 SD3R.n125 SD3R.t108 0.551
R256 SD3R.n126 SD3R.t26 0.551
R257 SD3R.n126 SD3R.t80 0.551
R258 SD3R.n127 SD3R.t25 0.551
R259 SD3R.n127 SD3R.t21 0.551
R260 SD3R.n128 SD3R.t83 0.551
R261 SD3R.n128 SD3R.t96 0.551
R262 SD3R.n129 SD3R.t102 0.551
R263 SD3R.n129 SD3R.t37 0.551
R264 SD3R.n130 SD3R.t35 0.551
R265 SD3R.n130 SD3R.t67 0.551
R266 SD3R.n36 SD3R.t16 0.551
R267 SD3R.n36 SD3R.t116 0.551
R268 SD3R.n37 SD3R.t64 0.551
R269 SD3R.n37 SD3R.t20 0.551
R270 SD3R.n38 SD3R.t77 0.551
R271 SD3R.n38 SD3R.t86 0.551
R272 SD3R.n39 SD3R.t72 0.551
R273 SD3R.n39 SD3R.t93 0.551
R274 SD3R.n40 SD3R.t45 0.551
R275 SD3R.n40 SD3R.t32 0.551
R276 SD3R.n35 SD3R.t89 0.551
R277 SD3R.n35 SD3R.t13 0.551
R278 SD3R.n34 SD3R.t74 0.551
R279 SD3R.n34 SD3R.t95 0.551
R280 SD3R.n33 SD3R.t110 0.551
R281 SD3R.n33 SD3R.t3 0.551
R282 SD3R.n32 SD3R.t9 0.551
R283 SD3R.n32 SD3R.t39 0.551
R284 SD3R.n31 SD3R.t107 0.551
R285 SD3R.n31 SD3R.t6 0.551
R286 SD3R.n30 SD3R.t84 0.551
R287 SD3R.n30 SD3R.t29 0.551
R288 SD3R.n41 SD3R.t18 0.551
R289 SD3R.n41 SD3R.t46 0.551
R290 SD3R.n42 SD3R.t58 0.551
R291 SD3R.n42 SD3R.t54 0.551
R292 SD3R.n43 SD3R.t85 0.551
R293 SD3R.n43 SD3R.t52 0.551
R294 SD3R.n44 SD3R.t44 0.551
R295 SD3R.n44 SD3R.t70 0.551
R296 SD3R.n45 SD3R.t128 0.551
R297 SD3R.n45 SD3R.t219 0.551
R298 SD3R.n46 SD3R.t133 0.551
R299 SD3R.n46 SD3R.t232 0.551
R300 SD3R.n47 SD3R.t195 0.551
R301 SD3R.n47 SD3R.t123 0.551
R302 SD3R.n48 SD3R.t198 0.551
R303 SD3R.n48 SD3R.t144 0.551
R304 SD3R.n49 SD3R.t138 0.551
R305 SD3R.n49 SD3R.t184 0.551
R306 SD3R.n50 SD3R.t125 0.551
R307 SD3R.n50 SD3R.t205 0.551
R308 SD3R.n51 SD3R.t137 0.551
R309 SD3R.n51 SD3R.t166 0.551
R310 SD3R.n52 SD3R.t189 0.551
R311 SD3R.n52 SD3R.t204 0.551
R312 SD3R.n53 SD3R.t183 0.551
R313 SD3R.n53 SD3R.t130 0.551
R314 SD3R.n54 SD3R.t153 0.551
R315 SD3R.n54 SD3R.t191 0.551
R316 SD3R.n55 SD3R.t161 0.551
R317 SD3R.n55 SD3R.t237 0.551
R318 SD3R.n56 SD3R.t224 0.551
R319 SD3R.n56 SD3R.t221 0.551
R320 SD3R.n57 SD3R.t158 0.551
R321 SD3R.n57 SD3R.t229 0.551
R322 SD3R.n58 SD3R.t176 0.551
R323 SD3R.n58 SD3R.t120 0.551
R324 SD3R.n59 SD3R.t181 0.551
R325 SD3R.n59 SD3R.t235 0.551
R326 SD3R.n60 SD3R.t233 0.551
R327 SD3R.n60 SD3R.t239 0.551
R328 SD3R.n61 SD3R.t143 0.551
R329 SD3R.n61 SD3R.t132 0.551
R330 SD3R.n62 SD3R.t162 0.551
R331 SD3R.n62 SD3R.t168 0.551
R332 SD3R.n63 SD3R.t177 0.551
R333 SD3R.n63 SD3R.t121 0.551
R334 SD3R.n64 SD3R.t187 0.551
R335 SD3R.n64 SD3R.t201 0.551
R336 SD3R.n65 SD3R.t225 0.551
R337 SD3R.n65 SD3R.t178 0.551
R338 SD3R.n66 SD3R.t197 0.551
R339 SD3R.n66 SD3R.t135 0.551
R340 SD3R.n67 SD3R.t223 0.551
R341 SD3R.n67 SD3R.t150 0.551
R342 SD3R.n68 SD3R.t140 0.551
R343 SD3R.n68 SD3R.t171 0.551
R344 SD3R.n69 SD3R.t164 0.551
R345 SD3R.n69 SD3R.t151 0.551
R346 SD3R.n70 SD3R.t212 0.551
R347 SD3R.n70 SD3R.t159 0.551
R348 SD3R.n71 SD3R.t192 0.551
R349 SD3R.n71 SD3R.t217 0.551
R350 SD3R.n73 SD3R.t203 0.551
R351 SD3R.n73 SD3R.t207 0.551
R352 SD3R.n72 SD3R.t211 0.551
R353 SD3R.n72 SD3R.t163 0.551
R354 SD3R.n146 SD3R.t0 0.551
R355 SD3R.n146 SD3R.t24 0.551
R356 SD3R.n21 SD3R.n28 0.43
R357 SD3R.n148 SD3R.n26 0.35
R358 SD3R.n131 SD3R.n27 0.347
R359 SD3R.n149 SD3R.n29 0.347
R360 SD3R.n150 SD3R.n25 0.224
R361 SD3R.n147 SD3R.n23 0.224
R362 SD3R.n148 SD3R.n147 0.091
R363 SD3R.n19 SD3R.n148 0.08
R364 SD3R SD3R.n150 0.054
R365 SD3R.n131 SD3R.n21 0.05
R366 SD3R.n149 SD3R.n19 0.05
R367 SD3R.n147 SD3R.n131 0.039
R368 SD3R.n150 SD3R.n149 0.039
R369 SD3R.n25 SD3R.n6 0.037
R370 SD3R.n23 SD3R.n0 0.037
R371 SD3R.n17 SD3R.n16 0.028
R372 SD3R.n16 SD3R.n15 0.028
R373 SD3R.n14 SD3R.n13 0.028
R374 SD3R.n13 SD3R.n12 0.028
R375 SD3R.n20 SD3R.n11 0.028
R376 SD3R.n9 SD3R.n8 0.028
R377 SD3R.n8 SD3R.n7 0.028
R378 SD3R.n5 SD3R.n4 0.028
R379 SD3R.n4 SD3R.n3 0.028
R380 SD3R.n18 SD3R.n2 0.028
R381 SD3R.n21 SD3R.n20 0.025
R382 SD3R.n19 SD3R.n18 0.025
R383 SD3R.n26 SD3R.n17 0.022
R384 SD3R.n23 SD3R.n22 0.021
R385 SD3R.n2 SD3R.n1 0.021
R386 SD3R.n25 SD3R.n24 0.021
R387 SD3R.n11 SD3R.n10 0.021
R388 SD3R.n29 SD3R.n5 0.02
R389 SD3R.n28 SD3R.n9 0.02
R390 SD3R.n27 SD3R.n14 0.02
R391 SD4R.n36 SD4R.t31 1.972
R392 SD4R.n11 SD4R.t99 1.972
R393 SD4R.n25 SD4R.t93 1.963
R394 SD4R.n51 SD4R.t65 1.963
R395 SD4R.n91 SD4R.n90 1.435
R396 SD4R.n63 SD4R.n62 1.435
R397 SD4R.n100 SD4R.n80 1.428
R398 SD4R.n99 SD4R.n81 1.428
R399 SD4R.n98 SD4R.n82 1.428
R400 SD4R.n97 SD4R.n83 1.428
R401 SD4R.n96 SD4R.n84 1.428
R402 SD4R.n95 SD4R.n85 1.428
R403 SD4R.n94 SD4R.n86 1.428
R404 SD4R.n93 SD4R.n87 1.428
R405 SD4R.n92 SD4R.n88 1.428
R406 SD4R.n91 SD4R.n89 1.428
R407 SD4R.n72 SD4R.n52 1.428
R408 SD4R.n71 SD4R.n53 1.428
R409 SD4R.n70 SD4R.n54 1.428
R410 SD4R.n69 SD4R.n55 1.428
R411 SD4R.n68 SD4R.n56 1.428
R412 SD4R.n67 SD4R.n57 1.428
R413 SD4R.n66 SD4R.n58 1.428
R414 SD4R.n65 SD4R.n59 1.428
R415 SD4R.n64 SD4R.n60 1.428
R416 SD4R.n63 SD4R.n61 1.428
R417 SD4R.n47 SD4R.n26 1.414
R418 SD4R.n46 SD4R.n27 1.414
R419 SD4R.n45 SD4R.n28 1.414
R420 SD4R.n44 SD4R.n29 1.414
R421 SD4R.n43 SD4R.n30 1.414
R422 SD4R.n42 SD4R.n31 1.414
R423 SD4R.n41 SD4R.n32 1.414
R424 SD4R.n40 SD4R.n33 1.414
R425 SD4R.n39 SD4R.n34 1.414
R426 SD4R.n36 SD4R.n35 1.414
R427 SD4R.n21 SD4R.n0 1.414
R428 SD4R.n20 SD4R.n1 1.414
R429 SD4R.n19 SD4R.n2 1.414
R430 SD4R.n18 SD4R.n3 1.414
R431 SD4R.n17 SD4R.n4 1.414
R432 SD4R.n16 SD4R.n5 1.414
R433 SD4R.n15 SD4R.n6 1.414
R434 SD4R.n14 SD4R.n7 1.414
R435 SD4R.n13 SD4R.n8 1.414
R436 SD4R.n12 SD4R.n9 1.414
R437 SD4R.n11 SD4R.n10 1.414
R438 SD4R.n38 SD4R.n37 1.413
R439 SD4R.n25 SD4R.n24 1.412
R440 SD4R.n25 SD4R.n23 1.412
R441 SD4R.n25 SD4R.n22 1.412
R442 SD4R.n51 SD4R.n50 1.412
R443 SD4R.n51 SD4R.n49 1.412
R444 SD4R.n51 SD4R.n48 1.412
R445 SD4R.n102 SD4R.n101 1.282
R446 SD4R.n106 SD4R.n103 1.28
R447 SD4R.n106 SD4R.n105 1.28
R448 SD4R.n106 SD4R.n104 1.28
R449 SD4R.n78 SD4R.n77 1.279
R450 SD4R.n78 SD4R.n76 1.279
R451 SD4R.n78 SD4R.n75 1.278
R452 SD4R.n74 SD4R.n73 1.278
R453 SD4R.n26 SD4R.t86 0.551
R454 SD4R.n26 SD4R.t40 0.551
R455 SD4R.n27 SD4R.t74 0.551
R456 SD4R.n27 SD4R.t42 0.551
R457 SD4R.n28 SD4R.t116 0.551
R458 SD4R.n28 SD4R.t110 0.551
R459 SD4R.n29 SD4R.t60 0.551
R460 SD4R.n29 SD4R.t19 0.551
R461 SD4R.n30 SD4R.t98 0.551
R462 SD4R.n30 SD4R.t64 0.551
R463 SD4R.n31 SD4R.t58 0.551
R464 SD4R.n31 SD4R.t18 0.551
R465 SD4R.n32 SD4R.t9 0.551
R466 SD4R.n32 SD4R.t49 0.551
R467 SD4R.n33 SD4R.t6 0.551
R468 SD4R.n33 SD4R.t15 0.551
R469 SD4R.n34 SD4R.t85 0.551
R470 SD4R.n34 SD4R.t76 0.551
R471 SD4R.n35 SD4R.t69 0.551
R472 SD4R.n35 SD4R.t37 0.551
R473 SD4R.n48 SD4R.t26 0.551
R474 SD4R.n48 SD4R.t94 0.551
R475 SD4R.n49 SD4R.t101 0.551
R476 SD4R.n49 SD4R.t51 0.551
R477 SD4R.n50 SD4R.t24 0.551
R478 SD4R.n50 SD4R.t92 0.551
R479 SD4R.n0 SD4R.t59 0.551
R480 SD4R.n0 SD4R.t108 0.551
R481 SD4R.n1 SD4R.t33 0.551
R482 SD4R.n1 SD4R.t68 0.551
R483 SD4R.n2 SD4R.t117 0.551
R484 SD4R.n2 SD4R.t2 0.551
R485 SD4R.n3 SD4R.t34 0.551
R486 SD4R.n3 SD4R.t78 0.551
R487 SD4R.n4 SD4R.t0 0.551
R488 SD4R.n4 SD4R.t43 0.551
R489 SD4R.n5 SD4R.t48 0.551
R490 SD4R.n5 SD4R.t97 0.551
R491 SD4R.n6 SD4R.t103 0.551
R492 SD4R.n6 SD4R.t38 0.551
R493 SD4R.n7 SD4R.t81 0.551
R494 SD4R.n7 SD4R.t90 0.551
R495 SD4R.n8 SD4R.t21 0.551
R496 SD4R.n8 SD4R.t28 0.551
R497 SD4R.n9 SD4R.t52 0.551
R498 SD4R.n9 SD4R.t44 0.551
R499 SD4R.n10 SD4R.t32 0.551
R500 SD4R.n10 SD4R.t107 0.551
R501 SD4R.n22 SD4R.t8 0.551
R502 SD4R.n22 SD4R.t50 0.551
R503 SD4R.n23 SD4R.t56 0.551
R504 SD4R.n23 SD4R.t106 0.551
R505 SD4R.n24 SD4R.t27 0.551
R506 SD4R.n24 SD4R.t67 0.551
R507 SD4R.n80 SD4R.t71 0.551
R508 SD4R.n80 SD4R.t109 0.551
R509 SD4R.n81 SD4R.t113 0.551
R510 SD4R.n81 SD4R.t119 0.551
R511 SD4R.n82 SD4R.t57 0.551
R512 SD4R.n82 SD4R.t62 0.551
R513 SD4R.n83 SD4R.t112 0.551
R514 SD4R.n83 SD4R.t16 0.551
R515 SD4R.n84 SD4R.t22 0.551
R516 SD4R.n84 SD4R.t61 0.551
R517 SD4R.n85 SD4R.t83 0.551
R518 SD4R.n85 SD4R.t14 0.551
R519 SD4R.n86 SD4R.t20 0.551
R520 SD4R.n86 SD4R.t47 0.551
R521 SD4R.n87 SD4R.t79 0.551
R522 SD4R.n87 SD4R.t88 0.551
R523 SD4R.n88 SD4R.t1 0.551
R524 SD4R.n88 SD4R.t35 0.551
R525 SD4R.n89 SD4R.t66 0.551
R526 SD4R.n89 SD4R.t70 0.551
R527 SD4R.n90 SD4R.t82 0.551
R528 SD4R.n90 SD4R.t13 0.551
R529 SD4R.n101 SD4R.t114 0.551
R530 SD4R.n101 SD4R.t41 0.551
R531 SD4R.n103 SD4R.t46 0.551
R532 SD4R.n103 SD4R.t4 0.551
R533 SD4R.n105 SD4R.t10 0.551
R534 SD4R.n105 SD4R.t53 0.551
R535 SD4R.n104 SD4R.t87 0.551
R536 SD4R.n104 SD4R.t96 0.551
R537 SD4R.n75 SD4R.t111 0.551
R538 SD4R.n75 SD4R.t104 0.551
R539 SD4R.n77 SD4R.t80 0.551
R540 SD4R.n77 SD4R.t36 0.551
R541 SD4R.n76 SD4R.t45 0.551
R542 SD4R.n76 SD4R.t89 0.551
R543 SD4R.n52 SD4R.t23 0.551
R544 SD4R.n52 SD4R.t91 0.551
R545 SD4R.n53 SD4R.t100 0.551
R546 SD4R.n53 SD4R.t95 0.551
R547 SD4R.n54 SD4R.t25 0.551
R548 SD4R.n54 SD4R.t17 0.551
R549 SD4R.n55 SD4R.t102 0.551
R550 SD4R.n55 SD4R.t63 0.551
R551 SD4R.n56 SD4R.t72 0.551
R552 SD4R.n56 SD4R.t29 0.551
R553 SD4R.n57 SD4R.t115 0.551
R554 SD4R.n57 SD4R.t77 0.551
R555 SD4R.n58 SD4R.t73 0.551
R556 SD4R.n58 SD4R.t30 0.551
R557 SD4R.n59 SD4R.t11 0.551
R558 SD4R.n59 SD4R.t5 0.551
R559 SD4R.n60 SD4R.t75 0.551
R560 SD4R.n60 SD4R.t54 0.551
R561 SD4R.n61 SD4R.t12 0.551
R562 SD4R.n61 SD4R.t7 0.551
R563 SD4R.n62 SD4R.t105 0.551
R564 SD4R.n62 SD4R.t55 0.551
R565 SD4R.n73 SD4R.t84 0.551
R566 SD4R.n73 SD4R.t39 0.551
R567 SD4R.n37 SD4R.t3 0.551
R568 SD4R.n37 SD4R.t118 0.551
R569 SD4R.n78 SD4R.n51 0.399
R570 SD4R.n79 SD4R.n25 0.347
R571 SD4R.n79 SD4R.n78 0.21
R572 SD4R SD4R.n106 0.112
R573 SD4R.n106 SD4R.n79 0.05
R574 SD4R.n74 SD4R.n72 0.008
R575 SD4R.n21 SD4R.n20 0.007
R576 SD4R.n20 SD4R.n19 0.007
R577 SD4R.n19 SD4R.n18 0.007
R578 SD4R.n18 SD4R.n17 0.007
R579 SD4R.n17 SD4R.n16 0.007
R580 SD4R.n16 SD4R.n15 0.007
R581 SD4R.n15 SD4R.n14 0.007
R582 SD4R.n14 SD4R.n13 0.007
R583 SD4R.n13 SD4R.n12 0.007
R584 SD4R.n12 SD4R.n11 0.007
R585 SD4R.n92 SD4R.n91 0.007
R586 SD4R.n93 SD4R.n92 0.007
R587 SD4R.n94 SD4R.n93 0.007
R588 SD4R.n95 SD4R.n94 0.007
R589 SD4R.n96 SD4R.n95 0.007
R590 SD4R.n97 SD4R.n96 0.007
R591 SD4R.n98 SD4R.n97 0.007
R592 SD4R.n99 SD4R.n98 0.007
R593 SD4R.n100 SD4R.n99 0.007
R594 SD4R.n102 SD4R.n100 0.007
R595 SD4R.n64 SD4R.n63 0.007
R596 SD4R.n65 SD4R.n64 0.007
R597 SD4R.n66 SD4R.n65 0.007
R598 SD4R.n67 SD4R.n66 0.007
R599 SD4R.n68 SD4R.n67 0.007
R600 SD4R.n69 SD4R.n68 0.007
R601 SD4R.n70 SD4R.n69 0.007
R602 SD4R.n71 SD4R.n70 0.007
R603 SD4R.n72 SD4R.n71 0.007
R604 SD4R.n47 SD4R.n46 0.007
R605 SD4R.n46 SD4R.n45 0.007
R606 SD4R.n45 SD4R.n44 0.007
R607 SD4R.n44 SD4R.n43 0.007
R608 SD4R.n43 SD4R.n42 0.007
R609 SD4R.n42 SD4R.n41 0.007
R610 SD4R.n41 SD4R.n40 0.007
R611 SD4R.n40 SD4R.n39 0.007
R612 SD4R.n39 SD4R.n38 0.007
R613 SD4R.n38 SD4R.n36 0.007
R614 SD4R.n25 SD4R.n21 0.006
R615 SD4R.n51 SD4R.n47 0.006
R616 SD4R.n78 SD4R.n74 0.005
R617 SD4R.n106 SD4R.n102 0.004
R618 SD2L.n14 SD2L.t90 1.972
R619 SD2L.n11 SD2L.t171 1.972
R620 SD2L.n9 SD2L.t144 1.972
R621 SD2L.n5 SD2L.t48 1.972
R622 SD2L.n4 SD2L.t187 1.972
R623 SD2L.n2 SD2L.t165 1.972
R624 SD2L.n19 SD2L.t31 1.963
R625 SD2L.n21 SD2L.t105 1.962
R626 SD2L.n0 SD2L.n144 1.435
R627 SD2L.n16 SD2L.n40 1.435
R628 SD2L.n12 SD2L.n69 1.435
R629 SD2L.n7 SD2L.n98 1.435
R630 SD2L.n23 SD2L.n135 1.428
R631 SD2L.n22 SD2L.n136 1.428
R632 SD2L.n22 SD2L.n137 1.428
R633 SD2L.n1 SD2L.n138 1.428
R634 SD2L.n1 SD2L.n139 1.428
R635 SD2L.n1 SD2L.n140 1.428
R636 SD2L.n1 SD2L.n141 1.428
R637 SD2L.n0 SD2L.n142 1.428
R638 SD2L.n0 SD2L.n143 1.428
R639 SD2L.n29 SD2L.n30 1.428
R640 SD2L.n29 SD2L.n31 1.428
R641 SD2L.n28 SD2L.n32 1.428
R642 SD2L.n28 SD2L.n33 1.428
R643 SD2L.n17 SD2L.n34 1.428
R644 SD2L.n17 SD2L.n35 1.428
R645 SD2L.n17 SD2L.n36 1.428
R646 SD2L.n17 SD2L.n37 1.428
R647 SD2L.n16 SD2L.n38 1.428
R648 SD2L.n16 SD2L.n39 1.428
R649 SD2L.n27 SD2L.n59 1.428
R650 SD2L.n27 SD2L.n60 1.428
R651 SD2L.n26 SD2L.n61 1.428
R652 SD2L.n26 SD2L.n62 1.428
R653 SD2L.n13 SD2L.n63 1.428
R654 SD2L.n13 SD2L.n64 1.428
R655 SD2L.n13 SD2L.n65 1.428
R656 SD2L.n13 SD2L.n66 1.428
R657 SD2L.n12 SD2L.n67 1.428
R658 SD2L.n12 SD2L.n68 1.428
R659 SD2L.n25 SD2L.n88 1.428
R660 SD2L.n25 SD2L.n89 1.428
R661 SD2L.n24 SD2L.n90 1.428
R662 SD2L.n24 SD2L.n91 1.428
R663 SD2L.n8 SD2L.n92 1.428
R664 SD2L.n8 SD2L.n93 1.428
R665 SD2L.n8 SD2L.n94 1.428
R666 SD2L.n8 SD2L.n95 1.428
R667 SD2L.n7 SD2L.n96 1.428
R668 SD2L.n7 SD2L.n97 1.428
R669 SD2L.n23 SD2L.n145 1.427
R670 SD2L.n21 SD2L.n45 1.414
R671 SD2L.n21 SD2L.n46 1.414
R672 SD2L.n21 SD2L.n47 1.414
R673 SD2L.n20 SD2L.n48 1.414
R674 SD2L.n20 SD2L.n49 1.414
R675 SD2L.n15 SD2L.n50 1.414
R676 SD2L.n15 SD2L.n51 1.414
R677 SD2L.n15 SD2L.n52 1.414
R678 SD2L.n15 SD2L.n53 1.414
R679 SD2L.n14 SD2L.n54 1.414
R680 SD2L.n14 SD2L.n55 1.414
R681 SD2L.n10 SD2L.n79 1.414
R682 SD2L.n10 SD2L.n80 1.414
R683 SD2L.n11 SD2L.n81 1.414
R684 SD2L.n11 SD2L.n82 1.414
R685 SD2L.n11 SD2L.n83 1.414
R686 SD2L.n9 SD2L.n78 1.414
R687 SD2L.n9 SD2L.n77 1.414
R688 SD2L.n10 SD2L.n76 1.414
R689 SD2L.n10 SD2L.n75 1.414
R690 SD2L.n10 SD2L.n74 1.414
R691 SD2L.n19 SD2L.n103 1.414
R692 SD2L.n19 SD2L.n104 1.414
R693 SD2L.n19 SD2L.n105 1.414
R694 SD2L.n18 SD2L.n106 1.414
R695 SD2L.n18 SD2L.n107 1.414
R696 SD2L.n6 SD2L.n108 1.414
R697 SD2L.n6 SD2L.n109 1.414
R698 SD2L.n6 SD2L.n110 1.414
R699 SD2L.n6 SD2L.n111 1.414
R700 SD2L.n5 SD2L.n112 1.414
R701 SD2L.n5 SD2L.n113 1.414
R702 SD2L.n3 SD2L.n122 1.414
R703 SD2L.n3 SD2L.n123 1.414
R704 SD2L.n4 SD2L.n124 1.414
R705 SD2L.n4 SD2L.n125 1.414
R706 SD2L.n4 SD2L.n126 1.414
R707 SD2L.n2 SD2L.n121 1.414
R708 SD2L.n2 SD2L.n120 1.414
R709 SD2L.n3 SD2L.n119 1.414
R710 SD2L.n3 SD2L.n118 1.414
R711 SD2L.n3 SD2L.n117 1.414
R712 SD2L.n10 SD2L.n87 1.412
R713 SD2L.n10 SD2L.n86 1.412
R714 SD2L.n10 SD2L.n85 1.412
R715 SD2L.n10 SD2L.n84 1.412
R716 SD2L.n19 SD2L.n116 1.412
R717 SD2L.n19 SD2L.n115 1.412
R718 SD2L.n19 SD2L.n114 1.412
R719 SD2L.n3 SD2L.n130 1.412
R720 SD2L.n3 SD2L.n129 1.412
R721 SD2L.n3 SD2L.n128 1.412
R722 SD2L.n3 SD2L.n127 1.412
R723 SD2L.n21 SD2L.n58 1.409
R724 SD2L.n21 SD2L.n57 1.409
R725 SD2L.n21 SD2L.n56 1.409
R726 SD2L.n29 SD2L.n41 1.281
R727 SD2L.n27 SD2L.n70 1.281
R728 SD2L.n25 SD2L.n99 1.281
R729 SD2L.n23 SD2L.n134 1.281
R730 SD2L.n29 SD2L.n42 1.28
R731 SD2L.n29 SD2L.n43 1.28
R732 SD2L.n29 SD2L.n44 1.28
R733 SD2L.n27 SD2L.n71 1.28
R734 SD2L.n27 SD2L.n72 1.28
R735 SD2L.n27 SD2L.n73 1.28
R736 SD2L.n25 SD2L.n100 1.28
R737 SD2L.n25 SD2L.n101 1.28
R738 SD2L.n25 SD2L.n102 1.28
R739 SD2L.n23 SD2L.n133 1.28
R740 SD2L.n23 SD2L.n132 1.28
R741 SD2L.n23 SD2L.n131 1.28
R742 SD2L.n135 SD2L.t76 0.551
R743 SD2L.n135 SD2L.t6 0.551
R744 SD2L.n136 SD2L.t12 0.551
R745 SD2L.n136 SD2L.t98 0.551
R746 SD2L.n137 SD2L.t114 0.551
R747 SD2L.n137 SD2L.t20 0.551
R748 SD2L.n138 SD2L.t41 0.551
R749 SD2L.n138 SD2L.t91 0.551
R750 SD2L.n139 SD2L.t109 0.551
R751 SD2L.n139 SD2L.t63 0.551
R752 SD2L.n140 SD2L.t50 0.551
R753 SD2L.n140 SD2L.t19 0.551
R754 SD2L.n141 SD2L.t27 0.551
R755 SD2L.n141 SD2L.t3 0.551
R756 SD2L.n142 SD2L.t53 0.551
R757 SD2L.n142 SD2L.t83 0.551
R758 SD2L.n143 SD2L.t103 0.551
R759 SD2L.n143 SD2L.t81 0.551
R760 SD2L.n144 SD2L.t10 0.551
R761 SD2L.n144 SD2L.t85 0.551
R762 SD2L.n134 SD2L.t112 0.551
R763 SD2L.n134 SD2L.t94 0.551
R764 SD2L.n133 SD2L.t14 0.551
R765 SD2L.n133 SD2L.t23 0.551
R766 SD2L.n132 SD2L.t106 0.551
R767 SD2L.n132 SD2L.t69 0.551
R768 SD2L.n131 SD2L.t87 0.551
R769 SD2L.n131 SD2L.t47 0.551
R770 SD2L.n30 SD2L.t123 0.551
R771 SD2L.n30 SD2L.t194 0.551
R772 SD2L.n31 SD2L.t143 0.551
R773 SD2L.n31 SD2L.t208 0.551
R774 SD2L.n32 SD2L.t149 0.551
R775 SD2L.n32 SD2L.t181 0.551
R776 SD2L.n33 SD2L.t126 0.551
R777 SD2L.n33 SD2L.t191 0.551
R778 SD2L.n34 SD2L.t134 0.551
R779 SD2L.n34 SD2L.t188 0.551
R780 SD2L.n35 SD2L.t186 0.551
R781 SD2L.n35 SD2L.t157 0.551
R782 SD2L.n36 SD2L.t185 0.551
R783 SD2L.n36 SD2L.t214 0.551
R784 SD2L.n37 SD2L.t132 0.551
R785 SD2L.n37 SD2L.t170 0.551
R786 SD2L.n38 SD2L.t200 0.551
R787 SD2L.n38 SD2L.t164 0.551
R788 SD2L.n39 SD2L.t136 0.551
R789 SD2L.n39 SD2L.t206 0.551
R790 SD2L.n40 SD2L.t130 0.551
R791 SD2L.n40 SD2L.t235 0.551
R792 SD2L.n41 SD2L.t178 0.551
R793 SD2L.n41 SD2L.t151 0.551
R794 SD2L.n42 SD2L.t167 0.551
R795 SD2L.n42 SD2L.t193 0.551
R796 SD2L.n43 SD2L.t153 0.551
R797 SD2L.n43 SD2L.t150 0.551
R798 SD2L.n44 SD2L.t237 0.551
R799 SD2L.n44 SD2L.t195 0.551
R800 SD2L.n58 SD2L.t102 0.551
R801 SD2L.n58 SD2L.t17 0.551
R802 SD2L.n57 SD2L.t52 0.551
R803 SD2L.n57 SD2L.t28 0.551
R804 SD2L.n56 SD2L.t96 0.551
R805 SD2L.n56 SD2L.t38 0.551
R806 SD2L.n45 SD2L.t42 0.551
R807 SD2L.n45 SD2L.t4 0.551
R808 SD2L.n46 SD2L.t74 0.551
R809 SD2L.n46 SD2L.t18 0.551
R810 SD2L.n47 SD2L.t70 0.551
R811 SD2L.n47 SD2L.t107 0.551
R812 SD2L.n48 SD2L.t30 0.551
R813 SD2L.n48 SD2L.t13 0.551
R814 SD2L.n49 SD2L.t101 0.551
R815 SD2L.n49 SD2L.t62 0.551
R816 SD2L.n50 SD2L.t115 0.551
R817 SD2L.n50 SD2L.t45 0.551
R818 SD2L.n51 SD2L.t80 0.551
R819 SD2L.n51 SD2L.t88 0.551
R820 SD2L.n52 SD2L.t97 0.551
R821 SD2L.n52 SD2L.t33 0.551
R822 SD2L.n53 SD2L.t21 0.551
R823 SD2L.n53 SD2L.t86 0.551
R824 SD2L.n54 SD2L.t24 0.551
R825 SD2L.n54 SD2L.t79 0.551
R826 SD2L.n55 SD2L.t51 0.551
R827 SD2L.n55 SD2L.t49 0.551
R828 SD2L.n59 SD2L.t40 0.551
R829 SD2L.n59 SD2L.t56 0.551
R830 SD2L.n60 SD2L.t8 0.551
R831 SD2L.n60 SD2L.t46 0.551
R832 SD2L.n61 SD2L.t104 0.551
R833 SD2L.n61 SD2L.t35 0.551
R834 SD2L.n62 SD2L.t116 0.551
R835 SD2L.n62 SD2L.t119 0.551
R836 SD2L.n63 SD2L.t58 0.551
R837 SD2L.n63 SD2L.t110 0.551
R838 SD2L.n64 SD2L.t29 0.551
R839 SD2L.n64 SD2L.t37 0.551
R840 SD2L.n65 SD2L.t39 0.551
R841 SD2L.n65 SD2L.t73 0.551
R842 SD2L.n66 SD2L.t5 0.551
R843 SD2L.n66 SD2L.t22 0.551
R844 SD2L.n67 SD2L.t65 0.551
R845 SD2L.n67 SD2L.t68 0.551
R846 SD2L.n68 SD2L.t84 0.551
R847 SD2L.n68 SD2L.t75 0.551
R848 SD2L.n69 SD2L.t44 0.551
R849 SD2L.n69 SD2L.t100 0.551
R850 SD2L.n70 SD2L.t108 0.551
R851 SD2L.n70 SD2L.t89 0.551
R852 SD2L.n71 SD2L.t93 0.551
R853 SD2L.n71 SD2L.t2 0.551
R854 SD2L.n72 SD2L.t26 0.551
R855 SD2L.n72 SD2L.t82 0.551
R856 SD2L.n73 SD2L.t1 0.551
R857 SD2L.n73 SD2L.t55 0.551
R858 SD2L.n79 SD2L.t135 0.551
R859 SD2L.n79 SD2L.t159 0.551
R860 SD2L.n80 SD2L.t146 0.551
R861 SD2L.n80 SD2L.t219 0.551
R862 SD2L.n81 SD2L.t177 0.551
R863 SD2L.n81 SD2L.t175 0.551
R864 SD2L.n82 SD2L.t205 0.551
R865 SD2L.n82 SD2L.t173 0.551
R866 SD2L.n83 SD2L.t148 0.551
R867 SD2L.n83 SD2L.t232 0.551
R868 SD2L.n78 SD2L.t226 0.551
R869 SD2L.n78 SD2L.t160 0.551
R870 SD2L.n77 SD2L.t215 0.551
R871 SD2L.n77 SD2L.t234 0.551
R872 SD2L.n76 SD2L.t222 0.551
R873 SD2L.n76 SD2L.t233 0.551
R874 SD2L.n75 SD2L.t183 0.551
R875 SD2L.n75 SD2L.t174 0.551
R876 SD2L.n74 SD2L.t180 0.551
R877 SD2L.n74 SD2L.t210 0.551
R878 SD2L.n84 SD2L.t220 0.551
R879 SD2L.n84 SD2L.t168 0.551
R880 SD2L.n85 SD2L.t128 0.551
R881 SD2L.n85 SD2L.t166 0.551
R882 SD2L.n86 SD2L.t155 0.551
R883 SD2L.n86 SD2L.t137 0.551
R884 SD2L.n87 SD2L.t209 0.551
R885 SD2L.n87 SD2L.t121 0.551
R886 SD2L.n88 SD2L.t231 0.551
R887 SD2L.n88 SD2L.t162 0.551
R888 SD2L.n89 SD2L.t204 0.551
R889 SD2L.n89 SD2L.t138 0.551
R890 SD2L.n90 SD2L.t147 0.551
R891 SD2L.n90 SD2L.t122 0.551
R892 SD2L.n91 SD2L.t161 0.551
R893 SD2L.n91 SD2L.t154 0.551
R894 SD2L.n92 SD2L.t156 0.551
R895 SD2L.n92 SD2L.t236 0.551
R896 SD2L.n93 SD2L.t223 0.551
R897 SD2L.n93 SD2L.t158 0.551
R898 SD2L.n94 SD2L.t125 0.551
R899 SD2L.n94 SD2L.t179 0.551
R900 SD2L.n95 SD2L.t131 0.551
R901 SD2L.n95 SD2L.t182 0.551
R902 SD2L.n96 SD2L.t139 0.551
R903 SD2L.n96 SD2L.t229 0.551
R904 SD2L.n97 SD2L.t199 0.551
R905 SD2L.n97 SD2L.t202 0.551
R906 SD2L.n98 SD2L.t133 0.551
R907 SD2L.n98 SD2L.t207 0.551
R908 SD2L.n99 SD2L.t120 0.551
R909 SD2L.n99 SD2L.t127 0.551
R910 SD2L.n100 SD2L.t230 0.551
R911 SD2L.n100 SD2L.t201 0.551
R912 SD2L.n101 SD2L.t221 0.551
R913 SD2L.n101 SD2L.t196 0.551
R914 SD2L.n102 SD2L.t124 0.551
R915 SD2L.n102 SD2L.t192 0.551
R916 SD2L.n103 SD2L.t36 0.551
R917 SD2L.n103 SD2L.t11 0.551
R918 SD2L.n104 SD2L.t25 0.551
R919 SD2L.n104 SD2L.t32 0.551
R920 SD2L.n105 SD2L.t15 0.551
R921 SD2L.n105 SD2L.t57 0.551
R922 SD2L.n106 SD2L.t113 0.551
R923 SD2L.n106 SD2L.t95 0.551
R924 SD2L.n107 SD2L.t16 0.551
R925 SD2L.n107 SD2L.t64 0.551
R926 SD2L.n108 SD2L.t77 0.551
R927 SD2L.n108 SD2L.t7 0.551
R928 SD2L.n109 SD2L.t72 0.551
R929 SD2L.n109 SD2L.t99 0.551
R930 SD2L.n110 SD2L.t71 0.551
R931 SD2L.n110 SD2L.t54 0.551
R932 SD2L.n111 SD2L.t60 0.551
R933 SD2L.n111 SD2L.t118 0.551
R934 SD2L.n112 SD2L.t67 0.551
R935 SD2L.n112 SD2L.t9 0.551
R936 SD2L.n113 SD2L.t43 0.551
R937 SD2L.n113 SD2L.t78 0.551
R938 SD2L.n114 SD2L.t34 0.551
R939 SD2L.n114 SD2L.t61 0.551
R940 SD2L.n115 SD2L.t66 0.551
R941 SD2L.n115 SD2L.t92 0.551
R942 SD2L.n116 SD2L.t111 0.551
R943 SD2L.n116 SD2L.t117 0.551
R944 SD2L.n122 SD2L.t212 0.551
R945 SD2L.n122 SD2L.t152 0.551
R946 SD2L.n123 SD2L.t217 0.551
R947 SD2L.n123 SD2L.t228 0.551
R948 SD2L.n124 SD2L.t140 0.551
R949 SD2L.n124 SD2L.t145 0.551
R950 SD2L.n125 SD2L.t224 0.551
R951 SD2L.n125 SD2L.t203 0.551
R952 SD2L.n126 SD2L.t218 0.551
R953 SD2L.n126 SD2L.t142 0.551
R954 SD2L.n121 SD2L.t163 0.551
R955 SD2L.n121 SD2L.t169 0.551
R956 SD2L.n120 SD2L.t129 0.551
R957 SD2L.n120 SD2L.t225 0.551
R958 SD2L.n119 SD2L.t141 0.551
R959 SD2L.n119 SD2L.t211 0.551
R960 SD2L.n118 SD2L.t239 0.551
R961 SD2L.n118 SD2L.t189 0.551
R962 SD2L.n117 SD2L.t190 0.551
R963 SD2L.n117 SD2L.t172 0.551
R964 SD2L.n127 SD2L.t227 0.551
R965 SD2L.n127 SD2L.t198 0.551
R966 SD2L.n128 SD2L.t213 0.551
R967 SD2L.n128 SD2L.t176 0.551
R968 SD2L.n129 SD2L.t197 0.551
R969 SD2L.n129 SD2L.t216 0.551
R970 SD2L.n130 SD2L.t184 0.551
R971 SD2L.n130 SD2L.t238 0.551
R972 SD2L.n145 SD2L.t59 0.551
R973 SD2L.n145 SD2L.t0 0.551
R974 SD2L.n146 SD2L.n3 0.455
R975 SD2L.n148 SD2L.n10 0.416
R976 SD2L SD2L.n21 0.281
R977 SD2L.n147 SD2L.n19 0.281
R978 SD2L.n149 SD2L.n27 0.155
R979 SD2L.n146 SD2L.n23 0.155
R980 SD2L.n147 SD2L.n146 0.13
R981 SD2L SD2L.n149 0.13
R982 SD2L.n147 SD2L.n25 0.103
R983 SD2L SD2L.n29 0.103
R984 SD2L.n148 SD2L.n147 0.091
R985 SD2L.n149 SD2L.n148 0.039
R986 SD2L.n10 SD2L.n11 0.038
R987 SD2L.n3 SD2L.n4 0.038
R988 SD2L.n28 SD2L.n17 0.028
R989 SD2L.n20 SD2L.n15 0.028
R990 SD2L.n26 SD2L.n13 0.028
R991 SD2L.n10 SD2L.n9 0.028
R992 SD2L.n24 SD2L.n8 0.028
R993 SD2L.n18 SD2L.n6 0.028
R994 SD2L.n3 SD2L.n2 0.028
R995 SD2L.n22 SD2L.n1 0.028
R996 SD2L.n21 SD2L.n20 0.025
R997 SD2L.n19 SD2L.n18 0.025
R998 SD2L.n29 SD2L.n28 0.022
R999 SD2L.n27 SD2L.n26 0.022
R1000 SD2L.n25 SD2L.n24 0.022
R1001 SD2L.n23 SD2L.n22 0.022
R1002 SD2L.n1 SD2L.n0 0.021
R1003 SD2L.n6 SD2L.n5 0.021
R1004 SD2L.n8 SD2L.n7 0.021
R1005 SD2L.n13 SD2L.n12 0.021
R1006 SD2L.n15 SD2L.n14 0.021
R1007 SD2L.n17 SD2L.n16 0.021
R1008 SD1L.n93 SD1L.t25 1.972
R1009 SD1L.n11 SD1L.t116 1.972
R1010 SD1L.n105 SD1L.t33 1.963
R1011 SD1L.n25 SD1L.t80 1.962
R1012 SD1L.n37 SD1L.n36 1.435
R1013 SD1L.n64 SD1L.n63 1.435
R1014 SD1L.n46 SD1L.n26 1.428
R1015 SD1L.n45 SD1L.n27 1.428
R1016 SD1L.n44 SD1L.n28 1.428
R1017 SD1L.n43 SD1L.n29 1.428
R1018 SD1L.n42 SD1L.n30 1.428
R1019 SD1L.n41 SD1L.n31 1.428
R1020 SD1L.n40 SD1L.n32 1.428
R1021 SD1L.n39 SD1L.n33 1.428
R1022 SD1L.n38 SD1L.n34 1.428
R1023 SD1L.n37 SD1L.n35 1.428
R1024 SD1L.n73 SD1L.n53 1.428
R1025 SD1L.n72 SD1L.n54 1.428
R1026 SD1L.n71 SD1L.n55 1.428
R1027 SD1L.n70 SD1L.n56 1.428
R1028 SD1L.n69 SD1L.n57 1.428
R1029 SD1L.n68 SD1L.n58 1.428
R1030 SD1L.n67 SD1L.n59 1.428
R1031 SD1L.n66 SD1L.n60 1.428
R1032 SD1L.n65 SD1L.n61 1.428
R1033 SD1L.n64 SD1L.n62 1.428
R1034 SD1L.n104 SD1L.n83 1.414
R1035 SD1L.n103 SD1L.n84 1.414
R1036 SD1L.n102 SD1L.n85 1.414
R1037 SD1L.n101 SD1L.n86 1.414
R1038 SD1L.n100 SD1L.n87 1.414
R1039 SD1L.n99 SD1L.n88 1.414
R1040 SD1L.n96 SD1L.n89 1.414
R1041 SD1L.n95 SD1L.n90 1.414
R1042 SD1L.n94 SD1L.n91 1.414
R1043 SD1L.n93 SD1L.n92 1.414
R1044 SD1L.n21 SD1L.n0 1.414
R1045 SD1L.n20 SD1L.n1 1.414
R1046 SD1L.n19 SD1L.n2 1.414
R1047 SD1L.n18 SD1L.n3 1.414
R1048 SD1L.n17 SD1L.n4 1.414
R1049 SD1L.n16 SD1L.n5 1.414
R1050 SD1L.n15 SD1L.n6 1.414
R1051 SD1L.n14 SD1L.n7 1.414
R1052 SD1L.n13 SD1L.n8 1.414
R1053 SD1L.n12 SD1L.n9 1.414
R1054 SD1L.n11 SD1L.n10 1.414
R1055 SD1L.n98 SD1L.n97 1.413
R1056 SD1L.n105 SD1L.n80 1.412
R1057 SD1L.n105 SD1L.n81 1.412
R1058 SD1L.n105 SD1L.n82 1.412
R1059 SD1L.n25 SD1L.n24 1.409
R1060 SD1L.n25 SD1L.n23 1.409
R1061 SD1L.n25 SD1L.n22 1.409
R1062 SD1L.n48 SD1L.n47 1.281
R1063 SD1L.n75 SD1L.n74 1.281
R1064 SD1L.n52 SD1L.n49 1.28
R1065 SD1L.n52 SD1L.n50 1.28
R1066 SD1L.n52 SD1L.n51 1.28
R1067 SD1L.n79 SD1L.n76 1.28
R1068 SD1L.n79 SD1L.n77 1.28
R1069 SD1L.n79 SD1L.n78 1.28
R1070 SD1L.n83 SD1L.t11 0.551
R1071 SD1L.n83 SD1L.t20 0.551
R1072 SD1L.n84 SD1L.t38 0.551
R1073 SD1L.n84 SD1L.t86 0.551
R1074 SD1L.n85 SD1L.t100 0.551
R1075 SD1L.n85 SD1L.t31 0.551
R1076 SD1L.n86 SD1L.t51 0.551
R1077 SD1L.n86 SD1L.t95 0.551
R1078 SD1L.n87 SD1L.t84 0.551
R1079 SD1L.n87 SD1L.t10 0.551
R1080 SD1L.n88 SD1L.t49 0.551
R1081 SD1L.n88 SD1L.t53 0.551
R1082 SD1L.n89 SD1L.t111 0.551
R1083 SD1L.n89 SD1L.t41 0.551
R1084 SD1L.n90 SD1L.t74 0.551
R1085 SD1L.n90 SD1L.t117 0.551
R1086 SD1L.n91 SD1L.t107 0.551
R1087 SD1L.n91 SD1L.t39 0.551
R1088 SD1L.n92 SD1L.t58 0.551
R1089 SD1L.n92 SD1L.t102 0.551
R1090 SD1L.n82 SD1L.t67 0.551
R1091 SD1L.n82 SD1L.t75 0.551
R1092 SD1L.n81 SD1L.t106 0.551
R1093 SD1L.n81 SD1L.t96 0.551
R1094 SD1L.n80 SD1L.t81 0.551
R1095 SD1L.n80 SD1L.t40 0.551
R1096 SD1L.n26 SD1L.t89 0.551
R1097 SD1L.n26 SD1L.t62 0.551
R1098 SD1L.n27 SD1L.t21 0.551
R1099 SD1L.n27 SD1L.t83 0.551
R1100 SD1L.n28 SD1L.t27 0.551
R1101 SD1L.n28 SD1L.t88 0.551
R1102 SD1L.n29 SD1L.t77 0.551
R1103 SD1L.n29 SD1L.t52 0.551
R1104 SD1L.n30 SD1L.t9 0.551
R1105 SD1L.n30 SD1L.t104 0.551
R1106 SD1L.n31 SD1L.t12 0.551
R1107 SD1L.n31 SD1L.t69 0.551
R1108 SD1L.n32 SD1L.t68 0.551
R1109 SD1L.n32 SD1L.t43 0.551
R1110 SD1L.n33 SD1L.t36 0.551
R1111 SD1L.n33 SD1L.t94 0.551
R1112 SD1L.n34 SD1L.t2 0.551
R1113 SD1L.n34 SD1L.t60 0.551
R1114 SD1L.n35 SD1L.t87 0.551
R1115 SD1L.n35 SD1L.t34 0.551
R1116 SD1L.n36 SD1L.t22 0.551
R1117 SD1L.n36 SD1L.t114 0.551
R1118 SD1L.n47 SD1L.t3 0.551
R1119 SD1L.n47 SD1L.t97 0.551
R1120 SD1L.n49 SD1L.t1 0.551
R1121 SD1L.n49 SD1L.t4 0.551
R1122 SD1L.n50 SD1L.t72 0.551
R1123 SD1L.n50 SD1L.t45 0.551
R1124 SD1L.n51 SD1L.t13 0.551
R1125 SD1L.n51 SD1L.t78 0.551
R1126 SD1L.n53 SD1L.t23 0.551
R1127 SD1L.n53 SD1L.t91 0.551
R1128 SD1L.n54 SD1L.t90 0.551
R1129 SD1L.n54 SD1L.t29 0.551
R1130 SD1L.n55 SD1L.t5 0.551
R1131 SD1L.n55 SD1L.t63 0.551
R1132 SD1L.n56 SD1L.t37 0.551
R1133 SD1L.n56 SD1L.t98 0.551
R1134 SD1L.n57 SD1L.t99 0.551
R1135 SD1L.n57 SD1L.t6 0.551
R1136 SD1L.n58 SD1L.t15 0.551
R1137 SD1L.n58 SD1L.t46 0.551
R1138 SD1L.n59 SD1L.t47 0.551
R1139 SD1L.n59 SD1L.t109 0.551
R1140 SD1L.n60 SD1L.t79 0.551
R1141 SD1L.n60 SD1L.t18 0.551
R1142 SD1L.n61 SD1L.t30 0.551
R1143 SD1L.n61 SD1L.t54 0.551
R1144 SD1L.n62 SD1L.t64 0.551
R1145 SD1L.n62 SD1L.t119 0.551
R1146 SD1L.n63 SD1L.t112 0.551
R1147 SD1L.n63 SD1L.t19 0.551
R1148 SD1L.n74 SD1L.t28 0.551
R1149 SD1L.n74 SD1L.t55 0.551
R1150 SD1L.n76 SD1L.t108 0.551
R1151 SD1L.n76 SD1L.t105 0.551
R1152 SD1L.n77 SD1L.t44 0.551
R1153 SD1L.n77 SD1L.t70 0.551
R1154 SD1L.n78 SD1L.t16 0.551
R1155 SD1L.n78 SD1L.t76 0.551
R1156 SD1L.n24 SD1L.t0 0.551
R1157 SD1L.n24 SD1L.t85 0.551
R1158 SD1L.n23 SD1L.t56 0.551
R1159 SD1L.n23 SD1L.t50 0.551
R1160 SD1L.n22 SD1L.t14 0.551
R1161 SD1L.n22 SD1L.t8 0.551
R1162 SD1L.n0 SD1L.t57 0.551
R1163 SD1L.n0 SD1L.t61 0.551
R1164 SD1L.n1 SD1L.t59 0.551
R1165 SD1L.n1 SD1L.t101 0.551
R1166 SD1L.n2 SD1L.t110 0.551
R1167 SD1L.n2 SD1L.t65 0.551
R1168 SD1L.n3 SD1L.t32 0.551
R1169 SD1L.n3 SD1L.t115 0.551
R1170 SD1L.n4 SD1L.t113 0.551
R1171 SD1L.n4 SD1L.t66 0.551
R1172 SD1L.n5 SD1L.t48 0.551
R1173 SD1L.n5 SD1L.t42 0.551
R1174 SD1L.n6 SD1L.t7 0.551
R1175 SD1L.n6 SD1L.t93 0.551
R1176 SD1L.n7 SD1L.t17 0.551
R1177 SD1L.n7 SD1L.t92 0.551
R1178 SD1L.n8 SD1L.t71 0.551
R1179 SD1L.n8 SD1L.t24 0.551
R1180 SD1L.n9 SD1L.t35 0.551
R1181 SD1L.n9 SD1L.t103 0.551
R1182 SD1L.n10 SD1L.t73 0.551
R1183 SD1L.n10 SD1L.t26 0.551
R1184 SD1L.n97 SD1L.t82 0.551
R1185 SD1L.n97 SD1L.t118 0.551
R1186 SD1L.n106 SD1L.n79 0.254
R1187 SD1L.n108 SD1L.n25 0.249
R1188 SD1L.n106 SD1L.n105 0.249
R1189 SD1L.n107 SD1L.n106 0.13
R1190 SD1L.n107 SD1L.n52 0.124
R1191 SD1L.n108 SD1L.n107 0.114
R1192 SD1L SD1L.n108 0.056
R1193 SD1L.n48 SD1L.n46 0.007
R1194 SD1L.n75 SD1L.n73 0.007
R1195 SD1L.n38 SD1L.n37 0.007
R1196 SD1L.n39 SD1L.n38 0.007
R1197 SD1L.n40 SD1L.n39 0.007
R1198 SD1L.n41 SD1L.n40 0.007
R1199 SD1L.n42 SD1L.n41 0.007
R1200 SD1L.n43 SD1L.n42 0.007
R1201 SD1L.n44 SD1L.n43 0.007
R1202 SD1L.n45 SD1L.n44 0.007
R1203 SD1L.n46 SD1L.n45 0.007
R1204 SD1L.n65 SD1L.n64 0.007
R1205 SD1L.n66 SD1L.n65 0.007
R1206 SD1L.n67 SD1L.n66 0.007
R1207 SD1L.n68 SD1L.n67 0.007
R1208 SD1L.n69 SD1L.n68 0.007
R1209 SD1L.n70 SD1L.n69 0.007
R1210 SD1L.n71 SD1L.n70 0.007
R1211 SD1L.n72 SD1L.n71 0.007
R1212 SD1L.n73 SD1L.n72 0.007
R1213 SD1L.n12 SD1L.n11 0.007
R1214 SD1L.n13 SD1L.n12 0.007
R1215 SD1L.n14 SD1L.n13 0.007
R1216 SD1L.n15 SD1L.n14 0.007
R1217 SD1L.n16 SD1L.n15 0.007
R1218 SD1L.n17 SD1L.n16 0.007
R1219 SD1L.n18 SD1L.n17 0.007
R1220 SD1L.n19 SD1L.n18 0.007
R1221 SD1L.n20 SD1L.n19 0.007
R1222 SD1L.n21 SD1L.n20 0.007
R1223 SD1L.n94 SD1L.n93 0.007
R1224 SD1L.n95 SD1L.n94 0.007
R1225 SD1L.n96 SD1L.n95 0.007
R1226 SD1L.n98 SD1L.n96 0.007
R1227 SD1L.n99 SD1L.n98 0.007
R1228 SD1L.n100 SD1L.n99 0.007
R1229 SD1L.n101 SD1L.n100 0.007
R1230 SD1L.n102 SD1L.n101 0.007
R1231 SD1L.n103 SD1L.n102 0.007
R1232 SD1L.n104 SD1L.n103 0.007
R1233 SD1L.n25 SD1L.n21 0.004
R1234 SD1L.n105 SD1L.n104 0.004
R1235 SD1L.n52 SD1L.n48 0.001
R1236 SD1L.n79 SD1L.n75 0.001
R1237 SD2R.n115 SD2R.t146 1.972
R1238 SD2R.n167 SD2R.t50 1.972
R1239 SD2R.n11 SD2R.t237 1.972
R1240 SD2R.n63 SD2R.t57 1.972
R1241 SD2R.n129 SD2R.t140 1.963
R1242 SD2R.n181 SD2R.t36 1.963
R1243 SD2R.n25 SD2R.t148 1.963
R1244 SD2R.n78 SD2R.t58 1.96
R1245 SD2R.n193 SD2R.n192 1.435
R1246 SD2R.n206 SD2R.n205 1.435
R1247 SD2R.n95 SD2R.n94 1.435
R1248 SD2R.n85 SD2R.n84 1.435
R1249 SD2R.n141 SD2R.n140 1.435
R1250 SD2R.n37 SD2R.n36 1.435
R1251 SD2R.n196 SD2R.n188 1.428
R1252 SD2R.n195 SD2R.n189 1.428
R1253 SD2R.n194 SD2R.n190 1.428
R1254 SD2R.n193 SD2R.n191 1.428
R1255 SD2R.n206 SD2R.n204 1.428
R1256 SD2R.n207 SD2R.n203 1.428
R1257 SD2R.n208 SD2R.n202 1.428
R1258 SD2R.n209 SD2R.n201 1.428
R1259 SD2R.n210 SD2R.n200 1.428
R1260 SD2R.n98 SD2R.n90 1.428
R1261 SD2R.n97 SD2R.n91 1.428
R1262 SD2R.n96 SD2R.n92 1.428
R1263 SD2R.n95 SD2R.n93 1.428
R1264 SD2R.n85 SD2R.n83 1.428
R1265 SD2R.n86 SD2R.n82 1.428
R1266 SD2R.n87 SD2R.n81 1.428
R1267 SD2R.n88 SD2R.n80 1.428
R1268 SD2R.n89 SD2R.n79 1.428
R1269 SD2R.n150 SD2R.n130 1.428
R1270 SD2R.n149 SD2R.n131 1.428
R1271 SD2R.n148 SD2R.n132 1.428
R1272 SD2R.n147 SD2R.n133 1.428
R1273 SD2R.n146 SD2R.n134 1.428
R1274 SD2R.n145 SD2R.n135 1.428
R1275 SD2R.n144 SD2R.n136 1.428
R1276 SD2R.n143 SD2R.n137 1.428
R1277 SD2R.n142 SD2R.n138 1.428
R1278 SD2R.n141 SD2R.n139 1.428
R1279 SD2R.n46 SD2R.n26 1.428
R1280 SD2R.n45 SD2R.n27 1.428
R1281 SD2R.n44 SD2R.n28 1.428
R1282 SD2R.n43 SD2R.n29 1.428
R1283 SD2R.n42 SD2R.n30 1.428
R1284 SD2R.n41 SD2R.n31 1.428
R1285 SD2R.n40 SD2R.n32 1.428
R1286 SD2R.n39 SD2R.n33 1.428
R1287 SD2R.n38 SD2R.n34 1.428
R1288 SD2R.n37 SD2R.n35 1.428
R1289 SD2R.n63 SD2R.n62 1.414
R1290 SD2R.n64 SD2R.n61 1.414
R1291 SD2R.n65 SD2R.n60 1.414
R1292 SD2R.n66 SD2R.n59 1.414
R1293 SD2R.n67 SD2R.n58 1.414
R1294 SD2R.n68 SD2R.n57 1.414
R1295 SD2R.n69 SD2R.n56 1.414
R1296 SD2R.n70 SD2R.n55 1.414
R1297 SD2R.n71 SD2R.n54 1.414
R1298 SD2R.n72 SD2R.n53 1.414
R1299 SD2R.n73 SD2R.n52 1.414
R1300 SD2R.n125 SD2R.n104 1.414
R1301 SD2R.n124 SD2R.n105 1.414
R1302 SD2R.n123 SD2R.n106 1.414
R1303 SD2R.n122 SD2R.n107 1.414
R1304 SD2R.n121 SD2R.n108 1.414
R1305 SD2R.n120 SD2R.n109 1.414
R1306 SD2R.n119 SD2R.n110 1.414
R1307 SD2R.n118 SD2R.n111 1.414
R1308 SD2R.n117 SD2R.n112 1.414
R1309 SD2R.n116 SD2R.n113 1.414
R1310 SD2R.n115 SD2R.n114 1.414
R1311 SD2R.n177 SD2R.n156 1.414
R1312 SD2R.n176 SD2R.n157 1.414
R1313 SD2R.n175 SD2R.n158 1.414
R1314 SD2R.n174 SD2R.n159 1.414
R1315 SD2R.n173 SD2R.n160 1.414
R1316 SD2R.n172 SD2R.n161 1.414
R1317 SD2R.n171 SD2R.n162 1.414
R1318 SD2R.n170 SD2R.n163 1.414
R1319 SD2R.n169 SD2R.n164 1.414
R1320 SD2R.n168 SD2R.n165 1.414
R1321 SD2R.n167 SD2R.n166 1.414
R1322 SD2R.n21 SD2R.n0 1.414
R1323 SD2R.n20 SD2R.n1 1.414
R1324 SD2R.n19 SD2R.n2 1.414
R1325 SD2R.n18 SD2R.n3 1.414
R1326 SD2R.n17 SD2R.n4 1.414
R1327 SD2R.n16 SD2R.n5 1.414
R1328 SD2R.n15 SD2R.n6 1.414
R1329 SD2R.n14 SD2R.n7 1.414
R1330 SD2R.n13 SD2R.n8 1.414
R1331 SD2R.n12 SD2R.n9 1.414
R1332 SD2R.n11 SD2R.n10 1.414
R1333 SD2R.n129 SD2R.n128 1.412
R1334 SD2R.n129 SD2R.n127 1.412
R1335 SD2R.n129 SD2R.n126 1.412
R1336 SD2R.n181 SD2R.n180 1.412
R1337 SD2R.n181 SD2R.n179 1.412
R1338 SD2R.n181 SD2R.n178 1.412
R1339 SD2R.n25 SD2R.n24 1.412
R1340 SD2R.n25 SD2R.n23 1.412
R1341 SD2R.n25 SD2R.n22 1.412
R1342 SD2R.n75 SD2R.n74 1.41
R1343 SD2R.n78 SD2R.n76 1.409
R1344 SD2R.n78 SD2R.n77 1.409
R1345 SD2R.n152 SD2R.n151 1.282
R1346 SD2R.n48 SD2R.n47 1.282
R1347 SD2R.n103 SD2R.n99 1.28
R1348 SD2R.n103 SD2R.n100 1.28
R1349 SD2R.n103 SD2R.n101 1.28
R1350 SD2R.n103 SD2R.n102 1.28
R1351 SD2R.n182 SD2R.n153 1.28
R1352 SD2R.n182 SD2R.n155 1.28
R1353 SD2R.n182 SD2R.n154 1.28
R1354 SD2R.n186 SD2R.n49 1.28
R1355 SD2R.n186 SD2R.n51 1.28
R1356 SD2R.n186 SD2R.n50 1.28
R1357 SD2R.n212 SD2R.n197 1.28
R1358 SD2R.n212 SD2R.n198 1.28
R1359 SD2R.n212 SD2R.n199 1.28
R1360 SD2R.n212 SD2R.n211 1.278
R1361 SD2R.n188 SD2R.t51 0.551
R1362 SD2R.n188 SD2R.t91 0.551
R1363 SD2R.n189 SD2R.t102 0.551
R1364 SD2R.n189 SD2R.t100 0.551
R1365 SD2R.n190 SD2R.t65 0.551
R1366 SD2R.n190 SD2R.t26 0.551
R1367 SD2R.n191 SD2R.t105 0.551
R1368 SD2R.n191 SD2R.t112 0.551
R1369 SD2R.n192 SD2R.t77 0.551
R1370 SD2R.n192 SD2R.t28 0.551
R1371 SD2R.n205 SD2R.t47 0.551
R1372 SD2R.n205 SD2R.t39 0.551
R1373 SD2R.n204 SD2R.t5 0.551
R1374 SD2R.n204 SD2R.t83 0.551
R1375 SD2R.n203 SD2R.t92 0.551
R1376 SD2R.n203 SD2R.t11 0.551
R1377 SD2R.n202 SD2R.t20 0.551
R1378 SD2R.n202 SD2R.t99 0.551
R1379 SD2R.n201 SD2R.t60 0.551
R1380 SD2R.n201 SD2R.t13 0.551
R1381 SD2R.n200 SD2R.t21 0.551
R1382 SD2R.n200 SD2R.t15 0.551
R1383 SD2R.n197 SD2R.t52 0.551
R1384 SD2R.n197 SD2R.t3 0.551
R1385 SD2R.n198 SD2R.t22 0.551
R1386 SD2R.n198 SD2R.t108 0.551
R1387 SD2R.n199 SD2R.t76 0.551
R1388 SD2R.n199 SD2R.t71 0.551
R1389 SD2R.n62 SD2R.t111 0.551
R1390 SD2R.n62 SD2R.t63 0.551
R1391 SD2R.n61 SD2R.t43 0.551
R1392 SD2R.n61 SD2R.t35 0.551
R1393 SD2R.n60 SD2R.t113 0.551
R1394 SD2R.n60 SD2R.t0 0.551
R1395 SD2R.n59 SD2R.t45 0.551
R1396 SD2R.n59 SD2R.t38 0.551
R1397 SD2R.n58 SD2R.t49 0.551
R1398 SD2R.n58 SD2R.t95 0.551
R1399 SD2R.n57 SD2R.t90 0.551
R1400 SD2R.n57 SD2R.t53 0.551
R1401 SD2R.n56 SD2R.t18 0.551
R1402 SD2R.n56 SD2R.t97 0.551
R1403 SD2R.n55 SD2R.t103 0.551
R1404 SD2R.n55 SD2R.t56 0.551
R1405 SD2R.n54 SD2R.t33 0.551
R1406 SD2R.n54 SD2R.t27 0.551
R1407 SD2R.n53 SD2R.t106 0.551
R1408 SD2R.n53 SD2R.t69 0.551
R1409 SD2R.n52 SD2R.t79 0.551
R1410 SD2R.n52 SD2R.t29 0.551
R1411 SD2R.n74 SD2R.t8 0.551
R1412 SD2R.n74 SD2R.t85 0.551
R1413 SD2R.n76 SD2R.t81 0.551
R1414 SD2R.n76 SD2R.t31 0.551
R1415 SD2R.n77 SD2R.t9 0.551
R1416 SD2R.n77 SD2R.t86 0.551
R1417 SD2R.n90 SD2R.t118 0.551
R1418 SD2R.n90 SD2R.t44 0.551
R1419 SD2R.n91 SD2R.t80 0.551
R1420 SD2R.n91 SD2R.t72 0.551
R1421 SD2R.n92 SD2R.t116 0.551
R1422 SD2R.n92 SD2R.t30 0.551
R1423 SD2R.n93 SD2R.t62 0.551
R1424 SD2R.n93 SD2R.t70 0.551
R1425 SD2R.n94 SD2R.t104 0.551
R1426 SD2R.n94 SD2R.t14 0.551
R1427 SD2R.n84 SD2R.t117 0.551
R1428 SD2R.n84 SD2R.t109 0.551
R1429 SD2R.n83 SD2R.t55 0.551
R1430 SD2R.n83 SD2R.t40 0.551
R1431 SD2R.n82 SD2R.t32 0.551
R1432 SD2R.n82 SD2R.t66 0.551
R1433 SD2R.n81 SD2R.t101 0.551
R1434 SD2R.n81 SD2R.t23 0.551
R1435 SD2R.n80 SD2R.t48 0.551
R1436 SD2R.n80 SD2R.t98 0.551
R1437 SD2R.n79 SD2R.t107 0.551
R1438 SD2R.n79 SD2R.t114 0.551
R1439 SD2R.n99 SD2R.t82 0.551
R1440 SD2R.n99 SD2R.t4 0.551
R1441 SD2R.n100 SD2R.t10 0.551
R1442 SD2R.n100 SD2R.t46 0.551
R1443 SD2R.n101 SD2R.t96 0.551
R1444 SD2R.n101 SD2R.t6 0.551
R1445 SD2R.n102 SD2R.t54 0.551
R1446 SD2R.n102 SD2R.t59 0.551
R1447 SD2R.n104 SD2R.t143 0.551
R1448 SD2R.n104 SD2R.t152 0.551
R1449 SD2R.n105 SD2R.t187 0.551
R1450 SD2R.n105 SD2R.t180 0.551
R1451 SD2R.n106 SD2R.t189 0.551
R1452 SD2R.n106 SD2R.t201 0.551
R1453 SD2R.n107 SD2R.t184 0.551
R1454 SD2R.n107 SD2R.t218 0.551
R1455 SD2R.n108 SD2R.t215 0.551
R1456 SD2R.n108 SD2R.t176 0.551
R1457 SD2R.n109 SD2R.t126 0.551
R1458 SD2R.n109 SD2R.t128 0.551
R1459 SD2R.n110 SD2R.t160 0.551
R1460 SD2R.n110 SD2R.t163 0.551
R1461 SD2R.n111 SD2R.t194 0.551
R1462 SD2R.n111 SD2R.t174 0.551
R1463 SD2R.n112 SD2R.t191 0.551
R1464 SD2R.n112 SD2R.t188 0.551
R1465 SD2R.n113 SD2R.t229 0.551
R1466 SD2R.n113 SD2R.t144 0.551
R1467 SD2R.n114 SD2R.t205 0.551
R1468 SD2R.n114 SD2R.t177 0.551
R1469 SD2R.n126 SD2R.t147 0.551
R1470 SD2R.n126 SD2R.t159 0.551
R1471 SD2R.n127 SD2R.t135 0.551
R1472 SD2R.n127 SD2R.t219 0.551
R1473 SD2R.n128 SD2R.t150 0.551
R1474 SD2R.n128 SD2R.t214 0.551
R1475 SD2R.n130 SD2R.t186 0.551
R1476 SD2R.n130 SD2R.t210 0.551
R1477 SD2R.n131 SD2R.t134 0.551
R1478 SD2R.n131 SD2R.t158 0.551
R1479 SD2R.n132 SD2R.t141 0.551
R1480 SD2R.n132 SD2R.t171 0.551
R1481 SD2R.n133 SD2R.t203 0.551
R1482 SD2R.n133 SD2R.t129 0.551
R1483 SD2R.n134 SD2R.t197 0.551
R1484 SD2R.n134 SD2R.t234 0.551
R1485 SD2R.n135 SD2R.t193 0.551
R1486 SD2R.n135 SD2R.t231 0.551
R1487 SD2R.n136 SD2R.t202 0.551
R1488 SD2R.n136 SD2R.t156 0.551
R1489 SD2R.n137 SD2R.t222 0.551
R1490 SD2R.n137 SD2R.t137 0.551
R1491 SD2R.n138 SD2R.t216 0.551
R1492 SD2R.n138 SD2R.t179 0.551
R1493 SD2R.n139 SD2R.t175 0.551
R1494 SD2R.n139 SD2R.t157 0.551
R1495 SD2R.n140 SD2R.t220 0.551
R1496 SD2R.n140 SD2R.t226 0.551
R1497 SD2R.n151 SD2R.t120 0.551
R1498 SD2R.n151 SD2R.t154 0.551
R1499 SD2R.n153 SD2R.t195 0.551
R1500 SD2R.n153 SD2R.t221 0.551
R1501 SD2R.n155 SD2R.t178 0.551
R1502 SD2R.n155 SD2R.t131 0.551
R1503 SD2R.n154 SD2R.t192 0.551
R1504 SD2R.n154 SD2R.t173 0.551
R1505 SD2R.n156 SD2R.t42 0.551
R1506 SD2R.n156 SD2R.t93 0.551
R1507 SD2R.n157 SD2R.t2 0.551
R1508 SD2R.n157 SD2R.t37 0.551
R1509 SD2R.n158 SD2R.t87 0.551
R1510 SD2R.n158 SD2R.t94 0.551
R1511 SD2R.n159 SD2R.t16 0.551
R1512 SD2R.n159 SD2R.t64 0.551
R1513 SD2R.n160 SD2R.t89 0.551
R1514 SD2R.n160 SD2R.t12 0.551
R1515 SD2R.n161 SD2R.t17 0.551
R1516 SD2R.n161 SD2R.t67 0.551
R1517 SD2R.n162 SD2R.t73 0.551
R1518 SD2R.n162 SD2R.t25 0.551
R1519 SD2R.n163 SD2R.t61 0.551
R1520 SD2R.n163 SD2R.t68 0.551
R1521 SD2R.n164 SD2R.t115 0.551
R1522 SD2R.n164 SD2R.t1 0.551
R1523 SD2R.n165 SD2R.t78 0.551
R1524 SD2R.n165 SD2R.t84 0.551
R1525 SD2R.n166 SD2R.t7 0.551
R1526 SD2R.n166 SD2R.t41 0.551
R1527 SD2R.n178 SD2R.t88 0.551
R1528 SD2R.n178 SD2R.t19 0.551
R1529 SD2R.n179 SD2R.t24 0.551
R1530 SD2R.n179 SD2R.t75 0.551
R1531 SD2R.n180 SD2R.t110 0.551
R1532 SD2R.n180 SD2R.t34 0.551
R1533 SD2R.n0 SD2R.t164 0.551
R1534 SD2R.n0 SD2R.t167 0.551
R1535 SD2R.n1 SD2R.t125 0.551
R1536 SD2R.n1 SD2R.t227 0.551
R1537 SD2R.n2 SD2R.t213 0.551
R1538 SD2R.n2 SD2R.t238 0.551
R1539 SD2R.n3 SD2R.t142 0.551
R1540 SD2R.n3 SD2R.t236 0.551
R1541 SD2R.n4 SD2R.t185 0.551
R1542 SD2R.n4 SD2R.t230 0.551
R1543 SD2R.n5 SD2R.t209 0.551
R1544 SD2R.n5 SD2R.t133 0.551
R1545 SD2R.n6 SD2R.t155 0.551
R1546 SD2R.n6 SD2R.t130 0.551
R1547 SD2R.n7 SD2R.t235 0.551
R1548 SD2R.n7 SD2R.t132 0.551
R1549 SD2R.n8 SD2R.t225 0.551
R1550 SD2R.n8 SD2R.t151 0.551
R1551 SD2R.n9 SD2R.t224 0.551
R1552 SD2R.n9 SD2R.t232 0.551
R1553 SD2R.n10 SD2R.t139 0.551
R1554 SD2R.n10 SD2R.t145 0.551
R1555 SD2R.n22 SD2R.t196 0.551
R1556 SD2R.n22 SD2R.t121 0.551
R1557 SD2R.n23 SD2R.t127 0.551
R1558 SD2R.n23 SD2R.t138 0.551
R1559 SD2R.n24 SD2R.t207 0.551
R1560 SD2R.n24 SD2R.t198 0.551
R1561 SD2R.n26 SD2R.t169 0.551
R1562 SD2R.n26 SD2R.t172 0.551
R1563 SD2R.n27 SD2R.t123 0.551
R1564 SD2R.n27 SD2R.t206 0.551
R1565 SD2R.n28 SD2R.t168 0.551
R1566 SD2R.n28 SD2R.t233 0.551
R1567 SD2R.n29 SD2R.t122 0.551
R1568 SD2R.n29 SD2R.t181 0.551
R1569 SD2R.n30 SD2R.t162 0.551
R1570 SD2R.n30 SD2R.t161 0.551
R1571 SD2R.n31 SD2R.t208 0.551
R1572 SD2R.n31 SD2R.t228 0.551
R1573 SD2R.n32 SD2R.t124 0.551
R1574 SD2R.n32 SD2R.t182 0.551
R1575 SD2R.n33 SD2R.t217 0.551
R1576 SD2R.n33 SD2R.t165 0.551
R1577 SD2R.n34 SD2R.t204 0.551
R1578 SD2R.n34 SD2R.t183 0.551
R1579 SD2R.n35 SD2R.t149 0.551
R1580 SD2R.n35 SD2R.t200 0.551
R1581 SD2R.n36 SD2R.t190 0.551
R1582 SD2R.n36 SD2R.t239 0.551
R1583 SD2R.n47 SD2R.t223 0.551
R1584 SD2R.n47 SD2R.t170 0.551
R1585 SD2R.n49 SD2R.t166 0.551
R1586 SD2R.n49 SD2R.t211 0.551
R1587 SD2R.n51 SD2R.t212 0.551
R1588 SD2R.n51 SD2R.t153 0.551
R1589 SD2R.n50 SD2R.t199 0.551
R1590 SD2R.n50 SD2R.t136 0.551
R1591 SD2R.n211 SD2R.t119 0.551
R1592 SD2R.n211 SD2R.t74 0.551
R1593 SD2R.n182 SD2R.n181 0.43
R1594 SD2R.n185 SD2R.n78 0.35
R1595 SD2R.n183 SD2R.n129 0.347
R1596 SD2R.n187 SD2R.n25 0.347
R1597 SD2R.n184 SD2R.n103 0.224
R1598 SD2R.n213 SD2R.n212 0.224
R1599 SD2R.n185 SD2R.n184 0.091
R1600 SD2R.n186 SD2R.n185 0.08
R1601 SD2R SD2R.n213 0.054
R1602 SD2R.n183 SD2R.n182 0.05
R1603 SD2R.n187 SD2R.n186 0.05
R1604 SD2R.n184 SD2R.n183 0.039
R1605 SD2R.n213 SD2R.n187 0.039
R1606 SD2R.n75 SD2R.n73 0.007
R1607 SD2R.n73 SD2R.n72 0.007
R1608 SD2R.n72 SD2R.n71 0.007
R1609 SD2R.n71 SD2R.n70 0.007
R1610 SD2R.n70 SD2R.n69 0.007
R1611 SD2R.n69 SD2R.n68 0.007
R1612 SD2R.n68 SD2R.n67 0.007
R1613 SD2R.n67 SD2R.n66 0.007
R1614 SD2R.n66 SD2R.n65 0.007
R1615 SD2R.n65 SD2R.n64 0.007
R1616 SD2R.n64 SD2R.n63 0.007
R1617 SD2R.n96 SD2R.n95 0.007
R1618 SD2R.n97 SD2R.n96 0.007
R1619 SD2R.n98 SD2R.n97 0.007
R1620 SD2R.n89 SD2R.n88 0.007
R1621 SD2R.n88 SD2R.n87 0.007
R1622 SD2R.n87 SD2R.n86 0.007
R1623 SD2R.n86 SD2R.n85 0.007
R1624 SD2R.n125 SD2R.n124 0.007
R1625 SD2R.n124 SD2R.n123 0.007
R1626 SD2R.n123 SD2R.n122 0.007
R1627 SD2R.n122 SD2R.n121 0.007
R1628 SD2R.n121 SD2R.n120 0.007
R1629 SD2R.n120 SD2R.n119 0.007
R1630 SD2R.n119 SD2R.n118 0.007
R1631 SD2R.n118 SD2R.n117 0.007
R1632 SD2R.n117 SD2R.n116 0.007
R1633 SD2R.n116 SD2R.n115 0.007
R1634 SD2R.n142 SD2R.n141 0.007
R1635 SD2R.n143 SD2R.n142 0.007
R1636 SD2R.n144 SD2R.n143 0.007
R1637 SD2R.n145 SD2R.n144 0.007
R1638 SD2R.n146 SD2R.n145 0.007
R1639 SD2R.n147 SD2R.n146 0.007
R1640 SD2R.n148 SD2R.n147 0.007
R1641 SD2R.n149 SD2R.n148 0.007
R1642 SD2R.n150 SD2R.n149 0.007
R1643 SD2R.n152 SD2R.n150 0.007
R1644 SD2R.n177 SD2R.n176 0.007
R1645 SD2R.n176 SD2R.n175 0.007
R1646 SD2R.n175 SD2R.n174 0.007
R1647 SD2R.n174 SD2R.n173 0.007
R1648 SD2R.n173 SD2R.n172 0.007
R1649 SD2R.n172 SD2R.n171 0.007
R1650 SD2R.n171 SD2R.n170 0.007
R1651 SD2R.n170 SD2R.n169 0.007
R1652 SD2R.n169 SD2R.n168 0.007
R1653 SD2R.n168 SD2R.n167 0.007
R1654 SD2R.n21 SD2R.n20 0.007
R1655 SD2R.n20 SD2R.n19 0.007
R1656 SD2R.n19 SD2R.n18 0.007
R1657 SD2R.n18 SD2R.n17 0.007
R1658 SD2R.n17 SD2R.n16 0.007
R1659 SD2R.n16 SD2R.n15 0.007
R1660 SD2R.n15 SD2R.n14 0.007
R1661 SD2R.n14 SD2R.n13 0.007
R1662 SD2R.n13 SD2R.n12 0.007
R1663 SD2R.n12 SD2R.n11 0.007
R1664 SD2R.n38 SD2R.n37 0.007
R1665 SD2R.n39 SD2R.n38 0.007
R1666 SD2R.n40 SD2R.n39 0.007
R1667 SD2R.n41 SD2R.n40 0.007
R1668 SD2R.n42 SD2R.n41 0.007
R1669 SD2R.n43 SD2R.n42 0.007
R1670 SD2R.n44 SD2R.n43 0.007
R1671 SD2R.n45 SD2R.n44 0.007
R1672 SD2R.n46 SD2R.n45 0.007
R1673 SD2R.n48 SD2R.n46 0.007
R1674 SD2R.n194 SD2R.n193 0.007
R1675 SD2R.n195 SD2R.n194 0.007
R1676 SD2R.n196 SD2R.n195 0.007
R1677 SD2R.n210 SD2R.n209 0.007
R1678 SD2R.n209 SD2R.n208 0.007
R1679 SD2R.n208 SD2R.n207 0.007
R1680 SD2R.n207 SD2R.n206 0.007
R1681 SD2R.n129 SD2R.n125 0.006
R1682 SD2R.n181 SD2R.n177 0.006
R1683 SD2R.n25 SD2R.n21 0.006
R1684 SD2R.n103 SD2R.n98 0.005
R1685 SD2R.n212 SD2R.n196 0.005
R1686 SD2R.n103 SD2R.n89 0.004
R1687 SD2R.n212 SD2R.n210 0.004
R1688 SD2R.n182 SD2R.n152 0.004
R1689 SD2R.n186 SD2R.n48 0.004
R1690 SD2R.n78 SD2R.n75 0.001
R1691 SD1R.n11 SD1R.t63 1.972
R1692 SD1R.n62 SD1R.t69 1.972
R1693 SD1R.n25 SD1R.t50 1.963
R1694 SD1R.n77 SD1R.t70 1.96
R1695 SD1R.n86 SD1R.n85 1.435
R1696 SD1R.n97 SD1R.n96 1.435
R1697 SD1R.n42 SD1R.n41 1.435
R1698 SD1R.n32 SD1R.n31 1.435
R1699 SD1R.n90 SD1R.n82 1.428
R1700 SD1R.n89 SD1R.n83 1.428
R1701 SD1R.n86 SD1R.n84 1.428
R1702 SD1R.n97 SD1R.n95 1.428
R1703 SD1R.n98 SD1R.n94 1.428
R1704 SD1R.n99 SD1R.n93 1.428
R1705 SD1R.n100 SD1R.n92 1.428
R1706 SD1R.n101 SD1R.n91 1.428
R1707 SD1R.n45 SD1R.n37 1.428
R1708 SD1R.n44 SD1R.n38 1.428
R1709 SD1R.n43 SD1R.n39 1.428
R1710 SD1R.n42 SD1R.n40 1.428
R1711 SD1R.n32 SD1R.n30 1.428
R1712 SD1R.n33 SD1R.n29 1.428
R1713 SD1R.n34 SD1R.n28 1.428
R1714 SD1R.n35 SD1R.n27 1.428
R1715 SD1R.n36 SD1R.n26 1.428
R1716 SD1R.n88 SD1R.n87 1.427
R1717 SD1R.n62 SD1R.n61 1.414
R1718 SD1R.n63 SD1R.n60 1.414
R1719 SD1R.n64 SD1R.n59 1.414
R1720 SD1R.n65 SD1R.n58 1.414
R1721 SD1R.n66 SD1R.n57 1.414
R1722 SD1R.n67 SD1R.n56 1.414
R1723 SD1R.n68 SD1R.n55 1.414
R1724 SD1R.n69 SD1R.n54 1.414
R1725 SD1R.n70 SD1R.n53 1.414
R1726 SD1R.n71 SD1R.n52 1.414
R1727 SD1R.n72 SD1R.n51 1.414
R1728 SD1R.n21 SD1R.n0 1.414
R1729 SD1R.n20 SD1R.n1 1.414
R1730 SD1R.n19 SD1R.n2 1.414
R1731 SD1R.n18 SD1R.n3 1.414
R1732 SD1R.n17 SD1R.n4 1.414
R1733 SD1R.n16 SD1R.n5 1.414
R1734 SD1R.n15 SD1R.n6 1.414
R1735 SD1R.n14 SD1R.n7 1.414
R1736 SD1R.n13 SD1R.n8 1.414
R1737 SD1R.n12 SD1R.n9 1.414
R1738 SD1R.n11 SD1R.n10 1.414
R1739 SD1R.n25 SD1R.n24 1.412
R1740 SD1R.n25 SD1R.n23 1.412
R1741 SD1R.n25 SD1R.n22 1.412
R1742 SD1R.n74 SD1R.n73 1.41
R1743 SD1R.n77 SD1R.n75 1.409
R1744 SD1R.n77 SD1R.n76 1.409
R1745 SD1R.n50 SD1R.n46 1.28
R1746 SD1R.n50 SD1R.n47 1.28
R1747 SD1R.n50 SD1R.n48 1.28
R1748 SD1R.n50 SD1R.n49 1.28
R1749 SD1R.n102 SD1R.n81 1.28
R1750 SD1R.n102 SD1R.n80 1.28
R1751 SD1R.n102 SD1R.n79 1.28
R1752 SD1R.n102 SD1R.n78 1.28
R1753 SD1R.n82 SD1R.t105 0.551
R1754 SD1R.n82 SD1R.t36 0.551
R1755 SD1R.n83 SD1R.t65 0.551
R1756 SD1R.n83 SD1R.t8 0.551
R1757 SD1R.n84 SD1R.t3 0.551
R1758 SD1R.n84 SD1R.t25 0.551
R1759 SD1R.n85 SD1R.t57 0.551
R1760 SD1R.n85 SD1R.t28 0.551
R1761 SD1R.n96 SD1R.t11 0.551
R1762 SD1R.n96 SD1R.t75 0.551
R1763 SD1R.n95 SD1R.t111 0.551
R1764 SD1R.n95 SD1R.t80 0.551
R1765 SD1R.n94 SD1R.t37 0.551
R1766 SD1R.n94 SD1R.t43 0.551
R1767 SD1R.n93 SD1R.t0 0.551
R1768 SD1R.n93 SD1R.t95 0.551
R1769 SD1R.n92 SD1R.t7 0.551
R1770 SD1R.n92 SD1R.t103 0.551
R1771 SD1R.n91 SD1R.t61 0.551
R1772 SD1R.n91 SD1R.t119 0.551
R1773 SD1R.n81 SD1R.t13 0.551
R1774 SD1R.n81 SD1R.t110 0.551
R1775 SD1R.n80 SD1R.t47 0.551
R1776 SD1R.n80 SD1R.t21 0.551
R1777 SD1R.n79 SD1R.t115 0.551
R1778 SD1R.n79 SD1R.t89 0.551
R1779 SD1R.n78 SD1R.t22 0.551
R1780 SD1R.n78 SD1R.t84 0.551
R1781 SD1R.n61 SD1R.t1 0.551
R1782 SD1R.n61 SD1R.t76 0.551
R1783 SD1R.n60 SD1R.t55 0.551
R1784 SD1R.n60 SD1R.t48 0.551
R1785 SD1R.n59 SD1R.t4 0.551
R1786 SD1R.n59 SD1R.t10 0.551
R1787 SD1R.n58 SD1R.t58 0.551
R1788 SD1R.n58 SD1R.t51 0.551
R1789 SD1R.n57 SD1R.t62 0.551
R1790 SD1R.n57 SD1R.t106 0.551
R1791 SD1R.n56 SD1R.t101 0.551
R1792 SD1R.n56 SD1R.t64 0.551
R1793 SD1R.n55 SD1R.t30 0.551
R1794 SD1R.n55 SD1R.t109 0.551
R1795 SD1R.n54 SD1R.t113 0.551
R1796 SD1R.n54 SD1R.t66 0.551
R1797 SD1R.n53 SD1R.t45 0.551
R1798 SD1R.n53 SD1R.t39 0.551
R1799 SD1R.n52 SD1R.t117 0.551
R1800 SD1R.n52 SD1R.t81 0.551
R1801 SD1R.n51 SD1R.t87 0.551
R1802 SD1R.n51 SD1R.t42 0.551
R1803 SD1R.n73 SD1R.t19 0.551
R1804 SD1R.n73 SD1R.t93 0.551
R1805 SD1R.n75 SD1R.t90 0.551
R1806 SD1R.n75 SD1R.t44 0.551
R1807 SD1R.n76 SD1R.t23 0.551
R1808 SD1R.n76 SD1R.t96 0.551
R1809 SD1R.n37 SD1R.t53 0.551
R1810 SD1R.n37 SD1R.t79 0.551
R1811 SD1R.n38 SD1R.t46 0.551
R1812 SD1R.n38 SD1R.t27 0.551
R1813 SD1R.n39 SD1R.t116 0.551
R1814 SD1R.n39 SD1R.t18 0.551
R1815 SD1R.n40 SD1R.t33 0.551
R1816 SD1R.n40 SD1R.t86 0.551
R1817 SD1R.n41 SD1R.t59 0.551
R1818 SD1R.n41 SD1R.t5 0.551
R1819 SD1R.n31 SD1R.t72 0.551
R1820 SD1R.n31 SD1R.t14 0.551
R1821 SD1R.n30 SD1R.t24 0.551
R1822 SD1R.n30 SD1R.t98 0.551
R1823 SD1R.n29 SD1R.t35 0.551
R1824 SD1R.n29 SD1R.t71 0.551
R1825 SD1R.n28 SD1R.t73 0.551
R1826 SD1R.n28 SD1R.t100 0.551
R1827 SD1R.n27 SD1R.t112 0.551
R1828 SD1R.n27 SD1R.t15 0.551
R1829 SD1R.n26 SD1R.t60 0.551
R1830 SD1R.n26 SD1R.t114 0.551
R1831 SD1R.n46 SD1R.t108 0.551
R1832 SD1R.n46 SD1R.t9 0.551
R1833 SD1R.n47 SD1R.t67 0.551
R1834 SD1R.n47 SD1R.t17 0.551
R1835 SD1R.n48 SD1R.t41 0.551
R1836 SD1R.n48 SD1R.t68 0.551
R1837 SD1R.n49 SD1R.t92 0.551
R1838 SD1R.n49 SD1R.t32 0.551
R1839 SD1R.n0 SD1R.t56 0.551
R1840 SD1R.n0 SD1R.t104 0.551
R1841 SD1R.n1 SD1R.t16 0.551
R1842 SD1R.n1 SD1R.t52 0.551
R1843 SD1R.n2 SD1R.t99 0.551
R1844 SD1R.n2 SD1R.t107 0.551
R1845 SD1R.n3 SD1R.t29 0.551
R1846 SD1R.n3 SD1R.t77 0.551
R1847 SD1R.n4 SD1R.t102 0.551
R1848 SD1R.n4 SD1R.t26 0.551
R1849 SD1R.n5 SD1R.t31 0.551
R1850 SD1R.n5 SD1R.t78 0.551
R1851 SD1R.n6 SD1R.t83 0.551
R1852 SD1R.n6 SD1R.t40 0.551
R1853 SD1R.n7 SD1R.t74 0.551
R1854 SD1R.n7 SD1R.t82 0.551
R1855 SD1R.n8 SD1R.t6 0.551
R1856 SD1R.n8 SD1R.t12 0.551
R1857 SD1R.n9 SD1R.t88 0.551
R1858 SD1R.n9 SD1R.t94 0.551
R1859 SD1R.n10 SD1R.t20 0.551
R1860 SD1R.n10 SD1R.t54 0.551
R1861 SD1R.n22 SD1R.t97 0.551
R1862 SD1R.n22 SD1R.t34 0.551
R1863 SD1R.n23 SD1R.t38 0.551
R1864 SD1R.n23 SD1R.t85 0.551
R1865 SD1R.n24 SD1R.t2 0.551
R1866 SD1R.n24 SD1R.t49 0.551
R1867 SD1R.n87 SD1R.t118 0.551
R1868 SD1R.n87 SD1R.t91 0.551
R1869 SD1R.n103 SD1R.n102 0.349
R1870 SD1R.n103 SD1R.n77 0.306
R1871 SD1R.n105 SD1R.n25 0.306
R1872 SD1R.n104 SD1R.n50 0.18
R1873 SD1R.n105 SD1R.n104 0.154
R1874 SD1R.n104 SD1R.n103 0.091
R1875 SD1R SD1R.n105 0.021
R1876 SD1R.n74 SD1R.n72 0.007
R1877 SD1R.n72 SD1R.n71 0.007
R1878 SD1R.n71 SD1R.n70 0.007
R1879 SD1R.n70 SD1R.n69 0.007
R1880 SD1R.n69 SD1R.n68 0.007
R1881 SD1R.n68 SD1R.n67 0.007
R1882 SD1R.n67 SD1R.n66 0.007
R1883 SD1R.n66 SD1R.n65 0.007
R1884 SD1R.n65 SD1R.n64 0.007
R1885 SD1R.n64 SD1R.n63 0.007
R1886 SD1R.n63 SD1R.n62 0.007
R1887 SD1R.n43 SD1R.n42 0.007
R1888 SD1R.n44 SD1R.n43 0.007
R1889 SD1R.n45 SD1R.n44 0.007
R1890 SD1R.n36 SD1R.n35 0.007
R1891 SD1R.n35 SD1R.n34 0.007
R1892 SD1R.n34 SD1R.n33 0.007
R1893 SD1R.n33 SD1R.n32 0.007
R1894 SD1R.n21 SD1R.n20 0.007
R1895 SD1R.n20 SD1R.n19 0.007
R1896 SD1R.n19 SD1R.n18 0.007
R1897 SD1R.n18 SD1R.n17 0.007
R1898 SD1R.n17 SD1R.n16 0.007
R1899 SD1R.n16 SD1R.n15 0.007
R1900 SD1R.n15 SD1R.n14 0.007
R1901 SD1R.n14 SD1R.n13 0.007
R1902 SD1R.n13 SD1R.n12 0.007
R1903 SD1R.n12 SD1R.n11 0.007
R1904 SD1R.n88 SD1R.n86 0.007
R1905 SD1R.n89 SD1R.n88 0.007
R1906 SD1R.n90 SD1R.n89 0.007
R1907 SD1R.n101 SD1R.n100 0.007
R1908 SD1R.n100 SD1R.n99 0.007
R1909 SD1R.n99 SD1R.n98 0.007
R1910 SD1R.n98 SD1R.n97 0.007
R1911 SD1R.n25 SD1R.n21 0.006
R1912 SD1R.n50 SD1R.n45 0.005
R1913 SD1R.n102 SD1R.n90 0.005
R1914 SD1R.n50 SD1R.n36 0.004
R1915 SD1R.n102 SD1R.n101 0.004
R1916 SD1R.n77 SD1R.n74 0.001
R1917 SD3L.n203 SD3L.t154 1.972
R1918 SD3L.n193 SD3L.t153 1.972
R1919 SD3L.n38 SD3L.t105 1.972
R1920 SD3L.n118 SD3L.t52 1.972
R1921 SD3L.n175 SD3L.t132 1.972
R1922 SD3L.n165 SD3L.t143 1.972
R1923 SD3L.n132 SD3L.t6 1.963
R1924 SD3L.n52 SD3L.t86 1.962
R1925 SD3L.n11 SD3L.n10 1.435
R1926 SD3L.n64 SD3L.n63 1.435
R1927 SD3L.n91 SD3L.n90 1.435
R1928 SD3L.n144 SD3L.n143 1.435
R1929 SD3L.n20 SD3L.n0 1.428
R1930 SD3L.n19 SD3L.n1 1.428
R1931 SD3L.n18 SD3L.n2 1.428
R1932 SD3L.n17 SD3L.n3 1.428
R1933 SD3L.n16 SD3L.n4 1.428
R1934 SD3L.n15 SD3L.n5 1.428
R1935 SD3L.n14 SD3L.n6 1.428
R1936 SD3L.n13 SD3L.n7 1.428
R1937 SD3L.n12 SD3L.n8 1.428
R1938 SD3L.n11 SD3L.n9 1.428
R1939 SD3L.n73 SD3L.n53 1.428
R1940 SD3L.n72 SD3L.n54 1.428
R1941 SD3L.n71 SD3L.n55 1.428
R1942 SD3L.n70 SD3L.n56 1.428
R1943 SD3L.n69 SD3L.n57 1.428
R1944 SD3L.n68 SD3L.n58 1.428
R1945 SD3L.n67 SD3L.n59 1.428
R1946 SD3L.n66 SD3L.n60 1.428
R1947 SD3L.n65 SD3L.n61 1.428
R1948 SD3L.n64 SD3L.n62 1.428
R1949 SD3L.n100 SD3L.n80 1.428
R1950 SD3L.n99 SD3L.n81 1.428
R1951 SD3L.n98 SD3L.n82 1.428
R1952 SD3L.n97 SD3L.n83 1.428
R1953 SD3L.n96 SD3L.n84 1.428
R1954 SD3L.n95 SD3L.n85 1.428
R1955 SD3L.n94 SD3L.n86 1.428
R1956 SD3L.n93 SD3L.n87 1.428
R1957 SD3L.n92 SD3L.n88 1.428
R1958 SD3L.n91 SD3L.n89 1.428
R1959 SD3L.n153 SD3L.n133 1.428
R1960 SD3L.n152 SD3L.n134 1.428
R1961 SD3L.n151 SD3L.n135 1.428
R1962 SD3L.n150 SD3L.n136 1.428
R1963 SD3L.n149 SD3L.n137 1.428
R1964 SD3L.n148 SD3L.n138 1.428
R1965 SD3L.n147 SD3L.n139 1.428
R1966 SD3L.n146 SD3L.n140 1.428
R1967 SD3L.n145 SD3L.n141 1.428
R1968 SD3L.n144 SD3L.n142 1.428
R1969 SD3L.n207 SD3L.n198 1.414
R1970 SD3L.n206 SD3L.n199 1.414
R1971 SD3L.n205 SD3L.n200 1.414
R1972 SD3L.n204 SD3L.n201 1.414
R1973 SD3L.n203 SD3L.n202 1.414
R1974 SD3L.n193 SD3L.n192 1.414
R1975 SD3L.n194 SD3L.n191 1.414
R1976 SD3L.n195 SD3L.n190 1.414
R1977 SD3L.n196 SD3L.n189 1.414
R1978 SD3L.n197 SD3L.n188 1.414
R1979 SD3L.n48 SD3L.n27 1.414
R1980 SD3L.n47 SD3L.n28 1.414
R1981 SD3L.n46 SD3L.n29 1.414
R1982 SD3L.n45 SD3L.n30 1.414
R1983 SD3L.n44 SD3L.n31 1.414
R1984 SD3L.n43 SD3L.n32 1.414
R1985 SD3L.n42 SD3L.n33 1.414
R1986 SD3L.n41 SD3L.n34 1.414
R1987 SD3L.n40 SD3L.n35 1.414
R1988 SD3L.n39 SD3L.n36 1.414
R1989 SD3L.n38 SD3L.n37 1.414
R1990 SD3L.n128 SD3L.n107 1.414
R1991 SD3L.n127 SD3L.n108 1.414
R1992 SD3L.n126 SD3L.n109 1.414
R1993 SD3L.n125 SD3L.n110 1.414
R1994 SD3L.n124 SD3L.n111 1.414
R1995 SD3L.n123 SD3L.n112 1.414
R1996 SD3L.n122 SD3L.n113 1.414
R1997 SD3L.n121 SD3L.n114 1.414
R1998 SD3L.n120 SD3L.n115 1.414
R1999 SD3L.n119 SD3L.n116 1.414
R2000 SD3L.n118 SD3L.n117 1.414
R2001 SD3L.n179 SD3L.n170 1.414
R2002 SD3L.n178 SD3L.n171 1.414
R2003 SD3L.n177 SD3L.n172 1.414
R2004 SD3L.n176 SD3L.n173 1.414
R2005 SD3L.n175 SD3L.n174 1.414
R2006 SD3L.n165 SD3L.n164 1.414
R2007 SD3L.n166 SD3L.n163 1.414
R2008 SD3L.n167 SD3L.n162 1.414
R2009 SD3L.n168 SD3L.n161 1.414
R2010 SD3L.n169 SD3L.n160 1.414
R2011 SD3L.n132 SD3L.n131 1.412
R2012 SD3L.n132 SD3L.n130 1.412
R2013 SD3L.n132 SD3L.n129 1.412
R2014 SD3L.n184 SD3L.n183 1.412
R2015 SD3L.n184 SD3L.n182 1.412
R2016 SD3L.n184 SD3L.n181 1.412
R2017 SD3L.n184 SD3L.n180 1.412
R2018 SD3L.n211 SD3L.n210 1.412
R2019 SD3L.n211 SD3L.n209 1.412
R2020 SD3L.n211 SD3L.n208 1.412
R2021 SD3L.n211 SD3L.n187 1.41
R2022 SD3L.n52 SD3L.n51 1.409
R2023 SD3L.n52 SD3L.n50 1.409
R2024 SD3L.n52 SD3L.n49 1.409
R2025 SD3L.n22 SD3L.n21 1.281
R2026 SD3L.n75 SD3L.n74 1.281
R2027 SD3L.n102 SD3L.n101 1.281
R2028 SD3L.n155 SD3L.n154 1.281
R2029 SD3L.n26 SD3L.n23 1.28
R2030 SD3L.n26 SD3L.n24 1.28
R2031 SD3L.n26 SD3L.n25 1.28
R2032 SD3L.n79 SD3L.n76 1.28
R2033 SD3L.n79 SD3L.n77 1.28
R2034 SD3L.n79 SD3L.n78 1.28
R2035 SD3L.n106 SD3L.n103 1.28
R2036 SD3L.n106 SD3L.n104 1.28
R2037 SD3L.n106 SD3L.n105 1.28
R2038 SD3L.n159 SD3L.n156 1.28
R2039 SD3L.n159 SD3L.n157 1.28
R2040 SD3L.n159 SD3L.n158 1.28
R2041 SD3L.n198 SD3L.t199 0.551
R2042 SD3L.n198 SD3L.t163 0.551
R2043 SD3L.n199 SD3L.t172 0.551
R2044 SD3L.n199 SD3L.t121 0.551
R2045 SD3L.n200 SD3L.t220 0.551
R2046 SD3L.n200 SD3L.t177 0.551
R2047 SD3L.n201 SD3L.t175 0.551
R2048 SD3L.n201 SD3L.t123 0.551
R2049 SD3L.n202 SD3L.t224 0.551
R2050 SD3L.n202 SD3L.t180 0.551
R2051 SD3L.n192 SD3L.t204 0.551
R2052 SD3L.n192 SD3L.t157 0.551
R2053 SD3L.n191 SD3L.t136 0.551
R2054 SD3L.n191 SD3L.t128 0.551
R2055 SD3L.n190 SD3L.t207 0.551
R2056 SD3L.n190 SD3L.t211 0.551
R2057 SD3L.n189 SD3L.t140 0.551
R2058 SD3L.n189 SD3L.t130 0.551
R2059 SD3L.n188 SD3L.t142 0.551
R2060 SD3L.n188 SD3L.t190 0.551
R2061 SD3L.n208 SD3L.t196 0.551
R2062 SD3L.n208 SD3L.t150 0.551
R2063 SD3L.n209 SD3L.t231 0.551
R2064 SD3L.n209 SD3L.t194 0.551
R2065 SD3L.n210 SD3L.t185 0.551
R2066 SD3L.n210 SD3L.t148 0.551
R2067 SD3L.n0 SD3L.t214 0.551
R2068 SD3L.n0 SD3L.t170 0.551
R2069 SD3L.n1 SD3L.t179 0.551
R2070 SD3L.n1 SD3L.t174 0.551
R2071 SD3L.n2 SD3L.t227 0.551
R2072 SD3L.n2 SD3L.t222 0.551
R2073 SD3L.n3 SD3L.t182 0.551
R2074 SD3L.n3 SD3L.t144 0.551
R2075 SD3L.n4 SD3L.t155 0.551
R2076 SD3L.n4 SD3L.t225 0.551
R2077 SD3L.n5 SD3L.t206 0.551
R2078 SD3L.n5 SD3L.t159 0.551
R2079 SD3L.n6 SD3L.t203 0.551
R2080 SD3L.n6 SD3L.t236 0.551
R2081 SD3L.n7 SD3L.t134 0.551
R2082 SD3L.n7 SD3L.t127 0.551
R2083 SD3L.n8 SD3L.t217 0.551
R2084 SD3L.n8 SD3L.t187 0.551
R2085 SD3L.n9 SD3L.t139 0.551
R2086 SD3L.n9 SD3L.t146 0.551
R2087 SD3L.n10 SD3L.t228 0.551
R2088 SD3L.n10 SD3L.t189 0.551
R2089 SD3L.n21 SD3L.t176 0.551
R2090 SD3L.n21 SD3L.t126 0.551
R2091 SD3L.n23 SD3L.t120 0.551
R2092 SD3L.n23 SD3L.t168 0.551
R2093 SD3L.n24 SD3L.t162 0.551
R2094 SD3L.n24 SD3L.t234 0.551
R2095 SD3L.n25 SD3L.t201 0.551
R2096 SD3L.n25 SD3L.t195 0.551
R2097 SD3L.n51 SD3L.t84 0.551
R2098 SD3L.n51 SD3L.t10 0.551
R2099 SD3L.n50 SD3L.t62 0.551
R2100 SD3L.n50 SD3L.t17 0.551
R2101 SD3L.n49 SD3L.t23 0.551
R2102 SD3L.n49 SD3L.t70 0.551
R2103 SD3L.n27 SD3L.t51 0.551
R2104 SD3L.n27 SD3L.t60 0.551
R2105 SD3L.n28 SD3L.t15 0.551
R2106 SD3L.n28 SD3L.t118 0.551
R2107 SD3L.n29 SD3L.t12 0.551
R2108 SD3L.n29 SD3L.t44 0.551
R2109 SD3L.n30 SD3L.t32 0.551
R2110 SD3L.n30 SD3L.t34 0.551
R2111 SD3L.n31 SD3L.t5 0.551
R2112 SD3L.n31 SD3L.t106 0.551
R2113 SD3L.n32 SD3L.t47 0.551
R2114 SD3L.n32 SD3L.t13 0.551
R2115 SD3L.n33 SD3L.t111 0.551
R2116 SD3L.n33 SD3L.t42 0.551
R2117 SD3L.n34 SD3L.t110 0.551
R2118 SD3L.n34 SD3L.t80 0.551
R2119 SD3L.n35 SD3L.t115 0.551
R2120 SD3L.n35 SD3L.t78 0.551
R2121 SD3L.n36 SD3L.t4 0.551
R2122 SD3L.n36 SD3L.t91 0.551
R2123 SD3L.n37 SD3L.t103 0.551
R2124 SD3L.n37 SD3L.t24 0.551
R2125 SD3L.n53 SD3L.t114 0.551
R2126 SD3L.n53 SD3L.t85 0.551
R2127 SD3L.n54 SD3L.t39 0.551
R2128 SD3L.n54 SD3L.t35 0.551
R2129 SD3L.n55 SD3L.t100 0.551
R2130 SD3L.n55 SD3L.t33 0.551
R2131 SD3L.n56 SD3L.t45 0.551
R2132 SD3L.n56 SD3L.t50 0.551
R2133 SD3L.n57 SD3L.t69 0.551
R2134 SD3L.n57 SD3L.t43 0.551
R2135 SD3L.n58 SD3L.t119 0.551
R2136 SD3L.n58 SD3L.t107 0.551
R2137 SD3L.n59 SD3L.t0 0.551
R2138 SD3L.n59 SD3L.t59 0.551
R2139 SD3L.n60 SD3L.t22 0.551
R2140 SD3L.n60 SD3L.t82 0.551
R2141 SD3L.n61 SD3L.t49 0.551
R2142 SD3L.n61 SD3L.t57 0.551
R2143 SD3L.n62 SD3L.t37 0.551
R2144 SD3L.n62 SD3L.t113 0.551
R2145 SD3L.n63 SD3L.t31 0.551
R2146 SD3L.n63 SD3L.t2 0.551
R2147 SD3L.n74 SD3L.t56 0.551
R2148 SD3L.n74 SD3L.t1 0.551
R2149 SD3L.n76 SD3L.t46 0.551
R2150 SD3L.n76 SD3L.t87 0.551
R2151 SD3L.n77 SD3L.t19 0.551
R2152 SD3L.n77 SD3L.t99 0.551
R2153 SD3L.n78 SD3L.t95 0.551
R2154 SD3L.n78 SD3L.t64 0.551
R2155 SD3L.n80 SD3L.t202 0.551
R2156 SD3L.n80 SD3L.t124 0.551
R2157 SD3L.n81 SD3L.t141 0.551
R2158 SD3L.n81 SD3L.t147 0.551
R2159 SD3L.n82 SD3L.t209 0.551
R2160 SD3L.n82 SD3L.t213 0.551
R2161 SD3L.n83 SD3L.t122 0.551
R2162 SD3L.n83 SD3L.t165 0.551
R2163 SD3L.n84 SD3L.t167 0.551
R2164 SD3L.n84 SD3L.t200 0.551
R2165 SD3L.n85 SD3L.t233 0.551
R2166 SD3L.n85 SD3L.t161 0.551
R2167 SD3L.n86 SD3L.t152 0.551
R2168 SD3L.n86 SD3L.t198 0.551
R2169 SD3L.n87 SD3L.t230 0.551
R2170 SD3L.n87 SD3L.t223 0.551
R2171 SD3L.n88 SD3L.t149 0.551
R2172 SD3L.n88 SD3L.t192 0.551
R2173 SD3L.n89 SD3L.t216 0.551
R2174 SD3L.n89 SD3L.t219 0.551
R2175 SD3L.n90 SD3L.t138 0.551
R2176 SD3L.n90 SD3L.t171 0.551
R2177 SD3L.n101 SD3L.t133 0.551
R2178 SD3L.n101 SD3L.t184 0.551
R2179 SD3L.n103 SD3L.t193 0.551
R2180 SD3L.n103 SD3L.t218 0.551
R2181 SD3L.n104 SD3L.t210 0.551
R2182 SD3L.n104 SD3L.t197 0.551
R2183 SD3L.n105 SD3L.t151 0.551
R2184 SD3L.n105 SD3L.t145 0.551
R2185 SD3L.n107 SD3L.t9 0.551
R2186 SD3L.n107 SD3L.t83 0.551
R2187 SD3L.n108 SD3L.t18 0.551
R2188 SD3L.n108 SD3L.t66 0.551
R2189 SD3L.n109 SD3L.t94 0.551
R2190 SD3L.n109 SD3L.t26 0.551
R2191 SD3L.n110 SD3L.t20 0.551
R2192 SD3L.n110 SD3L.t53 0.551
R2193 SD3L.n111 SD3L.t72 0.551
R2194 SD3L.n111 SD3L.t36 0.551
R2195 SD3L.n112 SD3L.t65 0.551
R2196 SD3L.n112 SD3L.t90 0.551
R2197 SD3L.n113 SD3L.t93 0.551
R2198 SD3L.n113 SD3L.t67 0.551
R2199 SD3L.n114 SD3L.t71 0.551
R2200 SD3L.n114 SD3L.t28 0.551
R2201 SD3L.n115 SD3L.t79 0.551
R2202 SD3L.n115 SD3L.t116 0.551
R2203 SD3L.n116 SD3L.t16 0.551
R2204 SD3L.n116 SD3L.t92 0.551
R2205 SD3L.n117 SD3L.t97 0.551
R2206 SD3L.n117 SD3L.t77 0.551
R2207 SD3L.n129 SD3L.t98 0.551
R2208 SD3L.n129 SD3L.t63 0.551
R2209 SD3L.n130 SD3L.t96 0.551
R2210 SD3L.n130 SD3L.t112 0.551
R2211 SD3L.n131 SD3L.t21 0.551
R2212 SD3L.n131 SD3L.t30 0.551
R2213 SD3L.n133 SD3L.t61 0.551
R2214 SD3L.n133 SD3L.t108 0.551
R2215 SD3L.n134 SD3L.t81 0.551
R2216 SD3L.n134 SD3L.t55 0.551
R2217 SD3L.n135 SD3L.t76 0.551
R2218 SD3L.n135 SD3L.t117 0.551
R2219 SD3L.n136 SD3L.t74 0.551
R2220 SD3L.n136 SD3L.t89 0.551
R2221 SD3L.n137 SD3L.t109 0.551
R2222 SD3L.n137 SD3L.t14 0.551
R2223 SD3L.n138 SD3L.t68 0.551
R2224 SD3L.n138 SD3L.t41 0.551
R2225 SD3L.n139 SD3L.t54 0.551
R2226 SD3L.n139 SD3L.t25 0.551
R2227 SD3L.n140 SD3L.t27 0.551
R2228 SD3L.n140 SD3L.t75 0.551
R2229 SD3L.n141 SD3L.t11 0.551
R2230 SD3L.n141 SD3L.t102 0.551
R2231 SD3L.n142 SD3L.t38 0.551
R2232 SD3L.n142 SD3L.t73 0.551
R2233 SD3L.n143 SD3L.t40 0.551
R2234 SD3L.n143 SD3L.t48 0.551
R2235 SD3L.n154 SD3L.t104 0.551
R2236 SD3L.n154 SD3L.t101 0.551
R2237 SD3L.n156 SD3L.t88 0.551
R2238 SD3L.n156 SD3L.t29 0.551
R2239 SD3L.n157 SD3L.t58 0.551
R2240 SD3L.n157 SD3L.t3 0.551
R2241 SD3L.n158 SD3L.t8 0.551
R2242 SD3L.n158 SD3L.t7 0.551
R2243 SD3L.n170 SD3L.t215 0.551
R2244 SD3L.n170 SD3L.t131 0.551
R2245 SD3L.n171 SD3L.t137 0.551
R2246 SD3L.n171 SD3L.t188 0.551
R2247 SD3L.n172 SD3L.t205 0.551
R2248 SD3L.n172 SD3L.t129 0.551
R2249 SD3L.n173 SD3L.t237 0.551
R2250 SD3L.n173 SD3L.t169 0.551
R2251 SD3L.n174 SD3L.t181 0.551
R2252 SD3L.n174 SD3L.t235 0.551
R2253 SD3L.n164 SD3L.t221 0.551
R2254 SD3L.n164 SD3L.t135 0.551
R2255 SD3L.n163 SD3L.t173 0.551
R2256 SD3L.n163 SD3L.t178 0.551
R2257 SD3L.n162 SD3L.t208 0.551
R2258 SD3L.n162 SD3L.t212 0.551
R2259 SD3L.n161 SD3L.t156 0.551
R2260 SD3L.n161 SD3L.t164 0.551
R2261 SD3L.n160 SD3L.t166 0.551
R2262 SD3L.n160 SD3L.t239 0.551
R2263 SD3L.n180 SD3L.t183 0.551
R2264 SD3L.n180 SD3L.t191 0.551
R2265 SD3L.n181 SD3L.t229 0.551
R2266 SD3L.n181 SD3L.t158 0.551
R2267 SD3L.n182 SD3L.t186 0.551
R2268 SD3L.n182 SD3L.t226 0.551
R2269 SD3L.n183 SD3L.t232 0.551
R2270 SD3L.n183 SD3L.t160 0.551
R2271 SD3L.n187 SD3L.t125 0.551
R2272 SD3L.n187 SD3L.t238 0.551
R2273 SD3L.n185 SD3L.n184 0.455
R2274 SD3L.n212 SD3L.n211 0.417
R2275 SD3L.n214 SD3L.n52 0.281
R2276 SD3L.n186 SD3L.n132 0.281
R2277 SD3L.n213 SD3L.n79 0.155
R2278 SD3L.n185 SD3L.n159 0.155
R2279 SD3L.n186 SD3L.n185 0.13
R2280 SD3L.n214 SD3L.n213 0.13
R2281 SD3L.n214 SD3L.n26 0.103
R2282 SD3L.n186 SD3L.n106 0.103
R2283 SD3L.n212 SD3L.n186 0.091
R2284 SD3L.n213 SD3L.n212 0.039
R2285 SD3L SD3L.n214 0.015
R2286 SD3L.n22 SD3L.n20 0.007
R2287 SD3L.n75 SD3L.n73 0.007
R2288 SD3L.n102 SD3L.n100 0.007
R2289 SD3L.n155 SD3L.n153 0.007
R2290 SD3L.n12 SD3L.n11 0.007
R2291 SD3L.n13 SD3L.n12 0.007
R2292 SD3L.n14 SD3L.n13 0.007
R2293 SD3L.n15 SD3L.n14 0.007
R2294 SD3L.n16 SD3L.n15 0.007
R2295 SD3L.n17 SD3L.n16 0.007
R2296 SD3L.n18 SD3L.n17 0.007
R2297 SD3L.n19 SD3L.n18 0.007
R2298 SD3L.n20 SD3L.n19 0.007
R2299 SD3L.n39 SD3L.n38 0.007
R2300 SD3L.n40 SD3L.n39 0.007
R2301 SD3L.n41 SD3L.n40 0.007
R2302 SD3L.n42 SD3L.n41 0.007
R2303 SD3L.n43 SD3L.n42 0.007
R2304 SD3L.n44 SD3L.n43 0.007
R2305 SD3L.n45 SD3L.n44 0.007
R2306 SD3L.n46 SD3L.n45 0.007
R2307 SD3L.n47 SD3L.n46 0.007
R2308 SD3L.n48 SD3L.n47 0.007
R2309 SD3L.n65 SD3L.n64 0.007
R2310 SD3L.n66 SD3L.n65 0.007
R2311 SD3L.n67 SD3L.n66 0.007
R2312 SD3L.n68 SD3L.n67 0.007
R2313 SD3L.n69 SD3L.n68 0.007
R2314 SD3L.n70 SD3L.n69 0.007
R2315 SD3L.n71 SD3L.n70 0.007
R2316 SD3L.n72 SD3L.n71 0.007
R2317 SD3L.n73 SD3L.n72 0.007
R2318 SD3L.n92 SD3L.n91 0.007
R2319 SD3L.n93 SD3L.n92 0.007
R2320 SD3L.n94 SD3L.n93 0.007
R2321 SD3L.n95 SD3L.n94 0.007
R2322 SD3L.n96 SD3L.n95 0.007
R2323 SD3L.n97 SD3L.n96 0.007
R2324 SD3L.n98 SD3L.n97 0.007
R2325 SD3L.n99 SD3L.n98 0.007
R2326 SD3L.n100 SD3L.n99 0.007
R2327 SD3L.n119 SD3L.n118 0.007
R2328 SD3L.n120 SD3L.n119 0.007
R2329 SD3L.n121 SD3L.n120 0.007
R2330 SD3L.n122 SD3L.n121 0.007
R2331 SD3L.n123 SD3L.n122 0.007
R2332 SD3L.n124 SD3L.n123 0.007
R2333 SD3L.n125 SD3L.n124 0.007
R2334 SD3L.n126 SD3L.n125 0.007
R2335 SD3L.n127 SD3L.n126 0.007
R2336 SD3L.n128 SD3L.n127 0.007
R2337 SD3L.n145 SD3L.n144 0.007
R2338 SD3L.n146 SD3L.n145 0.007
R2339 SD3L.n147 SD3L.n146 0.007
R2340 SD3L.n148 SD3L.n147 0.007
R2341 SD3L.n149 SD3L.n148 0.007
R2342 SD3L.n150 SD3L.n149 0.007
R2343 SD3L.n151 SD3L.n150 0.007
R2344 SD3L.n152 SD3L.n151 0.007
R2345 SD3L.n153 SD3L.n152 0.007
R2346 SD3L.n176 SD3L.n175 0.007
R2347 SD3L.n177 SD3L.n176 0.007
R2348 SD3L.n178 SD3L.n177 0.007
R2349 SD3L.n179 SD3L.n178 0.007
R2350 SD3L.n169 SD3L.n168 0.007
R2351 SD3L.n168 SD3L.n167 0.007
R2352 SD3L.n167 SD3L.n166 0.007
R2353 SD3L.n166 SD3L.n165 0.007
R2354 SD3L.n204 SD3L.n203 0.007
R2355 SD3L.n205 SD3L.n204 0.007
R2356 SD3L.n206 SD3L.n205 0.007
R2357 SD3L.n207 SD3L.n206 0.007
R2358 SD3L.n197 SD3L.n196 0.007
R2359 SD3L.n196 SD3L.n195 0.007
R2360 SD3L.n195 SD3L.n194 0.007
R2361 SD3L.n194 SD3L.n193 0.007
R2362 SD3L.n184 SD3L.n169 0.006
R2363 SD3L.n211 SD3L.n197 0.006
R2364 SD3L.n52 SD3L.n48 0.004
R2365 SD3L.n132 SD3L.n128 0.004
R2366 SD3L.n184 SD3L.n179 0.004
R2367 SD3L.n211 SD3L.n207 0.004
R2368 SD3L.n26 SD3L.n22 0.001
R2369 SD3L.n79 SD3L.n75 0.001
R2370 SD3L.n106 SD3L.n102 0.001
R2371 SD3L.n159 SD3L.n155 0.001
R2372 SD4L.n15 SD4L.t23 1.972
R2373 SD4L.n5 SD4L.t22 1.972
R2374 SD4L.n67 SD4L.t1 1.972
R2375 SD4L.n57 SD4L.t15 1.972
R2376 SD4L.n36 SD4L.n35 1.435
R2377 SD4L.n91 SD4L.n90 1.435
R2378 SD4L.n45 SD4L.n25 1.428
R2379 SD4L.n44 SD4L.n26 1.428
R2380 SD4L.n43 SD4L.n27 1.428
R2381 SD4L.n42 SD4L.n28 1.428
R2382 SD4L.n41 SD4L.n29 1.428
R2383 SD4L.n40 SD4L.n30 1.428
R2384 SD4L.n39 SD4L.n31 1.428
R2385 SD4L.n38 SD4L.n32 1.428
R2386 SD4L.n37 SD4L.n33 1.428
R2387 SD4L.n36 SD4L.n34 1.428
R2388 SD4L.n100 SD4L.n80 1.428
R2389 SD4L.n99 SD4L.n81 1.428
R2390 SD4L.n98 SD4L.n82 1.428
R2391 SD4L.n97 SD4L.n83 1.428
R2392 SD4L.n96 SD4L.n84 1.428
R2393 SD4L.n95 SD4L.n85 1.428
R2394 SD4L.n94 SD4L.n86 1.428
R2395 SD4L.n93 SD4L.n87 1.428
R2396 SD4L.n92 SD4L.n88 1.428
R2397 SD4L.n91 SD4L.n89 1.428
R2398 SD4L.n19 SD4L.n10 1.414
R2399 SD4L.n18 SD4L.n11 1.414
R2400 SD4L.n17 SD4L.n12 1.414
R2401 SD4L.n16 SD4L.n13 1.414
R2402 SD4L.n15 SD4L.n14 1.414
R2403 SD4L.n5 SD4L.n4 1.414
R2404 SD4L.n6 SD4L.n3 1.414
R2405 SD4L.n7 SD4L.n2 1.414
R2406 SD4L.n8 SD4L.n1 1.414
R2407 SD4L.n9 SD4L.n0 1.414
R2408 SD4L.n71 SD4L.n62 1.414
R2409 SD4L.n70 SD4L.n63 1.414
R2410 SD4L.n69 SD4L.n64 1.414
R2411 SD4L.n68 SD4L.n65 1.414
R2412 SD4L.n67 SD4L.n66 1.414
R2413 SD4L.n57 SD4L.n56 1.414
R2414 SD4L.n58 SD4L.n55 1.414
R2415 SD4L.n59 SD4L.n54 1.414
R2416 SD4L.n60 SD4L.n53 1.414
R2417 SD4L.n61 SD4L.n52 1.414
R2418 SD4L.n24 SD4L.n23 1.412
R2419 SD4L.n24 SD4L.n22 1.412
R2420 SD4L.n24 SD4L.n21 1.412
R2421 SD4L.n24 SD4L.n20 1.412
R2422 SD4L.n76 SD4L.n75 1.412
R2423 SD4L.n76 SD4L.n74 1.412
R2424 SD4L.n76 SD4L.n73 1.412
R2425 SD4L.n76 SD4L.n72 1.412
R2426 SD4L.n47 SD4L.n46 1.281
R2427 SD4L.n51 SD4L.n48 1.28
R2428 SD4L.n51 SD4L.n49 1.28
R2429 SD4L.n51 SD4L.n50 1.28
R2430 SD4L.n104 SD4L.n79 1.279
R2431 SD4L.n104 SD4L.n101 1.279
R2432 SD4L.n104 SD4L.n102 1.279
R2433 SD4L.n104 SD4L.n103 1.279
R2434 SD4L.n77 SD4L.n76 0.572
R2435 SD4L.n10 SD4L.t70 0.551
R2436 SD4L.n10 SD4L.t35 0.551
R2437 SD4L.n11 SD4L.t45 0.551
R2438 SD4L.n11 SD4L.t114 0.551
R2439 SD4L.n12 SD4L.t93 0.551
R2440 SD4L.n12 SD4L.t49 0.551
R2441 SD4L.n13 SD4L.t46 0.551
R2442 SD4L.n13 SD4L.t115 0.551
R2443 SD4L.n14 SD4L.t95 0.551
R2444 SD4L.n14 SD4L.t50 0.551
R2445 SD4L.n4 SD4L.t76 0.551
R2446 SD4L.n4 SD4L.t28 0.551
R2447 SD4L.n3 SD4L.t9 0.551
R2448 SD4L.n3 SD4L.t119 0.551
R2449 SD4L.n2 SD4L.t79 0.551
R2450 SD4L.n2 SD4L.t83 0.551
R2451 SD4L.n1 SD4L.t11 0.551
R2452 SD4L.n1 SD4L.t3 0.551
R2453 SD4L.n0 SD4L.t14 0.551
R2454 SD4L.n0 SD4L.t61 0.551
R2455 SD4L.n20 SD4L.t116 0.551
R2456 SD4L.n20 SD4L.t113 0.551
R2457 SD4L.n21 SD4L.t68 0.551
R2458 SD4L.n21 SD4L.t19 0.551
R2459 SD4L.n22 SD4L.t103 0.551
R2460 SD4L.n22 SD4L.t63 0.551
R2461 SD4L.n23 SD4L.t55 0.551
R2462 SD4L.n23 SD4L.t18 0.551
R2463 SD4L.n25 SD4L.t10 0.551
R2464 SD4L.n25 SD4L.t58 0.551
R2465 SD4L.n26 SD4L.t69 0.551
R2466 SD4L.n26 SD4L.t74 0.551
R2467 SD4L.n27 SD4L.t16 0.551
R2468 SD4L.n27 SD4L.t20 0.551
R2469 SD4L.n28 SD4L.t56 0.551
R2470 SD4L.n28 SD4L.t89 0.551
R2471 SD4L.n29 SD4L.t90 0.551
R2472 SD4L.n29 SD4L.t5 0.551
R2473 SD4L.n30 SD4L.t42 0.551
R2474 SD4L.n30 SD4L.t86 0.551
R2475 SD4L.n31 SD4L.t80 0.551
R2476 SD4L.n31 SD4L.t4 0.551
R2477 SD4L.n32 SD4L.t40 0.551
R2478 SD4L.n32 SD4L.t33 0.551
R2479 SD4L.n33 SD4L.t77 0.551
R2480 SD4L.n33 SD4L.t109 0.551
R2481 SD4L.n34 SD4L.t24 0.551
R2482 SD4L.n34 SD4L.t30 0.551
R2483 SD4L.n35 SD4L.t66 0.551
R2484 SD4L.n35 SD4L.t96 0.551
R2485 SD4L.n46 SD4L.t64 0.551
R2486 SD4L.n46 SD4L.t106 0.551
R2487 SD4L.n48 SD4L.t111 0.551
R2488 SD4L.n48 SD4L.t26 0.551
R2489 SD4L.n49 SD4L.t17 0.551
R2490 SD4L.n49 SD4L.t0 0.551
R2491 SD4L.n50 SD4L.t78 0.551
R2492 SD4L.n50 SD4L.t72 0.551
R2493 SD4L.n62 SD4L.t88 0.551
R2494 SD4L.n62 SD4L.t2 0.551
R2495 SD4L.n63 SD4L.t8 0.551
R2496 SD4L.n63 SD4L.t57 0.551
R2497 SD4L.n64 SD4L.t75 0.551
R2498 SD4L.n64 SD4L.t117 0.551
R2499 SD4L.n65 SD4L.t110 0.551
R2500 SD4L.n65 SD4L.t41 0.551
R2501 SD4L.n66 SD4L.t51 0.551
R2502 SD4L.n66 SD4L.t105 0.551
R2503 SD4L.n56 SD4L.t92 0.551
R2504 SD4L.n56 SD4L.t6 0.551
R2505 SD4L.n55 SD4L.t44 0.551
R2506 SD4L.n55 SD4L.t48 0.551
R2507 SD4L.n54 SD4L.t82 0.551
R2508 SD4L.n54 SD4L.t84 0.551
R2509 SD4L.n53 SD4L.t27 0.551
R2510 SD4L.n53 SD4L.t34 0.551
R2511 SD4L.n52 SD4L.t37 0.551
R2512 SD4L.n52 SD4L.t112 0.551
R2513 SD4L.n72 SD4L.t53 0.551
R2514 SD4L.n72 SD4L.t60 0.551
R2515 SD4L.n73 SD4L.t100 0.551
R2516 SD4L.n73 SD4L.t29 0.551
R2517 SD4L.n74 SD4L.t54 0.551
R2518 SD4L.n74 SD4L.t98 0.551
R2519 SD4L.n75 SD4L.t102 0.551
R2520 SD4L.n75 SD4L.t32 0.551
R2521 SD4L.n101 SD4L.t87 0.551
R2522 SD4L.n101 SD4L.t43 0.551
R2523 SD4L.n102 SD4L.t52 0.551
R2524 SD4L.n102 SD4L.t91 0.551
R2525 SD4L.n103 SD4L.t99 0.551
R2526 SD4L.n103 SD4L.t59 0.551
R2527 SD4L.n80 SD4L.t21 0.551
R2528 SD4L.n80 SD4L.t94 0.551
R2529 SD4L.n81 SD4L.t101 0.551
R2530 SD4L.n81 SD4L.t97 0.551
R2531 SD4L.n82 SD4L.t38 0.551
R2532 SD4L.n82 SD4L.t31 0.551
R2533 SD4L.n83 SD4L.t104 0.551
R2534 SD4L.n83 SD4L.t71 0.551
R2535 SD4L.n84 SD4L.t81 0.551
R2536 SD4L.n84 SD4L.t36 0.551
R2537 SD4L.n85 SD4L.t13 0.551
R2538 SD4L.n85 SD4L.t85 0.551
R2539 SD4L.n86 SD4L.t12 0.551
R2540 SD4L.n86 SD4L.t47 0.551
R2541 SD4L.n87 SD4L.t65 0.551
R2542 SD4L.n87 SD4L.t62 0.551
R2543 SD4L.n88 SD4L.t25 0.551
R2544 SD4L.n88 SD4L.t107 0.551
R2545 SD4L.n89 SD4L.t67 0.551
R2546 SD4L.n89 SD4L.t73 0.551
R2547 SD4L.n90 SD4L.t39 0.551
R2548 SD4L.n90 SD4L.t108 0.551
R2549 SD4L.n79 SD4L.t7 0.551
R2550 SD4L.n79 SD4L.t118 0.551
R2551 SD4L.n78 SD4L.n24 0.403
R2552 SD4L.n105 SD4L.n78 0.166
R2553 SD4L.n78 SD4L.n77 0.091
R2554 SD4L.n105 SD4L.n104 0.091
R2555 SD4L.n77 SD4L.n51 0.09
R2556 SD4L SD4L.n105 0.012
R2557 SD4L.n47 SD4L.n45 0.007
R2558 SD4L.n16 SD4L.n15 0.007
R2559 SD4L.n17 SD4L.n16 0.007
R2560 SD4L.n18 SD4L.n17 0.007
R2561 SD4L.n19 SD4L.n18 0.007
R2562 SD4L.n9 SD4L.n8 0.007
R2563 SD4L.n8 SD4L.n7 0.007
R2564 SD4L.n7 SD4L.n6 0.007
R2565 SD4L.n6 SD4L.n5 0.007
R2566 SD4L.n37 SD4L.n36 0.007
R2567 SD4L.n38 SD4L.n37 0.007
R2568 SD4L.n39 SD4L.n38 0.007
R2569 SD4L.n40 SD4L.n39 0.007
R2570 SD4L.n41 SD4L.n40 0.007
R2571 SD4L.n42 SD4L.n41 0.007
R2572 SD4L.n43 SD4L.n42 0.007
R2573 SD4L.n44 SD4L.n43 0.007
R2574 SD4L.n45 SD4L.n44 0.007
R2575 SD4L.n68 SD4L.n67 0.007
R2576 SD4L.n69 SD4L.n68 0.007
R2577 SD4L.n70 SD4L.n69 0.007
R2578 SD4L.n71 SD4L.n70 0.007
R2579 SD4L.n61 SD4L.n60 0.007
R2580 SD4L.n60 SD4L.n59 0.007
R2581 SD4L.n59 SD4L.n58 0.007
R2582 SD4L.n58 SD4L.n57 0.007
R2583 SD4L.n92 SD4L.n91 0.007
R2584 SD4L.n93 SD4L.n92 0.007
R2585 SD4L.n94 SD4L.n93 0.007
R2586 SD4L.n95 SD4L.n94 0.007
R2587 SD4L.n96 SD4L.n95 0.007
R2588 SD4L.n97 SD4L.n96 0.007
R2589 SD4L.n98 SD4L.n97 0.007
R2590 SD4L.n99 SD4L.n98 0.007
R2591 SD4L.n100 SD4L.n99 0.007
R2592 SD4L.n24 SD4L.n9 0.006
R2593 SD4L.n76 SD4L.n61 0.006
R2594 SD4L.n104 SD4L.n100 0.006
R2595 SD4L.n24 SD4L.n19 0.004
R2596 SD4L.n76 SD4L.n71 0.004
R2597 SD4L.n51 SD4L.n47 0.001
C43 SD1R a_n13364_5836# 59.49fF
C44 G12R a_n13364_5836# 99.81fF $ **FLOATING
C45 SD1L a_n13364_5836# 56.70fF
C46 G12L a_n13364_5836# 100.76fF $ **FLOATING
C47 SD2R a_n13364_5836# 103.45fF
C48 G23R a_n13364_5836# 99.81fF $ **FLOATING
C49 SD2L a_n13364_5836# 164.83fF
C50 G23L a_n13364_5836# 100.76fF $ **FLOATING
C51 SD4R a_n13364_5836# 77.75fF
C52 SD3R a_n13364_5836# 103.42fF
C53 G34R a_n13364_5836# 99.81fF $ **FLOATING
C54 SD4L a_n13364_5836# 50.00fF
C55 SD3L a_n13364_5836# 85.71fF
C56 G34L a_n13364_5836# 100.76fF $ **FLOATING
C57 SD4L.n0 a_n13364_5836# 4.21fF
C58 SD4L.n1 a_n13364_5836# 4.21fF
C59 SD4L.n2 a_n13364_5836# 4.21fF
C60 SD4L.n3 a_n13364_5836# 4.21fF
C61 SD4L.n4 a_n13364_5836# 4.21fF
C62 SD4L.t22 a_n13364_5836# 3.82fF $ **FLOATING
C63 SD4L.n5 a_n13364_5836# 11.42fF
C64 SD4L.n6 a_n13364_5836# 5.02fF
C65 SD4L.n7 a_n13364_5836# 5.02fF
C66 SD4L.n8 a_n13364_5836# 5.02fF
C67 SD4L.n9 a_n13364_5836# 4.96fF
C68 SD4L.n10 a_n13364_5836# 4.21fF
C69 SD4L.n11 a_n13364_5836# 4.21fF
C70 SD4L.n12 a_n13364_5836# 4.21fF
C71 SD4L.n13 a_n13364_5836# 4.21fF
C72 SD4L.n14 a_n13364_5836# 4.21fF
C73 SD4L.t23 a_n13364_5836# 3.82fF $ **FLOATING
C74 SD4L.n15 a_n13364_5836# 11.46fF
C75 SD4L.n16 a_n13364_5836# 5.02fF
C76 SD4L.n17 a_n13364_5836# 5.02fF
C77 SD4L.n18 a_n13364_5836# 5.02fF
C78 SD4L.n19 a_n13364_5836# 4.28fF
C79 SD4L.n20 a_n13364_5836# 4.21fF
C80 SD4L.n21 a_n13364_5836# 4.21fF
C81 SD4L.n22 a_n13364_5836# 4.21fF
C82 SD4L.n23 a_n13364_5836# 4.21fF
C83 SD4L.n24 a_n13364_5836# 78.13fF
C84 SD4L.n25 a_n13364_5836# 4.21fF
C85 SD4L.n26 a_n13364_5836# 4.21fF
C86 SD4L.n27 a_n13364_5836# 4.21fF
C87 SD4L.n28 a_n13364_5836# 4.21fF
C88 SD4L.n29 a_n13364_5836# 4.21fF
C89 SD4L.n30 a_n13364_5836# 4.21fF
C90 SD4L.n31 a_n13364_5836# 4.21fF
C91 SD4L.n32 a_n13364_5836# 4.21fF
C92 SD4L.n33 a_n13364_5836# 4.21fF
C93 SD4L.n34 a_n13364_5836# 4.21fF
C94 SD4L.n35 a_n13364_5836# 4.24fF
C95 SD4L.n36 a_n13364_5836# 11.76fF
C96 SD4L.n37 a_n13364_5836# 5.01fF
C97 SD4L.n38 a_n13364_5836# 5.01fF
C98 SD4L.n39 a_n13364_5836# 5.01fF
C99 SD4L.n40 a_n13364_5836# 5.01fF
C100 SD4L.n41 a_n13364_5836# 5.01fF
C101 SD4L.n42 a_n13364_5836# 5.01fF
C102 SD4L.n43 a_n13364_5836# 5.01fF
C103 SD4L.n44 a_n13364_5836# 5.01fF
C104 SD4L.n45 a_n13364_5836# 5.16fF
C105 SD4L.n46 a_n13364_5836# 4.19fF
C106 SD4L.n47 a_n13364_5836# 4.08fF
C107 SD4L.n48 a_n13364_5836# 4.19fF
C108 SD4L.n49 a_n13364_5836# 4.19fF
C109 SD4L.n50 a_n13364_5836# 4.19fF
C110 SD4L.n51 a_n13364_5836# 36.79fF
C111 SD4L.n52 a_n13364_5836# 4.21fF
C112 SD4L.n53 a_n13364_5836# 4.21fF
C113 SD4L.n54 a_n13364_5836# 4.21fF
C114 SD4L.n55 a_n13364_5836# 4.21fF
C115 SD4L.n56 a_n13364_5836# 4.21fF
C116 SD4L.t15 a_n13364_5836# 3.82fF $ **FLOATING
C117 SD4L.n57 a_n13364_5836# 11.72fF
C118 SD4L.n58 a_n13364_5836# 5.02fF
C119 SD4L.n59 a_n13364_5836# 5.02fF
C120 SD4L.n60 a_n13364_5836# 5.02fF
C121 SD4L.n61 a_n13364_5836# 4.96fF
C122 SD4L.n62 a_n13364_5836# 4.21fF
C123 SD4L.n63 a_n13364_5836# 4.21fF
C124 SD4L.n64 a_n13364_5836# 4.21fF
C125 SD4L.n65 a_n13364_5836# 4.21fF
C126 SD4L.n66 a_n13364_5836# 4.21fF
C127 SD4L.t1 a_n13364_5836# 3.82fF $ **FLOATING
C128 SD4L.n67 a_n13364_5836# 13.40fF
C129 SD4L.n68 a_n13364_5836# 5.02fF
C130 SD4L.n69 a_n13364_5836# 5.02fF
C131 SD4L.n70 a_n13364_5836# 5.02fF
C132 SD4L.n71 a_n13364_5836# 4.28fF
C133 SD4L.n72 a_n13364_5836# 4.21fF
C134 SD4L.n73 a_n13364_5836# 4.21fF
C135 SD4L.n74 a_n13364_5836# 4.21fF
C136 SD4L.n75 a_n13364_5836# 4.21fF
C137 SD4L.n76 a_n13364_5836# 104.61fF
C138 SD4L.n77 a_n13364_5836# 124.74fF
C139 SD4L.n78 a_n13364_5836# 99.48fF
C140 SD4L.n79 a_n13364_5836# 4.19fF
C141 SD4L.n80 a_n13364_5836# 4.21fF
C142 SD4L.n81 a_n13364_5836# 4.21fF
C143 SD4L.n82 a_n13364_5836# 4.21fF
C144 SD4L.n83 a_n13364_5836# 4.21fF
C145 SD4L.n84 a_n13364_5836# 4.21fF
C146 SD4L.n85 a_n13364_5836# 4.21fF
C147 SD4L.n86 a_n13364_5836# 4.21fF
C148 SD4L.n87 a_n13364_5836# 4.21fF
C149 SD4L.n88 a_n13364_5836# 4.21fF
C150 SD4L.n89 a_n13364_5836# 4.21fF
C151 SD4L.n90 a_n13364_5836# 4.24fF
C152 SD4L.n91 a_n13364_5836# 11.76fF
C153 SD4L.n92 a_n13364_5836# 5.01fF
C154 SD4L.n93 a_n13364_5836# 5.01fF
C155 SD4L.n94 a_n13364_5836# 5.01fF
C156 SD4L.n95 a_n13364_5836# 5.01fF
C157 SD4L.n96 a_n13364_5836# 5.01fF
C158 SD4L.n97 a_n13364_5836# 5.01fF
C159 SD4L.n98 a_n13364_5836# 5.01fF
C160 SD4L.n99 a_n13364_5836# 5.01fF
C161 SD4L.n100 a_n13364_5836# 4.96fF
C162 SD4L.n101 a_n13364_5836# 4.18fF
C163 SD4L.n102 a_n13364_5836# 4.18fF
C164 SD4L.n103 a_n13364_5836# 4.18fF
C165 SD4L.n104 a_n13364_5836# 41.00fF
C166 SD4L.n105 a_n13364_5836# 51.43fF
C167 SD3L.n0 a_n13364_5836# 4.61fF
C168 SD3L.n1 a_n13364_5836# 4.61fF
C169 SD3L.n2 a_n13364_5836# 4.61fF
C170 SD3L.n3 a_n13364_5836# 4.61fF
C171 SD3L.n4 a_n13364_5836# 4.61fF
C172 SD3L.n5 a_n13364_5836# 4.61fF
C173 SD3L.n6 a_n13364_5836# 4.61fF
C174 SD3L.n7 a_n13364_5836# 4.61fF
C175 SD3L.n8 a_n13364_5836# 4.61fF
C176 SD3L.n9 a_n13364_5836# 4.61fF
C177 SD3L.n10 a_n13364_5836# 4.64fF
C178 SD3L.n11 a_n13364_5836# 12.86fF
C179 SD3L.n12 a_n13364_5836# 5.49fF
C180 SD3L.n13 a_n13364_5836# 5.49fF
C181 SD3L.n14 a_n13364_5836# 5.49fF
C182 SD3L.n15 a_n13364_5836# 5.49fF
C183 SD3L.n16 a_n13364_5836# 5.49fF
C184 SD3L.n17 a_n13364_5836# 5.49fF
C185 SD3L.n18 a_n13364_5836# 5.49fF
C186 SD3L.n19 a_n13364_5836# 5.49fF
C187 SD3L.n20 a_n13364_5836# 5.64fF
C188 SD3L.n21 a_n13364_5836# 4.58fF
C189 SD3L.n22 a_n13364_5836# 4.47fF
C190 SD3L.n23 a_n13364_5836# 4.58fF
C191 SD3L.n24 a_n13364_5836# 4.58fF
C192 SD3L.n25 a_n13364_5836# 4.58fF
C193 SD3L.n26 a_n13364_5836# 41.95fF
C194 SD3L.n27 a_n13364_5836# 4.60fF
C195 SD3L.n28 a_n13364_5836# 4.60fF
C196 SD3L.n29 a_n13364_5836# 4.60fF
C197 SD3L.n30 a_n13364_5836# 4.60fF
C198 SD3L.n31 a_n13364_5836# 4.60fF
C199 SD3L.n32 a_n13364_5836# 4.60fF
C200 SD3L.n33 a_n13364_5836# 4.60fF
C201 SD3L.n34 a_n13364_5836# 4.60fF
C202 SD3L.n35 a_n13364_5836# 4.60fF
C203 SD3L.n36 a_n13364_5836# 4.60fF
C204 SD3L.n37 a_n13364_5836# 4.60fF
C205 SD3L.t105 a_n13364_5836# 4.18fF $ **FLOATING
C206 SD3L.n38 a_n13364_5836# 12.54fF
C207 SD3L.n39 a_n13364_5836# 5.49fF
C208 SD3L.n40 a_n13364_5836# 5.49fF
C209 SD3L.n41 a_n13364_5836# 5.49fF
C210 SD3L.n42 a_n13364_5836# 5.49fF
C211 SD3L.n43 a_n13364_5836# 5.49fF
C212 SD3L.n44 a_n13364_5836# 5.49fF
C213 SD3L.n45 a_n13364_5836# 5.49fF
C214 SD3L.n46 a_n13364_5836# 5.49fF
C215 SD3L.n47 a_n13364_5836# 5.49fF
C216 SD3L.n48 a_n13364_5836# 4.69fF
C217 SD3L.n49 a_n13364_5836# 4.60fF
C218 SD3L.n50 a_n13364_5836# 4.60fF
C219 SD3L.n51 a_n13364_5836# 4.60fF
C220 SD3L.t86 a_n13364_5836# 4.15fF $ **FLOATING
C221 SD3L.n52 a_n13364_5836# 70.96fF
C222 SD3L.n53 a_n13364_5836# 4.61fF
C223 SD3L.n54 a_n13364_5836# 4.61fF
C224 SD3L.n55 a_n13364_5836# 4.61fF
C225 SD3L.n56 a_n13364_5836# 4.61fF
C226 SD3L.n57 a_n13364_5836# 4.61fF
C227 SD3L.n58 a_n13364_5836# 4.61fF
C228 SD3L.n59 a_n13364_5836# 4.61fF
C229 SD3L.n60 a_n13364_5836# 4.61fF
C230 SD3L.n61 a_n13364_5836# 4.61fF
C231 SD3L.n62 a_n13364_5836# 4.61fF
C232 SD3L.n63 a_n13364_5836# 4.64fF
C233 SD3L.n64 a_n13364_5836# 12.86fF
C234 SD3L.n65 a_n13364_5836# 5.49fF
C235 SD3L.n66 a_n13364_5836# 5.49fF
C236 SD3L.n67 a_n13364_5836# 5.49fF
C237 SD3L.n68 a_n13364_5836# 5.49fF
C238 SD3L.n69 a_n13364_5836# 5.49fF
C239 SD3L.n70 a_n13364_5836# 5.49fF
C240 SD3L.n71 a_n13364_5836# 5.49fF
C241 SD3L.n72 a_n13364_5836# 5.49fF
C242 SD3L.n73 a_n13364_5836# 5.64fF
C243 SD3L.n74 a_n13364_5836# 4.58fF
C244 SD3L.n75 a_n13364_5836# 4.47fF
C245 SD3L.n76 a_n13364_5836# 4.58fF
C246 SD3L.n77 a_n13364_5836# 4.58fF
C247 SD3L.n78 a_n13364_5836# 4.58fF
C248 SD3L.n79 a_n13364_5836# 49.16fF
C249 SD3L.n80 a_n13364_5836# 4.61fF
C250 SD3L.n81 a_n13364_5836# 4.61fF
C251 SD3L.n82 a_n13364_5836# 4.61fF
C252 SD3L.n83 a_n13364_5836# 4.61fF
C253 SD3L.n84 a_n13364_5836# 4.61fF
C254 SD3L.n85 a_n13364_5836# 4.61fF
C255 SD3L.n86 a_n13364_5836# 4.61fF
C256 SD3L.n87 a_n13364_5836# 4.61fF
C257 SD3L.n88 a_n13364_5836# 4.61fF
C258 SD3L.n89 a_n13364_5836# 4.61fF
C259 SD3L.n90 a_n13364_5836# 4.64fF
C260 SD3L.n91 a_n13364_5836# 12.86fF
C261 SD3L.n92 a_n13364_5836# 5.49fF
C262 SD3L.n93 a_n13364_5836# 5.49fF
C263 SD3L.n94 a_n13364_5836# 5.49fF
C264 SD3L.n95 a_n13364_5836# 5.49fF
C265 SD3L.n96 a_n13364_5836# 5.49fF
C266 SD3L.n97 a_n13364_5836# 5.49fF
C267 SD3L.n98 a_n13364_5836# 5.49fF
C268 SD3L.n99 a_n13364_5836# 5.49fF
C269 SD3L.n100 a_n13364_5836# 5.64fF
C270 SD3L.n101 a_n13364_5836# 4.58fF
C271 SD3L.n102 a_n13364_5836# 4.47fF
C272 SD3L.n103 a_n13364_5836# 4.58fF
C273 SD3L.n104 a_n13364_5836# 4.58fF
C274 SD3L.n105 a_n13364_5836# 4.58fF
C275 SD3L.n106 a_n13364_5836# 41.95fF
C276 SD3L.n107 a_n13364_5836# 4.60fF
C277 SD3L.n108 a_n13364_5836# 4.60fF
C278 SD3L.n109 a_n13364_5836# 4.60fF
C279 SD3L.n110 a_n13364_5836# 4.60fF
C280 SD3L.n111 a_n13364_5836# 4.60fF
C281 SD3L.n112 a_n13364_5836# 4.60fF
C282 SD3L.n113 a_n13364_5836# 4.60fF
C283 SD3L.n114 a_n13364_5836# 4.60fF
C284 SD3L.n115 a_n13364_5836# 4.60fF
C285 SD3L.n116 a_n13364_5836# 4.60fF
C286 SD3L.n117 a_n13364_5836# 4.60fF
C287 SD3L.t52 a_n13364_5836# 4.18fF $ **FLOATING
C288 SD3L.n118 a_n13364_5836# 12.54fF
C289 SD3L.n119 a_n13364_5836# 5.49fF
C290 SD3L.n120 a_n13364_5836# 5.49fF
C291 SD3L.n121 a_n13364_5836# 5.49fF
C292 SD3L.n122 a_n13364_5836# 5.49fF
C293 SD3L.n123 a_n13364_5836# 5.49fF
C294 SD3L.n124 a_n13364_5836# 5.49fF
C295 SD3L.n125 a_n13364_5836# 5.49fF
C296 SD3L.n126 a_n13364_5836# 5.49fF
C297 SD3L.n127 a_n13364_5836# 5.49fF
C298 SD3L.n128 a_n13364_5836# 4.69fF
C299 SD3L.n129 a_n13364_5836# 4.60fF
C300 SD3L.n130 a_n13364_5836# 4.60fF
C301 SD3L.n131 a_n13364_5836# 4.60fF
C302 SD3L.t6 a_n13364_5836# 4.15fF $ **FLOATING
C303 SD3L.n132 a_n13364_5836# 70.96fF
C304 SD3L.n133 a_n13364_5836# 4.61fF
C305 SD3L.n134 a_n13364_5836# 4.61fF
C306 SD3L.n135 a_n13364_5836# 4.61fF
C307 SD3L.n136 a_n13364_5836# 4.61fF
C308 SD3L.n137 a_n13364_5836# 4.61fF
C309 SD3L.n138 a_n13364_5836# 4.61fF
C310 SD3L.n139 a_n13364_5836# 4.61fF
C311 SD3L.n140 a_n13364_5836# 4.61fF
C312 SD3L.n141 a_n13364_5836# 4.61fF
C313 SD3L.n142 a_n13364_5836# 4.61fF
C314 SD3L.n143 a_n13364_5836# 4.64fF
C315 SD3L.n144 a_n13364_5836# 12.86fF
C316 SD3L.n145 a_n13364_5836# 5.49fF
C317 SD3L.n146 a_n13364_5836# 5.49fF
C318 SD3L.n147 a_n13364_5836# 5.49fF
C319 SD3L.n148 a_n13364_5836# 5.49fF
C320 SD3L.n149 a_n13364_5836# 5.49fF
C321 SD3L.n150 a_n13364_5836# 5.49fF
C322 SD3L.n151 a_n13364_5836# 5.49fF
C323 SD3L.n152 a_n13364_5836# 5.49fF
C324 SD3L.n153 a_n13364_5836# 5.64fF
C325 SD3L.n154 a_n13364_5836# 4.58fF
C326 SD3L.n155 a_n13364_5836# 4.47fF
C327 SD3L.n156 a_n13364_5836# 4.58fF
C328 SD3L.n157 a_n13364_5836# 4.58fF
C329 SD3L.n158 a_n13364_5836# 4.58fF
C330 SD3L.n159 a_n13364_5836# 49.16fF
C331 SD3L.n160 a_n13364_5836# 4.60fF
C332 SD3L.n161 a_n13364_5836# 4.60fF
C333 SD3L.n162 a_n13364_5836# 4.60fF
C334 SD3L.n163 a_n13364_5836# 4.60fF
C335 SD3L.n164 a_n13364_5836# 4.60fF
C336 SD3L.t143 a_n13364_5836# 4.18fF $ **FLOATING
C337 SD3L.n165 a_n13364_5836# 12.83fF
C338 SD3L.n166 a_n13364_5836# 5.49fF
C339 SD3L.n167 a_n13364_5836# 5.49fF
C340 SD3L.n168 a_n13364_5836# 5.49fF
C341 SD3L.n169 a_n13364_5836# 5.43fF
C342 SD3L.n170 a_n13364_5836# 4.60fF
C343 SD3L.n171 a_n13364_5836# 4.60fF
C344 SD3L.n172 a_n13364_5836# 4.60fF
C345 SD3L.n173 a_n13364_5836# 4.60fF
C346 SD3L.n174 a_n13364_5836# 4.60fF
C347 SD3L.t132 a_n13364_5836# 4.18fF $ **FLOATING
C348 SD3L.n175 a_n13364_5836# 14.66fF
C349 SD3L.n176 a_n13364_5836# 5.49fF
C350 SD3L.n177 a_n13364_5836# 5.49fF
C351 SD3L.n178 a_n13364_5836# 5.49fF
C352 SD3L.n179 a_n13364_5836# 4.68fF
C353 SD3L.n180 a_n13364_5836# 4.60fF
C354 SD3L.n181 a_n13364_5836# 4.60fF
C355 SD3L.n182 a_n13364_5836# 4.60fF
C356 SD3L.n183 a_n13364_5836# 4.60fF
C357 SD3L.n184 a_n13364_5836# 94.87fF
C358 SD3L.n185 a_n13364_5836# 141.09fF
C359 SD3L.n186 a_n13364_5836# 93.43fF
C360 SD3L.n187 a_n13364_5836# 4.60fF
C361 SD3L.n188 a_n13364_5836# 4.60fF
C362 SD3L.n189 a_n13364_5836# 4.60fF
C363 SD3L.n190 a_n13364_5836# 4.60fF
C364 SD3L.n191 a_n13364_5836# 4.60fF
C365 SD3L.n192 a_n13364_5836# 4.60fF
C366 SD3L.t153 a_n13364_5836# 4.18fF $ **FLOATING
C367 SD3L.n193 a_n13364_5836# 12.49fF
C368 SD3L.n194 a_n13364_5836# 5.49fF
C369 SD3L.n195 a_n13364_5836# 5.49fF
C370 SD3L.n196 a_n13364_5836# 5.49fF
C371 SD3L.n197 a_n13364_5836# 5.43fF
C372 SD3L.n198 a_n13364_5836# 4.60fF
C373 SD3L.n199 a_n13364_5836# 4.60fF
C374 SD3L.n200 a_n13364_5836# 4.60fF
C375 SD3L.n201 a_n13364_5836# 4.60fF
C376 SD3L.n202 a_n13364_5836# 4.60fF
C377 SD3L.t154 a_n13364_5836# 4.18fF $ **FLOATING
C378 SD3L.n203 a_n13364_5836# 12.54fF
C379 SD3L.n204 a_n13364_5836# 5.49fF
C380 SD3L.n205 a_n13364_5836# 5.49fF
C381 SD3L.n206 a_n13364_5836# 5.49fF
C382 SD3L.n207 a_n13364_5836# 4.68fF
C383 SD3L.n208 a_n13364_5836# 4.60fF
C384 SD3L.n209 a_n13364_5836# 4.60fF
C385 SD3L.n210 a_n13364_5836# 4.60fF
C386 SD3L.n211 a_n13364_5836# 87.05fF
C387 SD3L.n212 a_n13364_5836# 86.47fF
C388 SD3L.n213 a_n13364_5836# 58.90fF
C389 SD3L.n214 a_n13364_5836# 79.13fF
C390 SD1R.n0 a_n13364_5836# 4.22fF
C391 SD1R.n1 a_n13364_5836# 4.22fF
C392 SD1R.n2 a_n13364_5836# 4.22fF
C393 SD1R.n3 a_n13364_5836# 4.22fF
C394 SD1R.n4 a_n13364_5836# 4.22fF
C395 SD1R.n5 a_n13364_5836# 4.22fF
C396 SD1R.n6 a_n13364_5836# 4.22fF
C397 SD1R.n7 a_n13364_5836# 4.22fF
C398 SD1R.n8 a_n13364_5836# 4.22fF
C399 SD1R.n9 a_n13364_5836# 4.22fF
C400 SD1R.n10 a_n13364_5836# 4.22fF
C401 SD1R.t63 a_n13364_5836# 3.82fF $ **FLOATING
C402 SD1R.n11 a_n13364_5836# 11.44fF
C403 SD1R.n12 a_n13364_5836# 5.03fF
C404 SD1R.n13 a_n13364_5836# 5.03fF
C405 SD1R.n14 a_n13364_5836# 5.03fF
C406 SD1R.n15 a_n13364_5836# 5.03fF
C407 SD1R.n16 a_n13364_5836# 5.03fF
C408 SD1R.n17 a_n13364_5836# 5.03fF
C409 SD1R.n18 a_n13364_5836# 5.03fF
C410 SD1R.n19 a_n13364_5836# 5.03fF
C411 SD1R.n20 a_n13364_5836# 5.03fF
C412 SD1R.n21 a_n13364_5836# 4.98fF
C413 SD1R.t50 a_n13364_5836# 3.80fF $ **FLOATING
C414 SD1R.n22 a_n13364_5836# 4.22fF
C415 SD1R.n23 a_n13364_5836# 4.22fF
C416 SD1R.n24 a_n13364_5836# 4.22fF
C417 SD1R.n25 a_n13364_5836# 69.07fF
C418 SD1R.n26 a_n13364_5836# 4.22fF
C419 SD1R.n27 a_n13364_5836# 4.22fF
C420 SD1R.n28 a_n13364_5836# 4.22fF
C421 SD1R.n29 a_n13364_5836# 4.22fF
C422 SD1R.n30 a_n13364_5836# 4.22fF
C423 SD1R.n31 a_n13364_5836# 4.25fF
C424 SD1R.n32 a_n13364_5836# 11.74fF
C425 SD1R.n33 a_n13364_5836# 5.02fF
C426 SD1R.n34 a_n13364_5836# 5.02fF
C427 SD1R.n35 a_n13364_5836# 5.02fF
C428 SD1R.n36 a_n13364_5836# 4.29fF
C429 SD1R.n37 a_n13364_5836# 4.22fF
C430 SD1R.n38 a_n13364_5836# 4.22fF
C431 SD1R.n39 a_n13364_5836# 4.22fF
C432 SD1R.n40 a_n13364_5836# 4.22fF
C433 SD1R.n41 a_n13364_5836# 4.25fF
C434 SD1R.n42 a_n13364_5836# 11.78fF
C435 SD1R.n43 a_n13364_5836# 5.02fF
C436 SD1R.n44 a_n13364_5836# 5.02fF
C437 SD1R.n45 a_n13364_5836# 4.69fF
C438 SD1R.n46 a_n13364_5836# 4.20fF
C439 SD1R.n47 a_n13364_5836# 4.20fF
C440 SD1R.n48 a_n13364_5836# 4.20fF
C441 SD1R.n49 a_n13364_5836# 4.20fF
C442 SD1R.n50 a_n13364_5836# 51.38fF
C443 SD1R.n51 a_n13364_5836# 4.22fF
C444 SD1R.n52 a_n13364_5836# 4.22fF
C445 SD1R.n53 a_n13364_5836# 4.22fF
C446 SD1R.n54 a_n13364_5836# 4.22fF
C447 SD1R.n55 a_n13364_5836# 4.22fF
C448 SD1R.n56 a_n13364_5836# 4.22fF
C449 SD1R.n57 a_n13364_5836# 4.22fF
C450 SD1R.n58 a_n13364_5836# 4.22fF
C451 SD1R.n59 a_n13364_5836# 4.22fF
C452 SD1R.n60 a_n13364_5836# 4.22fF
C453 SD1R.n61 a_n13364_5836# 4.22fF
C454 SD1R.t69 a_n13364_5836# 3.83fF $ **FLOATING
C455 SD1R.n62 a_n13364_5836# 11.44fF
C456 SD1R.n63 a_n13364_5836# 5.03fF
C457 SD1R.n64 a_n13364_5836# 5.03fF
C458 SD1R.n65 a_n13364_5836# 5.03fF
C459 SD1R.n66 a_n13364_5836# 5.03fF
C460 SD1R.n67 a_n13364_5836# 5.03fF
C461 SD1R.n68 a_n13364_5836# 5.03fF
C462 SD1R.n69 a_n13364_5836# 5.03fF
C463 SD1R.n70 a_n13364_5836# 5.03fF
C464 SD1R.n71 a_n13364_5836# 5.03fF
C465 SD1R.n72 a_n13364_5836# 5.18fF
C466 SD1R.n73 a_n13364_5836# 4.22fF
C467 SD1R.n74 a_n13364_5836# 4.06fF
C468 SD1R.n75 a_n13364_5836# 4.21fF
C469 SD1R.n76 a_n13364_5836# 4.21fF
C470 SD1R.t70 a_n13364_5836# 3.80fF $ **FLOATING
C471 SD1R.n77 a_n13364_5836# 64.81fF
C472 SD1R.n78 a_n13364_5836# 4.20fF
C473 SD1R.n79 a_n13364_5836# 4.20fF
C474 SD1R.n80 a_n13364_5836# 4.20fF
C475 SD1R.n81 a_n13364_5836# 4.20fF
C476 SD1R.n82 a_n13364_5836# 4.22fF
C477 SD1R.n83 a_n13364_5836# 4.22fF
C478 SD1R.n84 a_n13364_5836# 4.22fF
C479 SD1R.n85 a_n13364_5836# 4.25fF
C480 SD1R.n86 a_n13364_5836# 11.78fF
C481 SD1R.n87 a_n13364_5836# 4.22fF
C482 SD1R.n88 a_n13364_5836# 5.02fF
C483 SD1R.n89 a_n13364_5836# 5.02fF
C484 SD1R.n90 a_n13364_5836# 4.69fF
C485 SD1R.n91 a_n13364_5836# 4.22fF
C486 SD1R.n92 a_n13364_5836# 4.22fF
C487 SD1R.n93 a_n13364_5836# 4.22fF
C488 SD1R.n94 a_n13364_5836# 4.22fF
C489 SD1R.n95 a_n13364_5836# 4.22fF
C490 SD1R.n96 a_n13364_5836# 4.25fF
C491 SD1R.n97 a_n13364_5836# 11.74fF
C492 SD1R.n98 a_n13364_5836# 5.02fF
C493 SD1R.n99 a_n13364_5836# 5.02fF
C494 SD1R.n100 a_n13364_5836# 5.02fF
C495 SD1R.n101 a_n13364_5836# 4.29fF
C496 SD1R.n102 a_n13364_5836# 81.61fF
C497 SD1R.n103 a_n13364_5836# 120.41fF
C498 SD1R.n104 a_n13364_5836# 70.14fF
C499 SD1R.n105 a_n13364_5836# 79.35fF
C500 SD2R.n0 a_n13364_5836# 4.55fF
C501 SD2R.n1 a_n13364_5836# 4.55fF
C502 SD2R.n2 a_n13364_5836# 4.55fF
C503 SD2R.n3 a_n13364_5836# 4.55fF
C504 SD2R.n4 a_n13364_5836# 4.55fF
C505 SD2R.n5 a_n13364_5836# 4.55fF
C506 SD2R.n6 a_n13364_5836# 4.55fF
C507 SD2R.n7 a_n13364_5836# 4.55fF
C508 SD2R.n8 a_n13364_5836# 4.55fF
C509 SD2R.n9 a_n13364_5836# 4.55fF
C510 SD2R.n10 a_n13364_5836# 4.55fF
C511 SD2R.t237 a_n13364_5836# 4.13fF $ **FLOATING
C512 SD2R.n11 a_n13364_5836# 12.35fF
C513 SD2R.n12 a_n13364_5836# 5.43fF
C514 SD2R.n13 a_n13364_5836# 5.43fF
C515 SD2R.n14 a_n13364_5836# 5.43fF
C516 SD2R.n15 a_n13364_5836# 5.43fF
C517 SD2R.n16 a_n13364_5836# 5.43fF
C518 SD2R.n17 a_n13364_5836# 5.43fF
C519 SD2R.n18 a_n13364_5836# 5.43fF
C520 SD2R.n19 a_n13364_5836# 5.43fF
C521 SD2R.n20 a_n13364_5836# 5.43fF
C522 SD2R.n21 a_n13364_5836# 5.37fF
C523 SD2R.t148 a_n13364_5836# 4.10fF $ **FLOATING
C524 SD2R.n22 a_n13364_5836# 4.55fF
C525 SD2R.n23 a_n13364_5836# 4.55fF
C526 SD2R.n24 a_n13364_5836# 4.55fF
C527 SD2R.n25 a_n13364_5836# 79.87fF
C528 SD2R.n26 a_n13364_5836# 4.55fF
C529 SD2R.n27 a_n13364_5836# 4.55fF
C530 SD2R.n28 a_n13364_5836# 4.55fF
C531 SD2R.n29 a_n13364_5836# 4.55fF
C532 SD2R.n30 a_n13364_5836# 4.55fF
C533 SD2R.n31 a_n13364_5836# 4.55fF
C534 SD2R.n32 a_n13364_5836# 4.55fF
C535 SD2R.n33 a_n13364_5836# 4.55fF
C536 SD2R.n34 a_n13364_5836# 4.55fF
C537 SD2R.n35 a_n13364_5836# 4.55fF
C538 SD2R.n36 a_n13364_5836# 4.59fF
C539 SD2R.n37 a_n13364_5836# 12.71fF
C540 SD2R.n38 a_n13364_5836# 5.42fF
C541 SD2R.n39 a_n13364_5836# 5.42fF
C542 SD2R.n40 a_n13364_5836# 5.42fF
C543 SD2R.n41 a_n13364_5836# 5.42fF
C544 SD2R.n42 a_n13364_5836# 5.42fF
C545 SD2R.n43 a_n13364_5836# 5.42fF
C546 SD2R.n44 a_n13364_5836# 5.42fF
C547 SD2R.n45 a_n13364_5836# 5.42fF
C548 SD2R.n46 a_n13364_5836# 5.34fF
C549 SD2R.n47 a_n13364_5836# 4.53fF
C550 SD2R.n48 a_n13364_5836# 4.91fF
C551 SD2R.n49 a_n13364_5836# 4.53fF
C552 SD2R.n50 a_n13364_5836# 4.53fF
C553 SD2R.n51 a_n13364_5836# 4.53fF
C554 SD2R.n52 a_n13364_5836# 4.55fF
C555 SD2R.n53 a_n13364_5836# 4.55fF
C556 SD2R.n54 a_n13364_5836# 4.55fF
C557 SD2R.n55 a_n13364_5836# 4.55fF
C558 SD2R.n56 a_n13364_5836# 4.55fF
C559 SD2R.n57 a_n13364_5836# 4.55fF
C560 SD2R.n58 a_n13364_5836# 4.55fF
C561 SD2R.n59 a_n13364_5836# 4.55fF
C562 SD2R.n60 a_n13364_5836# 4.55fF
C563 SD2R.n61 a_n13364_5836# 4.55fF
C564 SD2R.n62 a_n13364_5836# 4.55fF
C565 SD2R.t57 a_n13364_5836# 4.13fF $ **FLOATING
C566 SD2R.n63 a_n13364_5836# 12.35fF
C567 SD2R.n64 a_n13364_5836# 5.43fF
C568 SD2R.n65 a_n13364_5836# 5.43fF
C569 SD2R.n66 a_n13364_5836# 5.43fF
C570 SD2R.n67 a_n13364_5836# 5.43fF
C571 SD2R.n68 a_n13364_5836# 5.43fF
C572 SD2R.n69 a_n13364_5836# 5.43fF
C573 SD2R.n70 a_n13364_5836# 5.43fF
C574 SD2R.n71 a_n13364_5836# 5.43fF
C575 SD2R.n72 a_n13364_5836# 5.43fF
C576 SD2R.n73 a_n13364_5836# 5.59fF
C577 SD2R.n74 a_n13364_5836# 4.55fF
C578 SD2R.n75 a_n13364_5836# 4.38fF
C579 SD2R.n76 a_n13364_5836# 4.55fF
C580 SD2R.n77 a_n13364_5836# 4.55fF
C581 SD2R.t58 a_n13364_5836# 4.10fF $ **FLOATING
C582 SD2R.n78 a_n13364_5836# 75.74fF
C583 SD2R.n79 a_n13364_5836# 4.55fF
C584 SD2R.n80 a_n13364_5836# 4.55fF
C585 SD2R.n81 a_n13364_5836# 4.55fF
C586 SD2R.n82 a_n13364_5836# 4.55fF
C587 SD2R.n83 a_n13364_5836# 4.55fF
C588 SD2R.n84 a_n13364_5836# 4.59fF
C589 SD2R.n85 a_n13364_5836# 12.67fF
C590 SD2R.n86 a_n13364_5836# 5.42fF
C591 SD2R.n87 a_n13364_5836# 5.42fF
C592 SD2R.n88 a_n13364_5836# 5.42fF
C593 SD2R.n89 a_n13364_5836# 4.63fF
C594 SD2R.n90 a_n13364_5836# 4.55fF
C595 SD2R.n91 a_n13364_5836# 4.55fF
C596 SD2R.n92 a_n13364_5836# 4.55fF
C597 SD2R.n93 a_n13364_5836# 4.55fF
C598 SD2R.n94 a_n13364_5836# 4.59fF
C599 SD2R.n95 a_n13364_5836# 12.71fF
C600 SD2R.n96 a_n13364_5836# 5.42fF
C601 SD2R.n97 a_n13364_5836# 5.42fF
C602 SD2R.n98 a_n13364_5836# 5.06fF
C603 SD2R.n99 a_n13364_5836# 4.53fF
C604 SD2R.n100 a_n13364_5836# 4.53fF
C605 SD2R.n101 a_n13364_5836# 4.53fF
C606 SD2R.n102 a_n13364_5836# 4.53fF
C607 SD2R.n103 a_n13364_5836# 61.26fF
C608 SD2R.n104 a_n13364_5836# 4.55fF
C609 SD2R.n105 a_n13364_5836# 4.55fF
C610 SD2R.n106 a_n13364_5836# 4.55fF
C611 SD2R.n107 a_n13364_5836# 4.55fF
C612 SD2R.n108 a_n13364_5836# 4.55fF
C613 SD2R.n109 a_n13364_5836# 4.55fF
C614 SD2R.n110 a_n13364_5836# 4.55fF
C615 SD2R.n111 a_n13364_5836# 4.55fF
C616 SD2R.n112 a_n13364_5836# 4.55fF
C617 SD2R.n113 a_n13364_5836# 4.55fF
C618 SD2R.n114 a_n13364_5836# 4.55fF
C619 SD2R.t146 a_n13364_5836# 4.13fF $ **FLOATING
C620 SD2R.n115 a_n13364_5836# 12.35fF
C621 SD2R.n116 a_n13364_5836# 5.43fF
C622 SD2R.n117 a_n13364_5836# 5.43fF
C623 SD2R.n118 a_n13364_5836# 5.43fF
C624 SD2R.n119 a_n13364_5836# 5.43fF
C625 SD2R.n120 a_n13364_5836# 5.43fF
C626 SD2R.n121 a_n13364_5836# 5.43fF
C627 SD2R.n122 a_n13364_5836# 5.43fF
C628 SD2R.n123 a_n13364_5836# 5.43fF
C629 SD2R.n124 a_n13364_5836# 5.43fF
C630 SD2R.n125 a_n13364_5836# 5.37fF
C631 SD2R.t140 a_n13364_5836# 4.10fF $ **FLOATING
C632 SD2R.n126 a_n13364_5836# 4.55fF
C633 SD2R.n127 a_n13364_5836# 4.55fF
C634 SD2R.n128 a_n13364_5836# 4.55fF
C635 SD2R.n129 a_n13364_5836# 79.87fF
C636 SD2R.n130 a_n13364_5836# 4.55fF
C637 SD2R.n131 a_n13364_5836# 4.55fF
C638 SD2R.n132 a_n13364_5836# 4.55fF
C639 SD2R.n133 a_n13364_5836# 4.55fF
C640 SD2R.n134 a_n13364_5836# 4.55fF
C641 SD2R.n135 a_n13364_5836# 4.55fF
C642 SD2R.n136 a_n13364_5836# 4.55fF
C643 SD2R.n137 a_n13364_5836# 4.55fF
C644 SD2R.n138 a_n13364_5836# 4.55fF
C645 SD2R.n139 a_n13364_5836# 4.55fF
C646 SD2R.n140 a_n13364_5836# 4.59fF
C647 SD2R.n141 a_n13364_5836# 12.71fF
C648 SD2R.n142 a_n13364_5836# 5.42fF
C649 SD2R.n143 a_n13364_5836# 5.42fF
C650 SD2R.n144 a_n13364_5836# 5.42fF
C651 SD2R.n145 a_n13364_5836# 5.42fF
C652 SD2R.n146 a_n13364_5836# 5.42fF
C653 SD2R.n147 a_n13364_5836# 5.42fF
C654 SD2R.n148 a_n13364_5836# 5.42fF
C655 SD2R.n149 a_n13364_5836# 5.42fF
C656 SD2R.n150 a_n13364_5836# 5.34fF
C657 SD2R.n151 a_n13364_5836# 4.53fF
C658 SD2R.n152 a_n13364_5836# 4.91fF
C659 SD2R.n153 a_n13364_5836# 4.53fF
C660 SD2R.n154 a_n13364_5836# 4.53fF
C661 SD2R.n155 a_n13364_5836# 4.53fF
C662 SD2R.n156 a_n13364_5836# 4.55fF
C663 SD2R.n157 a_n13364_5836# 4.55fF
C664 SD2R.n158 a_n13364_5836# 4.55fF
C665 SD2R.n159 a_n13364_5836# 4.55fF
C666 SD2R.n160 a_n13364_5836# 4.55fF
C667 SD2R.n161 a_n13364_5836# 4.55fF
C668 SD2R.n162 a_n13364_5836# 4.55fF
C669 SD2R.n163 a_n13364_5836# 4.55fF
C670 SD2R.n164 a_n13364_5836# 4.55fF
C671 SD2R.n165 a_n13364_5836# 4.55fF
C672 SD2R.n166 a_n13364_5836# 4.55fF
C673 SD2R.t50 a_n13364_5836# 4.13fF $ **FLOATING
C674 SD2R.n167 a_n13364_5836# 12.35fF
C675 SD2R.n168 a_n13364_5836# 5.43fF
C676 SD2R.n169 a_n13364_5836# 5.43fF
C677 SD2R.n170 a_n13364_5836# 5.43fF
C678 SD2R.n171 a_n13364_5836# 5.43fF
C679 SD2R.n172 a_n13364_5836# 5.43fF
C680 SD2R.n173 a_n13364_5836# 5.43fF
C681 SD2R.n174 a_n13364_5836# 5.43fF
C682 SD2R.n175 a_n13364_5836# 5.43fF
C683 SD2R.n176 a_n13364_5836# 5.43fF
C684 SD2R.n177 a_n13364_5836# 5.37fF
C685 SD2R.t36 a_n13364_5836# 4.10fF $ **FLOATING
C686 SD2R.n178 a_n13364_5836# 4.55fF
C687 SD2R.n179 a_n13364_5836# 4.55fF
C688 SD2R.n180 a_n13364_5836# 4.55fF
C689 SD2R.n181 a_n13364_5836# 94.03fF
C690 SD2R.n182 a_n13364_5836# 126.04fF
C691 SD2R.n183 a_n13364_5836# 68.68fF
C692 SD2R.n184 a_n13364_5836# 59.99fF
C693 SD2R.n185 a_n13364_5836# 84.54fF
C694 SD2R.n186 a_n13364_5836# 66.41fF
C695 SD2R.n187 a_n13364_5836# 68.68fF
C696 SD2R.n188 a_n13364_5836# 4.55fF
C697 SD2R.n189 a_n13364_5836# 4.55fF
C698 SD2R.n190 a_n13364_5836# 4.55fF
C699 SD2R.n191 a_n13364_5836# 4.55fF
C700 SD2R.n192 a_n13364_5836# 4.59fF
C701 SD2R.n193 a_n13364_5836# 12.71fF
C702 SD2R.n194 a_n13364_5836# 5.42fF
C703 SD2R.n195 a_n13364_5836# 5.42fF
C704 SD2R.n196 a_n13364_5836# 5.06fF
C705 SD2R.n197 a_n13364_5836# 4.53fF
C706 SD2R.n198 a_n13364_5836# 4.53fF
C707 SD2R.n199 a_n13364_5836# 4.53fF
C708 SD2R.n200 a_n13364_5836# 4.55fF
C709 SD2R.n201 a_n13364_5836# 4.55fF
C710 SD2R.n202 a_n13364_5836# 4.55fF
C711 SD2R.n203 a_n13364_5836# 4.55fF
C712 SD2R.n204 a_n13364_5836# 4.55fF
C713 SD2R.n205 a_n13364_5836# 4.59fF
C714 SD2R.n206 a_n13364_5836# 12.67fF
C715 SD2R.n207 a_n13364_5836# 5.42fF
C716 SD2R.n208 a_n13364_5836# 5.42fF
C717 SD2R.n209 a_n13364_5836# 5.42fF
C718 SD2R.n210 a_n13364_5836# 4.63fF
C719 SD2R.n211 a_n13364_5836# 4.53fF
C720 SD2R.n212 a_n13364_5836# 61.26fF
C721 SD2R.n213 a_n13364_5836# 53.21fF
C722 SD1L.n0 a_n13364_5836# 4.45fF
C723 SD1L.n1 a_n13364_5836# 4.45fF
C724 SD1L.n2 a_n13364_5836# 4.45fF
C725 SD1L.n3 a_n13364_5836# 4.45fF
C726 SD1L.n4 a_n13364_5836# 4.45fF
C727 SD1L.n5 a_n13364_5836# 4.45fF
C728 SD1L.n6 a_n13364_5836# 4.45fF
C729 SD1L.n7 a_n13364_5836# 4.45fF
C730 SD1L.n8 a_n13364_5836# 4.45fF
C731 SD1L.n9 a_n13364_5836# 4.45fF
C732 SD1L.n10 a_n13364_5836# 4.45fF
C733 SD1L.t116 a_n13364_5836# 4.04fF $ **FLOATING
C734 SD1L.n11 a_n13364_5836# 12.12fF
C735 SD1L.n12 a_n13364_5836# 5.31fF
C736 SD1L.n13 a_n13364_5836# 5.31fF
C737 SD1L.n14 a_n13364_5836# 5.31fF
C738 SD1L.n15 a_n13364_5836# 5.31fF
C739 SD1L.n16 a_n13364_5836# 5.31fF
C740 SD1L.n17 a_n13364_5836# 5.31fF
C741 SD1L.n18 a_n13364_5836# 5.31fF
C742 SD1L.n19 a_n13364_5836# 5.31fF
C743 SD1L.n20 a_n13364_5836# 5.31fF
C744 SD1L.n21 a_n13364_5836# 4.53fF
C745 SD1L.n22 a_n13364_5836# 4.45fF
C746 SD1L.n23 a_n13364_5836# 4.45fF
C747 SD1L.n24 a_n13364_5836# 4.45fF
C748 SD1L.t80 a_n13364_5836# 4.01fF $ **FLOATING
C749 SD1L.n25 a_n13364_5836# 64.52fF
C750 SD1L.n26 a_n13364_5836# 4.45fF
C751 SD1L.n27 a_n13364_5836# 4.45fF
C752 SD1L.n28 a_n13364_5836# 4.45fF
C753 SD1L.n29 a_n13364_5836# 4.45fF
C754 SD1L.n30 a_n13364_5836# 4.45fF
C755 SD1L.n31 a_n13364_5836# 4.45fF
C756 SD1L.n32 a_n13364_5836# 4.45fF
C757 SD1L.n33 a_n13364_5836# 4.45fF
C758 SD1L.n34 a_n13364_5836# 4.45fF
C759 SD1L.n35 a_n13364_5836# 4.45fF
C760 SD1L.n36 a_n13364_5836# 4.49fF
C761 SD1L.n37 a_n13364_5836# 12.43fF
C762 SD1L.n38 a_n13364_5836# 5.30fF
C763 SD1L.n39 a_n13364_5836# 5.30fF
C764 SD1L.n40 a_n13364_5836# 5.30fF
C765 SD1L.n41 a_n13364_5836# 5.30fF
C766 SD1L.n42 a_n13364_5836# 5.30fF
C767 SD1L.n43 a_n13364_5836# 5.30fF
C768 SD1L.n44 a_n13364_5836# 5.30fF
C769 SD1L.n45 a_n13364_5836# 5.30fF
C770 SD1L.n46 a_n13364_5836# 5.45fF
C771 SD1L.n47 a_n13364_5836# 4.43fF
C772 SD1L.n48 a_n13364_5836# 4.32fF
C773 SD1L.n49 a_n13364_5836# 4.43fF
C774 SD1L.n50 a_n13364_5836# 4.43fF
C775 SD1L.n51 a_n13364_5836# 4.43fF
C776 SD1L.n52 a_n13364_5836# 43.45fF
C777 SD1L.n53 a_n13364_5836# 4.45fF
C778 SD1L.n54 a_n13364_5836# 4.45fF
C779 SD1L.n55 a_n13364_5836# 4.45fF
C780 SD1L.n56 a_n13364_5836# 4.45fF
C781 SD1L.n57 a_n13364_5836# 4.45fF
C782 SD1L.n58 a_n13364_5836# 4.45fF
C783 SD1L.n59 a_n13364_5836# 4.45fF
C784 SD1L.n60 a_n13364_5836# 4.45fF
C785 SD1L.n61 a_n13364_5836# 4.45fF
C786 SD1L.n62 a_n13364_5836# 4.45fF
C787 SD1L.n63 a_n13364_5836# 4.49fF
C788 SD1L.n64 a_n13364_5836# 12.43fF
C789 SD1L.n65 a_n13364_5836# 5.30fF
C790 SD1L.n66 a_n13364_5836# 5.30fF
C791 SD1L.n67 a_n13364_5836# 5.30fF
C792 SD1L.n68 a_n13364_5836# 5.30fF
C793 SD1L.n69 a_n13364_5836# 5.30fF
C794 SD1L.n70 a_n13364_5836# 5.30fF
C795 SD1L.n71 a_n13364_5836# 5.30fF
C796 SD1L.n72 a_n13364_5836# 5.30fF
C797 SD1L.n73 a_n13364_5836# 5.45fF
C798 SD1L.n74 a_n13364_5836# 4.43fF
C799 SD1L.n75 a_n13364_5836# 4.32fF
C800 SD1L.n76 a_n13364_5836# 4.43fF
C801 SD1L.n77 a_n13364_5836# 4.43fF
C802 SD1L.n78 a_n13364_5836# 4.43fF
C803 SD1L.n79 a_n13364_5836# 69.73fF
C804 SD1L.t33 a_n13364_5836# 4.01fF $ **FLOATING
C805 SD1L.n80 a_n13364_5836# 4.45fF
C806 SD1L.n81 a_n13364_5836# 4.45fF
C807 SD1L.n82 a_n13364_5836# 4.45fF
C808 SD1L.n83 a_n13364_5836# 4.45fF
C809 SD1L.n84 a_n13364_5836# 4.45fF
C810 SD1L.n85 a_n13364_5836# 4.45fF
C811 SD1L.n86 a_n13364_5836# 4.45fF
C812 SD1L.n87 a_n13364_5836# 4.45fF
C813 SD1L.n88 a_n13364_5836# 4.45fF
C814 SD1L.n89 a_n13364_5836# 4.45fF
C815 SD1L.n90 a_n13364_5836# 4.45fF
C816 SD1L.n91 a_n13364_5836# 4.45fF
C817 SD1L.n92 a_n13364_5836# 4.45fF
C818 SD1L.t25 a_n13364_5836# 4.04fF $ **FLOATING
C819 SD1L.n93 a_n13364_5836# 12.12fF
C820 SD1L.n94 a_n13364_5836# 5.31fF
C821 SD1L.n95 a_n13364_5836# 5.31fF
C822 SD1L.n96 a_n13364_5836# 5.31fF
C823 SD1L.n97 a_n13364_5836# 4.45fF
C824 SD1L.n98 a_n13364_5836# 5.30fF
C825 SD1L.n99 a_n13364_5836# 5.31fF
C826 SD1L.n100 a_n13364_5836# 5.31fF
C827 SD1L.n101 a_n13364_5836# 5.31fF
C828 SD1L.n102 a_n13364_5836# 5.31fF
C829 SD1L.n103 a_n13364_5836# 5.31fF
C830 SD1L.n104 a_n13364_5836# 4.53fF
C831 SD1L.n105 a_n13364_5836# 64.52fF
C832 SD1L.n106 a_n13364_5836# 110.85fF
C833 SD1L.n107 a_n13364_5836# 66.70fF
C834 SD1L.n108 a_n13364_5836# 76.52fF
C835 SD2L.n0 a_n13364_5836# 18.37fF
C836 SD2L.n1 a_n13364_5836# 21.97fF
C837 SD2L.n2 a_n13364_5836# 18.34fF
C838 SD2L.n3 a_n13364_5836# 121.57fF
C839 SD2L.n4 a_n13364_5836# 25.66fF
C840 SD2L.n5 a_n13364_5836# 18.05fF
C841 SD2L.n6 a_n13364_5836# 21.98fF
C842 SD2L.n7 a_n13364_5836# 18.37fF
C843 SD2L.n8 a_n13364_5836# 21.97fF
C844 SD2L.n9 a_n13364_5836# 18.00fF
C845 SD2L.n10 a_n13364_5836# 113.86fF
C846 SD2L.n11 a_n13364_5836# 23.54fF
C847 SD2L.n12 a_n13364_5836# 18.37fF
C848 SD2L.n13 a_n13364_5836# 21.97fF
C849 SD2L.n14 a_n13364_5836# 18.05fF
C850 SD2L.n15 a_n13364_5836# 21.98fF
C851 SD2L.n16 a_n13364_5836# 18.37fF
C852 SD2L.n17 a_n13364_5836# 21.97fF
C853 SD2L.n18 a_n13364_5836# 10.99fF
C854 SD2L.n19 a_n13364_5836# 86.72fF
C855 SD2L.n20 a_n13364_5836# 10.99fF
C856 SD2L.n21 a_n13364_5836# 86.72fF
C857 SD2L.n22 a_n13364_5836# 10.98fF
C858 SD2L.n23 a_n13364_5836# 64.82fF
C859 SD2L.n24 a_n13364_5836# 10.98fF
C860 SD2L.n25 a_n13364_5836# 57.61fF
C861 SD2L.n26 a_n13364_5836# 10.98fF
C862 SD2L.n27 a_n13364_5836# 64.82fF
C863 SD2L.n28 a_n13364_5836# 10.98fF
C864 SD2L.n29 a_n13364_5836# 57.61fF
C865 SD2L.n30 a_n13364_5836# 4.61fF
C866 SD2L.n31 a_n13364_5836# 4.61fF
C867 SD2L.n32 a_n13364_5836# 4.61fF
C868 SD2L.n33 a_n13364_5836# 4.61fF
C869 SD2L.n34 a_n13364_5836# 4.61fF
C870 SD2L.n35 a_n13364_5836# 4.61fF
C871 SD2L.n36 a_n13364_5836# 4.61fF
C872 SD2L.n37 a_n13364_5836# 4.61fF
C873 SD2L.n38 a_n13364_5836# 4.61fF
C874 SD2L.n39 a_n13364_5836# 4.61fF
C875 SD2L.n40 a_n13364_5836# 4.65fF
C876 SD2L.n41 a_n13364_5836# 4.59fF
C877 SD2L.n42 a_n13364_5836# 4.59fF
C878 SD2L.n43 a_n13364_5836# 4.59fF
C879 SD2L.n44 a_n13364_5836# 4.59fF
C880 SD2L.n45 a_n13364_5836# 4.61fF
C881 SD2L.n46 a_n13364_5836# 4.61fF
C882 SD2L.n47 a_n13364_5836# 4.61fF
C883 SD2L.n48 a_n13364_5836# 4.61fF
C884 SD2L.n49 a_n13364_5836# 4.61fF
C885 SD2L.n50 a_n13364_5836# 4.61fF
C886 SD2L.n51 a_n13364_5836# 4.61fF
C887 SD2L.n52 a_n13364_5836# 4.61fF
C888 SD2L.n53 a_n13364_5836# 4.61fF
C889 SD2L.n54 a_n13364_5836# 4.61fF
C890 SD2L.n55 a_n13364_5836# 4.61fF
C891 SD2L.t90 a_n13364_5836# 4.18fF $ **FLOATING
C892 SD2L.n56 a_n13364_5836# 4.61fF
C893 SD2L.n57 a_n13364_5836# 4.61fF
C894 SD2L.n58 a_n13364_5836# 4.61fF
C895 SD2L.t105 a_n13364_5836# 4.15fF $ **FLOATING
C896 SD2L.n59 a_n13364_5836# 4.61fF
C897 SD2L.n60 a_n13364_5836# 4.61fF
C898 SD2L.n61 a_n13364_5836# 4.61fF
C899 SD2L.n62 a_n13364_5836# 4.61fF
C900 SD2L.n63 a_n13364_5836# 4.61fF
C901 SD2L.n64 a_n13364_5836# 4.61fF
C902 SD2L.n65 a_n13364_5836# 4.61fF
C903 SD2L.n66 a_n13364_5836# 4.61fF
C904 SD2L.n67 a_n13364_5836# 4.61fF
C905 SD2L.n68 a_n13364_5836# 4.61fF
C906 SD2L.n69 a_n13364_5836# 4.65fF
C907 SD2L.n70 a_n13364_5836# 4.59fF
C908 SD2L.n71 a_n13364_5836# 4.59fF
C909 SD2L.n72 a_n13364_5836# 4.59fF
C910 SD2L.n73 a_n13364_5836# 4.59fF
C911 SD2L.n74 a_n13364_5836# 4.61fF
C912 SD2L.n75 a_n13364_5836# 4.61fF
C913 SD2L.n76 a_n13364_5836# 4.61fF
C914 SD2L.n77 a_n13364_5836# 4.61fF
C915 SD2L.n78 a_n13364_5836# 4.61fF
C916 SD2L.t144 a_n13364_5836# 4.18fF $ **FLOATING
C917 SD2L.n79 a_n13364_5836# 4.61fF
C918 SD2L.n80 a_n13364_5836# 4.61fF
C919 SD2L.n81 a_n13364_5836# 4.61fF
C920 SD2L.n82 a_n13364_5836# 4.61fF
C921 SD2L.n83 a_n13364_5836# 4.61fF
C922 SD2L.t171 a_n13364_5836# 4.18fF $ **FLOATING
C923 SD2L.n84 a_n13364_5836# 4.61fF
C924 SD2L.n85 a_n13364_5836# 4.61fF
C925 SD2L.n86 a_n13364_5836# 4.61fF
C926 SD2L.n87 a_n13364_5836# 4.61fF
C927 SD2L.n88 a_n13364_5836# 4.61fF
C928 SD2L.n89 a_n13364_5836# 4.61fF
C929 SD2L.n90 a_n13364_5836# 4.61fF
C930 SD2L.n91 a_n13364_5836# 4.61fF
C931 SD2L.n92 a_n13364_5836# 4.61fF
C932 SD2L.n93 a_n13364_5836# 4.61fF
C933 SD2L.n94 a_n13364_5836# 4.61fF
C934 SD2L.n95 a_n13364_5836# 4.61fF
C935 SD2L.n96 a_n13364_5836# 4.61fF
C936 SD2L.n97 a_n13364_5836# 4.61fF
C937 SD2L.n98 a_n13364_5836# 4.65fF
C938 SD2L.n99 a_n13364_5836# 4.59fF
C939 SD2L.n100 a_n13364_5836# 4.59fF
C940 SD2L.n101 a_n13364_5836# 4.59fF
C941 SD2L.n102 a_n13364_5836# 4.59fF
C942 SD2L.n103 a_n13364_5836# 4.61fF
C943 SD2L.n104 a_n13364_5836# 4.61fF
C944 SD2L.n105 a_n13364_5836# 4.61fF
C945 SD2L.n106 a_n13364_5836# 4.61fF
C946 SD2L.n107 a_n13364_5836# 4.61fF
C947 SD2L.n108 a_n13364_5836# 4.61fF
C948 SD2L.n109 a_n13364_5836# 4.61fF
C949 SD2L.n110 a_n13364_5836# 4.61fF
C950 SD2L.n111 a_n13364_5836# 4.61fF
C951 SD2L.n112 a_n13364_5836# 4.61fF
C952 SD2L.n113 a_n13364_5836# 4.61fF
C953 SD2L.t48 a_n13364_5836# 4.18fF $ **FLOATING
C954 SD2L.n114 a_n13364_5836# 4.61fF
C955 SD2L.n115 a_n13364_5836# 4.61fF
C956 SD2L.n116 a_n13364_5836# 4.61fF
C957 SD2L.t31 a_n13364_5836# 4.15fF $ **FLOATING
C958 SD2L.n117 a_n13364_5836# 4.61fF
C959 SD2L.n118 a_n13364_5836# 4.61fF
C960 SD2L.n119 a_n13364_5836# 4.61fF
C961 SD2L.n120 a_n13364_5836# 4.61fF
C962 SD2L.n121 a_n13364_5836# 4.61fF
C963 SD2L.t165 a_n13364_5836# 4.18fF $ **FLOATING
C964 SD2L.n122 a_n13364_5836# 4.61fF
C965 SD2L.n123 a_n13364_5836# 4.61fF
C966 SD2L.n124 a_n13364_5836# 4.61fF
C967 SD2L.n125 a_n13364_5836# 4.61fF
C968 SD2L.n126 a_n13364_5836# 4.61fF
C969 SD2L.t187 a_n13364_5836# 4.19fF $ **FLOATING
C970 SD2L.n127 a_n13364_5836# 4.61fF
C971 SD2L.n128 a_n13364_5836# 4.61fF
C972 SD2L.n129 a_n13364_5836# 4.61fF
C973 SD2L.n130 a_n13364_5836# 4.61fF
C974 SD2L.n131 a_n13364_5836# 4.59fF
C975 SD2L.n132 a_n13364_5836# 4.59fF
C976 SD2L.n133 a_n13364_5836# 4.59fF
C977 SD2L.n134 a_n13364_5836# 4.59fF
C978 SD2L.n135 a_n13364_5836# 4.61fF
C979 SD2L.n136 a_n13364_5836# 4.61fF
C980 SD2L.n137 a_n13364_5836# 4.61fF
C981 SD2L.n138 a_n13364_5836# 4.61fF
C982 SD2L.n139 a_n13364_5836# 4.61fF
C983 SD2L.n140 a_n13364_5836# 4.61fF
C984 SD2L.n141 a_n13364_5836# 4.61fF
C985 SD2L.n142 a_n13364_5836# 4.61fF
C986 SD2L.n143 a_n13364_5836# 4.61fF
C987 SD2L.n144 a_n13364_5836# 4.65fF
C988 SD2L.n145 a_n13364_5836# 4.61fF
C989 SD2L.n146 a_n13364_5836# 141.25fF
C990 SD2L.n147 a_n13364_5836# 93.54fF
C991 SD2L.n148 a_n13364_5836# 86.46fF
C992 SD2L.n149 a_n13364_5836# 58.97fF
C993 SD4R.n0 a_n13364_5836# 4.40fF
C994 SD4R.n1 a_n13364_5836# 4.40fF
C995 SD4R.n2 a_n13364_5836# 4.40fF
C996 SD4R.n3 a_n13364_5836# 4.40fF
C997 SD4R.n4 a_n13364_5836# 4.40fF
C998 SD4R.n5 a_n13364_5836# 4.40fF
C999 SD4R.n6 a_n13364_5836# 4.40fF
C1000 SD4R.n7 a_n13364_5836# 4.40fF
C1001 SD4R.n8 a_n13364_5836# 4.40fF
C1002 SD4R.n9 a_n13364_5836# 4.40fF
C1003 SD4R.n10 a_n13364_5836# 4.40fF
C1004 SD4R.t99 a_n13364_5836# 3.99fF $ **FLOATING
C1005 SD4R.n11 a_n13364_5836# 11.94fF
C1006 SD4R.n12 a_n13364_5836# 5.25fF
C1007 SD4R.n13 a_n13364_5836# 5.25fF
C1008 SD4R.n14 a_n13364_5836# 5.25fF
C1009 SD4R.n15 a_n13364_5836# 5.25fF
C1010 SD4R.n16 a_n13364_5836# 5.25fF
C1011 SD4R.n17 a_n13364_5836# 5.25fF
C1012 SD4R.n18 a_n13364_5836# 5.25fF
C1013 SD4R.n19 a_n13364_5836# 5.25fF
C1014 SD4R.n20 a_n13364_5836# 5.25fF
C1015 SD4R.n21 a_n13364_5836# 5.20fF
C1016 SD4R.t93 a_n13364_5836# 3.96fF $ **FLOATING
C1017 SD4R.n22 a_n13364_5836# 4.40fF
C1018 SD4R.n23 a_n13364_5836# 4.40fF
C1019 SD4R.n24 a_n13364_5836# 4.40fF
C1020 SD4R.n25 a_n13364_5836# 77.21fF
C1021 SD4R.n26 a_n13364_5836# 4.40fF
C1022 SD4R.n27 a_n13364_5836# 4.40fF
C1023 SD4R.n28 a_n13364_5836# 4.40fF
C1024 SD4R.n29 a_n13364_5836# 4.40fF
C1025 SD4R.n30 a_n13364_5836# 4.40fF
C1026 SD4R.n31 a_n13364_5836# 4.40fF
C1027 SD4R.n32 a_n13364_5836# 4.40fF
C1028 SD4R.n33 a_n13364_5836# 4.40fF
C1029 SD4R.n34 a_n13364_5836# 4.40fF
C1030 SD4R.n35 a_n13364_5836# 4.40fF
C1031 SD4R.t31 a_n13364_5836# 3.99fF $ **FLOATING
C1032 SD4R.n36 a_n13364_5836# 11.94fF
C1033 SD4R.n37 a_n13364_5836# 4.40fF
C1034 SD4R.n38 a_n13364_5836# 5.24fF
C1035 SD4R.n39 a_n13364_5836# 5.25fF
C1036 SD4R.n40 a_n13364_5836# 5.25fF
C1037 SD4R.n41 a_n13364_5836# 5.25fF
C1038 SD4R.n42 a_n13364_5836# 5.25fF
C1039 SD4R.n43 a_n13364_5836# 5.25fF
C1040 SD4R.n44 a_n13364_5836# 5.25fF
C1041 SD4R.n45 a_n13364_5836# 5.25fF
C1042 SD4R.n46 a_n13364_5836# 5.25fF
C1043 SD4R.n47 a_n13364_5836# 5.20fF
C1044 SD4R.t65 a_n13364_5836# 3.96fF $ **FLOATING
C1045 SD4R.n48 a_n13364_5836# 4.40fF
C1046 SD4R.n49 a_n13364_5836# 4.40fF
C1047 SD4R.n50 a_n13364_5836# 4.40fF
C1048 SD4R.n51 a_n13364_5836# 85.16fF
C1049 SD4R.n52 a_n13364_5836# 4.40fF
C1050 SD4R.n53 a_n13364_5836# 4.40fF
C1051 SD4R.n54 a_n13364_5836# 4.40fF
C1052 SD4R.n55 a_n13364_5836# 4.40fF
C1053 SD4R.n56 a_n13364_5836# 4.40fF
C1054 SD4R.n57 a_n13364_5836# 4.40fF
C1055 SD4R.n58 a_n13364_5836# 4.40fF
C1056 SD4R.n59 a_n13364_5836# 4.40fF
C1057 SD4R.n60 a_n13364_5836# 4.40fF
C1058 SD4R.n61 a_n13364_5836# 4.40fF
C1059 SD4R.n62 a_n13364_5836# 4.44fF
C1060 SD4R.n63 a_n13364_5836# 12.29fF
C1061 SD4R.n64 a_n13364_5836# 5.24fF
C1062 SD4R.n65 a_n13364_5836# 5.24fF
C1063 SD4R.n66 a_n13364_5836# 5.24fF
C1064 SD4R.n67 a_n13364_5836# 5.24fF
C1065 SD4R.n68 a_n13364_5836# 5.24fF
C1066 SD4R.n69 a_n13364_5836# 5.24fF
C1067 SD4R.n70 a_n13364_5836# 5.24fF
C1068 SD4R.n71 a_n13364_5836# 5.24fF
C1069 SD4R.n72 a_n13364_5836# 5.41fF
C1070 SD4R.n73 a_n13364_5836# 4.38fF
C1071 SD4R.n74 a_n13364_5836# 3.82fF
C1072 SD4R.n75 a_n13364_5836# 4.38fF
C1073 SD4R.n76 a_n13364_5836# 4.37fF
C1074 SD4R.n77 a_n13364_5836# 4.37fF
C1075 SD4R.n78 a_n13364_5836# 145.55fF
C1076 SD4R.n79 a_n13364_5836# 97.56fF
C1077 SD4R.n80 a_n13364_5836# 4.40fF
C1078 SD4R.n81 a_n13364_5836# 4.40fF
C1079 SD4R.n82 a_n13364_5836# 4.40fF
C1080 SD4R.n83 a_n13364_5836# 4.40fF
C1081 SD4R.n84 a_n13364_5836# 4.40fF
C1082 SD4R.n85 a_n13364_5836# 4.40fF
C1083 SD4R.n86 a_n13364_5836# 4.40fF
C1084 SD4R.n87 a_n13364_5836# 4.40fF
C1085 SD4R.n88 a_n13364_5836# 4.40fF
C1086 SD4R.n89 a_n13364_5836# 4.40fF
C1087 SD4R.n90 a_n13364_5836# 4.44fF
C1088 SD4R.n91 a_n13364_5836# 12.29fF
C1089 SD4R.n92 a_n13364_5836# 5.24fF
C1090 SD4R.n93 a_n13364_5836# 5.24fF
C1091 SD4R.n94 a_n13364_5836# 5.24fF
C1092 SD4R.n95 a_n13364_5836# 5.24fF
C1093 SD4R.n96 a_n13364_5836# 5.24fF
C1094 SD4R.n97 a_n13364_5836# 5.24fF
C1095 SD4R.n98 a_n13364_5836# 5.24fF
C1096 SD4R.n99 a_n13364_5836# 5.24fF
C1097 SD4R.n100 a_n13364_5836# 5.17fF
C1098 SD4R.n101 a_n13364_5836# 4.38fF
C1099 SD4R.n102 a_n13364_5836# 4.75fF
C1100 SD4R.n103 a_n13364_5836# 4.38fF
C1101 SD4R.n104 a_n13364_5836# 4.38fF
C1102 SD4R.n105 a_n13364_5836# 4.38fF
C1103 SD4R.n106 a_n13364_5836# 73.16fF
C1104 SD3R.n0 a_n13364_5836# 28.85fF
C1105 SD3R.n1 a_n13364_5836# 18.08fF
C1106 SD3R.n2 a_n13364_5836# 21.62fF
C1107 SD3R.n3 a_n13364_5836# 17.72fF
C1108 SD3R.n4 a_n13364_5836# 21.64fF
C1109 SD3R.n5 a_n13364_5836# 21.64fF
C1110 SD3R.n6 a_n13364_5836# 28.85fF
C1111 SD3R.n7 a_n13364_5836# 17.72fF
C1112 SD3R.n8 a_n13364_5836# 21.64fF
C1113 SD3R.n9 a_n13364_5836# 21.64fF
C1114 SD3R.n10 a_n13364_5836# 18.08fF
C1115 SD3R.n11 a_n13364_5836# 21.62fF
C1116 SD3R.n12 a_n13364_5836# 17.72fF
C1117 SD3R.n13 a_n13364_5836# 21.64fF
C1118 SD3R.n14 a_n13364_5836# 21.64fF
C1119 SD3R.n15 a_n13364_5836# 17.72fF
C1120 SD3R.n16 a_n13364_5836# 21.64fF
C1121 SD3R.n17 a_n13364_5836# 21.64fF
C1122 SD3R.n18 a_n13364_5836# 10.81fF
C1123 SD3R.n19 a_n13364_5836# 81.85fF
C1124 SD3R.n20 a_n13364_5836# 10.81fF
C1125 SD3R.n21 a_n13364_5836# 141.30fF
C1126 SD3R.n22 a_n13364_5836# 18.08fF
C1127 SD3R.n23 a_n13364_5836# 76.14fF
C1128 SD3R.n24 a_n13364_5836# 18.08fF
C1129 SD3R.n25 a_n13364_5836# 76.14fF
C1130 SD3R.n26 a_n13364_5836# 85.47fF
C1131 SD3R.n27 a_n13364_5836# 84.99fF
C1132 SD3R.n28 a_n13364_5836# 99.11fF
C1133 SD3R.n29 a_n13364_5836# 84.99fF
C1134 SD3R.n30 a_n13364_5836# 4.54fF
C1135 SD3R.n31 a_n13364_5836# 4.54fF
C1136 SD3R.n32 a_n13364_5836# 4.54fF
C1137 SD3R.n33 a_n13364_5836# 4.54fF
C1138 SD3R.n34 a_n13364_5836# 4.54fF
C1139 SD3R.n35 a_n13364_5836# 4.58fF
C1140 SD3R.n36 a_n13364_5836# 4.54fF
C1141 SD3R.n37 a_n13364_5836# 4.54fF
C1142 SD3R.n38 a_n13364_5836# 4.54fF
C1143 SD3R.n39 a_n13364_5836# 4.54fF
C1144 SD3R.n40 a_n13364_5836# 4.58fF
C1145 SD3R.n41 a_n13364_5836# 4.51fF
C1146 SD3R.n42 a_n13364_5836# 4.51fF
C1147 SD3R.n43 a_n13364_5836# 4.51fF
C1148 SD3R.n44 a_n13364_5836# 4.51fF
C1149 SD3R.n45 a_n13364_5836# 4.54fF
C1150 SD3R.n46 a_n13364_5836# 4.54fF
C1151 SD3R.n47 a_n13364_5836# 4.54fF
C1152 SD3R.n48 a_n13364_5836# 4.54fF
C1153 SD3R.n49 a_n13364_5836# 4.54fF
C1154 SD3R.n50 a_n13364_5836# 4.54fF
C1155 SD3R.n51 a_n13364_5836# 4.54fF
C1156 SD3R.n52 a_n13364_5836# 4.54fF
C1157 SD3R.n53 a_n13364_5836# 4.54fF
C1158 SD3R.n54 a_n13364_5836# 4.54fF
C1159 SD3R.n55 a_n13364_5836# 4.54fF
C1160 SD3R.t213 a_n13364_5836# 4.11fF $ **FLOATING
C1161 SD3R.t185 a_n13364_5836# 4.09fF $ **FLOATING
C1162 SD3R.n56 a_n13364_5836# 4.54fF
C1163 SD3R.n57 a_n13364_5836# 4.54fF
C1164 SD3R.n58 a_n13364_5836# 4.54fF
C1165 SD3R.n59 a_n13364_5836# 4.54fF
C1166 SD3R.n60 a_n13364_5836# 4.54fF
C1167 SD3R.n61 a_n13364_5836# 4.54fF
C1168 SD3R.n62 a_n13364_5836# 4.54fF
C1169 SD3R.n63 a_n13364_5836# 4.54fF
C1170 SD3R.n64 a_n13364_5836# 4.54fF
C1171 SD3R.n65 a_n13364_5836# 4.54fF
C1172 SD3R.n66 a_n13364_5836# 4.54fF
C1173 SD3R.n67 a_n13364_5836# 4.54fF
C1174 SD3R.n68 a_n13364_5836# 4.54fF
C1175 SD3R.n69 a_n13364_5836# 4.58fF
C1176 SD3R.n70 a_n13364_5836# 4.52fF
C1177 SD3R.n71 a_n13364_5836# 4.51fF
C1178 SD3R.n72 a_n13364_5836# 4.51fF
C1179 SD3R.n73 a_n13364_5836# 4.51fF
C1180 SD3R.n74 a_n13364_5836# 4.54fF
C1181 SD3R.n75 a_n13364_5836# 4.54fF
C1182 SD3R.n76 a_n13364_5836# 4.54fF
C1183 SD3R.n77 a_n13364_5836# 4.54fF
C1184 SD3R.n78 a_n13364_5836# 4.54fF
C1185 SD3R.n79 a_n13364_5836# 4.54fF
C1186 SD3R.n80 a_n13364_5836# 4.54fF
C1187 SD3R.n81 a_n13364_5836# 4.54fF
C1188 SD3R.n82 a_n13364_5836# 4.54fF
C1189 SD3R.n83 a_n13364_5836# 4.54fF
C1190 SD3R.n84 a_n13364_5836# 4.54fF
C1191 SD3R.t22 a_n13364_5836# 4.12fF $ **FLOATING
C1192 SD3R.n85 a_n13364_5836# 4.54fF
C1193 SD3R.n86 a_n13364_5836# 4.53fF
C1194 SD3R.n87 a_n13364_5836# 4.53fF
C1195 SD3R.t23 a_n13364_5836# 4.08fF $ **FLOATING
C1196 SD3R.n88 a_n13364_5836# 4.54fF
C1197 SD3R.n89 a_n13364_5836# 4.54fF
C1198 SD3R.n90 a_n13364_5836# 4.54fF
C1199 SD3R.n91 a_n13364_5836# 4.54fF
C1200 SD3R.n92 a_n13364_5836# 4.54fF
C1201 SD3R.n93 a_n13364_5836# 4.54fF
C1202 SD3R.n94 a_n13364_5836# 4.54fF
C1203 SD3R.n95 a_n13364_5836# 4.54fF
C1204 SD3R.n96 a_n13364_5836# 4.54fF
C1205 SD3R.n97 a_n13364_5836# 4.54fF
C1206 SD3R.n98 a_n13364_5836# 4.54fF
C1207 SD3R.t139 a_n13364_5836# 4.11fF $ **FLOATING
C1208 SD3R.t220 a_n13364_5836# 4.09fF $ **FLOATING
C1209 SD3R.n99 a_n13364_5836# 4.54fF
C1210 SD3R.n100 a_n13364_5836# 4.54fF
C1211 SD3R.n101 a_n13364_5836# 4.54fF
C1212 SD3R.n102 a_n13364_5836# 4.54fF
C1213 SD3R.n103 a_n13364_5836# 4.54fF
C1214 SD3R.n104 a_n13364_5836# 4.54fF
C1215 SD3R.n105 a_n13364_5836# 4.54fF
C1216 SD3R.n106 a_n13364_5836# 4.54fF
C1217 SD3R.n107 a_n13364_5836# 4.54fF
C1218 SD3R.n108 a_n13364_5836# 4.54fF
C1219 SD3R.n109 a_n13364_5836# 4.54fF
C1220 SD3R.n110 a_n13364_5836# 4.54fF
C1221 SD3R.n111 a_n13364_5836# 4.54fF
C1222 SD3R.n112 a_n13364_5836# 4.58fF
C1223 SD3R.n113 a_n13364_5836# 4.52fF
C1224 SD3R.n114 a_n13364_5836# 4.51fF
C1225 SD3R.n115 a_n13364_5836# 4.51fF
C1226 SD3R.n116 a_n13364_5836# 4.51fF
C1227 SD3R.n117 a_n13364_5836# 4.54fF
C1228 SD3R.n118 a_n13364_5836# 4.54fF
C1229 SD3R.n119 a_n13364_5836# 4.54fF
C1230 SD3R.n120 a_n13364_5836# 4.54fF
C1231 SD3R.n121 a_n13364_5836# 4.54fF
C1232 SD3R.n122 a_n13364_5836# 4.54fF
C1233 SD3R.n123 a_n13364_5836# 4.54fF
C1234 SD3R.n124 a_n13364_5836# 4.54fF
C1235 SD3R.n125 a_n13364_5836# 4.54fF
C1236 SD3R.n126 a_n13364_5836# 4.54fF
C1237 SD3R.n127 a_n13364_5836# 4.54fF
C1238 SD3R.t48 a_n13364_5836# 4.11fF $ **FLOATING
C1239 SD3R.t42 a_n13364_5836# 4.09fF $ **FLOATING
C1240 SD3R.n128 a_n13364_5836# 4.54fF
C1241 SD3R.n129 a_n13364_5836# 4.54fF
C1242 SD3R.n130 a_n13364_5836# 4.54fF
C1243 SD3R.n131 a_n13364_5836# 68.48fF
C1244 SD3R.n132 a_n13364_5836# 4.51fF
C1245 SD3R.n133 a_n13364_5836# 4.51fF
C1246 SD3R.n134 a_n13364_5836# 4.51fF
C1247 SD3R.n135 a_n13364_5836# 4.51fF
C1248 SD3R.n136 a_n13364_5836# 4.54fF
C1249 SD3R.n137 a_n13364_5836# 4.54fF
C1250 SD3R.n138 a_n13364_5836# 4.54fF
C1251 SD3R.n139 a_n13364_5836# 4.54fF
C1252 SD3R.n140 a_n13364_5836# 4.58fF
C1253 SD3R.n141 a_n13364_5836# 4.54fF
C1254 SD3R.n142 a_n13364_5836# 4.54fF
C1255 SD3R.n143 a_n13364_5836# 4.54fF
C1256 SD3R.n144 a_n13364_5836# 4.54fF
C1257 SD3R.n145 a_n13364_5836# 4.58fF
C1258 SD3R.n146 a_n13364_5836# 4.54fF
C1259 SD3R.n147 a_n13364_5836# 59.82fF
C1260 SD3R.n148 a_n13364_5836# 84.30fF
C1261 SD3R.n149 a_n13364_5836# 68.48fF
C1262 SD3R.n150 a_n13364_5836# 53.06fF
