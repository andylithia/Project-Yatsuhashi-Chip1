** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/LNAs.sch
**.subckt LNAs
XM1 n_ds1 vgate1 net1 GND sky130_fd_pr__nfet_01v8 L=L W=W nf=NF ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=M m=M
Ldeg1 net1 GND 1n m=1
V1 net2 GND 1.8
V2 net3 GND dc 0 ac 0 portnum 1 z0 50
C2 net5 net3 1u m=1
V3 net4 GND dc 0 ac 0 portnum 2 z0 50
C4 net4 net6 1u m=1
Ldeg2 vgate1 net5 0 m=1
XM2 vbias1 vbias1 GND GND sky130_fd_pr__nfet_01v8 L=L W=W nf=NF ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=M m=M
R1 vbias1 vgate1 10k m=1
C1 vbias1 GND 100p m=1
I0 net2 vbias1 2m
Lload1 net2 n_ds1 5n m=1
V4 __UNCONNECTED_PIN__0 GND 1.8
XM3 net2 n_ds1 net6 GND sky130_fd_pr__nfet_01v8 L=L W=W nf=NF ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=M m=M
I1 net7 GND 2m
Lload2 net6 net7 100n m=1
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.param L=2
.param W=40
.param W2=20
.param NF=1
.param M=1
.op
.dc V4 0 1.8 0.01
.plot @m.xm1.msky130_fd_pr__nfet_01v8[vgs]
.plot @m.xm1.msky130_fd_pr__nfet_01v8[vds]
.print @m.xm3.msky130_fd_pr__nfet_01v8[vgs]
.print @m.xm3.msky130_fd_pr__nfet_01v8[vds]
.sp dec 100 1e9 100e9 0
.control
run
display
plot db(S_1_1) db(S_1_2) db(S_2_2) db(S_2_1)
plot S_1_1 smithgrid
print @m.xm1.msky130_fd_pr__nfet_01v8[id]
print @m.xm1.msky130_fd_pr__nfet_01v8[vgs]
print @m.xm1.msky130_fd_pr__nfet_01v8[vds]
print @m.xm3.msky130_fd_pr__nfet_01v8[vgs]
print @m.xm3.msky130_fd_pr__nfet_01v8[vds]
print @m.xm3.msky130_fd_pr__nfet_01v8[id]
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
