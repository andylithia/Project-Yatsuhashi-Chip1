.subckt NMOS_30_0p5_30_diff4x_2 SD1L SD2L GL SD1R SD2R GR SUB
X0 SD2L.t119 GL SD1L.t47 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X1 SD1L.t33 GL SD2L.t118 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X2 SD2L.t117 GL SD1L.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X3 SD2L.t116 GL SD1L.t22 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X4 SD2R.t119 GR SD1R.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X5 SD1L.t29 GL SD2L.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X6 SD1R.t6 GR SD2R.t118 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X7 SD1R.t48 GR SD2R.t117 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X8 SD2L.t114 GL SD1L.t68 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X9 SD1L.t46 GL SD2L.t113 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X10 SD2R.t116 GR SD1R.t89 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X11 SD1L.t113 GL SD2L.t112 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X12 SD1R.t72 GR SD2R.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X13 SD1L.t32 GL SD2L.t111 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X14 SD1L.t27 GL SD2L.t110 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X15 SD2R.t114 GR SD1R.t93 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X16 SD1L.t100 GL SD2L.t109 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X17 SD2R.t113 GR SD1R.t90 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X18 SD2R.t112 GR SD1R.t70 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X19 SD1L.t19 GL SD2L.t108 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X20 SD1L.t112 GL SD2L.t107 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X21 SD2R.t111 GR SD1R.t71 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X22 SD2L.t106 GL SD1L.t17 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X23 SD1R.t29 GR SD2R.t110 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X24 SD1L.t110 GL SD2L.t105 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X25 SD2R.t109 GR SD1R.t7 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X26 SD2L.t104 GL SD1L.t108 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X27 SD1R.t2 GR SD2R.t108 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X28 SD1L.t36 GL SD2L.t103 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X29 SD2L.t102 GL SD1L.t31 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X30 SD1R.t14 GR SD2R.t107 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X31 SD2R.t106 GR SD1R.t99 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X32 SD2L.t101 GL SD1L.t111 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X33 SD2R.t105 GR SD1R.t57 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X34 SD2L.t100 GL SD1L.t34 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X35 SD1R.t52 GR SD2R.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X36 SD2L.t99 GL SD1L.t35 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X37 SD1R.t105 GR SD2R.t103 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X38 SD2R.t102 GR SD1R.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X39 SD1L.t23 GL SD2L.t98 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X40 SD1L.t93 GL SD2L.t97 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X41 SD2R.t101 GR SD1R.t19 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X42 SD1L.t28 GL SD2L.t96 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X43 SD1L.t69 GL SD2L.t95 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X44 SD2L.t94 GL SD1L.t38 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X45 SD2R.t100 GR SD1R.t34 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X46 SD2L.t93 GL SD1L.t73 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X47 SD1R.t41 GR SD2R.t99 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X48 SD1R.t30 GR SD2R.t98 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X49 SD1L.t99 GL SD2L.t92 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X50 SD2L.t91 GL SD1L.t50 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X51 SD1L.t98 GL SD2L.t90 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X52 SD2R.t97 GR SD1R.t58 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X53 SD1L.t13 GL SD2L.t89 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X54 SD1L.t30 GL SD2L.t88 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X55 SD2L.t87 GL SD1L.t18 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X56 SD2L.t86 GL SD1L.t37 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X57 SD2R.t96 GR SD1R.t73 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X58 SD2L.t85 GL SD1L.t5 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X59 SD2L.t84 GL SD1L.t8 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X60 SD1L.t105 GL SD2L.t83 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X61 SD1R.t94 GR SD2R.t95 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X62 SD1R.t16 GR SD2R.t94 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X63 SD2R.t93 GR SD1R.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X64 SD1R.t95 GR SD2R.t92 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X65 SD2R.t91 GR SD1R.t84 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X66 SD2R.t90 GR SD1R.t85 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X67 SD1L.t51 GL SD2L.t82 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X68 SD2R.t89 GR SD1R.t112 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X69 SD1R.t74 GR SD2R.t88 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X70 SD2R.t87 GR SD1R.t82 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X71 SD2L.t81 GL SD1L.t52 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X72 SD1R.t33 GR SD2R.t86 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X73 SD1L.t53 GL SD2L.t80 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X74 SD2L.t79 GL SD1L.t54 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X75 SD2R.t85 GR SD1R.t83 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X76 SD2R.t84 GR SD1R.t0 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X77 SD1L.t55 GL SD2L.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X78 SD2L.t77 GL SD1L.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X79 SD2R.t83 GR SD1R.t86 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X80 SD2R.t82 GR SD1R.t8 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X81 SD1R.t1 GR SD2R.t81 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X82 SD2R.t80 GR SD1R.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X83 SD1L.t57 GL SD2L.t76 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X84 SD1R.t113 GR SD2R.t79 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X85 SD2L.t75 GL SD1L.t58 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X86 SD2R.t78 GR SD1R.t75 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X87 SD2L.t74 GL SD1L.t59 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X88 SD2R.t77 GR SD1R.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X89 SD1L.t60 GL SD2L.t73 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X90 SD2R.t76 GR SD1R.t5 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X91 SD2R.t75 GR SD1R.t96 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X92 SD1L.t61 GL SD2L.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X93 SD1R.t59 GR SD2R.t74 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X94 SD2L.t71 GL SD1L.t62 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X95 SD1R.t53 GR SD2R.t73 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X96 SD1R.t35 GR SD2R.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X97 SD2R.t71 GR SD1R.t114 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X98 SD2R.t70 GR SD1R.t42 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X99 SD2L.t70 GL SD1L.t63 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X100 SD2L.t69 GL SD1L.t64 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X101 SD1R.t76 GR SD2R.t69 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X102 SD2L.t68 GL SD1L.t65 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X103 SD2R.t68 GR SD1R.t97 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X104 SD2R.t67 GR SD1R.t60 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X105 SD2L.t67 GL SD1L.t66 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X106 SD2L.t66 GL SD1L.t67 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X107 SD1R.t54 GR SD2R.t66 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X108 SD2L.t65 GL SD1L.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X109 SD2L.t64 GL SD1L.t0 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X110 SD1R.t106 GR SD2R.t65 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X111 SD1R.t36 GR SD2R.t64 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X112 SD2L.t63 GL SD1L.t1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X113 SD1L.t6 GL SD2L.t62 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X114 SD2R.t63 GR SD1R.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X115 SD1R.t43 GR SD2R.t62 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X116 SD2R.t61 GR SD1R.t77 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X117 SD1L.t70 GL SD2L.t61 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X118 SD1L.t20 GL SD2L.t60 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X119 SD2R.t60 GR SD1R.t98 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X120 SD1L.t71 GL SD2L.t59 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X121 SD1L.t21 GL SD2L.t58 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X122 SD1R.t61 GR SD2R.t59 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X123 SD2L.t57 GL SD1L.t7 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X124 SD1L.t114 GL SD2L.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X125 SD2R.t58 GR SD1R.t55 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X126 SD2R.t57 GR SD1R.t107 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X127 SD2L.t55 GL SD1L.t116 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X128 SD1L.t118 GL SD2L.t54 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X129 SD2L.t53 GL SD1L.t109 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X130 SD2L.t52 GL SD1L.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X131 SD2R.t56 GR SD1R.t62 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X132 SD2L.t51 GL SD1L.t117 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X133 SD1R.t37 GR SD2R.t55 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X134 SD2L.t50 GL SD1L.t106 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X135 SD1L.t74 GL SD2L.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X136 SD2L.t48 GL SD1L.t75 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X137 SD2R.t54 GR SD1R.t116 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X138 SD1R.t44 GR SD2R.t53 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X139 SD1L.t76 GL SD2L.t47 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X140 SD2L.t46 GL SD1L.t77 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X141 SD2R.t52 GR SD1R.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X142 SD1L.t78 GL SD2L.t45 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X143 SD1R.t100 GR SD2R.t51 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X144 SD2L.t44 GL SD1L.t79 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X145 SD1R.t63 GR SD2R.t50 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X146 SD1R.t108 GR SD2R.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X147 SD1L.t2 GL SD2L.t43 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X148 SD2L.t42 GL SD1L.t80 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X149 SD1L.t81 GL SD2L.t41 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X150 SD1L.t82 GL SD2L.t40 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X151 SD1L.t83 GL SD2L.t39 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X152 SD2R.t48 GR SD1R.t20 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X153 SD1L.t84 GL SD2L.t38 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X154 SD2R.t47 GR SD1R.t32 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X155 SD2L.t37 GL SD1L.t85 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X156 SD2R.t46 GR SD1R.t25 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X157 SD1R.t11 GR SD2R.t45 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X158 SD2L.t36 GL SD1L.t86 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X159 SD1R.t91 GR SD2R.t44 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X160 SD2L.t35 GL SD1L.t87 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X161 SD1R.t3 GR SD2R.t43 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X162 SD2L.t34 GL SD1L.t88 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X163 SD1R.t92 GR SD2R.t42 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X164 SD2R.t41 GR SD1R.t31 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X165 SD2L.t33 GL SD1L.t89 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X166 SD2L.t32 GL SD1L.t90 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X167 SD2L.t31 GL SD1L.t91 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X168 SD1L.t48 GL SD2L.t30 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X169 SD1R.t12 GR SD2R.t40 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X170 SD2L.t29 GL SD1L.t92 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X171 SD1L.t94 GL SD2L.t28 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X172 SD1R.t117 GR SD2R.t39 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X173 SD1R.t79 GR SD2R.t38 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X174 SD1L.t97 GL SD2L.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X175 SD1L.t96 GL SD2L.t26 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X176 SD1R.t13 GR SD2R.t37 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X177 SD1R.t15 GR SD2R.t36 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X178 SD2L.t25 GL SD1L.t101 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X179 SD1R.t101 GR SD2R.t35 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X180 SD2L.t24 GL SD1L.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X181 SD1L.t103 GL SD2L.t23 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X182 SD1L.t95 GL SD2L.t22 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X183 SD2R.t34 GR SD1R.t64 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X184 SD1R.t21 GR SD2R.t33 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X185 SD2L.t21 GL SD1L.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X186 SD1R.t38 GR SD2R.t32 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X187 SD1L.t119 GL SD2L.t20 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X188 SD1R.t45 GR SD2R.t31 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X189 SD1L.t107 GL SD2L.t19 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X190 SD2R.t30 GR SD1R.t109 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X191 SD2R.t29 GR SD1R.t39 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X192 SD1R.t118 GR SD2R.t28 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X193 SD1L.t42 GL SD2L.t18 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X194 SD2R.t27 GR SD1R.t26 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X195 SD2R.t26 GR SD1R.t46 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X196 SD1R.t80 GR SD2R.t25 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X197 SD2L.t17 GL SD1L.t14 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X198 SD1L.t25 GL SD2L.t16 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X199 SD2R.t24 GR SD1R.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X200 SD2R.t23 GR SD1R.t65 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X201 SD2R.t22 GR SD1R.t110 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X202 SD1L.t43 GL SD2L.t15 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X203 SD1R.t22 GR SD2R.t21 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X204 SD1L.t3 GL SD2L.t14 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X205 SD1R.t40 GR SD2R.t20 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X206 SD1R.t119 GR SD2R.t19 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X207 SD2R.t18 GR SD1R.t47 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X208 SD1R.t81 GR SD2R.t17 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X209 SD2R.t16 GR SD1R.t103 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X210 SD1R.t66 GR SD2R.t15 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X211 SD1R.t111 GR SD2R.t14 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X212 SD2R.t13 GR SD1R.t23 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X213 SD1L.t15 GL SD2L.t13 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X214 SD1R.t4 GR SD2R.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X215 SD2R.t11 GR SD1R.t67 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X216 SD2R.t10 GR SD1R.t24 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X217 SD1R.t50 GR SD2R.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X218 SD2L.t12 GL SD1L.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X219 SD1L.t26 GL SD2L.t11 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X220 SD2L.t10 GL SD1L.t41 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X221 SD1L.t24 GL SD2L.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X222 SD1R.t17 GR SD2R.t8 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X223 SD2L.t8 GL SD1L.t44 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X224 SD2L.t7 GL SD1L.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X225 SD1L.t40 GL SD2L.t6 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X226 SD1R.t68 GR SD2R.t7 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X227 SD1L.t45 GL SD2L.t5 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X228 SD2R.t6 GR SD1R.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X229 SD1R.t51 GR SD2R.t5 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X230 SD2R.t4 GR SD1R.t18 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X231 SD1L.t4 GL SD2L.t4 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X232 SD1R.t69 GR SD2R.t3 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X233 SD2L.t3 GL SD1L.t39 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X234 SD1L.t16 GL SD2L.t2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X235 SD1R.t28 GR SD2R.t2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X236 SD2R.t1 GR SD1R.t87 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X237 SD1R.t88 GR SD2R.t0 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X238 SD2L.t1 GL SD1L.t11 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X239 SD2L.t0 GL SD1L.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
C0 SD1L SD1R 68.17fF
C1 GR SD2L 15.75fF
C2 SD1R GL 13.75fF
C3 SD1R SD2R 832.35fF
C4 SD1L GL 97.85fF
C5 SD1L SD2R 39.99fF
C6 SD2R GL 16.59fF
C7 m4_11500_n11600# SD2L 2.89fF
C8 SD1R GR 93.48fF
C9 SD1L GR 16.95fF
C10 GR GL 28.25fF
C11 SD2R GR 99.27fF
C12 SD1R SD2L 34.60fF
C13 SD1L SD2L 832.59fF
C14 SD2L GL 97.33fF
C15 SD2R SD2L 57.01fF
R0 SD1L.n13 SD1L.t53 1.972
R1 SD1L.n0 SD1L.t5 1.972
R2 SD1L.n8 SD1L.t42 1.972
R3 SD1L.n6 SD1L.t44 1.972
R4 SD1L.n4 SD1L.n39 1.435
R5 SD1L.n2 SD1L.n28 1.435
R6 SD1L.n11 SD1L.n29 1.428
R7 SD1L.n11 SD1L.n30 1.428
R8 SD1L.n10 SD1L.n31 1.428
R9 SD1L.n10 SD1L.n32 1.428
R10 SD1L.n5 SD1L.n33 1.428
R11 SD1L.n5 SD1L.n34 1.428
R12 SD1L.n5 SD1L.n35 1.428
R13 SD1L.n5 SD1L.n36 1.428
R14 SD1L.n4 SD1L.n37 1.428
R15 SD1L.n4 SD1L.n38 1.428
R16 SD1L.n9 SD1L.n18 1.428
R17 SD1L.n9 SD1L.n19 1.428
R18 SD1L.n9 SD1L.n20 1.428
R19 SD1L.n3 SD1L.n21 1.428
R20 SD1L.n3 SD1L.n22 1.428
R21 SD1L.n3 SD1L.n23 1.428
R22 SD1L.n3 SD1L.n24 1.428
R23 SD1L.n2 SD1L.n25 1.428
R24 SD1L.n2 SD1L.n26 1.428
R25 SD1L.n2 SD1L.n27 1.428
R26 SD1L.n1 SD1L.n62 1.414
R27 SD1L.n12 SD1L.n63 1.414
R28 SD1L.n12 SD1L.n64 1.414
R29 SD1L.n13 SD1L.n65 1.414
R30 SD1L.n13 SD1L.n66 1.414
R31 SD1L.n0 SD1L.n72 1.414
R32 SD1L.n0 SD1L.n71 1.414
R33 SD1L.n1 SD1L.n70 1.414
R34 SD1L.n1 SD1L.n69 1.414
R35 SD1L.n1 SD1L.n68 1.414
R36 SD1L.n7 SD1L.n49 1.414
R37 SD1L.n7 SD1L.n50 1.414
R38 SD1L.n8 SD1L.n51 1.414
R39 SD1L.n8 SD1L.n52 1.414
R40 SD1L.n8 SD1L.n53 1.414
R41 SD1L.n6 SD1L.n48 1.414
R42 SD1L.n6 SD1L.n47 1.414
R43 SD1L.n7 SD1L.n46 1.414
R44 SD1L.n7 SD1L.n45 1.414
R45 SD1L.n7 SD1L.n44 1.414
R46 SD1L.n7 SD1L.n57 1.412
R47 SD1L.n7 SD1L.n56 1.412
R48 SD1L.n7 SD1L.n55 1.412
R49 SD1L.n7 SD1L.n54 1.412
R50 SD1L.n1 SD1L.n59 1.412
R51 SD1L.n1 SD1L.n60 1.412
R52 SD1L.n1 SD1L.n61 1.412
R53 SD1L.n1 SD1L.n67 1.41
R54 SD1L.n11 SD1L.n40 1.281
R55 SD1L.n11 SD1L.n41 1.28
R56 SD1L.n11 SD1L.n42 1.28
R57 SD1L.n11 SD1L.n43 1.28
R58 SD1L.n9 SD1L.n16 1.279
R59 SD1L.n9 SD1L.n15 1.279
R60 SD1L.n9 SD1L.n14 1.279
R61 SD1L.n9 SD1L.n17 1.278
R62 SD1L.n62 SD1L.t92 0.551
R63 SD1L.n62 SD1L.t70 0.551
R64 SD1L.n63 SD1L.t72 0.551
R65 SD1L.n63 SD1L.t19 0.551
R66 SD1L.n64 SD1L.t12 0.551
R67 SD1L.n64 SD1L.t71 0.551
R68 SD1L.n65 SD1L.t1 0.551
R69 SD1L.n65 SD1L.t13 0.551
R70 SD1L.n66 SD1L.t10 0.551
R71 SD1L.n66 SD1L.t118 0.551
R72 SD1L.n72 SD1L.t117 0.551
R73 SD1L.n72 SD1L.t69 0.551
R74 SD1L.n71 SD1L.t9 0.551
R75 SD1L.n71 SD1L.t45 0.551
R76 SD1L.n70 SD1L.t87 0.551
R77 SD1L.n70 SD1L.t83 0.551
R78 SD1L.n69 SD1L.t115 0.551
R79 SD1L.n69 SD1L.t4 0.551
R80 SD1L.n68 SD1L.t68 0.551
R81 SD1L.n68 SD1L.t61 0.551
R82 SD1L.n61 SD1L.t111 0.551
R83 SD1L.n61 SD1L.t100 0.551
R84 SD1L.n60 SD1L.t90 0.551
R85 SD1L.n60 SD1L.t51 0.551
R86 SD1L.n59 SD1L.t11 0.551
R87 SD1L.n59 SD1L.t21 0.551
R88 SD1L.n49 SD1L.t52 0.551
R89 SD1L.n49 SD1L.t33 0.551
R90 SD1L.n50 SD1L.t39 0.551
R91 SD1L.n50 SD1L.t48 0.551
R92 SD1L.n51 SD1L.t62 0.551
R93 SD1L.n51 SD1L.t29 0.551
R94 SD1L.n52 SD1L.t17 0.551
R95 SD1L.n52 SD1L.t94 0.551
R96 SD1L.n53 SD1L.t116 0.551
R97 SD1L.n53 SD1L.t93 0.551
R98 SD1L.n48 SD1L.t58 0.551
R99 SD1L.n48 SD1L.t16 0.551
R100 SD1L.n47 SD1L.t89 0.551
R101 SD1L.n47 SD1L.t84 0.551
R102 SD1L.n46 SD1L.t59 0.551
R103 SD1L.n46 SD1L.t55 0.551
R104 SD1L.n45 SD1L.t14 0.551
R105 SD1L.n45 SD1L.t119 0.551
R106 SD1L.n44 SD1L.t101 0.551
R107 SD1L.n44 SD1L.t99 0.551
R108 SD1L.n54 SD1L.t80 0.551
R109 SD1L.n54 SD1L.t74 0.551
R110 SD1L.n55 SD1L.t73 0.551
R111 SD1L.n55 SD1L.t15 0.551
R112 SD1L.n56 SD1L.t79 0.551
R113 SD1L.n56 SD1L.t30 0.551
R114 SD1L.n57 SD1L.t38 0.551
R115 SD1L.n57 SD1L.t107 0.551
R116 SD1L.n29 SD1L.t47 0.551
R117 SD1L.n29 SD1L.t24 0.551
R118 SD1L.n30 SD1L.t41 0.551
R119 SD1L.n30 SD1L.t110 0.551
R120 SD1L.n31 SD1L.t49 0.551
R121 SD1L.n31 SD1L.t96 0.551
R122 SD1L.n32 SD1L.t67 0.551
R123 SD1L.n32 SD1L.t78 0.551
R124 SD1L.n33 SD1L.t77 0.551
R125 SD1L.n33 SD1L.t114 0.551
R126 SD1L.n34 SD1L.t18 0.551
R127 SD1L.n34 SD1L.t28 0.551
R128 SD1L.n35 SD1L.t35 0.551
R129 SD1L.n35 SD1L.t27 0.551
R130 SD1L.n36 SD1L.t22 0.551
R131 SD1L.n36 SD1L.t98 0.551
R132 SD1L.n37 SD1L.t88 0.551
R133 SD1L.n37 SD1L.t43 0.551
R134 SD1L.n38 SD1L.t106 0.551
R135 SD1L.n38 SD1L.t95 0.551
R136 SD1L.n39 SD1L.t91 0.551
R137 SD1L.n39 SD1L.t82 0.551
R138 SD1L.n40 SD1L.t31 0.551
R139 SD1L.n40 SD1L.t113 0.551
R140 SD1L.n41 SD1L.t8 0.551
R141 SD1L.n41 SD1L.t60 0.551
R142 SD1L.n42 SD1L.t75 0.551
R143 SD1L.n42 SD1L.t20 0.551
R144 SD1L.n43 SD1L.t65 0.551
R145 SD1L.n43 SD1L.t81 0.551
R146 SD1L.n17 SD1L.t63 0.551
R147 SD1L.n17 SD1L.t2 0.551
R148 SD1L.n16 SD1L.t54 0.551
R149 SD1L.n16 SD1L.t6 0.551
R150 SD1L.n15 SD1L.t37 0.551
R151 SD1L.n15 SD1L.t36 0.551
R152 SD1L.n14 SD1L.t108 0.551
R153 SD1L.n14 SD1L.t46 0.551
R154 SD1L.n18 SD1L.t104 0.551
R155 SD1L.n18 SD1L.t26 0.551
R156 SD1L.n19 SD1L.t85 0.551
R157 SD1L.n19 SD1L.t3 0.551
R158 SD1L.n20 SD1L.t7 0.551
R159 SD1L.n20 SD1L.t97 0.551
R160 SD1L.n21 SD1L.t66 0.551
R161 SD1L.n21 SD1L.t76 0.551
R162 SD1L.n22 SD1L.t56 0.551
R163 SD1L.n22 SD1L.t105 0.551
R164 SD1L.n23 SD1L.t50 0.551
R165 SD1L.n23 SD1L.t23 0.551
R166 SD1L.n24 SD1L.t34 0.551
R167 SD1L.n24 SD1L.t32 0.551
R168 SD1L.n25 SD1L.t102 0.551
R169 SD1L.n25 SD1L.t40 0.551
R170 SD1L.n26 SD1L.t86 0.551
R171 SD1L.n26 SD1L.t25 0.551
R172 SD1L.n27 SD1L.t109 0.551
R173 SD1L.n27 SD1L.t103 0.551
R174 SD1L.n28 SD1L.t64 0.551
R175 SD1L.n28 SD1L.t57 0.551
R176 SD1L.n67 SD1L.t0 0.551
R177 SD1L.n67 SD1L.t112 0.551
R178 SD1L.n58 SD1L.n7 0.523
R179 SD1L.n73 SD1L.n1 0.392
R180 SD1L.n74 SD1L.n73 0.099
R181 SD1L.n58 SD1L.n11 0.078
R182 SD1L.n74 SD1L.n9 0.078
R183 SD1L.n73 SD1L.n58 0.07
R184 SD1L.n9 SD1L.n3 0.041
R185 SD1L SD1L.n74 0.04
R186 SD1L.n7 SD1L.n8 0.038
R187 SD1L.n7 SD1L.n6 0.028
R188 SD1L.n10 SD1L.n5 0.028
R189 SD1L.n3 SD1L.n2 0.028
R190 SD1L.n1 SD1L.n0 0.028
R191 SD1L.n11 SD1L.n10 0.022
R192 SD1L.n12 SD1L.n13 0.021
R193 SD1L.n5 SD1L.n4 0.021
R194 SD1L.n1 SD1L.n12 0.019
R195 SD2L.n64 SD2L.t31 1.972
R196 SD2L.n11 SD2L.t69 1.972
R197 SD2L.n78 SD2L.t41 1.963
R198 SD2L.n25 SD2L.t43 1.962
R199 SD2L.n93 SD2L.n92 1.435
R200 SD2L.n37 SD2L.n36 1.435
R201 SD2L.n103 SD2L.n83 1.428
R202 SD2L.n102 SD2L.n84 1.428
R203 SD2L.n101 SD2L.n85 1.428
R204 SD2L.n100 SD2L.n86 1.428
R205 SD2L.n99 SD2L.n87 1.428
R206 SD2L.n96 SD2L.n88 1.428
R207 SD2L.n95 SD2L.n89 1.428
R208 SD2L.n94 SD2L.n90 1.428
R209 SD2L.n93 SD2L.n91 1.428
R210 SD2L.n46 SD2L.n26 1.428
R211 SD2L.n45 SD2L.n27 1.428
R212 SD2L.n44 SD2L.n28 1.428
R213 SD2L.n43 SD2L.n29 1.428
R214 SD2L.n42 SD2L.n30 1.428
R215 SD2L.n41 SD2L.n31 1.428
R216 SD2L.n40 SD2L.n32 1.428
R217 SD2L.n39 SD2L.n33 1.428
R218 SD2L.n38 SD2L.n34 1.428
R219 SD2L.n37 SD2L.n35 1.428
R220 SD2L.n98 SD2L.n97 1.427
R221 SD2L.n74 SD2L.n53 1.414
R222 SD2L.n73 SD2L.n54 1.414
R223 SD2L.n72 SD2L.n55 1.414
R224 SD2L.n71 SD2L.n56 1.414
R225 SD2L.n70 SD2L.n57 1.414
R226 SD2L.n69 SD2L.n58 1.414
R227 SD2L.n68 SD2L.n59 1.414
R228 SD2L.n67 SD2L.n60 1.414
R229 SD2L.n66 SD2L.n61 1.414
R230 SD2L.n65 SD2L.n62 1.414
R231 SD2L.n64 SD2L.n63 1.414
R232 SD2L.n21 SD2L.n0 1.414
R233 SD2L.n20 SD2L.n1 1.414
R234 SD2L.n19 SD2L.n2 1.414
R235 SD2L.n18 SD2L.n3 1.414
R236 SD2L.n17 SD2L.n4 1.414
R237 SD2L.n16 SD2L.n5 1.414
R238 SD2L.n15 SD2L.n6 1.414
R239 SD2L.n14 SD2L.n7 1.414
R240 SD2L.n13 SD2L.n8 1.414
R241 SD2L.n12 SD2L.n9 1.414
R242 SD2L.n11 SD2L.n10 1.414
R243 SD2L.n78 SD2L.n77 1.412
R244 SD2L.n78 SD2L.n76 1.412
R245 SD2L.n78 SD2L.n75 1.412
R246 SD2L.n25 SD2L.n24 1.409
R247 SD2L.n25 SD2L.n23 1.409
R248 SD2L.n25 SD2L.n22 1.409
R249 SD2L.n48 SD2L.n47 1.281
R250 SD2L.n104 SD2L.n82 1.281
R251 SD2L.n52 SD2L.n49 1.28
R252 SD2L.n52 SD2L.n50 1.28
R253 SD2L.n52 SD2L.n51 1.28
R254 SD2L.n105 SD2L.n81 1.28
R255 SD2L.n105 SD2L.n80 1.28
R256 SD2L.n105 SD2L.n79 1.28
R257 SD2L.n83 SD2L.t92 0.551
R258 SD2L.n83 SD2L.t17 0.551
R259 SD2L.n84 SD2L.t19 0.551
R260 SD2L.n84 SD2L.t25 0.551
R261 SD2L.n85 SD2L.t88 0.551
R262 SD2L.n85 SD2L.t94 0.551
R263 SD2L.n86 SD2L.t13 0.551
R264 SD2L.n86 SD2L.t44 0.551
R265 SD2L.n87 SD2L.t49 0.551
R266 SD2L.n87 SD2L.t93 0.551
R267 SD2L.n88 SD2L.t30 0.551
R268 SD2L.n88 SD2L.t81 0.551
R269 SD2L.n89 SD2L.t115 0.551
R270 SD2L.n89 SD2L.t3 0.551
R271 SD2L.n90 SD2L.t28 0.551
R272 SD2L.n90 SD2L.t71 0.551
R273 SD2L.n91 SD2L.t97 0.551
R274 SD2L.n91 SD2L.t106 0.551
R275 SD2L.n92 SD2L.t18 0.551
R276 SD2L.n92 SD2L.t55 0.551
R277 SD2L.n82 SD2L.t20 0.551
R278 SD2L.n82 SD2L.t74 0.551
R279 SD2L.n81 SD2L.t78 0.551
R280 SD2L.n81 SD2L.t33 0.551
R281 SD2L.n80 SD2L.t38 0.551
R282 SD2L.n80 SD2L.t75 0.551
R283 SD2L.n79 SD2L.t2 0.551
R284 SD2L.n79 SD2L.t8 0.551
R285 SD2L.n26 SD2L.t72 0.551
R286 SD2L.n26 SD2L.t117 0.551
R287 SD2L.n27 SD2L.t107 0.551
R288 SD2L.n27 SD2L.t114 0.551
R289 SD2L.n28 SD2L.t58 0.551
R290 SD2L.n28 SD2L.t64 0.551
R291 SD2L.n29 SD2L.t82 0.551
R292 SD2L.n29 SD2L.t1 0.551
R293 SD2L.n30 SD2L.t109 0.551
R294 SD2L.n30 SD2L.t32 0.551
R295 SD2L.n31 SD2L.t61 0.551
R296 SD2L.n31 SD2L.t101 0.551
R297 SD2L.n32 SD2L.t108 0.551
R298 SD2L.n32 SD2L.t29 0.551
R299 SD2L.n33 SD2L.t59 0.551
R300 SD2L.n33 SD2L.t65 0.551
R301 SD2L.n34 SD2L.t89 0.551
R302 SD2L.n34 SD2L.t12 0.551
R303 SD2L.n35 SD2L.t54 0.551
R304 SD2L.n35 SD2L.t63 0.551
R305 SD2L.n36 SD2L.t80 0.551
R306 SD2L.n36 SD2L.t7 0.551
R307 SD2L.n47 SD2L.t4 0.551
R308 SD2L.n47 SD2L.t35 0.551
R309 SD2L.n49 SD2L.t39 0.551
R310 SD2L.n49 SD2L.t0 0.551
R311 SD2L.n50 SD2L.t5 0.551
R312 SD2L.n50 SD2L.t51 0.551
R313 SD2L.n51 SD2L.t95 0.551
R314 SD2L.n51 SD2L.t85 0.551
R315 SD2L.n53 SD2L.t9 0.551
R316 SD2L.n53 SD2L.t102 0.551
R317 SD2L.n54 SD2L.t105 0.551
R318 SD2L.n54 SD2L.t119 0.551
R319 SD2L.n55 SD2L.t26 0.551
R320 SD2L.n55 SD2L.t10 0.551
R321 SD2L.n56 SD2L.t45 0.551
R322 SD2L.n56 SD2L.t52 0.551
R323 SD2L.n57 SD2L.t56 0.551
R324 SD2L.n57 SD2L.t66 0.551
R325 SD2L.n58 SD2L.t96 0.551
R326 SD2L.n58 SD2L.t46 0.551
R327 SD2L.n59 SD2L.t110 0.551
R328 SD2L.n59 SD2L.t87 0.551
R329 SD2L.n60 SD2L.t90 0.551
R330 SD2L.n60 SD2L.t99 0.551
R331 SD2L.n61 SD2L.t15 0.551
R332 SD2L.n61 SD2L.t116 0.551
R333 SD2L.n62 SD2L.t22 0.551
R334 SD2L.n62 SD2L.t34 0.551
R335 SD2L.n63 SD2L.t40 0.551
R336 SD2L.n63 SD2L.t50 0.551
R337 SD2L.n75 SD2L.t112 0.551
R338 SD2L.n75 SD2L.t84 0.551
R339 SD2L.n76 SD2L.t73 0.551
R340 SD2L.n76 SD2L.t48 0.551
R341 SD2L.n77 SD2L.t60 0.551
R342 SD2L.n77 SD2L.t68 0.551
R343 SD2L.n24 SD2L.t62 0.551
R344 SD2L.n24 SD2L.t70 0.551
R345 SD2L.n23 SD2L.t103 0.551
R346 SD2L.n23 SD2L.t79 0.551
R347 SD2L.n22 SD2L.t113 0.551
R348 SD2L.n22 SD2L.t86 0.551
R349 SD2L.n0 SD2L.t11 0.551
R350 SD2L.n0 SD2L.t104 0.551
R351 SD2L.n1 SD2L.t14 0.551
R352 SD2L.n1 SD2L.t24 0.551
R353 SD2L.n2 SD2L.t27 0.551
R354 SD2L.n2 SD2L.t37 0.551
R355 SD2L.n3 SD2L.t47 0.551
R356 SD2L.n3 SD2L.t57 0.551
R357 SD2L.n4 SD2L.t83 0.551
R358 SD2L.n4 SD2L.t67 0.551
R359 SD2L.n5 SD2L.t98 0.551
R360 SD2L.n5 SD2L.t77 0.551
R361 SD2L.n6 SD2L.t111 0.551
R362 SD2L.n6 SD2L.t91 0.551
R363 SD2L.n7 SD2L.t6 0.551
R364 SD2L.n7 SD2L.t100 0.551
R365 SD2L.n8 SD2L.t16 0.551
R366 SD2L.n8 SD2L.t21 0.551
R367 SD2L.n9 SD2L.t23 0.551
R368 SD2L.n9 SD2L.t36 0.551
R369 SD2L.n10 SD2L.t76 0.551
R370 SD2L.n10 SD2L.t53 0.551
R371 SD2L.n97 SD2L.t118 0.551
R372 SD2L.n97 SD2L.t42 0.551
R373 SD2L.n106 SD2L.n78 0.39
R374 SD2L.n108 SD2L.n25 0.39
R375 SD2L.n106 SD2L.n105 0.366
R376 SD2L.n107 SD2L.n52 0.265
R377 SD2L.n107 SD2L.n106 0.101
R378 SD2L.n108 SD2L.n107 0.097
R379 SD2L SD2L.n108 0.01
R380 SD2L.n48 SD2L.n46 0.007
R381 SD2L.n104 SD2L.n103 0.007
R382 SD2L.n38 SD2L.n37 0.007
R383 SD2L.n39 SD2L.n38 0.007
R384 SD2L.n40 SD2L.n39 0.007
R385 SD2L.n41 SD2L.n40 0.007
R386 SD2L.n42 SD2L.n41 0.007
R387 SD2L.n43 SD2L.n42 0.007
R388 SD2L.n44 SD2L.n43 0.007
R389 SD2L.n45 SD2L.n44 0.007
R390 SD2L.n46 SD2L.n45 0.007
R391 SD2L.n65 SD2L.n64 0.007
R392 SD2L.n66 SD2L.n65 0.007
R393 SD2L.n67 SD2L.n66 0.007
R394 SD2L.n68 SD2L.n67 0.007
R395 SD2L.n69 SD2L.n68 0.007
R396 SD2L.n70 SD2L.n69 0.007
R397 SD2L.n71 SD2L.n70 0.007
R398 SD2L.n72 SD2L.n71 0.007
R399 SD2L.n73 SD2L.n72 0.007
R400 SD2L.n74 SD2L.n73 0.007
R401 SD2L.n12 SD2L.n11 0.007
R402 SD2L.n13 SD2L.n12 0.007
R403 SD2L.n14 SD2L.n13 0.007
R404 SD2L.n15 SD2L.n14 0.007
R405 SD2L.n16 SD2L.n15 0.007
R406 SD2L.n17 SD2L.n16 0.007
R407 SD2L.n18 SD2L.n17 0.007
R408 SD2L.n19 SD2L.n18 0.007
R409 SD2L.n20 SD2L.n19 0.007
R410 SD2L.n21 SD2L.n20 0.007
R411 SD2L.n94 SD2L.n93 0.007
R412 SD2L.n95 SD2L.n94 0.007
R413 SD2L.n96 SD2L.n95 0.007
R414 SD2L.n98 SD2L.n96 0.007
R415 SD2L.n99 SD2L.n98 0.007
R416 SD2L.n100 SD2L.n99 0.007
R417 SD2L.n101 SD2L.n100 0.007
R418 SD2L.n102 SD2L.n101 0.007
R419 SD2L.n103 SD2L.n102 0.007
R420 SD2L.n78 SD2L.n74 0.004
R421 SD2L.n25 SD2L.n21 0.004
R422 SD2L.n52 SD2L.n48 0.001
R423 SD2L.n105 SD2L.n104 0.001
R424 SD1R.n5 SD1R.t67 1.972
R425 SD1R.n2 SD1R.t20 1.972
R426 SD1R.n14 SD1R.t4 1.963
R427 SD1R.n15 SD1R.t61 1.963
R428 SD1R.n0 SD1R.n72 1.435
R429 SD1R.n8 SD1R.n42 1.435
R430 SD1R.n13 SD1R.n63 1.428
R431 SD1R.n13 SD1R.n64 1.428
R432 SD1R.n12 SD1R.n65 1.428
R433 SD1R.n12 SD1R.n66 1.428
R434 SD1R.n1 SD1R.n67 1.428
R435 SD1R.n1 SD1R.n68 1.428
R436 SD1R.n1 SD1R.n69 1.428
R437 SD1R.n0 SD1R.n70 1.428
R438 SD1R.n0 SD1R.n71 1.428
R439 SD1R.n11 SD1R.n32 1.428
R440 SD1R.n11 SD1R.n33 1.428
R441 SD1R.n10 SD1R.n34 1.428
R442 SD1R.n10 SD1R.n35 1.428
R443 SD1R.n9 SD1R.n36 1.428
R444 SD1R.n9 SD1R.n37 1.428
R445 SD1R.n9 SD1R.n38 1.428
R446 SD1R.n9 SD1R.n39 1.428
R447 SD1R.n8 SD1R.n40 1.428
R448 SD1R.n8 SD1R.n41 1.428
R449 SD1R.n1 SD1R.n73 1.427
R450 SD1R.n14 SD1R.n16 1.414
R451 SD1R.n7 SD1R.n17 1.414
R452 SD1R.n7 SD1R.n18 1.414
R453 SD1R.n7 SD1R.n19 1.414
R454 SD1R.n7 SD1R.n20 1.414
R455 SD1R.n6 SD1R.n21 1.414
R456 SD1R.n6 SD1R.n22 1.414
R457 SD1R.n6 SD1R.n23 1.414
R458 SD1R.n6 SD1R.n24 1.414
R459 SD1R.n5 SD1R.n25 1.414
R460 SD1R.n5 SD1R.n26 1.414
R461 SD1R.n15 SD1R.n45 1.414
R462 SD1R.n4 SD1R.n46 1.414
R463 SD1R.n4 SD1R.n47 1.414
R464 SD1R.n4 SD1R.n48 1.414
R465 SD1R.n4 SD1R.n49 1.414
R466 SD1R.n3 SD1R.n50 1.414
R467 SD1R.n3 SD1R.n51 1.414
R468 SD1R.n3 SD1R.n52 1.414
R469 SD1R.n3 SD1R.n53 1.414
R470 SD1R.n2 SD1R.n54 1.414
R471 SD1R.n2 SD1R.n55 1.414
R472 SD1R.n14 SD1R.n29 1.412
R473 SD1R.n14 SD1R.n28 1.412
R474 SD1R.n14 SD1R.n27 1.412
R475 SD1R.n15 SD1R.n58 1.412
R476 SD1R.n15 SD1R.n57 1.412
R477 SD1R.n15 SD1R.n56 1.412
R478 SD1R.n13 SD1R.n74 1.282
R479 SD1R.n13 SD1R.n62 1.28
R480 SD1R.n13 SD1R.n75 1.28
R481 SD1R.n13 SD1R.n61 1.28
R482 SD1R.n11 SD1R.n44 1.279
R483 SD1R.n11 SD1R.n30 1.279
R484 SD1R.n11 SD1R.n31 1.278
R485 SD1R.n11 SD1R.n43 1.278
R486 SD1R.n63 SD1R.t87 0.551
R487 SD1R.n63 SD1R.t50 0.551
R488 SD1R.n64 SD1R.t32 0.551
R489 SD1R.n64 SD1R.t22 0.551
R490 SD1R.n65 SD1R.t55 0.551
R491 SD1R.n65 SD1R.t117 0.551
R492 SD1R.n66 SD1R.t97 0.551
R493 SD1R.n66 SD1R.t44 0.551
R494 SD1R.n67 SD1R.t58 0.551
R495 SD1R.n67 SD1R.t105 0.551
R496 SD1R.n68 SD1R.t99 0.551
R497 SD1R.n68 SD1R.t72 0.551
R498 SD1R.n69 SD1R.t64 0.551
R499 SD1R.n69 SD1R.t68 0.551
R500 SD1R.n70 SD1R.t25 0.551
R501 SD1R.n70 SD1R.t80 0.551
R502 SD1R.n71 SD1R.t62 0.551
R503 SD1R.n71 SD1R.t13 0.551
R504 SD1R.n72 SD1R.t42 0.551
R505 SD1R.n72 SD1R.t100 0.551
R506 SD1R.n74 SD1R.t7 0.551
R507 SD1R.n74 SD1R.t6 0.551
R508 SD1R.n62 SD1R.t73 0.551
R509 SD1R.n62 SD1R.t14 0.551
R510 SD1R.n75 SD1R.t82 0.551
R511 SD1R.n75 SD1R.t43 0.551
R512 SD1R.n61 SD1R.t114 0.551
R513 SD1R.n61 SD1R.t63 0.551
R514 SD1R.n31 SD1R.t102 0.551
R515 SD1R.n31 SD1R.t16 0.551
R516 SD1R.n44 SD1R.t18 0.551
R517 SD1R.n44 SD1R.t111 0.551
R518 SD1R.n30 SD1R.t47 0.551
R519 SD1R.n30 SD1R.t45 0.551
R520 SD1R.n32 SD1R.t10 0.551
R521 SD1R.n32 SD1R.t74 0.551
R522 SD1R.n33 SD1R.t112 0.551
R523 SD1R.n33 SD1R.t106 0.551
R524 SD1R.n34 SD1R.t34 0.551
R525 SD1R.n34 SD1R.t113 0.551
R526 SD1R.n35 SD1R.t46 0.551
R527 SD1R.n35 SD1R.t69 0.551
R528 SD1R.n36 SD1R.t27 0.551
R529 SD1R.n36 SD1R.t81 0.551
R530 SD1R.n37 SD1R.t65 0.551
R531 SD1R.n37 SD1R.t38 0.551
R532 SD1R.n38 SD1R.t115 0.551
R533 SD1R.n38 SD1R.t35 0.551
R534 SD1R.n39 SD1R.t75 0.551
R535 SD1R.n39 SD1R.t37 0.551
R536 SD1R.n40 SD1R.t84 0.551
R537 SD1R.n40 SD1R.t76 0.551
R538 SD1R.n41 SD1R.t24 0.551
R539 SD1R.n41 SD1R.t29 0.551
R540 SD1R.n42 SD1R.t89 0.551
R541 SD1R.n42 SD1R.t28 0.551
R542 SD1R.n43 SD1R.t77 0.551
R543 SD1R.n43 SD1R.t3 0.551
R544 SD1R.n16 SD1R.t93 0.551
R545 SD1R.n16 SD1R.t91 0.551
R546 SD1R.n17 SD1R.t85 0.551
R547 SD1R.n17 SD1R.t88 0.551
R548 SD1R.n18 SD1R.t78 0.551
R549 SD1R.n18 SD1R.t11 0.551
R550 SD1R.n19 SD1R.t49 0.551
R551 SD1R.n19 SD1R.t66 0.551
R552 SD1R.n20 SD1R.t116 0.551
R553 SD1R.n20 SD1R.t30 0.551
R554 SD1R.n21 SD1R.t19 0.551
R555 SD1R.n21 SD1R.t119 0.551
R556 SD1R.n22 SD1R.t110 0.551
R557 SD1R.n22 SD1R.t41 0.551
R558 SD1R.n23 SD1R.t39 0.551
R559 SD1R.n23 SD1R.t21 0.551
R560 SD1R.n24 SD1R.t9 0.551
R561 SD1R.n24 SD1R.t33 0.551
R562 SD1R.n25 SD1R.t109 0.551
R563 SD1R.n25 SD1R.t101 0.551
R564 SD1R.n26 SD1R.t8 0.551
R565 SD1R.n26 SD1R.t51 0.551
R566 SD1R.n27 SD1R.t98 0.551
R567 SD1R.n27 SD1R.t52 0.551
R568 SD1R.n28 SD1R.t70 0.551
R569 SD1R.n28 SD1R.t12 0.551
R570 SD1R.n29 SD1R.t5 0.551
R571 SD1R.n29 SD1R.t2 0.551
R572 SD1R.n45 SD1R.t31 0.551
R573 SD1R.n45 SD1R.t59 0.551
R574 SD1R.n46 SD1R.t56 0.551
R575 SD1R.n46 SD1R.t79 0.551
R576 SD1R.n47 SD1R.t86 0.551
R577 SD1R.n47 SD1R.t95 0.551
R578 SD1R.n48 SD1R.t23 0.551
R579 SD1R.n48 SD1R.t108 0.551
R580 SD1R.n49 SD1R.t83 0.551
R581 SD1R.n49 SD1R.t17 0.551
R582 SD1R.n50 SD1R.t103 0.551
R583 SD1R.n50 SD1R.t36 0.551
R584 SD1R.n51 SD1R.t60 0.551
R585 SD1R.n51 SD1R.t118 0.551
R586 SD1R.n52 SD1R.t107 0.551
R587 SD1R.n52 SD1R.t54 0.551
R588 SD1R.n53 SD1R.t71 0.551
R589 SD1R.n53 SD1R.t48 0.551
R590 SD1R.n54 SD1R.t96 0.551
R591 SD1R.n54 SD1R.t1 0.551
R592 SD1R.n55 SD1R.t90 0.551
R593 SD1R.n55 SD1R.t92 0.551
R594 SD1R.n56 SD1R.t104 0.551
R595 SD1R.n56 SD1R.t40 0.551
R596 SD1R.n57 SD1R.t26 0.551
R597 SD1R.n57 SD1R.t53 0.551
R598 SD1R.n58 SD1R.t57 0.551
R599 SD1R.n58 SD1R.t15 0.551
R600 SD1R.n73 SD1R.t0 0.551
R601 SD1R.n73 SD1R.t94 0.551
R602 SD1R.n59 SD1R.n15 0.525
R603 SD1R.n60 SD1R.n14 0.485
R604 SD1R.n59 SD1R.n11 0.172
R605 SD1R.n76 SD1R.n13 0.169
R606 SD1R.n60 SD1R.n59 0.162
R607 SD1R.n76 SD1R.n60 0.04
R608 SD1R SD1R.n76 0.037
R609 SD1R.n10 SD1R.n9 0.028
R610 SD1R.n7 SD1R.n6 0.028
R611 SD1R.n6 SD1R.n5 0.028
R612 SD1R.n4 SD1R.n3 0.028
R613 SD1R.n3 SD1R.n2 0.028
R614 SD1R.n12 SD1R.n1 0.028
R615 SD1R.n11 SD1R.n10 0.027
R616 SD1R.n13 SD1R.n12 0.025
R617 SD1R.n1 SD1R.n0 0.021
R618 SD1R.n9 SD1R.n8 0.021
R619 SD1R.n15 SD1R.n4 0.02
R620 SD1R.n14 SD1R.n7 0.02
R621 SD2R.n92 SD2R.t50 1.972
R622 SD2R.n36 SD2R.t94 1.972
R623 SD2R.n104 SD2R.t70 1.963
R624 SD2R.n51 SD2R.t116 1.96
R625 SD2R.n16 SD2R.n15 1.435
R626 SD2R.n6 SD2R.n5 1.435
R627 SD2R.n68 SD2R.n67 1.435
R628 SD2R.n58 SD2R.n57 1.435
R629 SD2R.n19 SD2R.n11 1.428
R630 SD2R.n18 SD2R.n12 1.428
R631 SD2R.n17 SD2R.n13 1.428
R632 SD2R.n16 SD2R.n14 1.428
R633 SD2R.n6 SD2R.n4 1.428
R634 SD2R.n7 SD2R.n3 1.428
R635 SD2R.n8 SD2R.n2 1.428
R636 SD2R.n9 SD2R.n1 1.428
R637 SD2R.n10 SD2R.n0 1.428
R638 SD2R.n71 SD2R.n63 1.428
R639 SD2R.n70 SD2R.n64 1.428
R640 SD2R.n69 SD2R.n65 1.428
R641 SD2R.n68 SD2R.n66 1.428
R642 SD2R.n58 SD2R.n56 1.428
R643 SD2R.n59 SD2R.n55 1.428
R644 SD2R.n60 SD2R.n54 1.428
R645 SD2R.n61 SD2R.n53 1.428
R646 SD2R.n62 SD2R.n52 1.428
R647 SD2R.n103 SD2R.n82 1.414
R648 SD2R.n102 SD2R.n83 1.414
R649 SD2R.n101 SD2R.n84 1.414
R650 SD2R.n100 SD2R.n85 1.414
R651 SD2R.n99 SD2R.n86 1.414
R652 SD2R.n98 SD2R.n87 1.414
R653 SD2R.n97 SD2R.n88 1.414
R654 SD2R.n96 SD2R.n89 1.414
R655 SD2R.n93 SD2R.n90 1.414
R656 SD2R.n92 SD2R.n91 1.414
R657 SD2R.n36 SD2R.n35 1.414
R658 SD2R.n37 SD2R.n34 1.414
R659 SD2R.n38 SD2R.n33 1.414
R660 SD2R.n39 SD2R.n32 1.414
R661 SD2R.n40 SD2R.n31 1.414
R662 SD2R.n41 SD2R.n30 1.414
R663 SD2R.n42 SD2R.n29 1.414
R664 SD2R.n43 SD2R.n28 1.414
R665 SD2R.n44 SD2R.n27 1.414
R666 SD2R.n45 SD2R.n26 1.414
R667 SD2R.n46 SD2R.n25 1.414
R668 SD2R.n95 SD2R.n94 1.413
R669 SD2R.n104 SD2R.n79 1.412
R670 SD2R.n104 SD2R.n80 1.412
R671 SD2R.n104 SD2R.n81 1.412
R672 SD2R.n48 SD2R.n47 1.41
R673 SD2R.n51 SD2R.n49 1.409
R674 SD2R.n51 SD2R.n50 1.409
R675 SD2R.n24 SD2R.n20 1.28
R676 SD2R.n24 SD2R.n21 1.28
R677 SD2R.n24 SD2R.n22 1.28
R678 SD2R.n24 SD2R.n23 1.28
R679 SD2R.n76 SD2R.n72 1.28
R680 SD2R.n76 SD2R.n73 1.28
R681 SD2R.n76 SD2R.n74 1.28
R682 SD2R.n76 SD2R.n75 1.28
R683 SD2R.n82 SD2R.t7 0.551
R684 SD2R.n82 SD2R.t106 0.551
R685 SD2R.n83 SD2R.t115 0.551
R686 SD2R.n83 SD2R.t97 0.551
R687 SD2R.n84 SD2R.t103 0.551
R688 SD2R.n84 SD2R.t84 0.551
R689 SD2R.n85 SD2R.t95 0.551
R690 SD2R.n85 SD2R.t68 0.551
R691 SD2R.n86 SD2R.t53 0.551
R692 SD2R.n86 SD2R.t58 0.551
R693 SD2R.n87 SD2R.t39 0.551
R694 SD2R.n87 SD2R.t47 0.551
R695 SD2R.n88 SD2R.t21 0.551
R696 SD2R.n88 SD2R.t1 0.551
R697 SD2R.n89 SD2R.t9 0.551
R698 SD2R.n89 SD2R.t109 0.551
R699 SD2R.n90 SD2R.t107 0.551
R700 SD2R.n90 SD2R.t87 0.551
R701 SD2R.n91 SD2R.t62 0.551
R702 SD2R.n91 SD2R.t71 0.551
R703 SD2R.n81 SD2R.t51 0.551
R704 SD2R.n81 SD2R.t56 0.551
R705 SD2R.n80 SD2R.t37 0.551
R706 SD2R.n80 SD2R.t46 0.551
R707 SD2R.n79 SD2R.t25 0.551
R708 SD2R.n79 SD2R.t34 0.551
R709 SD2R.n35 SD2R.t14 0.551
R710 SD2R.n35 SD2R.t24 0.551
R711 SD2R.n34 SD2R.t31 0.551
R712 SD2R.n34 SD2R.t4 0.551
R713 SD2R.n33 SD2R.t43 0.551
R714 SD2R.n33 SD2R.t18 0.551
R715 SD2R.n32 SD2R.t88 0.551
R716 SD2R.n32 SD2R.t61 0.551
R717 SD2R.n31 SD2R.t65 0.551
R718 SD2R.n31 SD2R.t77 0.551
R719 SD2R.n30 SD2R.t79 0.551
R720 SD2R.n30 SD2R.t89 0.551
R721 SD2R.n29 SD2R.t3 0.551
R722 SD2R.n29 SD2R.t100 0.551
R723 SD2R.n28 SD2R.t17 0.551
R724 SD2R.n28 SD2R.t26 0.551
R725 SD2R.n27 SD2R.t32 0.551
R726 SD2R.n27 SD2R.t6 0.551
R727 SD2R.n26 SD2R.t72 0.551
R728 SD2R.n26 SD2R.t23 0.551
R729 SD2R.n25 SD2R.t55 0.551
R730 SD2R.n25 SD2R.t63 0.551
R731 SD2R.n47 SD2R.t69 0.551
R732 SD2R.n47 SD2R.t78 0.551
R733 SD2R.n49 SD2R.t110 0.551
R734 SD2R.n49 SD2R.t91 0.551
R735 SD2R.n50 SD2R.t2 0.551
R736 SD2R.n50 SD2R.t10 0.551
R737 SD2R.n11 SD2R.t44 0.551
R738 SD2R.n11 SD2R.t90 0.551
R739 SD2R.n12 SD2R.t108 0.551
R740 SD2R.n12 SD2R.t114 0.551
R741 SD2R.n13 SD2R.t40 0.551
R742 SD2R.n13 SD2R.t76 0.551
R743 SD2R.n14 SD2R.t104 0.551
R744 SD2R.n14 SD2R.t112 0.551
R745 SD2R.n15 SD2R.t12 0.551
R746 SD2R.n15 SD2R.t60 0.551
R747 SD2R.n5 SD2R.t5 0.551
R748 SD2R.n5 SD2R.t11 0.551
R749 SD2R.n4 SD2R.t35 0.551
R750 SD2R.n4 SD2R.t82 0.551
R751 SD2R.n3 SD2R.t86 0.551
R752 SD2R.n3 SD2R.t30 0.551
R753 SD2R.n2 SD2R.t33 0.551
R754 SD2R.n2 SD2R.t80 0.551
R755 SD2R.n1 SD2R.t99 0.551
R756 SD2R.n1 SD2R.t29 0.551
R757 SD2R.n0 SD2R.t19 0.551
R758 SD2R.n0 SD2R.t22 0.551
R759 SD2R.n20 SD2R.t0 0.551
R760 SD2R.n20 SD2R.t52 0.551
R761 SD2R.n21 SD2R.t45 0.551
R762 SD2R.n21 SD2R.t93 0.551
R763 SD2R.n22 SD2R.t15 0.551
R764 SD2R.n22 SD2R.t54 0.551
R765 SD2R.n23 SD2R.t98 0.551
R766 SD2R.n23 SD2R.t101 0.551
R767 SD2R.n63 SD2R.t74 0.551
R768 SD2R.n63 SD2R.t119 0.551
R769 SD2R.n64 SD2R.t36 0.551
R770 SD2R.n64 SD2R.t41 0.551
R771 SD2R.n65 SD2R.t73 0.551
R772 SD2R.n65 SD2R.t105 0.551
R773 SD2R.n66 SD2R.t20 0.551
R774 SD2R.n66 SD2R.t27 0.551
R775 SD2R.n67 SD2R.t59 0.551
R776 SD2R.n67 SD2R.t102 0.551
R777 SD2R.n57 SD2R.t42 0.551
R778 SD2R.n57 SD2R.t48 0.551
R779 SD2R.n56 SD2R.t81 0.551
R780 SD2R.n56 SD2R.t113 0.551
R781 SD2R.n55 SD2R.t117 0.551
R782 SD2R.n55 SD2R.t75 0.551
R783 SD2R.n54 SD2R.t66 0.551
R784 SD2R.n54 SD2R.t111 0.551
R785 SD2R.n53 SD2R.t28 0.551
R786 SD2R.n53 SD2R.t57 0.551
R787 SD2R.n52 SD2R.t64 0.551
R788 SD2R.n52 SD2R.t67 0.551
R789 SD2R.n72 SD2R.t38 0.551
R790 SD2R.n72 SD2R.t83 0.551
R791 SD2R.n73 SD2R.t92 0.551
R792 SD2R.n73 SD2R.t13 0.551
R793 SD2R.n74 SD2R.t49 0.551
R794 SD2R.n74 SD2R.t85 0.551
R795 SD2R.n75 SD2R.t8 0.551
R796 SD2R.n75 SD2R.t16 0.551
R797 SD2R.n94 SD2R.t118 0.551
R798 SD2R.n94 SD2R.t96 0.551
R799 SD2R.n77 SD2R.n76 0.303
R800 SD2R.n77 SD2R.n51 0.296
R801 SD2R.n105 SD2R.n104 0.296
R802 SD2R.n78 SD2R.n24 0.171
R803 SD2R.n105 SD2R.n78 0.099
R804 SD2R.n78 SD2R.n77 0.07
R805 SD2R SD2R.n105 0.042
R806 SD2R.n48 SD2R.n46 0.007
R807 SD2R.n46 SD2R.n45 0.007
R808 SD2R.n45 SD2R.n44 0.007
R809 SD2R.n44 SD2R.n43 0.007
R810 SD2R.n43 SD2R.n42 0.007
R811 SD2R.n42 SD2R.n41 0.007
R812 SD2R.n41 SD2R.n40 0.007
R813 SD2R.n40 SD2R.n39 0.007
R814 SD2R.n39 SD2R.n38 0.007
R815 SD2R.n38 SD2R.n37 0.007
R816 SD2R.n37 SD2R.n36 0.007
R817 SD2R.n17 SD2R.n16 0.007
R818 SD2R.n18 SD2R.n17 0.007
R819 SD2R.n19 SD2R.n18 0.007
R820 SD2R.n10 SD2R.n9 0.007
R821 SD2R.n9 SD2R.n8 0.007
R822 SD2R.n8 SD2R.n7 0.007
R823 SD2R.n7 SD2R.n6 0.007
R824 SD2R.n69 SD2R.n68 0.007
R825 SD2R.n70 SD2R.n69 0.007
R826 SD2R.n71 SD2R.n70 0.007
R827 SD2R.n62 SD2R.n61 0.007
R828 SD2R.n61 SD2R.n60 0.007
R829 SD2R.n60 SD2R.n59 0.007
R830 SD2R.n59 SD2R.n58 0.007
R831 SD2R.n103 SD2R.n102 0.007
R832 SD2R.n102 SD2R.n101 0.007
R833 SD2R.n101 SD2R.n100 0.007
R834 SD2R.n100 SD2R.n99 0.007
R835 SD2R.n99 SD2R.n98 0.007
R836 SD2R.n98 SD2R.n97 0.007
R837 SD2R.n97 SD2R.n96 0.007
R838 SD2R.n96 SD2R.n95 0.007
R839 SD2R.n95 SD2R.n93 0.007
R840 SD2R.n93 SD2R.n92 0.007
R841 SD2R.n104 SD2R.n103 0.006
R842 SD2R.n24 SD2R.n19 0.005
R843 SD2R.n76 SD2R.n71 0.005
R844 SD2R.n24 SD2R.n10 0.004
R845 SD2R.n76 SD2R.n62 0.004
R846 SD2R.n51 SD2R.n48 0.001
C16 m4_11500_n11600# SUB 1.79fF
C17 SD1R SUB 94.98fF
C18 SD2R SUB 82.48fF
C19 GR SUB 99.81fF $ **FLOATING
C20 SD1L SUB 73.54fF
C21 SD2L SUB 69.08fF
C22 GL SUB 100.76fF $ **FLOATING
C23 SD2R.n0 SUB 3.93fF
C24 SD2R.n1 SUB 3.93fF
C25 SD2R.n2 SUB 3.93fF
C26 SD2R.n3 SUB 3.93fF
C27 SD2R.n4 SUB 3.93fF
C28 SD2R.n5 SUB 3.96fF
C29 SD2R.n6 SUB 10.94fF
C30 SD2R.n7 SUB 4.68fF
C31 SD2R.n8 SUB 4.68fF
C32 SD2R.n9 SUB 4.68fF
C33 SD2R.n10 SUB 4.00fF
C34 SD2R.n11 SUB 3.93fF
C35 SD2R.n12 SUB 3.93fF
C36 SD2R.n13 SUB 3.93fF
C37 SD2R.n14 SUB 3.93fF
C38 SD2R.n15 SUB 3.96fF
C39 SD2R.n16 SUB 10.98fF
C40 SD2R.n17 SUB 4.68fF
C41 SD2R.n18 SUB 4.68fF
C42 SD2R.n19 SUB 4.37fF
C43 SD2R.n20 SUB 3.91fF
C44 SD2R.n21 SUB 3.91fF
C45 SD2R.n22 SUB 3.91fF
C46 SD2R.n23 SUB 3.91fF
C47 SD2R.n24 SUB 46.79fF
C48 SD2R.n25 SUB 3.93fF
C49 SD2R.n26 SUB 3.93fF
C50 SD2R.n27 SUB 3.93fF
C51 SD2R.n28 SUB 3.93fF
C52 SD2R.n29 SUB 3.93fF
C53 SD2R.n30 SUB 3.93fF
C54 SD2R.n31 SUB 3.93fF
C55 SD2R.n32 SUB 3.93fF
C56 SD2R.n33 SUB 3.93fF
C57 SD2R.n34 SUB 3.93fF
C58 SD2R.n35 SUB 3.93fF
C59 SD2R.t94 SUB 3.56fF $ **FLOATING
C60 SD2R.n36 SUB 10.66fF
C61 SD2R.n37 SUB 4.68fF
C62 SD2R.n38 SUB 4.68fF
C63 SD2R.n39 SUB 4.68fF
C64 SD2R.n40 SUB 4.68fF
C65 SD2R.n41 SUB 4.68fF
C66 SD2R.n42 SUB 4.68fF
C67 SD2R.n43 SUB 4.68fF
C68 SD2R.n44 SUB 4.68fF
C69 SD2R.n45 SUB 4.68fF
C70 SD2R.n46 SUB 4.83fF
C71 SD2R.n47 SUB 3.93fF
C72 SD2R.n48 SUB 3.79fF
C73 SD2R.n49 SUB 3.93fF
C74 SD2R.n50 SUB 3.93fF
C75 SD2R.t116 SUB 3.54fF $ **FLOATING
C76 SD2R.n51 SUB 59.30fF
C77 SD2R.n52 SUB 3.93fF
C78 SD2R.n53 SUB 3.93fF
C79 SD2R.n54 SUB 3.93fF
C80 SD2R.n55 SUB 3.93fF
C81 SD2R.n56 SUB 3.93fF
C82 SD2R.n57 SUB 3.96fF
C83 SD2R.n58 SUB 10.94fF
C84 SD2R.n59 SUB 4.68fF
C85 SD2R.n60 SUB 4.68fF
C86 SD2R.n61 SUB 4.68fF
C87 SD2R.n62 SUB 4.00fF
C88 SD2R.n63 SUB 3.93fF
C89 SD2R.n64 SUB 3.93fF
C90 SD2R.n65 SUB 3.93fF
C91 SD2R.n66 SUB 3.93fF
C92 SD2R.n67 SUB 3.96fF
C93 SD2R.n68 SUB 10.98fF
C94 SD2R.n69 SUB 4.68fF
C95 SD2R.n70 SUB 4.68fF
C96 SD2R.n71 SUB 4.37fF
C97 SD2R.n72 SUB 3.91fF
C98 SD2R.n73 SUB 3.91fF
C99 SD2R.n74 SUB 3.91fF
C100 SD2R.n75 SUB 3.91fF
C101 SD2R.n76 SUB 76.32fF
C102 SD2R.n77 SUB 132.84fF
C103 SD2R.n78 SUB 71.44fF
C104 SD2R.n79 SUB 3.93fF
C105 SD2R.n80 SUB 3.93fF
C106 SD2R.n81 SUB 3.93fF
C107 SD2R.t70 SUB 3.54fF $ **FLOATING
C108 SD2R.n82 SUB 3.93fF
C109 SD2R.n83 SUB 3.93fF
C110 SD2R.n84 SUB 3.93fF
C111 SD2R.n85 SUB 3.93fF
C112 SD2R.n86 SUB 3.93fF
C113 SD2R.n87 SUB 3.93fF
C114 SD2R.n88 SUB 3.93fF
C115 SD2R.n89 SUB 3.93fF
C116 SD2R.n90 SUB 3.93fF
C117 SD2R.n91 SUB 3.93fF
C118 SD2R.t50 SUB 3.56fF $ **FLOATING
C119 SD2R.n92 SUB 10.66fF
C120 SD2R.n93 SUB 4.68fF
C121 SD2R.n94 SUB 3.93fF
C122 SD2R.n95 SUB 4.68fF
C123 SD2R.n96 SUB 4.68fF
C124 SD2R.n97 SUB 4.68fF
C125 SD2R.n98 SUB 4.68fF
C126 SD2R.n99 SUB 4.68fF
C127 SD2R.n100 SUB 4.68fF
C128 SD2R.n101 SUB 4.68fF
C129 SD2R.n102 SUB 4.68fF
C130 SD2R.n103 SUB 4.64fF
C131 SD2R.n104 SUB 63.27fF
C132 SD2R.n105 SUB 106.32fF
C133 SD1R.n0 SUB 15.36fF
C134 SD1R.n1 SUB 18.37fF
C135 SD1R.n2 SUB 15.06fF
C136 SD1R.n3 SUB 18.38fF
C137 SD1R.n4 SUB 18.38fF
C138 SD1R.n5 SUB 15.06fF
C139 SD1R.n6 SUB 18.38fF
C140 SD1R.n7 SUB 18.38fF
C141 SD1R.n8 SUB 15.36fF
C142 SD1R.n9 SUB 18.37fF
C143 SD1R.n10 SUB 9.19fF
C144 SD1R.n11 SUB 55.93fF
C145 SD1R.n12 SUB 9.19fF
C146 SD1R.n13 SUB 56.21fF
C147 SD1R.n14 SUB 87.68fF
C148 SD1R.n15 SUB 93.60fF
C149 SD1R.n16 SUB 3.85fF
C150 SD1R.n17 SUB 3.85fF
C151 SD1R.n18 SUB 3.85fF
C152 SD1R.n19 SUB 3.85fF
C153 SD1R.n20 SUB 3.85fF
C154 SD1R.n21 SUB 3.85fF
C155 SD1R.n22 SUB 3.85fF
C156 SD1R.n23 SUB 3.85fF
C157 SD1R.n24 SUB 3.85fF
C158 SD1R.n25 SUB 3.85fF
C159 SD1R.n26 SUB 3.85fF
C160 SD1R.t67 SUB 3.50fF $ **FLOATING
C161 SD1R.t4 SUB 3.47fF $ **FLOATING
C162 SD1R.n27 SUB 3.85fF
C163 SD1R.n28 SUB 3.85fF
C164 SD1R.n29 SUB 3.85fF
C165 SD1R.n30 SUB 3.83fF
C166 SD1R.n31 SUB 3.84fF
C167 SD1R.n32 SUB 3.86fF
C168 SD1R.n33 SUB 3.86fF
C169 SD1R.n34 SUB 3.86fF
C170 SD1R.n35 SUB 3.86fF
C171 SD1R.n36 SUB 3.86fF
C172 SD1R.n37 SUB 3.86fF
C173 SD1R.n38 SUB 3.86fF
C174 SD1R.n39 SUB 3.86fF
C175 SD1R.n40 SUB 3.86fF
C176 SD1R.n41 SUB 3.86fF
C177 SD1R.n42 SUB 3.89fF
C178 SD1R.n43 SUB 3.83fF
C179 SD1R.n44 SUB 3.83fF
C180 SD1R.n45 SUB 3.85fF
C181 SD1R.n46 SUB 3.85fF
C182 SD1R.n47 SUB 3.85fF
C183 SD1R.n48 SUB 3.85fF
C184 SD1R.n49 SUB 3.85fF
C185 SD1R.n50 SUB 3.85fF
C186 SD1R.n51 SUB 3.85fF
C187 SD1R.n52 SUB 3.85fF
C188 SD1R.n53 SUB 3.85fF
C189 SD1R.n54 SUB 3.85fF
C190 SD1R.n55 SUB 3.85fF
C191 SD1R.t20 SUB 3.50fF $ **FLOATING
C192 SD1R.t61 SUB 3.47fF $ **FLOATING
C193 SD1R.n56 SUB 3.85fF
C194 SD1R.n57 SUB 3.85fF
C195 SD1R.n58 SUB 3.85fF
C196 SD1R.n59 SUB 150.53fF
C197 SD1R.n60 SUB 113.95fF
C198 SD1R.n61 SUB 3.83fF
C199 SD1R.n62 SUB 3.83fF
C200 SD1R.n63 SUB 3.86fF
C201 SD1R.n64 SUB 3.86fF
C202 SD1R.n65 SUB 3.86fF
C203 SD1R.n66 SUB 3.86fF
C204 SD1R.n67 SUB 3.86fF
C205 SD1R.n68 SUB 3.86fF
C206 SD1R.n69 SUB 3.86fF
C207 SD1R.n70 SUB 3.86fF
C208 SD1R.n71 SUB 3.86fF
C209 SD1R.n72 SUB 3.89fF
C210 SD1R.n73 SUB 3.86fF
C211 SD1R.n74 SUB 3.84fF
C212 SD1R.n75 SUB 3.83fF
C213 SD1R.n76 SUB 50.12fF
C214 SD2L.n0 SUB 3.85fF
C215 SD2L.n1 SUB 3.85fF
C216 SD2L.n2 SUB 3.85fF
C217 SD2L.n3 SUB 3.85fF
C218 SD2L.n4 SUB 3.85fF
C219 SD2L.n5 SUB 3.85fF
C220 SD2L.n6 SUB 3.85fF
C221 SD2L.n7 SUB 3.85fF
C222 SD2L.n8 SUB 3.85fF
C223 SD2L.n9 SUB 3.85fF
C224 SD2L.n10 SUB 3.85fF
C225 SD2L.t69 SUB 3.50fF $ **FLOATING
C226 SD2L.n11 SUB 10.49fF
C227 SD2L.n12 SUB 4.59fF
C228 SD2L.n13 SUB 4.59fF
C229 SD2L.n14 SUB 4.59fF
C230 SD2L.n15 SUB 4.59fF
C231 SD2L.n16 SUB 4.59fF
C232 SD2L.n17 SUB 4.59fF
C233 SD2L.n18 SUB 4.59fF
C234 SD2L.n19 SUB 4.59fF
C235 SD2L.n20 SUB 4.59fF
C236 SD2L.n21 SUB 3.92fF
C237 SD2L.n22 SUB 3.85fF
C238 SD2L.n23 SUB 3.85fF
C239 SD2L.n24 SUB 3.85fF
C240 SD2L.t43 SUB 3.47fF $ **FLOATING
C241 SD2L.n25 SUB 71.70fF
C242 SD2L.n26 SUB 3.86fF
C243 SD2L.n27 SUB 3.86fF
C244 SD2L.n28 SUB 3.86fF
C245 SD2L.n29 SUB 3.86fF
C246 SD2L.n30 SUB 3.86fF
C247 SD2L.n31 SUB 3.86fF
C248 SD2L.n32 SUB 3.86fF
C249 SD2L.n33 SUB 3.86fF
C250 SD2L.n34 SUB 3.86fF
C251 SD2L.n35 SUB 3.86fF
C252 SD2L.n36 SUB 3.89fF
C253 SD2L.n37 SUB 10.77fF
C254 SD2L.n38 SUB 4.59fF
C255 SD2L.n39 SUB 4.59fF
C256 SD2L.n40 SUB 4.59fF
C257 SD2L.n41 SUB 4.59fF
C258 SD2L.n42 SUB 4.59fF
C259 SD2L.n43 SUB 4.59fF
C260 SD2L.n44 SUB 4.59fF
C261 SD2L.n45 SUB 4.59fF
C262 SD2L.n46 SUB 4.72fF
C263 SD2L.n47 SUB 3.84fF
C264 SD2L.n48 SUB 3.74fF
C265 SD2L.n49 SUB 3.83fF
C266 SD2L.n50 SUB 3.83fF
C267 SD2L.n51 SUB 3.83fF
C268 SD2L.n52 SUB 53.45fF
C269 SD2L.n53 SUB 3.85fF
C270 SD2L.n54 SUB 3.85fF
C271 SD2L.n55 SUB 3.85fF
C272 SD2L.n56 SUB 3.85fF
C273 SD2L.n57 SUB 3.85fF
C274 SD2L.n58 SUB 3.85fF
C275 SD2L.n59 SUB 3.85fF
C276 SD2L.n60 SUB 3.85fF
C277 SD2L.n61 SUB 3.85fF
C278 SD2L.n62 SUB 3.85fF
C279 SD2L.n63 SUB 3.85fF
C280 SD2L.t31 SUB 3.50fF $ **FLOATING
C281 SD2L.n64 SUB 10.49fF
C282 SD2L.n65 SUB 4.59fF
C283 SD2L.n66 SUB 4.59fF
C284 SD2L.n67 SUB 4.59fF
C285 SD2L.n68 SUB 4.59fF
C286 SD2L.n69 SUB 4.59fF
C287 SD2L.n70 SUB 4.59fF
C288 SD2L.n71 SUB 4.59fF
C289 SD2L.n72 SUB 4.59fF
C290 SD2L.n73 SUB 4.59fF
C291 SD2L.n74 SUB 3.92fF
C292 SD2L.n75 SUB 3.85fF
C293 SD2L.n76 SUB 3.85fF
C294 SD2L.n77 SUB 3.85fF
C295 SD2L.t41 SUB 3.47fF $ **FLOATING
C296 SD2L.n78 SUB 71.70fF
C297 SD2L.n79 SUB 3.83fF
C298 SD2L.n80 SUB 3.83fF
C299 SD2L.n81 SUB 3.83fF
C300 SD2L.n82 SUB 3.84fF
C301 SD2L.n83 SUB 3.86fF
C302 SD2L.n84 SUB 3.86fF
C303 SD2L.n85 SUB 3.86fF
C304 SD2L.n86 SUB 3.86fF
C305 SD2L.n87 SUB 3.86fF
C306 SD2L.n88 SUB 3.86fF
C307 SD2L.n89 SUB 3.86fF
C308 SD2L.n90 SUB 3.86fF
C309 SD2L.n91 SUB 3.86fF
C310 SD2L.n92 SUB 3.89fF
C311 SD2L.n93 SUB 10.77fF
C312 SD2L.n94 SUB 4.59fF
C313 SD2L.n95 SUB 4.59fF
C314 SD2L.n96 SUB 4.59fF
C315 SD2L.n97 SUB 3.86fF
C316 SD2L.n98 SUB 4.59fF
C317 SD2L.n99 SUB 4.59fF
C318 SD2L.n100 SUB 4.59fF
C319 SD2L.n101 SUB 4.59fF
C320 SD2L.n102 SUB 4.59fF
C321 SD2L.n103 SUB 4.72fF
C322 SD2L.n104 SUB 3.74fF
C323 SD2L.n105 SUB 72.49fF
C324 SD2L.n106 SUB 153.29fF
C325 SD2L.n107 SUB 88.85fF
C326 SD2L.n108 SUB 82.60fF
C327 SD1L.n0 SUB 15.36fF
C328 SD1L.n1 SUB 89.49fF
C329 SD1L.n2 SUB 20.36fF
C330 SD1L.n3 SUB 18.74fF
C331 SD1L.n4 SUB 15.67fF
C332 SD1L.n5 SUB 18.74fF
C333 SD1L.n6 SUB 15.64fF
C334 SD1L.n7 SUB 117.64fF
C335 SD1L.n8 SUB 21.90fF
C336 SD1L.n9 SUB 50.97fF
C337 SD1L.n10 SUB 9.37fF
C338 SD1L.n11 SUB 46.28fF
C339 SD1L.n12 SUB 9.38fF
C340 SD1L.n13 SUB 15.40fF
C341 SD1L.n14 SUB 3.91fF
C342 SD1L.n15 SUB 3.91fF
C343 SD1L.n16 SUB 3.91fF
C344 SD1L.n17 SUB 3.91fF
C345 SD1L.n18 SUB 3.93fF
C346 SD1L.n19 SUB 3.93fF
C347 SD1L.n20 SUB 3.93fF
C348 SD1L.n21 SUB 3.93fF
C349 SD1L.n22 SUB 3.93fF
C350 SD1L.n23 SUB 3.93fF
C351 SD1L.n24 SUB 3.93fF
C352 SD1L.n25 SUB 3.93fF
C353 SD1L.n26 SUB 3.93fF
C354 SD1L.n27 SUB 3.93fF
C355 SD1L.n28 SUB 3.97fF
C356 SD1L.n29 SUB 3.93fF
C357 SD1L.n30 SUB 3.93fF
C358 SD1L.n31 SUB 3.93fF
C359 SD1L.n32 SUB 3.93fF
C360 SD1L.n33 SUB 3.93fF
C361 SD1L.n34 SUB 3.93fF
C362 SD1L.n35 SUB 3.93fF
C363 SD1L.n36 SUB 3.93fF
C364 SD1L.n37 SUB 3.93fF
C365 SD1L.n38 SUB 3.93fF
C366 SD1L.n39 SUB 3.97fF
C367 SD1L.n40 SUB 3.91fF
C368 SD1L.n41 SUB 3.91fF
C369 SD1L.n42 SUB 3.91fF
C370 SD1L.n43 SUB 3.91fF
C371 SD1L.n44 SUB 3.93fF
C372 SD1L.n45 SUB 3.93fF
C373 SD1L.n46 SUB 3.93fF
C374 SD1L.n47 SUB 3.93fF
C375 SD1L.n48 SUB 3.93fF
C376 SD1L.t44 SUB 3.57fF $ **FLOATING
C377 SD1L.n49 SUB 3.93fF
C378 SD1L.n50 SUB 3.93fF
C379 SD1L.n51 SUB 3.93fF
C380 SD1L.n52 SUB 3.93fF
C381 SD1L.n53 SUB 3.93fF
C382 SD1L.t42 SUB 3.57fF $ **FLOATING
C383 SD1L.n54 SUB 3.93fF
C384 SD1L.n55 SUB 3.93fF
C385 SD1L.n56 SUB 3.93fF
C386 SD1L.n57 SUB 3.93fF
C387 SD1L.n58 SUB 138.82fF
C388 SD1L.n59 SUB 3.93fF
C389 SD1L.n60 SUB 3.93fF
C390 SD1L.n61 SUB 3.93fF
C391 SD1L.n62 SUB 3.93fF
C392 SD1L.n63 SUB 3.93fF
C393 SD1L.n64 SUB 3.93fF
C394 SD1L.n65 SUB 3.93fF
C395 SD1L.n66 SUB 3.93fF
C396 SD1L.t53 SUB 3.57fF $ **FLOATING
C397 SD1L.n67 SUB 3.93fF
C398 SD1L.n68 SUB 3.93fF
C399 SD1L.n69 SUB 3.93fF
C400 SD1L.n70 SUB 3.93fF
C401 SD1L.n71 SUB 3.93fF
C402 SD1L.n72 SUB 3.93fF
C403 SD1L.t5 SUB 3.57fF $ **FLOATING
C404 SD1L.n73 SUB 96.96fF
C405 SD1L.n74 SUB 80.24fF
.ends