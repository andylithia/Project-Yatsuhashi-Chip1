magic
tech sky130A
magscale 1 2
timestamp 1658291001
<< pwell >>
rect -812 -439 812 439
<< nmos >>
rect -616 109 -416 229
rect -358 109 -158 229
rect -100 109 100 229
rect 158 109 358 229
rect 416 109 616 229
rect -616 -229 -416 -109
rect -358 -229 -158 -109
rect -100 -229 100 -109
rect 158 -229 358 -109
rect 416 -229 616 -109
<< ndiff >>
rect -674 217 -616 229
rect -674 121 -662 217
rect -628 121 -616 217
rect -674 109 -616 121
rect -416 217 -358 229
rect -416 121 -404 217
rect -370 121 -358 217
rect -416 109 -358 121
rect -158 217 -100 229
rect -158 121 -146 217
rect -112 121 -100 217
rect -158 109 -100 121
rect 100 217 158 229
rect 100 121 112 217
rect 146 121 158 217
rect 100 109 158 121
rect 358 217 416 229
rect 358 121 370 217
rect 404 121 416 217
rect 358 109 416 121
rect 616 217 674 229
rect 616 121 628 217
rect 662 121 674 217
rect 616 109 674 121
rect -674 -121 -616 -109
rect -674 -217 -662 -121
rect -628 -217 -616 -121
rect -674 -229 -616 -217
rect -416 -121 -358 -109
rect -416 -217 -404 -121
rect -370 -217 -358 -121
rect -416 -229 -358 -217
rect -158 -121 -100 -109
rect -158 -217 -146 -121
rect -112 -217 -100 -121
rect -158 -229 -100 -217
rect 100 -121 158 -109
rect 100 -217 112 -121
rect 146 -217 158 -121
rect 100 -229 158 -217
rect 358 -121 416 -109
rect 358 -217 370 -121
rect 404 -217 416 -121
rect 358 -229 416 -217
rect 616 -121 674 -109
rect 616 -217 628 -121
rect 662 -217 674 -121
rect 616 -229 674 -217
<< ndiffc >>
rect -662 121 -628 217
rect -404 121 -370 217
rect -146 121 -112 217
rect 112 121 146 217
rect 370 121 404 217
rect 628 121 662 217
rect -662 -217 -628 -121
rect -404 -217 -370 -121
rect -146 -217 -112 -121
rect 112 -217 146 -121
rect 370 -217 404 -121
rect 628 -217 662 -121
<< psubdiff >>
rect -776 369 -680 403
rect 680 369 776 403
rect -776 307 -742 369
rect 742 307 776 369
rect -776 -369 -742 -307
rect 742 -369 776 -307
rect -776 -403 -680 -369
rect 680 -403 776 -369
<< psubdiffcont >>
rect -680 369 680 403
rect -776 -307 -742 307
rect 742 -307 776 307
rect -680 -403 680 -369
<< poly >>
rect -616 301 -416 317
rect -616 267 -600 301
rect -432 267 -416 301
rect -616 229 -416 267
rect -358 301 -158 317
rect -358 267 -342 301
rect -174 267 -158 301
rect -358 229 -158 267
rect -100 301 100 317
rect -100 267 -84 301
rect 84 267 100 301
rect -100 229 100 267
rect 158 301 358 317
rect 158 267 174 301
rect 342 267 358 301
rect 158 229 358 267
rect 416 301 616 317
rect 416 267 432 301
rect 600 267 616 301
rect 416 229 616 267
rect -616 71 -416 109
rect -616 37 -600 71
rect -432 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 109
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 109
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect 416 71 616 109
rect 416 37 432 71
rect 600 37 616 71
rect 416 21 616 37
rect -616 -37 -416 -21
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -616 -109 -416 -71
rect -358 -37 -158 -21
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -358 -109 -158 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect 158 -37 358 -21
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 158 -109 358 -71
rect 416 -37 616 -21
rect 416 -71 432 -37
rect 600 -71 616 -37
rect 416 -109 616 -71
rect -616 -267 -416 -229
rect -616 -301 -600 -267
rect -432 -301 -416 -267
rect -616 -317 -416 -301
rect -358 -267 -158 -229
rect -358 -301 -342 -267
rect -174 -301 -158 -267
rect -358 -317 -158 -301
rect -100 -267 100 -229
rect -100 -301 -84 -267
rect 84 -301 100 -267
rect -100 -317 100 -301
rect 158 -267 358 -229
rect 158 -301 174 -267
rect 342 -301 358 -267
rect 158 -317 358 -301
rect 416 -267 616 -229
rect 416 -301 432 -267
rect 600 -301 616 -267
rect 416 -317 616 -301
<< polycont >>
rect -600 267 -432 301
rect -342 267 -174 301
rect -84 267 84 301
rect 174 267 342 301
rect 432 267 600 301
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect -600 -301 -432 -267
rect -342 -301 -174 -267
rect -84 -301 84 -267
rect 174 -301 342 -267
rect 432 -301 600 -267
<< locali >>
rect -776 369 -680 403
rect 680 369 776 403
rect -776 307 -742 369
rect 742 307 776 369
rect -616 267 -600 301
rect -432 267 -416 301
rect -358 267 -342 301
rect -174 267 -158 301
rect -100 267 -84 301
rect 84 267 100 301
rect 158 267 174 301
rect 342 267 358 301
rect 416 267 432 301
rect 600 267 616 301
rect -662 217 -628 233
rect -662 105 -628 121
rect -404 217 -370 233
rect -404 105 -370 121
rect -146 217 -112 233
rect -146 105 -112 121
rect 112 217 146 233
rect 112 105 146 121
rect 370 217 404 233
rect 370 105 404 121
rect 628 217 662 233
rect 628 105 662 121
rect -616 37 -600 71
rect -432 37 -416 71
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect 416 37 432 71
rect 600 37 616 71
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 416 -71 432 -37
rect 600 -71 616 -37
rect -662 -121 -628 -105
rect -662 -233 -628 -217
rect -404 -121 -370 -105
rect -404 -233 -370 -217
rect -146 -121 -112 -105
rect -146 -233 -112 -217
rect 112 -121 146 -105
rect 112 -233 146 -217
rect 370 -121 404 -105
rect 370 -233 404 -217
rect 628 -121 662 -105
rect 628 -233 662 -217
rect -616 -301 -600 -267
rect -432 -301 -416 -267
rect -358 -301 -342 -267
rect -174 -301 -158 -267
rect -100 -301 -84 -267
rect 84 -301 100 -267
rect 158 -301 174 -267
rect 342 -301 358 -267
rect 416 -301 432 -267
rect 600 -301 616 -267
rect -776 -369 -742 -307
rect 742 -369 776 -307
rect -776 -403 -680 -369
rect 680 -403 776 -369
<< viali >>
rect -600 267 -432 301
rect -342 267 -174 301
rect -84 267 84 301
rect 174 267 342 301
rect 432 267 600 301
rect -662 121 -628 217
rect -404 121 -370 217
rect -146 121 -112 217
rect 112 121 146 217
rect 370 121 404 217
rect 628 121 662 217
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect -662 -217 -628 -121
rect -404 -217 -370 -121
rect -146 -217 -112 -121
rect 112 -217 146 -121
rect 370 -217 404 -121
rect 628 -217 662 -121
rect -600 -301 -432 -267
rect -342 -301 -174 -267
rect -84 -301 84 -267
rect 174 -301 342 -267
rect 432 -301 600 -267
<< metal1 >>
rect -612 301 -420 307
rect -612 267 -600 301
rect -432 267 -420 301
rect -612 261 -420 267
rect -354 301 -162 307
rect -354 267 -342 301
rect -174 267 -162 301
rect -354 261 -162 267
rect -96 301 96 307
rect -96 267 -84 301
rect 84 267 96 301
rect -96 261 96 267
rect 162 301 354 307
rect 162 267 174 301
rect 342 267 354 301
rect 162 261 354 267
rect 420 301 612 307
rect 420 267 432 301
rect 600 267 612 301
rect 420 261 612 267
rect -668 217 -622 229
rect -668 121 -662 217
rect -628 121 -622 217
rect -668 109 -622 121
rect -410 217 -364 229
rect -410 121 -404 217
rect -370 121 -364 217
rect -410 109 -364 121
rect -152 217 -106 229
rect -152 121 -146 217
rect -112 121 -106 217
rect -152 109 -106 121
rect 106 217 152 229
rect 106 121 112 217
rect 146 121 152 217
rect 106 109 152 121
rect 364 217 410 229
rect 364 121 370 217
rect 404 121 410 217
rect 364 109 410 121
rect 622 217 668 229
rect 622 121 628 217
rect 662 121 668 217
rect 622 109 668 121
rect -612 71 -420 77
rect -612 37 -600 71
rect -432 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 432 71
rect 600 37 612 71
rect 420 31 612 37
rect -612 -37 -420 -31
rect -612 -71 -600 -37
rect -432 -71 -420 -37
rect -612 -77 -420 -71
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect 420 -37 612 -31
rect 420 -71 432 -37
rect 600 -71 612 -37
rect 420 -77 612 -71
rect -668 -121 -622 -109
rect -668 -217 -662 -121
rect -628 -217 -622 -121
rect -668 -229 -622 -217
rect -410 -121 -364 -109
rect -410 -217 -404 -121
rect -370 -217 -364 -121
rect -410 -229 -364 -217
rect -152 -121 -106 -109
rect -152 -217 -146 -121
rect -112 -217 -106 -121
rect -152 -229 -106 -217
rect 106 -121 152 -109
rect 106 -217 112 -121
rect 146 -217 152 -121
rect 106 -229 152 -217
rect 364 -121 410 -109
rect 364 -217 370 -121
rect 404 -217 410 -121
rect 364 -229 410 -217
rect 622 -121 668 -109
rect 622 -217 628 -121
rect 662 -217 668 -121
rect 622 -229 668 -217
rect -612 -267 -420 -261
rect -612 -301 -600 -267
rect -432 -301 -420 -267
rect -612 -307 -420 -301
rect -354 -267 -162 -261
rect -354 -301 -342 -267
rect -174 -301 -162 -267
rect -354 -307 -162 -301
rect -96 -267 96 -261
rect -96 -301 -84 -267
rect 84 -301 96 -267
rect -96 -307 96 -301
rect 162 -267 354 -261
rect 162 -301 174 -267
rect 342 -301 354 -267
rect 162 -307 354 -301
rect 420 -267 612 -261
rect 420 -301 432 -267
rect 600 -301 612 -267
rect 420 -307 612 -301
<< properties >>
string FIXED_BBOX -759 -386 759 386
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.6 l 1 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
