.subckt NMOS_30_0p5_30_interdigital_diff4x SD1L SD2L GL SD1R SD2R GR SUB
X0 SD2L.t119 GL SD1L.t118 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X1 SD2R.t119 GR SD1R.t69 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X2 SD1R.t107 GR SD2R.t118 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X3 SD2L.t118 GL SD1L.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X4 SD2L.t117 GL SD1L.t13 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X5 SD1L.t28 GL SD2L.t116 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X6 SD2R.t117 GR SD1R.t33 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X7 SD1L.t95 GL SD2L.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X8 SD1L.t47 GL SD2L.t114 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X9 SD1R.t58 GR SD2R.t116 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X10 SD1R.t83 GR SD2R.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X11 SD1R.t114 GR SD2R.t114 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X12 SD2R.t113 GR SD1R.t55 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X13 SD1R.t24 GR SD2R.t112 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X14 SD2L.t113 GL SD1L.t61 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X15 SD2R.t111 GR SD1R.t43 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X16 SD1R.t63 GR SD2R.t110 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X17 SD2R.t109 GR SD1R.t92 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X18 SD2L.t112 GL SD1L.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X19 SD2L.t111 GL SD1L.t63 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X20 SD2R.t108 GR SD1R.t97 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X21 SD1L.t59 GL SD2L.t110 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X22 SD1R.t98 GR SD2R.t107 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X23 SD2L.t109 GL SD1L.t119 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X24 SD2L.t108 GL SD1L.t25 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X25 SD1R.t18 GR SD2R.t106 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X26 SD2R.t105 GR SD1R.t57 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X27 SD1L.t16 GL SD2L.t107 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X28 SD2L.t106 GL SD1L.t90 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X29 SD1R.t91 GR SD2R.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X30 SD1R.t100 GR SD2R.t103 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X31 SD2L.t105 GL SD1L.t93 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X32 SD1R.t111 GR SD2R.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X33 SD1L.t97 GL SD2L.t104 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X34 SD1R.t118 GR SD2R.t101 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X35 SD1R.t36 GR SD2R.t100 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X36 SD2R.t99 GR SD1R.t31 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X37 SD2R.t98 GR SD1R.t61 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X38 SD1L.t94 GL SD2L.t103 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X39 SD1L.t65 GL SD2L.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X40 SD1L.t62 GL SD2L.t101 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X41 SD2R.t97 GR SD1R.t77 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X42 SD2R.t96 GR SD1R.t99 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X43 SD1R.t7 GR SD2R.t95 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X44 SD1R.t113 GR SD2R.t94 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X45 SD2R.t93 GR SD1R.t17 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X46 SD2R.t92 GR SD1R.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X47 SD1L.t98 GL SD2L.t100 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X48 SD2R.t91 GR SD1R.t16 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X49 SD2L.t99 GL SD1L.t101 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X50 SD2L.t98 GL SD1L.t114 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X51 SD2L.t97 GL SD1L.t113 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X52 SD1R.t28 GR SD2R.t90 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X53 SD2L.t96 GL SD1L.t96 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X54 SD2R.t89 GR SD1R.t6 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X55 SD2R.t88 GR SD1R.t59 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X56 SD2L.t95 GL SD1L.t58 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X57 SD2L.t94 GL SD1L.t4 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X58 SD1R.t26 GR SD2R.t87 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X59 SD1R.t95 GR SD2R.t86 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X60 SD1R.t96 GR SD2R.t85 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X61 SD1L.t37 GL SD2L.t93 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X62 SD2R.t84 GR SD1R.t23 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X63 SD1R.t22 GR SD2R.t83 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X64 SD2R.t82 GR SD1R.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X65 SD2R.t81 GR SD1R.t66 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X66 SD1R.t38 GR SD2R.t80 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X67 SD1L.t11 GL SD2L.t92 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X68 SD2R.t79 GR SD1R.t52 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X69 SD1L.t52 GL SD2L.t91 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X70 SD1R.t81 GR SD2R.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X71 SD2R.t77 GR SD1R.t90 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X72 SD2L.t90 GL SD1L.t18 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X73 SD1L.t92 GL SD2L.t89 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X74 SD2R.t76 GR SD1R.t88 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X75 SD2L.t88 GL SD1L.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X76 SD2L.t87 GL SD1L.t105 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X77 SD2R.t75 GR SD1R.t29 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X78 SD1R.t104 GR SD2R.t74 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X79 SD2L.t86 GL SD1L.t115 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X80 SD2L.t85 GL SD1L.t60 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X81 SD2L.t84 GL SD1L.t81 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X82 SD1R.t39 GR SD2R.t73 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X83 SD2L.t83 GL SD1L.t41 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X84 SD1L.t44 GL SD2L.t82 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X85 SD1R.t44 GR SD2R.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X86 SD2L.t81 GL SD1L.t91 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X87 SD1L.t106 GL SD2L.t80 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X88 SD1R.t87 GR SD2R.t71 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X89 SD2L.t79 GL SD1L.t75 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X90 SD1L.t26 GL SD2L.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X91 SD1L.t89 GL SD2L.t77 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X92 SD2L.t76 GL SD1L.t29 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X93 SD1L.t57 GL SD2L.t75 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X94 SD1R.t34 GR SD2R.t70 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X95 SD1R.t51 GR SD2R.t69 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X96 SD2L.t74 GL SD1L.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X97 SD2L.t73 GL SD1L.t76 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X98 SD1R.t8 GR SD2R.t68 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X99 SD1L.t80 GL SD2L.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X100 SD1L.t85 GL SD2L.t71 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X101 SD2L.t70 GL SD1L.t36 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X102 SD1L.t67 GL SD2L.t69 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X103 SD1L.t112 GL SD2L.t68 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X104 SD2R.t67 GR SD1R.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X105 SD1L.t104 GL SD2L.t67 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X106 SD2R.t66 GR SD1R.t75 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X107 SD2L.t66 GL SD1L.t14 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X108 SD1R.t54 GR SD2R.t65 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X109 SD2L.t65 GL SD1L.t69 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X110 SD2R.t64 GR SD1R.t102 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X111 SD2L.t64 GL SD1L.t83 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X112 SD1R.t45 GR SD2R.t63 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X113 SD2L.t63 GL SD1L.t32 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X114 SD2R.t62 GR SD1R.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X115 SD1L.t116 GL SD2L.t62 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X116 SD2L.t61 GL SD1L.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X117 SD2R.t61 GR SD1R.t46 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X118 SD2R.t60 GR SD1R.t2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X119 SD1L.t24 GL SD2L.t60 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X120 SD1L.t9 GL SD2L.t59 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X121 SD2R.t59 GR SD1R.t47 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X122 SD1R.t4 GR SD2R.t58 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X123 SD2L.t58 GL SD1L.t3 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X124 SD1L.t68 GL SD2L.t57 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X125 SD1L.t21 GL SD2L.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X126 SD1R.t109 GR SD2R.t57 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X127 SD1R.t5 GR SD2R.t56 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X128 SD2L.t55 GL SD1L.t54 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X129 SD1L.t34 GL SD2L.t54 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X130 SD2L.t53 GL SD1L.t82 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X131 SD2R.t55 GR SD1R.t32 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X132 SD1L.t111 GL SD2L.t52 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X133 SD2R.t54 GR SD1R.t119 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X134 SD1R.t70 GR SD2R.t53 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X135 SD2L.t51 GL SD1L.t40 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X136 SD2R.t52 GR SD1R.t48 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X137 SD1R.t67 GR SD2R.t51 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X138 SD1L.t2 GL SD2L.t50 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X139 SD2R.t50 GR SD1R.t15 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X140 SD1R.t19 GR SD2R.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X141 SD1L.t27 GL SD2L.t49 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X142 SD2L.t48 GL SD1L.t74 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X143 SD2L.t47 GL SD1L.t71 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X144 SD1R.t13 GR SD2R.t48 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X145 SD1R.t89 GR SD2R.t47 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X146 SD2R.t46 GR SD1R.t117 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X147 SD1R.t80 GR SD2R.t45 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X148 SD1L.t23 GL SD2L.t46 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X149 SD1L.t53 GL SD2L.t45 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X150 SD2R.t44 GR SD1R.t94 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X151 SD2R.t43 GR SD1R.t93 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X152 SD1L.t39 GL SD2L.t44 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X153 SD1L.t84 GL SD2L.t43 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X154 SD1L.t88 GL SD2L.t42 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X155 SD1R.t105 GR SD2R.t42 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X156 SD1L.t17 GL SD2L.t41 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X157 SD2L.t40 GL SD1L.t73 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X158 SD2R.t41 GR SD1R.t40 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X159 SD1R.t115 GR SD2R.t40 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X160 SD2R.t39 GR SD1R.t101 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X161 SD1R.t50 GR SD2R.t38 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X162 SD1R.t27 GR SD2R.t37 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X163 SD2R.t36 GR SD1R.t76 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X164 SD2R.t35 GR SD1R.t3 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X165 SD1R.t62 GR SD2R.t34 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X166 SD1L.t66 GL SD2L.t39 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X167 SD1L.t51 GL SD2L.t38 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X168 SD2L.t37 GL SD1L.t7 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X169 SD2L.t36 GL SD1L.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X170 SD1R.t25 GR SD2R.t33 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X171 SD1L.t35 GL SD2L.t35 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X172 SD1L.t55 GL SD2L.t34 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X173 SD2R.t32 GR SD1R.t79 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X174 SD1L.t8 GL SD2L.t33 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X175 SD1R.t53 GR SD2R.t31 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X176 SD1L.t64 GL SD2L.t32 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X177 SD2R.t30 GR SD1R.t116 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X178 SD2R.t29 GR SD1R.t35 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X179 SD2R.t28 GR SD1R.t108 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X180 SD2R.t27 GR SD1R.t41 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X181 SD1R.t110 GR SD2R.t26 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X182 SD1R.t42 GR SD2R.t25 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X183 SD2R.t24 GR SD1R.t60 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X184 SD1R.t37 GR SD2R.t23 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X185 SD2R.t22 GR SD1R.t85 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X186 SD2L.t31 GL SD1L.t33 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X187 SD2L.t30 GL SD1L.t46 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X188 SD2L.t29 GL SD1L.t108 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X189 SD2R.t21 GR SD1R.t73 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X190 SD2L.t28 GL SD1L.t1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X191 SD2R.t20 GR SD1R.t71 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X192 SD1L.t19 GL SD2L.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X193 SD1R.t1 GR SD2R.t19 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X194 SD2L.t26 GL SD1L.t20 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X195 SD1R.t68 GR SD2R.t18 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X196 SD1R.t0 GR SD2R.t17 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X197 SD1L.t117 GL SD2L.t25 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X198 SD2R.t16 GR SD1R.t11 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X199 SD1L.t31 GL SD2L.t24 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X200 SD1R.t65 GR SD2R.t15 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X201 SD1L.t48 GL SD2L.t23 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X202 SD2R.t14 GR SD1R.t78 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X203 SD1L.t45 GL SD2L.t22 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X204 SD1R.t74 GR SD2R.t13 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X205 SD2L.t21 GL SD1L.t5 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X206 SD2L.t20 GL SD1L.t38 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X207 SD1R.t84 GR SD2R.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X208 SD1L.t86 GL SD2L.t19 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X209 SD2R.t11 GR SD1R.t86 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X210 SD1R.t106 GR SD2R.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X211 SD2L.t18 GL SD1L.t109 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X212 SD2L.t17 GL SD1L.t110 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X213 SD2L.t16 GL SD1L.t77 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X214 SD1R.t112 GR SD2R.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X215 SD2R.t8 GR SD1R.t64 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X216 SD1L.t99 GL SD2L.t15 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X217 SD1L.t0 GL SD2L.t14 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X218 SD2L.t13 GL SD1L.t107 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X219 SD2R.t7 GR SD1R.t103 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X220 SD2L.t12 GL SD1L.t30 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X221 SD1R.t20 GR SD2R.t6 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X222 SD1L.t49 GL SD2L.t11 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X223 SD1L.t6 GL SD2L.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X224 SD1R.t14 GR SD2R.t5 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X225 SD1L.t43 GL SD2L.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X226 SD2R.t4 GR SD1R.t72 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X227 SD1L.t70 GL SD2L.t8 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X228 SD2L.t7 GL SD1L.t42 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X229 SD1L.t15 GL SD2L.t6 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X230 SD2L.t5 GL SD1L.t22 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X231 SD2R.t3 GR SD1R.t30 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X232 SD1L.t103 GL SD2L.t4 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X233 SD2R.t2 GR SD1R.t21 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X234 SD2L.t3 GL SD1L.t79 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X235 SD1L.t50 GL SD2L.t2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X236 SD2R.t1 GR SD1R.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X237 SD2R.t0 GR SD1R.t82 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X238 SD2L.t1 GL SD1L.t87 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X239 SD2L.t0 GL SD1L.t100 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
C0 SD1L SD2R 36.54fF
C1 SD2L SD2R 50.41fF
C2 GR SD2R 116.25fF
C3 SD1L GL 112.81fF
C4 SD2L GL 112.76fF
C5 SD2R SD1R 1294.62fF
C6 GR GL 27.31fF
C7 SD1R GL 15.71fF
C8 SD1L SD2L 1294.36fF
C9 SD1L GR 20.74fF
C10 SD2L GR 17.10fF
C11 SD1L SD1R 63.14fF
C12 SD2L SD1R 28.64fF
C13 GR SD1R 107.41fF
C14 SD2R GL 16.51fF
R0 SD1L.n25 SD1L.t35 2.284
R1 SD1L.n11 SD1L.t73 2.284
R2 SD1L.n79 SD1L.t98 2.284
R3 SD1L.n65 SD1L.t115 2.284
R4 SD1L.n109 SD1L.n108 1.74
R5 SD1L.n50 SD1L.n49 1.739
R6 SD1L.n36 SD1L.n35 1.739
R7 SD1L.n97 SD1L.n96 1.739
R8 SD1L.n50 SD1L.n48 1.702
R9 SD1L.n51 SD1L.n47 1.702
R10 SD1L.n52 SD1L.n46 1.702
R11 SD1L.n53 SD1L.n45 1.702
R12 SD1L.n54 SD1L.n44 1.702
R13 SD1L.n55 SD1L.n43 1.702
R14 SD1L.n57 SD1L.n41 1.702
R15 SD1L.n2 SD1L.n40 1.702
R16 SD1L.n39 SD1L.n31 1.702
R17 SD1L.n38 SD1L.n32 1.702
R18 SD1L.n37 SD1L.n33 1.702
R19 SD1L.n36 SD1L.n34 1.702
R20 SD1L.n97 SD1L.n95 1.702
R21 SD1L.n98 SD1L.n94 1.702
R22 SD1L.n99 SD1L.n93 1.702
R23 SD1L.n100 SD1L.n92 1.702
R24 SD1L.n101 SD1L.n91 1.702
R25 SD1L.n102 SD1L.n90 1.702
R26 SD1L.n104 SD1L.n88 1.702
R27 SD1L.n3 SD1L.n87 1.702
R28 SD1L.n113 SD1L.n105 1.702
R29 SD1L.n112 SD1L.n106 1.702
R30 SD1L.n109 SD1L.n107 1.702
R31 SD1L.n111 SD1L.n110 1.701
R32 SD1L.n25 SD1L.n24 1.696
R33 SD1L.n26 SD1L.n23 1.696
R34 SD1L.n27 SD1L.n22 1.696
R35 SD1L.n28 SD1L.n21 1.696
R36 SD1L.n29 SD1L.n20 1.696
R37 SD1L.n30 SD1L.n19 1.696
R38 SD1L.n0 SD1L.n18 1.696
R39 SD1L.n17 SD1L.n4 1.696
R40 SD1L.n16 SD1L.n5 1.696
R41 SD1L.n15 SD1L.n6 1.696
R42 SD1L.n14 SD1L.n7 1.696
R43 SD1L.n13 SD1L.n8 1.696
R44 SD1L.n12 SD1L.n9 1.696
R45 SD1L.n11 SD1L.n10 1.696
R46 SD1L.n79 SD1L.n78 1.696
R47 SD1L.n80 SD1L.n77 1.696
R48 SD1L.n81 SD1L.n76 1.696
R49 SD1L.n82 SD1L.n75 1.696
R50 SD1L.n83 SD1L.n74 1.696
R51 SD1L.n84 SD1L.n73 1.696
R52 SD1L.n1 SD1L.n72 1.696
R53 SD1L.n71 SD1L.n58 1.696
R54 SD1L.n70 SD1L.n59 1.696
R55 SD1L.n69 SD1L.n60 1.696
R56 SD1L.n68 SD1L.n61 1.696
R57 SD1L.n67 SD1L.n62 1.696
R58 SD1L.n66 SD1L.n63 1.696
R59 SD1L.n65 SD1L.n64 1.696
R60 SD1L.n56 SD1L.n42 1.678
R61 SD1L.n103 SD1L.n89 1.678
R62 SD1L.n85 SD1L.n1 0.569
R63 SD1L.n24 SD1L.t60 0.551
R64 SD1L.n24 SD1L.t15 0.551
R65 SD1L.n23 SD1L.t109 0.551
R66 SD1L.n23 SD1L.t39 0.551
R67 SD1L.n22 SD1L.t102 0.551
R68 SD1L.n22 SD1L.t49 0.551
R69 SD1L.n21 SD1L.t5 0.551
R70 SD1L.n21 SD1L.t24 0.551
R71 SD1L.n20 SD1L.t119 0.551
R72 SD1L.n20 SD1L.t99 0.551
R73 SD1L.n19 SD1L.t82 0.551
R74 SD1L.n19 SD1L.t116 0.551
R75 SD1L.n18 SD1L.t63 0.551
R76 SD1L.n18 SD1L.t66 0.551
R77 SD1L.n4 SD1L.t78 0.551
R78 SD1L.n4 SD1L.t6 0.551
R79 SD1L.n5 SD1L.t38 0.551
R80 SD1L.n5 SD1L.t9 0.551
R81 SD1L.n6 SD1L.t69 0.551
R82 SD1L.n6 SD1L.t19 0.551
R83 SD1L.n7 SD1L.t36 0.551
R84 SD1L.n7 SD1L.t106 0.551
R85 SD1L.n8 SD1L.t61 0.551
R86 SD1L.n8 SD1L.t28 0.551
R87 SD1L.n9 SD1L.t76 0.551
R88 SD1L.n9 SD1L.t44 0.551
R89 SD1L.n10 SD1L.t22 0.551
R90 SD1L.n10 SD1L.t27 0.551
R91 SD1L.n78 SD1L.t42 0.551
R92 SD1L.n78 SD1L.t2 0.551
R93 SD1L.n77 SD1L.t3 0.551
R94 SD1L.n77 SD1L.t16 0.551
R95 SD1L.n76 SD1L.t20 0.551
R96 SD1L.n76 SD1L.t104 0.551
R97 SD1L.n75 SD1L.t75 0.551
R98 SD1L.n75 SD1L.t59 0.551
R99 SD1L.n74 SD1L.t72 0.551
R100 SD1L.n74 SD1L.t85 0.551
R101 SD1L.n73 SD1L.t10 0.551
R102 SD1L.n73 SD1L.t103 0.551
R103 SD1L.n72 SD1L.t71 0.551
R104 SD1L.n72 SD1L.t52 0.551
R105 SD1L.n58 SD1L.t100 0.551
R106 SD1L.n58 SD1L.t88 0.551
R107 SD1L.n59 SD1L.t74 0.551
R108 SD1L.n59 SD1L.t62 0.551
R109 SD1L.n60 SD1L.t93 0.551
R110 SD1L.n60 SD1L.t23 0.551
R111 SD1L.n61 SD1L.t113 0.551
R112 SD1L.n61 SD1L.t94 0.551
R113 SD1L.n62 SD1L.t46 0.551
R114 SD1L.n62 SD1L.t64 0.551
R115 SD1L.n63 SD1L.t12 0.551
R116 SD1L.n63 SD1L.t95 0.551
R117 SD1L.n64 SD1L.t33 0.551
R118 SD1L.n64 SD1L.t26 0.551
R119 SD1L.n49 SD1L.t56 0.551
R120 SD1L.n49 SD1L.t112 0.551
R121 SD1L.n48 SD1L.t41 0.551
R122 SD1L.n48 SD1L.t111 0.551
R123 SD1L.n47 SD1L.t32 0.551
R124 SD1L.n47 SD1L.t84 0.551
R125 SD1L.n46 SD1L.t1 0.551
R126 SD1L.n46 SD1L.t50 0.551
R127 SD1L.n45 SD1L.t30 0.551
R128 SD1L.n45 SD1L.t45 0.551
R129 SD1L.n44 SD1L.t87 0.551
R130 SD1L.n44 SD1L.t70 0.551
R131 SD1L.n43 SD1L.t29 0.551
R132 SD1L.n43 SD1L.t92 0.551
R133 SD1L.n42 SD1L.t4 0.551
R134 SD1L.n42 SD1L.t57 0.551
R135 SD1L.n41 SD1L.t105 0.551
R136 SD1L.n41 SD1L.t21 0.551
R137 SD1L.n40 SD1L.t7 0.551
R138 SD1L.n40 SD1L.t86 0.551
R139 SD1L.n31 SD1L.t108 0.551
R140 SD1L.n31 SD1L.t55 0.551
R141 SD1L.n32 SD1L.t77 0.551
R142 SD1L.n32 SD1L.t31 0.551
R143 SD1L.n33 SD1L.t13 0.551
R144 SD1L.n33 SD1L.t65 0.551
R145 SD1L.n34 SD1L.t91 0.551
R146 SD1L.n34 SD1L.t11 0.551
R147 SD1L.n35 SD1L.t96 0.551
R148 SD1L.n35 SD1L.t67 0.551
R149 SD1L.n96 SD1L.t114 0.551
R150 SD1L.n96 SD1L.t97 0.551
R151 SD1L.n95 SD1L.t81 0.551
R152 SD1L.n95 SD1L.t34 0.551
R153 SD1L.n94 SD1L.t83 0.551
R154 SD1L.n94 SD1L.t53 0.551
R155 SD1L.n93 SD1L.t40 0.551
R156 SD1L.n93 SD1L.t8 0.551
R157 SD1L.n92 SD1L.t107 0.551
R158 SD1L.n92 SD1L.t48 0.551
R159 SD1L.n91 SD1L.t79 0.551
R160 SD1L.n91 SD1L.t43 0.551
R161 SD1L.n90 SD1L.t90 0.551
R162 SD1L.n90 SD1L.t47 0.551
R163 SD1L.n89 SD1L.t58 0.551
R164 SD1L.n89 SD1L.t89 0.551
R165 SD1L.n88 SD1L.t18 0.551
R166 SD1L.n88 SD1L.t68 0.551
R167 SD1L.n87 SD1L.t14 0.551
R168 SD1L.n87 SD1L.t17 0.551
R169 SD1L.n105 SD1L.t54 0.551
R170 SD1L.n105 SD1L.t51 0.551
R171 SD1L.n106 SD1L.t110 0.551
R172 SD1L.n106 SD1L.t117 0.551
R173 SD1L.n107 SD1L.t25 0.551
R174 SD1L.n107 SD1L.t37 0.551
R175 SD1L.n108 SD1L.t101 0.551
R176 SD1L.n108 SD1L.t80 0.551
R177 SD1L.n110 SD1L.t118 0.551
R178 SD1L.n110 SD1L.t0 0.551
R179 SD1L.n86 SD1L.n0 0.437
R180 SD1L.n114 SD1L.n86 0.099
R181 SD1L.n85 SD1L.n2 0.075
R182 SD1L.n114 SD1L.n3 0.075
R183 SD1L.n86 SD1L.n85 0.07
R184 SD1L SD1L.n114 0.04
R185 SD1L.n26 SD1L.n25 0.037
R186 SD1L.n27 SD1L.n26 0.037
R187 SD1L.n28 SD1L.n27 0.037
R188 SD1L.n29 SD1L.n28 0.037
R189 SD1L.n30 SD1L.n29 0.037
R190 SD1L.n0 SD1L.n30 0.037
R191 SD1L.n17 SD1L.n16 0.037
R192 SD1L.n16 SD1L.n15 0.037
R193 SD1L.n15 SD1L.n14 0.037
R194 SD1L.n14 SD1L.n13 0.037
R195 SD1L.n13 SD1L.n12 0.037
R196 SD1L.n12 SD1L.n11 0.037
R197 SD1L.n80 SD1L.n79 0.037
R198 SD1L.n81 SD1L.n80 0.037
R199 SD1L.n82 SD1L.n81 0.037
R200 SD1L.n83 SD1L.n82 0.037
R201 SD1L.n84 SD1L.n83 0.037
R202 SD1L.n1 SD1L.n84 0.037
R203 SD1L.n71 SD1L.n70 0.037
R204 SD1L.n70 SD1L.n69 0.037
R205 SD1L.n69 SD1L.n68 0.037
R206 SD1L.n68 SD1L.n67 0.037
R207 SD1L.n67 SD1L.n66 0.037
R208 SD1L.n66 SD1L.n65 0.037
R209 SD1L.n51 SD1L.n50 0.037
R210 SD1L.n52 SD1L.n51 0.037
R211 SD1L.n53 SD1L.n52 0.037
R212 SD1L.n54 SD1L.n53 0.037
R213 SD1L.n55 SD1L.n54 0.037
R214 SD1L.n56 SD1L.n55 0.037
R215 SD1L.n57 SD1L.n56 0.037
R216 SD1L.n2 SD1L.n57 0.037
R217 SD1L.n39 SD1L.n38 0.037
R218 SD1L.n38 SD1L.n37 0.037
R219 SD1L.n37 SD1L.n36 0.037
R220 SD1L.n98 SD1L.n97 0.037
R221 SD1L.n99 SD1L.n98 0.037
R222 SD1L.n100 SD1L.n99 0.037
R223 SD1L.n101 SD1L.n100 0.037
R224 SD1L.n102 SD1L.n101 0.037
R225 SD1L.n103 SD1L.n102 0.037
R226 SD1L.n104 SD1L.n103 0.037
R227 SD1L.n3 SD1L.n104 0.037
R228 SD1L.n113 SD1L.n112 0.037
R229 SD1L.n112 SD1L.n111 0.037
R230 SD1L.n111 SD1L.n109 0.037
R231 SD1L.n3 SD1L.n113 0.037
R232 SD1L.n2 SD1L.n39 0.037
R233 SD1L.n1 SD1L.n71 0.036
R234 SD1L.n0 SD1L.n17 0.036
R235 SD2L.n5 SD2L.t72 2.285
R236 SD2L.n77 SD2L.t61 2.284
R237 SD2L.n63 SD2L.t69 2.284
R238 SD2L.n19 SD2L.t98 2.284
R239 SD2L.n45 SD2L.n44 1.739
R240 SD2L.n31 SD2L.n30 1.739
R241 SD2L.n99 SD2L.n98 1.739
R242 SD2L.n114 SD2L.n113 1.739
R243 SD2L.n45 SD2L.n43 1.702
R244 SD2L.n46 SD2L.n42 1.702
R245 SD2L.n47 SD2L.n41 1.702
R246 SD2L.n48 SD2L.n40 1.702
R247 SD2L.n49 SD2L.n39 1.702
R248 SD2L.n50 SD2L.n38 1.702
R249 SD2L.n52 SD2L.n36 1.702
R250 SD2L.n53 SD2L.n35 1.702
R251 SD2L.n54 SD2L.n34 1.702
R252 SD2L.n55 SD2L.n33 1.702
R253 SD2L.n56 SD2L.n32 1.702
R254 SD2L.n31 SD2L.n29 1.702
R255 SD2L.n99 SD2L.n97 1.702
R256 SD2L.n100 SD2L.n96 1.702
R257 SD2L.n101 SD2L.n95 1.702
R258 SD2L.n102 SD2L.n94 1.702
R259 SD2L.n105 SD2L.n93 1.702
R260 SD2L.n107 SD2L.n91 1.702
R261 SD2L.n108 SD2L.n90 1.702
R262 SD2L.n109 SD2L.n89 1.702
R263 SD2L.n110 SD2L.n88 1.702
R264 SD2L.n111 SD2L.n87 1.702
R265 SD2L.n114 SD2L.n112 1.702
R266 SD2L.n104 SD2L.n103 1.701
R267 SD2L.n77 SD2L.n76 1.696
R268 SD2L.n78 SD2L.n75 1.696
R269 SD2L.n79 SD2L.n74 1.696
R270 SD2L.n80 SD2L.n73 1.696
R271 SD2L.n81 SD2L.n72 1.696
R272 SD2L.n82 SD2L.n71 1.696
R273 SD2L.n83 SD2L.n70 1.696
R274 SD2L.n84 SD2L.n69 1.696
R275 SD2L.n85 SD2L.n68 1.696
R276 SD2L.n67 SD2L.n58 1.696
R277 SD2L.n66 SD2L.n59 1.696
R278 SD2L.n65 SD2L.n60 1.696
R279 SD2L.n64 SD2L.n61 1.696
R280 SD2L.n63 SD2L.n62 1.696
R281 SD2L.n19 SD2L.n18 1.696
R282 SD2L.n20 SD2L.n17 1.696
R283 SD2L.n21 SD2L.n16 1.696
R284 SD2L.n22 SD2L.n15 1.696
R285 SD2L.n23 SD2L.n14 1.696
R286 SD2L.n24 SD2L.n13 1.696
R287 SD2L.n25 SD2L.n12 1.696
R288 SD2L.n26 SD2L.n11 1.696
R289 SD2L.n27 SD2L.n10 1.696
R290 SD2L.n9 SD2L.n0 1.696
R291 SD2L.n8 SD2L.n1 1.696
R292 SD2L.n7 SD2L.n2 1.696
R293 SD2L.n6 SD2L.n3 1.696
R294 SD2L.n5 SD2L.n4 1.696
R295 SD2L.n51 SD2L.n37 1.678
R296 SD2L.n106 SD2L.n92 1.678
R297 SD2L.n44 SD2L.t35 0.551
R298 SD2L.n44 SD2L.t85 0.551
R299 SD2L.n43 SD2L.t6 0.551
R300 SD2L.n43 SD2L.t18 0.551
R301 SD2L.n42 SD2L.t44 0.551
R302 SD2L.n42 SD2L.t88 0.551
R303 SD2L.n41 SD2L.t11 0.551
R304 SD2L.n41 SD2L.t21 0.551
R305 SD2L.n40 SD2L.t60 0.551
R306 SD2L.n40 SD2L.t109 0.551
R307 SD2L.n39 SD2L.t15 0.551
R308 SD2L.n39 SD2L.t53 0.551
R309 SD2L.n38 SD2L.t62 0.551
R310 SD2L.n38 SD2L.t111 0.551
R311 SD2L.n37 SD2L.t39 0.551
R312 SD2L.n37 SD2L.t74 0.551
R313 SD2L.n36 SD2L.t10 0.551
R314 SD2L.n36 SD2L.t20 0.551
R315 SD2L.n35 SD2L.t59 0.551
R316 SD2L.n35 SD2L.t65 0.551
R317 SD2L.n34 SD2L.t27 0.551
R318 SD2L.n34 SD2L.t70 0.551
R319 SD2L.n33 SD2L.t80 0.551
R320 SD2L.n33 SD2L.t113 0.551
R321 SD2L.n32 SD2L.t116 0.551
R322 SD2L.n32 SD2L.t73 0.551
R323 SD2L.n29 SD2L.t82 0.551
R324 SD2L.n29 SD2L.t5 0.551
R325 SD2L.n30 SD2L.t49 0.551
R326 SD2L.n30 SD2L.t40 0.551
R327 SD2L.n76 SD2L.t68 0.551
R328 SD2L.n76 SD2L.t83 0.551
R329 SD2L.n75 SD2L.t52 0.551
R330 SD2L.n75 SD2L.t63 0.551
R331 SD2L.n74 SD2L.t43 0.551
R332 SD2L.n74 SD2L.t28 0.551
R333 SD2L.n73 SD2L.t2 0.551
R334 SD2L.n73 SD2L.t12 0.551
R335 SD2L.n72 SD2L.t22 0.551
R336 SD2L.n72 SD2L.t1 0.551
R337 SD2L.n71 SD2L.t8 0.551
R338 SD2L.n71 SD2L.t76 0.551
R339 SD2L.n70 SD2L.t89 0.551
R340 SD2L.n70 SD2L.t94 0.551
R341 SD2L.n69 SD2L.t75 0.551
R342 SD2L.n69 SD2L.t87 0.551
R343 SD2L.n68 SD2L.t56 0.551
R344 SD2L.n68 SD2L.t37 0.551
R345 SD2L.n58 SD2L.t19 0.551
R346 SD2L.n58 SD2L.t29 0.551
R347 SD2L.n59 SD2L.t34 0.551
R348 SD2L.n59 SD2L.t16 0.551
R349 SD2L.n60 SD2L.t24 0.551
R350 SD2L.n60 SD2L.t117 0.551
R351 SD2L.n61 SD2L.t102 0.551
R352 SD2L.n61 SD2L.t81 0.551
R353 SD2L.n62 SD2L.t92 0.551
R354 SD2L.n62 SD2L.t96 0.551
R355 SD2L.n18 SD2L.t104 0.551
R356 SD2L.n18 SD2L.t84 0.551
R357 SD2L.n17 SD2L.t54 0.551
R358 SD2L.n17 SD2L.t64 0.551
R359 SD2L.n16 SD2L.t45 0.551
R360 SD2L.n16 SD2L.t51 0.551
R361 SD2L.n15 SD2L.t33 0.551
R362 SD2L.n15 SD2L.t13 0.551
R363 SD2L.n14 SD2L.t23 0.551
R364 SD2L.n14 SD2L.t3 0.551
R365 SD2L.n13 SD2L.t9 0.551
R366 SD2L.n13 SD2L.t106 0.551
R367 SD2L.n12 SD2L.t114 0.551
R368 SD2L.n12 SD2L.t95 0.551
R369 SD2L.n11 SD2L.t77 0.551
R370 SD2L.n11 SD2L.t90 0.551
R371 SD2L.n10 SD2L.t57 0.551
R372 SD2L.n10 SD2L.t66 0.551
R373 SD2L.n0 SD2L.t41 0.551
R374 SD2L.n0 SD2L.t55 0.551
R375 SD2L.n1 SD2L.t38 0.551
R376 SD2L.n1 SD2L.t17 0.551
R377 SD2L.n2 SD2L.t25 0.551
R378 SD2L.n2 SD2L.t119 0.551
R379 SD2L.n3 SD2L.t14 0.551
R380 SD2L.n3 SD2L.t108 0.551
R381 SD2L.n4 SD2L.t93 0.551
R382 SD2L.n4 SD2L.t99 0.551
R383 SD2L.n98 SD2L.t100 0.551
R384 SD2L.n98 SD2L.t7 0.551
R385 SD2L.n97 SD2L.t50 0.551
R386 SD2L.n97 SD2L.t58 0.551
R387 SD2L.n96 SD2L.t107 0.551
R388 SD2L.n96 SD2L.t26 0.551
R389 SD2L.n95 SD2L.t67 0.551
R390 SD2L.n95 SD2L.t79 0.551
R391 SD2L.n94 SD2L.t110 0.551
R392 SD2L.n94 SD2L.t36 0.551
R393 SD2L.n93 SD2L.t4 0.551
R394 SD2L.n93 SD2L.t47 0.551
R395 SD2L.n92 SD2L.t91 0.551
R396 SD2L.n92 SD2L.t0 0.551
R397 SD2L.n91 SD2L.t42 0.551
R398 SD2L.n91 SD2L.t48 0.551
R399 SD2L.n90 SD2L.t101 0.551
R400 SD2L.n90 SD2L.t105 0.551
R401 SD2L.n89 SD2L.t46 0.551
R402 SD2L.n89 SD2L.t97 0.551
R403 SD2L.n88 SD2L.t103 0.551
R404 SD2L.n88 SD2L.t30 0.551
R405 SD2L.n87 SD2L.t32 0.551
R406 SD2L.n87 SD2L.t112 0.551
R407 SD2L.n112 SD2L.t115 0.551
R408 SD2L.n112 SD2L.t31 0.551
R409 SD2L.n113 SD2L.t78 0.551
R410 SD2L.n113 SD2L.t86 0.551
R411 SD2L.n103 SD2L.t71 0.551
R412 SD2L.n103 SD2L.t118 0.551
R413 SD2L.n116 SD2L.n86 0.406
R414 SD2L.n118 SD2L.n28 0.406
R415 SD2L.n116 SD2L.n115 0.398
R416 SD2L.n117 SD2L.n57 0.297
R417 SD2L.n117 SD2L.n116 0.101
R418 SD2L.n118 SD2L.n117 0.097
R419 SD2L.n46 SD2L.n45 0.037
R420 SD2L.n47 SD2L.n46 0.037
R421 SD2L.n48 SD2L.n47 0.037
R422 SD2L.n49 SD2L.n48 0.037
R423 SD2L.n50 SD2L.n49 0.037
R424 SD2L.n51 SD2L.n50 0.037
R425 SD2L.n52 SD2L.n51 0.037
R426 SD2L.n53 SD2L.n52 0.037
R427 SD2L.n54 SD2L.n53 0.037
R428 SD2L.n55 SD2L.n54 0.037
R429 SD2L.n56 SD2L.n55 0.037
R430 SD2L.n78 SD2L.n77 0.037
R431 SD2L.n79 SD2L.n78 0.037
R432 SD2L.n80 SD2L.n79 0.037
R433 SD2L.n81 SD2L.n80 0.037
R434 SD2L.n82 SD2L.n81 0.037
R435 SD2L.n83 SD2L.n82 0.037
R436 SD2L.n84 SD2L.n83 0.037
R437 SD2L.n85 SD2L.n84 0.037
R438 SD2L.n67 SD2L.n66 0.037
R439 SD2L.n66 SD2L.n65 0.037
R440 SD2L.n65 SD2L.n64 0.037
R441 SD2L.n64 SD2L.n63 0.037
R442 SD2L.n20 SD2L.n19 0.037
R443 SD2L.n21 SD2L.n20 0.037
R444 SD2L.n22 SD2L.n21 0.037
R445 SD2L.n23 SD2L.n22 0.037
R446 SD2L.n24 SD2L.n23 0.037
R447 SD2L.n25 SD2L.n24 0.037
R448 SD2L.n26 SD2L.n25 0.037
R449 SD2L.n27 SD2L.n26 0.037
R450 SD2L.n9 SD2L.n8 0.037
R451 SD2L.n8 SD2L.n7 0.037
R452 SD2L.n7 SD2L.n6 0.037
R453 SD2L.n6 SD2L.n5 0.037
R454 SD2L.n100 SD2L.n99 0.037
R455 SD2L.n101 SD2L.n100 0.037
R456 SD2L.n102 SD2L.n101 0.037
R457 SD2L.n104 SD2L.n102 0.037
R458 SD2L.n105 SD2L.n104 0.037
R459 SD2L.n106 SD2L.n105 0.037
R460 SD2L.n107 SD2L.n106 0.037
R461 SD2L.n108 SD2L.n107 0.037
R462 SD2L.n109 SD2L.n108 0.037
R463 SD2L.n110 SD2L.n109 0.037
R464 SD2L.n111 SD2L.n110 0.037
R465 SD2L.n57 SD2L.n31 0.024
R466 SD2L.n115 SD2L.n114 0.024
R467 SD2L.n86 SD2L.n85 0.023
R468 SD2L.n28 SD2L.n27 0.023
R469 SD2L.n86 SD2L.n67 0.014
R470 SD2L.n28 SD2L.n9 0.014
R471 SD2L.n57 SD2L.n56 0.012
R472 SD2L.n115 SD2L.n111 0.012
R473 SD2L SD2L.n118 0.01
R474 SD1R.n57 SD1R.t81 2.284
R475 SD1R.n44 SD1R.t90 2.284
R476 SD1R.n86 SD1R.t14 2.284
R477 SD1R.n99 SD1R.t33 2.284
R478 SD1R.n60 SD1R.n59 1.74
R479 SD1R.n74 SD1R.n73 1.739
R480 SD1R.n20 SD1R.n19 1.739
R481 SD1R.n6 SD1R.n5 1.739
R482 SD1R.n74 SD1R.n72 1.702
R483 SD1R.n75 SD1R.n71 1.702
R484 SD1R.n76 SD1R.n70 1.702
R485 SD1R.n77 SD1R.n69 1.702
R486 SD1R.n78 SD1R.n68 1.702
R487 SD1R.n79 SD1R.n67 1.702
R488 SD1R.n81 SD1R.n65 1.702
R489 SD1R.n82 SD1R.n64 1.702
R490 SD1R.n83 SD1R.n63 1.702
R491 SD1R.n84 SD1R.n62 1.702
R492 SD1R.n0 SD1R.n61 1.702
R493 SD1R.n60 SD1R.n58 1.702
R494 SD1R.n20 SD1R.n18 1.702
R495 SD1R.n21 SD1R.n17 1.702
R496 SD1R.n22 SD1R.n16 1.702
R497 SD1R.n23 SD1R.n15 1.702
R498 SD1R.n24 SD1R.n14 1.702
R499 SD1R.n25 SD1R.n13 1.702
R500 SD1R.n27 SD1R.n11 1.702
R501 SD1R.n28 SD1R.n10 1.702
R502 SD1R.n29 SD1R.n9 1.702
R503 SD1R.n30 SD1R.n8 1.702
R504 SD1R.n1 SD1R.n7 1.702
R505 SD1R.n6 SD1R.n4 1.702
R506 SD1R.n57 SD1R.n56 1.696
R507 SD1R.n2 SD1R.n31 1.696
R508 SD1R.n55 SD1R.n32 1.696
R509 SD1R.n54 SD1R.n33 1.696
R510 SD1R.n53 SD1R.n34 1.696
R511 SD1R.n52 SD1R.n35 1.696
R512 SD1R.n51 SD1R.n36 1.696
R513 SD1R.n50 SD1R.n37 1.696
R514 SD1R.n49 SD1R.n38 1.696
R515 SD1R.n48 SD1R.n39 1.696
R516 SD1R.n47 SD1R.n40 1.696
R517 SD1R.n46 SD1R.n41 1.696
R518 SD1R.n45 SD1R.n42 1.696
R519 SD1R.n44 SD1R.n43 1.696
R520 SD1R.n86 SD1R.n85 1.696
R521 SD1R.n110 SD1R.n87 1.696
R522 SD1R.n109 SD1R.n88 1.696
R523 SD1R.n108 SD1R.n89 1.696
R524 SD1R.n107 SD1R.n90 1.696
R525 SD1R.n106 SD1R.n91 1.696
R526 SD1R.n105 SD1R.n92 1.696
R527 SD1R.n104 SD1R.n93 1.696
R528 SD1R.n103 SD1R.n94 1.696
R529 SD1R.n102 SD1R.n95 1.696
R530 SD1R.n101 SD1R.n96 1.696
R531 SD1R.n100 SD1R.n97 1.696
R532 SD1R.n99 SD1R.n98 1.696
R533 SD1R.n3 SD1R.n111 1.695
R534 SD1R.n80 SD1R.n66 1.678
R535 SD1R.n26 SD1R.n12 1.678
R536 SD1R.n112 SD1R.n3 0.571
R537 SD1R.n73 SD1R.t11 0.551
R538 SD1R.n73 SD1R.t37 0.551
R539 SD1R.n72 SD1R.t3 0.551
R540 SD1R.n72 SD1R.t84 0.551
R541 SD1R.n71 SD1R.t55 0.551
R542 SD1R.n71 SD1R.t28 0.551
R543 SD1R.n70 SD1R.t31 0.551
R544 SD1R.n70 SD1R.t39 0.551
R545 SD1R.n69 SD1R.t23 0.551
R546 SD1R.n69 SD1R.t113 0.551
R547 SD1R.n68 SD1R.t93 0.551
R548 SD1R.n68 SD1R.t67 0.551
R549 SD1R.n67 SD1R.t116 0.551
R550 SD1R.n67 SD1R.t115 0.551
R551 SD1R.n66 SD1R.t117 0.551
R552 SD1R.n66 SD1R.t110 0.551
R553 SD1R.n65 SD1R.t30 0.551
R554 SD1R.n65 SD1R.t118 0.551
R555 SD1R.n64 SD1R.t43 0.551
R556 SD1R.n64 SD1R.t95 0.551
R557 SD1R.n63 SD1R.t61 0.551
R558 SD1R.n63 SD1R.t18 0.551
R559 SD1R.n62 SD1R.t66 0.551
R560 SD1R.n62 SD1R.t45 0.551
R561 SD1R.n61 SD1R.t40 0.551
R562 SD1R.n61 SD1R.t19 0.551
R563 SD1R.n58 SD1R.t108 0.551
R564 SD1R.n58 SD1R.t50 0.551
R565 SD1R.n59 SD1R.t94 0.551
R566 SD1R.n59 SD1R.t83 0.551
R567 SD1R.n56 SD1R.t103 0.551
R568 SD1R.n56 SD1R.t70 0.551
R569 SD1R.n31 SD1R.t2 0.551
R570 SD1R.n31 SD1R.t98 0.551
R571 SD1R.n32 SD1R.t73 0.551
R572 SD1R.n32 SD1R.t5 0.551
R573 SD1R.n33 SD1R.t12 0.551
R574 SD1R.n33 SD1R.t24 0.551
R575 SD1R.n34 SD1R.t76 0.551
R576 SD1R.n34 SD1R.t51 0.551
R577 SD1R.n35 SD1R.t82 0.551
R578 SD1R.n35 SD1R.t114 0.551
R579 SD1R.n36 SD1R.t101 0.551
R580 SD1R.n36 SD1R.t38 0.551
R581 SD1R.n37 SD1R.t21 0.551
R582 SD1R.n37 SD1R.t89 0.551
R583 SD1R.n38 SD1R.t15 0.551
R584 SD1R.n38 SD1R.t96 0.551
R585 SD1R.n39 SD1R.t59 0.551
R586 SD1R.n39 SD1R.t13 0.551
R587 SD1R.n40 SD1R.t99 0.551
R588 SD1R.n40 SD1R.t36 0.551
R589 SD1R.n41 SD1R.t60 0.551
R590 SD1R.n41 SD1R.t25 0.551
R591 SD1R.n42 SD1R.t77 0.551
R592 SD1R.n42 SD1R.t111 0.551
R593 SD1R.n43 SD1R.t41 0.551
R594 SD1R.n43 SD1R.t44 0.551
R595 SD1R.n19 SD1R.t10 0.551
R596 SD1R.n19 SD1R.t34 0.551
R597 SD1R.n18 SD1R.t29 0.551
R598 SD1R.n18 SD1R.t109 0.551
R599 SD1R.n17 SD1R.t102 0.551
R600 SD1R.n17 SD1R.t80 0.551
R601 SD1R.n16 SD1R.t119 0.551
R602 SD1R.n16 SD1R.t53 0.551
R603 SD1R.n15 SD1R.t64 0.551
R604 SD1R.n15 SD1R.t65 0.551
R605 SD1R.n14 SD1R.t9 0.551
R606 SD1R.n14 SD1R.t20 0.551
R607 SD1R.n13 SD1R.t57 0.551
R608 SD1R.n13 SD1R.t58 0.551
R609 SD1R.n12 SD1R.t6 0.551
R610 SD1R.n12 SD1R.t87 0.551
R611 SD1R.n11 SD1R.t88 0.551
R612 SD1R.n11 SD1R.t4 0.551
R613 SD1R.n10 SD1R.t75 0.551
R614 SD1R.n10 SD1R.t105 0.551
R615 SD1R.n9 SD1R.t85 0.551
R616 SD1R.n9 SD1R.t62 0.551
R617 SD1R.n8 SD1R.t86 0.551
R618 SD1R.n8 SD1R.t68 0.551
R619 SD1R.n7 SD1R.t69 0.551
R620 SD1R.n7 SD1R.t112 0.551
R621 SD1R.n4 SD1R.t97 0.551
R622 SD1R.n4 SD1R.t22 0.551
R623 SD1R.n5 SD1R.t17 0.551
R624 SD1R.n5 SD1R.t8 0.551
R625 SD1R.n85 SD1R.t48 0.551
R626 SD1R.n85 SD1R.t26 0.551
R627 SD1R.n87 SD1R.t32 0.551
R628 SD1R.n87 SD1R.t100 0.551
R629 SD1R.n88 SD1R.t92 0.551
R630 SD1R.n88 SD1R.t1 0.551
R631 SD1R.n89 SD1R.t56 0.551
R632 SD1R.n89 SD1R.t91 0.551
R633 SD1R.n90 SD1R.t35 0.551
R634 SD1R.n90 SD1R.t27 0.551
R635 SD1R.n91 SD1R.t52 0.551
R636 SD1R.n91 SD1R.t107 0.551
R637 SD1R.n92 SD1R.t79 0.551
R638 SD1R.n92 SD1R.t104 0.551
R639 SD1R.n93 SD1R.t49 0.551
R640 SD1R.n93 SD1R.t106 0.551
R641 SD1R.n94 SD1R.t78 0.551
R642 SD1R.n94 SD1R.t7 0.551
R643 SD1R.n95 SD1R.t72 0.551
R644 SD1R.n95 SD1R.t74 0.551
R645 SD1R.n96 SD1R.t47 0.551
R646 SD1R.n96 SD1R.t54 0.551
R647 SD1R.n97 SD1R.t71 0.551
R648 SD1R.n97 SD1R.t42 0.551
R649 SD1R.n98 SD1R.t46 0.551
R650 SD1R.n98 SD1R.t63 0.551
R651 SD1R.n111 SD1R.t16 0.551
R652 SD1R.n111 SD1R.t0 0.551
R653 SD1R.n113 SD1R.n2 0.531
R654 SD1R.n113 SD1R.n112 0.162
R655 SD1R.n112 SD1R.n0 0.122
R656 SD1R.n114 SD1R.n1 0.118
R657 SD1R.n114 SD1R.n113 0.04
R658 SD1R.n75 SD1R.n74 0.037
R659 SD1R.n76 SD1R.n75 0.037
R660 SD1R.n77 SD1R.n76 0.037
R661 SD1R.n78 SD1R.n77 0.037
R662 SD1R.n79 SD1R.n78 0.037
R663 SD1R.n80 SD1R.n79 0.037
R664 SD1R.n81 SD1R.n80 0.037
R665 SD1R.n82 SD1R.n81 0.037
R666 SD1R.n83 SD1R.n82 0.037
R667 SD1R.n84 SD1R.n83 0.037
R668 SD1R.n0 SD1R.n84 0.037
R669 SD1R.n2 SD1R.n55 0.037
R670 SD1R.n55 SD1R.n54 0.037
R671 SD1R.n54 SD1R.n53 0.037
R672 SD1R.n53 SD1R.n52 0.037
R673 SD1R.n52 SD1R.n51 0.037
R674 SD1R.n51 SD1R.n50 0.037
R675 SD1R.n50 SD1R.n49 0.037
R676 SD1R.n49 SD1R.n48 0.037
R677 SD1R.n48 SD1R.n47 0.037
R678 SD1R.n47 SD1R.n46 0.037
R679 SD1R.n46 SD1R.n45 0.037
R680 SD1R.n45 SD1R.n44 0.037
R681 SD1R.n21 SD1R.n20 0.037
R682 SD1R.n22 SD1R.n21 0.037
R683 SD1R.n23 SD1R.n22 0.037
R684 SD1R.n24 SD1R.n23 0.037
R685 SD1R.n25 SD1R.n24 0.037
R686 SD1R.n26 SD1R.n25 0.037
R687 SD1R.n27 SD1R.n26 0.037
R688 SD1R.n28 SD1R.n27 0.037
R689 SD1R.n29 SD1R.n28 0.037
R690 SD1R.n30 SD1R.n29 0.037
R691 SD1R.n1 SD1R.n30 0.037
R692 SD1R SD1R.n114 0.037
R693 SD1R.n3 SD1R.n110 0.037
R694 SD1R.n110 SD1R.n109 0.037
R695 SD1R.n109 SD1R.n108 0.037
R696 SD1R.n108 SD1R.n107 0.037
R697 SD1R.n107 SD1R.n106 0.037
R698 SD1R.n106 SD1R.n105 0.037
R699 SD1R.n105 SD1R.n104 0.037
R700 SD1R.n104 SD1R.n103 0.037
R701 SD1R.n103 SD1R.n102 0.037
R702 SD1R.n102 SD1R.n101 0.037
R703 SD1R.n101 SD1R.n100 0.037
R704 SD1R.n100 SD1R.n99 0.037
R705 SD1R.n1 SD1R.n6 0.037
R706 SD1R.n0 SD1R.n60 0.037
R707 SD1R.n3 SD1R.n86 0.036
R708 SD1R.n2 SD1R.n57 0.036
R709 SD2R.n71 SD2R.t115 2.285
R710 SD2R.n85 SD2R.t16 2.284
R711 SD2R.n27 SD2R.t92 2.284
R712 SD2R.n13 SD2R.t68 2.284
R713 SD2R.n51 SD2R.n50 1.739
R714 SD2R.n37 SD2R.n36 1.739
R715 SD2R.n94 SD2R.n93 1.739
R716 SD2R.n107 SD2R.n106 1.739
R717 SD2R.n51 SD2R.n49 1.702
R718 SD2R.n52 SD2R.n48 1.702
R719 SD2R.n53 SD2R.n47 1.702
R720 SD2R.n54 SD2R.n46 1.702
R721 SD2R.n55 SD2R.n45 1.702
R722 SD2R.n56 SD2R.n44 1.702
R723 SD2R.n42 SD2R.n30 1.702
R724 SD2R.n41 SD2R.n31 1.702
R725 SD2R.n40 SD2R.n32 1.702
R726 SD2R.n39 SD2R.n33 1.702
R727 SD2R.n38 SD2R.n34 1.702
R728 SD2R.n37 SD2R.n35 1.702
R729 SD2R.n94 SD2R.n92 1.702
R730 SD2R.n95 SD2R.n91 1.702
R731 SD2R.n96 SD2R.n90 1.702
R732 SD2R.n97 SD2R.n89 1.702
R733 SD2R.n98 SD2R.n88 1.702
R734 SD2R.n99 SD2R.n87 1.702
R735 SD2R.n112 SD2R.n100 1.702
R736 SD2R.n111 SD2R.n101 1.702
R737 SD2R.n110 SD2R.n102 1.702
R738 SD2R.n109 SD2R.n103 1.702
R739 SD2R.n108 SD2R.n104 1.702
R740 SD2R.n107 SD2R.n105 1.702
R741 SD2R.n85 SD2R.n84 1.696
R742 SD2R.n83 SD2R.n58 1.696
R743 SD2R.n82 SD2R.n59 1.696
R744 SD2R.n81 SD2R.n60 1.696
R745 SD2R.n80 SD2R.n61 1.696
R746 SD2R.n79 SD2R.n62 1.696
R747 SD2R.n78 SD2R.n63 1.696
R748 SD2R.n77 SD2R.n64 1.696
R749 SD2R.n76 SD2R.n65 1.696
R750 SD2R.n75 SD2R.n66 1.696
R751 SD2R.n74 SD2R.n67 1.696
R752 SD2R.n73 SD2R.n68 1.696
R753 SD2R.n72 SD2R.n69 1.696
R754 SD2R.n71 SD2R.n70 1.696
R755 SD2R.n27 SD2R.n26 1.696
R756 SD2R.n25 SD2R.n0 1.696
R757 SD2R.n24 SD2R.n1 1.696
R758 SD2R.n23 SD2R.n2 1.696
R759 SD2R.n22 SD2R.n3 1.696
R760 SD2R.n21 SD2R.n4 1.696
R761 SD2R.n20 SD2R.n5 1.696
R762 SD2R.n19 SD2R.n6 1.696
R763 SD2R.n18 SD2R.n7 1.696
R764 SD2R.n17 SD2R.n8 1.696
R765 SD2R.n16 SD2R.n9 1.696
R766 SD2R.n15 SD2R.n10 1.696
R767 SD2R.n14 SD2R.n11 1.696
R768 SD2R.n13 SD2R.n12 1.696
R769 SD2R.n43 SD2R.n29 1.678
R770 SD2R.n114 SD2R.n113 1.677
R771 SD2R.n84 SD2R.t23 0.551
R772 SD2R.n84 SD2R.t35 0.551
R773 SD2R.n58 SD2R.t12 0.551
R774 SD2R.n58 SD2R.t113 0.551
R775 SD2R.n59 SD2R.t90 0.551
R776 SD2R.n59 SD2R.t99 0.551
R777 SD2R.n60 SD2R.t73 0.551
R778 SD2R.n60 SD2R.t84 0.551
R779 SD2R.n61 SD2R.t94 0.551
R780 SD2R.n61 SD2R.t43 0.551
R781 SD2R.n62 SD2R.t51 0.551
R782 SD2R.n62 SD2R.t30 0.551
R783 SD2R.n63 SD2R.t40 0.551
R784 SD2R.n63 SD2R.t46 0.551
R785 SD2R.n64 SD2R.t26 0.551
R786 SD2R.n64 SD2R.t3 0.551
R787 SD2R.n65 SD2R.t101 0.551
R788 SD2R.n65 SD2R.t111 0.551
R789 SD2R.n66 SD2R.t86 0.551
R790 SD2R.n66 SD2R.t98 0.551
R791 SD2R.n67 SD2R.t106 0.551
R792 SD2R.n67 SD2R.t81 0.551
R793 SD2R.n68 SD2R.t63 0.551
R794 SD2R.n68 SD2R.t41 0.551
R795 SD2R.n69 SD2R.t49 0.551
R796 SD2R.n69 SD2R.t28 0.551
R797 SD2R.n70 SD2R.t38 0.551
R798 SD2R.n70 SD2R.t44 0.551
R799 SD2R.n50 SD2R.t78 0.551
R800 SD2R.n50 SD2R.t7 0.551
R801 SD2R.n49 SD2R.t53 0.551
R802 SD2R.n49 SD2R.t60 0.551
R803 SD2R.n48 SD2R.t107 0.551
R804 SD2R.n48 SD2R.t21 0.551
R805 SD2R.n47 SD2R.t56 0.551
R806 SD2R.n47 SD2R.t62 0.551
R807 SD2R.n46 SD2R.t112 0.551
R808 SD2R.n46 SD2R.t36 0.551
R809 SD2R.n45 SD2R.t69 0.551
R810 SD2R.n45 SD2R.t0 0.551
R811 SD2R.n44 SD2R.t114 0.551
R812 SD2R.n44 SD2R.t39 0.551
R813 SD2R.n29 SD2R.t80 0.551
R814 SD2R.n29 SD2R.t2 0.551
R815 SD2R.n30 SD2R.t47 0.551
R816 SD2R.n30 SD2R.t50 0.551
R817 SD2R.n31 SD2R.t85 0.551
R818 SD2R.n31 SD2R.t88 0.551
R819 SD2R.n32 SD2R.t48 0.551
R820 SD2R.n32 SD2R.t96 0.551
R821 SD2R.n33 SD2R.t100 0.551
R822 SD2R.n33 SD2R.t24 0.551
R823 SD2R.n34 SD2R.t33 0.551
R824 SD2R.n34 SD2R.t97 0.551
R825 SD2R.n35 SD2R.t102 0.551
R826 SD2R.n35 SD2R.t27 0.551
R827 SD2R.n36 SD2R.t72 0.551
R828 SD2R.n36 SD2R.t77 0.551
R829 SD2R.n26 SD2R.t70 0.551
R830 SD2R.n26 SD2R.t75 0.551
R831 SD2R.n0 SD2R.t57 0.551
R832 SD2R.n0 SD2R.t64 0.551
R833 SD2R.n1 SD2R.t45 0.551
R834 SD2R.n1 SD2R.t54 0.551
R835 SD2R.n2 SD2R.t31 0.551
R836 SD2R.n2 SD2R.t8 0.551
R837 SD2R.n3 SD2R.t15 0.551
R838 SD2R.n3 SD2R.t1 0.551
R839 SD2R.n4 SD2R.t6 0.551
R840 SD2R.n4 SD2R.t105 0.551
R841 SD2R.n5 SD2R.t116 0.551
R842 SD2R.n5 SD2R.t89 0.551
R843 SD2R.n6 SD2R.t71 0.551
R844 SD2R.n6 SD2R.t76 0.551
R845 SD2R.n7 SD2R.t58 0.551
R846 SD2R.n7 SD2R.t66 0.551
R847 SD2R.n8 SD2R.t42 0.551
R848 SD2R.n8 SD2R.t22 0.551
R849 SD2R.n9 SD2R.t34 0.551
R850 SD2R.n9 SD2R.t11 0.551
R851 SD2R.n10 SD2R.t18 0.551
R852 SD2R.n10 SD2R.t119 0.551
R853 SD2R.n11 SD2R.t9 0.551
R854 SD2R.n11 SD2R.t108 0.551
R855 SD2R.n12 SD2R.t83 0.551
R856 SD2R.n12 SD2R.t93 0.551
R857 SD2R.n93 SD2R.t5 0.551
R858 SD2R.n93 SD2R.t52 0.551
R859 SD2R.n92 SD2R.t87 0.551
R860 SD2R.n92 SD2R.t91 0.551
R861 SD2R.n91 SD2R.t17 0.551
R862 SD2R.n91 SD2R.t55 0.551
R863 SD2R.n90 SD2R.t103 0.551
R864 SD2R.n90 SD2R.t109 0.551
R865 SD2R.n89 SD2R.t19 0.551
R866 SD2R.n89 SD2R.t67 0.551
R867 SD2R.n88 SD2R.t104 0.551
R868 SD2R.n88 SD2R.t29 0.551
R869 SD2R.n87 SD2R.t37 0.551
R870 SD2R.n87 SD2R.t79 0.551
R871 SD2R.n100 SD2R.t74 0.551
R872 SD2R.n100 SD2R.t82 0.551
R873 SD2R.n101 SD2R.t10 0.551
R874 SD2R.n101 SD2R.t14 0.551
R875 SD2R.n102 SD2R.t95 0.551
R876 SD2R.n102 SD2R.t4 0.551
R877 SD2R.n103 SD2R.t13 0.551
R878 SD2R.n103 SD2R.t59 0.551
R879 SD2R.n104 SD2R.t65 0.551
R880 SD2R.n104 SD2R.t20 0.551
R881 SD2R.n105 SD2R.t25 0.551
R882 SD2R.n105 SD2R.t61 0.551
R883 SD2R.n106 SD2R.t110 0.551
R884 SD2R.n106 SD2R.t117 0.551
R885 SD2R.n113 SD2R.t118 0.551
R886 SD2R.n113 SD2R.t32 0.551
R887 SD2R.n116 SD2R.n115 0.335
R888 SD2R.n116 SD2R.n86 0.27
R889 SD2R.n118 SD2R.n28 0.27
R890 SD2R.n117 SD2R.n57 0.203
R891 SD2R.n118 SD2R.n117 0.099
R892 SD2R.n117 SD2R.n116 0.07
R893 SD2R SD2R.n118 0.042
R894 SD2R.n83 SD2R.n82 0.037
R895 SD2R.n82 SD2R.n81 0.037
R896 SD2R.n81 SD2R.n80 0.037
R897 SD2R.n80 SD2R.n79 0.037
R898 SD2R.n79 SD2R.n78 0.037
R899 SD2R.n78 SD2R.n77 0.037
R900 SD2R.n77 SD2R.n76 0.037
R901 SD2R.n76 SD2R.n75 0.037
R902 SD2R.n75 SD2R.n74 0.037
R903 SD2R.n74 SD2R.n73 0.037
R904 SD2R.n73 SD2R.n72 0.037
R905 SD2R.n72 SD2R.n71 0.037
R906 SD2R.n52 SD2R.n51 0.037
R907 SD2R.n53 SD2R.n52 0.037
R908 SD2R.n54 SD2R.n53 0.037
R909 SD2R.n55 SD2R.n54 0.037
R910 SD2R.n56 SD2R.n55 0.037
R911 SD2R.n43 SD2R.n42 0.037
R912 SD2R.n42 SD2R.n41 0.037
R913 SD2R.n41 SD2R.n40 0.037
R914 SD2R.n40 SD2R.n39 0.037
R915 SD2R.n39 SD2R.n38 0.037
R916 SD2R.n38 SD2R.n37 0.037
R917 SD2R.n25 SD2R.n24 0.037
R918 SD2R.n24 SD2R.n23 0.037
R919 SD2R.n23 SD2R.n22 0.037
R920 SD2R.n22 SD2R.n21 0.037
R921 SD2R.n21 SD2R.n20 0.037
R922 SD2R.n20 SD2R.n19 0.037
R923 SD2R.n19 SD2R.n18 0.037
R924 SD2R.n18 SD2R.n17 0.037
R925 SD2R.n17 SD2R.n16 0.037
R926 SD2R.n16 SD2R.n15 0.037
R927 SD2R.n15 SD2R.n14 0.037
R928 SD2R.n14 SD2R.n13 0.037
R929 SD2R.n95 SD2R.n94 0.037
R930 SD2R.n96 SD2R.n95 0.037
R931 SD2R.n97 SD2R.n96 0.037
R932 SD2R.n98 SD2R.n97 0.037
R933 SD2R.n99 SD2R.n98 0.037
R934 SD2R.n114 SD2R.n112 0.037
R935 SD2R.n112 SD2R.n111 0.037
R936 SD2R.n111 SD2R.n110 0.037
R937 SD2R.n110 SD2R.n109 0.037
R938 SD2R.n109 SD2R.n108 0.037
R939 SD2R.n108 SD2R.n107 0.037
R940 SD2R.n86 SD2R.n85 0.032
R941 SD2R.n28 SD2R.n27 0.032
R942 SD2R.n57 SD2R.n56 0.027
R943 SD2R.n115 SD2R.n99 0.027
R944 SD2R.n57 SD2R.n43 0.009
R945 SD2R.n115 SD2R.n114 0.009
R946 SD2R.n86 SD2R.n83 0.004
R947 SD2R.n28 SD2R.n25 0.004
C15 SD1R SUB 101.39fF
C16 SD2R SUB 87.52fF
C17 GR SUB 104.85fF $ **FLOATING
C18 SD1L SUB 80.03fF
C19 SD2L SUB 64.98fF
C20 GL SUB 104.15fF $ **FLOATING
C21 SD2R.n0 SUB 10.65fF
C22 SD2R.n1 SUB 10.65fF
C23 SD2R.n2 SUB 10.65fF
C24 SD2R.n3 SUB 10.65fF
C25 SD2R.n4 SUB 10.65fF
C26 SD2R.n5 SUB 10.65fF
C27 SD2R.n6 SUB 10.65fF
C28 SD2R.n7 SUB 10.65fF
C29 SD2R.n8 SUB 10.65fF
C30 SD2R.n9 SUB 10.65fF
C31 SD2R.n10 SUB 10.65fF
C32 SD2R.n11 SUB 10.65fF
C33 SD2R.n12 SUB 10.65fF
C34 SD2R.t68 SUB 9.20fF $ **FLOATING
C35 SD2R.n13 SUB 5.48fF
C36 SD2R.n14 SUB 1.56fF
C37 SD2R.n15 SUB 1.56fF
C38 SD2R.n16 SUB 1.56fF
C39 SD2R.n17 SUB 1.56fF
C40 SD2R.n18 SUB 1.56fF
C41 SD2R.n19 SUB 1.56fF
C42 SD2R.n20 SUB 1.56fF
C43 SD2R.n21 SUB 1.56fF
C44 SD2R.n22 SUB 1.56fF
C45 SD2R.n23 SUB 1.56fF
C46 SD2R.n24 SUB 1.56fF
C47 SD2R.n25 SUB 1.17fF
C48 SD2R.n26 SUB 10.65fF
C49 SD2R.t92 SUB 9.20fF $ **FLOATING
C50 SD2R.n27 SUB 5.42fF
C51 SD2R.n28 SUB 48.30fF
C52 SD2R.n29 SUB 10.68fF
C53 SD2R.n30 SUB 10.65fF
C54 SD2R.n31 SUB 10.65fF
C55 SD2R.n32 SUB 10.65fF
C56 SD2R.n33 SUB 10.65fF
C57 SD2R.n34 SUB 10.65fF
C58 SD2R.n35 SUB 10.65fF
C59 SD2R.n36 SUB 10.69fF
C60 SD2R.n37 SUB 3.20fF
C61 SD2R.n38 SUB 1.56fF
C62 SD2R.n39 SUB 1.56fF
C63 SD2R.n40 SUB 1.56fF
C64 SD2R.n41 SUB 1.56fF
C65 SD2R.n42 SUB 1.56fF
C66 SD2R.n43 SUB 1.23fF
C67 SD2R.n44 SUB 10.65fF
C68 SD2R.n45 SUB 10.65fF
C69 SD2R.n46 SUB 10.65fF
C70 SD2R.n47 SUB 10.65fF
C71 SD2R.n48 SUB 10.65fF
C72 SD2R.n49 SUB 10.65fF
C73 SD2R.n50 SUB 10.69fF
C74 SD2R.n51 SUB 3.20fF
C75 SD2R.n52 SUB 1.56fF
C76 SD2R.n53 SUB 1.56fF
C77 SD2R.n54 SUB 1.56fF
C78 SD2R.n55 SUB 1.56fF
C79 SD2R.n56 SUB 1.45fF
C80 SD2R.n57 SUB 37.17fF
C81 SD2R.n58 SUB 10.65fF
C82 SD2R.n59 SUB 10.65fF
C83 SD2R.n60 SUB 10.65fF
C84 SD2R.n61 SUB 10.65fF
C85 SD2R.n62 SUB 10.65fF
C86 SD2R.n63 SUB 10.65fF
C87 SD2R.n64 SUB 10.65fF
C88 SD2R.n65 SUB 10.65fF
C89 SD2R.n66 SUB 10.65fF
C90 SD2R.n67 SUB 10.65fF
C91 SD2R.n68 SUB 10.65fF
C92 SD2R.n69 SUB 10.65fF
C93 SD2R.n70 SUB 10.65fF
C94 SD2R.t115 SUB 9.21fF $ **FLOATING
C95 SD2R.n71 SUB 5.48fF
C96 SD2R.n72 SUB 1.56fF
C97 SD2R.n73 SUB 1.56fF
C98 SD2R.n74 SUB 1.56fF
C99 SD2R.n75 SUB 1.56fF
C100 SD2R.n76 SUB 1.56fF
C101 SD2R.n77 SUB 1.56fF
C102 SD2R.n78 SUB 1.56fF
C103 SD2R.n79 SUB 1.56fF
C104 SD2R.n80 SUB 1.56fF
C105 SD2R.n81 SUB 1.56fF
C106 SD2R.n82 SUB 1.56fF
C107 SD2R.n83 SUB 1.17fF
C108 SD2R.n84 SUB 10.65fF
C109 SD2R.t16 SUB 9.20fF $ **FLOATING
C110 SD2R.n85 SUB 5.42fF
C111 SD2R.n86 SUB 49.05fF
C112 SD2R.n87 SUB 10.65fF
C113 SD2R.n88 SUB 10.65fF
C114 SD2R.n89 SUB 10.65fF
C115 SD2R.n90 SUB 10.65fF
C116 SD2R.n91 SUB 10.65fF
C117 SD2R.n92 SUB 10.65fF
C118 SD2R.n93 SUB 10.69fF
C119 SD2R.n94 SUB 3.20fF
C120 SD2R.n95 SUB 1.56fF
C121 SD2R.n96 SUB 1.56fF
C122 SD2R.n97 SUB 1.56fF
C123 SD2R.n98 SUB 1.56fF
C124 SD2R.n99 SUB 1.45fF
C125 SD2R.n100 SUB 10.65fF
C126 SD2R.n101 SUB 10.65fF
C127 SD2R.n102 SUB 10.65fF
C128 SD2R.n103 SUB 10.65fF
C129 SD2R.n104 SUB 10.65fF
C130 SD2R.n105 SUB 10.65fF
C131 SD2R.n106 SUB 10.69fF
C132 SD2R.n107 SUB 3.20fF
C133 SD2R.n108 SUB 1.56fF
C134 SD2R.n109 SUB 1.56fF
C135 SD2R.n110 SUB 1.56fF
C136 SD2R.n111 SUB 1.56fF
C137 SD2R.n112 SUB 1.56fF
C138 SD2R.n113 SUB 10.68fF
C139 SD2R.n114 SUB 1.23fF
C140 SD2R.n115 SUB 79.64fF
C141 SD2R.n116 SUB 203.53fF
C142 SD2R.n117 SUB 113.29fF
C143 SD2R.n118 SUB 155.86fF
C144 SD1R.n0 SUB 24.36fF
C145 SD1R.n1 SUB 24.59fF
C146 SD1R.n2 SUB 93.32fF
C147 SD1R.n3 SUB 102.07fF
C148 SD1R.n4 SUB 10.44fF
C149 SD1R.n5 SUB 10.47fF
C150 SD1R.n6 SUB 2.97fF
C151 SD1R.n7 SUB 10.44fF
C152 SD1R.n8 SUB 10.44fF
C153 SD1R.n9 SUB 10.44fF
C154 SD1R.n10 SUB 10.44fF
C155 SD1R.n11 SUB 10.44fF
C156 SD1R.n12 SUB 10.47fF
C157 SD1R.n13 SUB 10.44fF
C158 SD1R.n14 SUB 10.44fF
C159 SD1R.n15 SUB 10.44fF
C160 SD1R.n16 SUB 10.44fF
C161 SD1R.n17 SUB 10.44fF
C162 SD1R.n18 SUB 10.44fF
C163 SD1R.n19 SUB 10.47fF
C164 SD1R.n20 SUB 3.14fF
C165 SD1R.n21 SUB 1.53fF
C166 SD1R.n22 SUB 1.53fF
C167 SD1R.n23 SUB 1.53fF
C168 SD1R.n24 SUB 1.53fF
C169 SD1R.n25 SUB 1.53fF
C170 SD1R.n26 SUB 1.54fF
C171 SD1R.n27 SUB 1.53fF
C172 SD1R.n28 SUB 1.53fF
C173 SD1R.n29 SUB 1.53fF
C174 SD1R.n30 SUB 1.53fF
C175 SD1R.n31 SUB 10.44fF
C176 SD1R.n32 SUB 10.44fF
C177 SD1R.n33 SUB 10.44fF
C178 SD1R.n34 SUB 10.44fF
C179 SD1R.n35 SUB 10.44fF
C180 SD1R.n36 SUB 10.44fF
C181 SD1R.n37 SUB 10.44fF
C182 SD1R.n38 SUB 10.44fF
C183 SD1R.n39 SUB 10.44fF
C184 SD1R.n40 SUB 10.44fF
C185 SD1R.n41 SUB 10.44fF
C186 SD1R.n42 SUB 10.44fF
C187 SD1R.n43 SUB 10.44fF
C188 SD1R.t90 SUB 9.02fF $ **FLOATING
C189 SD1R.n44 SUB 5.37fF
C190 SD1R.n45 SUB 1.53fF
C191 SD1R.n46 SUB 1.53fF
C192 SD1R.n47 SUB 1.53fF
C193 SD1R.n48 SUB 1.53fF
C194 SD1R.n49 SUB 1.53fF
C195 SD1R.n50 SUB 1.53fF
C196 SD1R.n51 SUB 1.53fF
C197 SD1R.n52 SUB 1.53fF
C198 SD1R.n53 SUB 1.53fF
C199 SD1R.n54 SUB 1.53fF
C200 SD1R.n55 SUB 1.53fF
C201 SD1R.n56 SUB 10.44fF
C202 SD1R.t81 SUB 9.02fF $ **FLOATING
C203 SD1R.n57 SUB 5.31fF
C204 SD1R.n58 SUB 10.44fF
C205 SD1R.n59 SUB 10.48fF
C206 SD1R.n60 SUB 2.97fF
C207 SD1R.n61 SUB 10.44fF
C208 SD1R.n62 SUB 10.44fF
C209 SD1R.n63 SUB 10.44fF
C210 SD1R.n64 SUB 10.44fF
C211 SD1R.n65 SUB 10.44fF
C212 SD1R.n66 SUB 10.47fF
C213 SD1R.n67 SUB 10.44fF
C214 SD1R.n68 SUB 10.44fF
C215 SD1R.n69 SUB 10.44fF
C216 SD1R.n70 SUB 10.44fF
C217 SD1R.n71 SUB 10.44fF
C218 SD1R.n72 SUB 10.44fF
C219 SD1R.n73 SUB 10.47fF
C220 SD1R.n74 SUB 3.14fF
C221 SD1R.n75 SUB 1.53fF
C222 SD1R.n76 SUB 1.53fF
C223 SD1R.n77 SUB 1.53fF
C224 SD1R.n78 SUB 1.53fF
C225 SD1R.n79 SUB 1.53fF
C226 SD1R.n80 SUB 1.54fF
C227 SD1R.n81 SUB 1.53fF
C228 SD1R.n82 SUB 1.53fF
C229 SD1R.n83 SUB 1.53fF
C230 SD1R.n84 SUB 1.53fF
C231 SD1R.n85 SUB 10.44fF
C232 SD1R.t14 SUB 9.02fF $ **FLOATING
C233 SD1R.n86 SUB 5.31fF
C234 SD1R.n87 SUB 10.44fF
C235 SD1R.n88 SUB 10.44fF
C236 SD1R.n89 SUB 10.44fF
C237 SD1R.n90 SUB 10.44fF
C238 SD1R.n91 SUB 10.44fF
C239 SD1R.n92 SUB 10.44fF
C240 SD1R.n93 SUB 10.44fF
C241 SD1R.n94 SUB 10.44fF
C242 SD1R.n95 SUB 10.44fF
C243 SD1R.n96 SUB 10.44fF
C244 SD1R.n97 SUB 10.44fF
C245 SD1R.n98 SUB 10.44fF
C246 SD1R.t33 SUB 9.02fF $ **FLOATING
C247 SD1R.n99 SUB 5.37fF
C248 SD1R.n100 SUB 1.53fF
C249 SD1R.n101 SUB 1.53fF
C250 SD1R.n102 SUB 1.53fF
C251 SD1R.n103 SUB 1.53fF
C252 SD1R.n104 SUB 1.53fF
C253 SD1R.n105 SUB 1.53fF
C254 SD1R.n106 SUB 1.53fF
C255 SD1R.n107 SUB 1.53fF
C256 SD1R.n108 SUB 1.53fF
C257 SD1R.n109 SUB 1.53fF
C258 SD1R.n110 SUB 1.53fF
C259 SD1R.n111 SUB 10.44fF
C260 SD1R.n112 SUB 226.54fF
C261 SD1R.n113 SUB 179.58fF
C262 SD1R.n114 SUB 66.51fF
C263 SD2L.n0 SUB 10.27fF
C264 SD2L.n1 SUB 10.27fF
C265 SD2L.n2 SUB 10.27fF
C266 SD2L.n3 SUB 10.27fF
C267 SD2L.n4 SUB 10.27fF
C268 SD2L.t72 SUB 8.88fF $ **FLOATING
C269 SD2L.n5 SUB 5.28fF
C270 SD2L.n6 SUB 1.51fF
C271 SD2L.n7 SUB 1.51fF
C272 SD2L.n8 SUB 1.51fF
C273 SD2L.n9 SUB 1.23fF
C274 SD2L.n10 SUB 10.27fF
C275 SD2L.n11 SUB 10.27fF
C276 SD2L.n12 SUB 10.27fF
C277 SD2L.n13 SUB 10.27fF
C278 SD2L.n14 SUB 10.27fF
C279 SD2L.n15 SUB 10.27fF
C280 SD2L.n16 SUB 10.27fF
C281 SD2L.n17 SUB 10.27fF
C282 SD2L.n18 SUB 10.27fF
C283 SD2L.t98 SUB 8.88fF $ **FLOATING
C284 SD2L.n19 SUB 5.29fF
C285 SD2L.n20 SUB 1.51fF
C286 SD2L.n21 SUB 1.51fF
C287 SD2L.n22 SUB 1.51fF
C288 SD2L.n23 SUB 1.51fF
C289 SD2L.n24 SUB 1.51fF
C290 SD2L.n25 SUB 1.51fF
C291 SD2L.n26 SUB 1.51fF
C292 SD2L.n27 SUB 1.34fF
C293 SD2L.n28 SUB 63.20fF
C294 SD2L.n29 SUB 10.27fF
C295 SD2L.n30 SUB 10.31fF
C296 SD2L.n31 SUB 2.94fF
C297 SD2L.n32 SUB 10.27fF
C298 SD2L.n33 SUB 10.27fF
C299 SD2L.n34 SUB 10.27fF
C300 SD2L.n35 SUB 10.27fF
C301 SD2L.n36 SUB 10.27fF
C302 SD2L.n37 SUB 10.30fF
C303 SD2L.n38 SUB 10.27fF
C304 SD2L.n39 SUB 10.27fF
C305 SD2L.n40 SUB 10.27fF
C306 SD2L.n41 SUB 10.27fF
C307 SD2L.n42 SUB 10.27fF
C308 SD2L.n43 SUB 10.27fF
C309 SD2L.n44 SUB 10.31fF
C310 SD2L.n45 SUB 3.09fF
C311 SD2L.n46 SUB 1.51fF
C312 SD2L.n47 SUB 1.51fF
C313 SD2L.n48 SUB 1.51fF
C314 SD2L.n49 SUB 1.51fF
C315 SD2L.n50 SUB 1.51fF
C316 SD2L.n51 SUB 1.52fF
C317 SD2L.n52 SUB 1.51fF
C318 SD2L.n53 SUB 1.51fF
C319 SD2L.n54 SUB 1.51fF
C320 SD2L.n55 SUB 1.51fF
C321 SD2L.n56 SUB 1.22fF
C322 SD2L.n57 SUB 51.84fF
C323 SD2L.n58 SUB 10.27fF
C324 SD2L.n59 SUB 10.27fF
C325 SD2L.n60 SUB 10.27fF
C326 SD2L.n61 SUB 10.27fF
C327 SD2L.n62 SUB 10.27fF
C328 SD2L.t69 SUB 8.88fF $ **FLOATING
C329 SD2L.n63 SUB 5.29fF
C330 SD2L.n64 SUB 1.51fF
C331 SD2L.n65 SUB 1.51fF
C332 SD2L.n66 SUB 1.51fF
C333 SD2L.n67 SUB 1.23fF
C334 SD2L.n68 SUB 10.27fF
C335 SD2L.n69 SUB 10.27fF
C336 SD2L.n70 SUB 10.27fF
C337 SD2L.n71 SUB 10.27fF
C338 SD2L.n72 SUB 10.27fF
C339 SD2L.n73 SUB 10.27fF
C340 SD2L.n74 SUB 10.27fF
C341 SD2L.n75 SUB 10.27fF
C342 SD2L.n76 SUB 10.27fF
C343 SD2L.t61 SUB 8.88fF $ **FLOATING
C344 SD2L.n77 SUB 5.29fF
C345 SD2L.n78 SUB 1.51fF
C346 SD2L.n79 SUB 1.51fF
C347 SD2L.n80 SUB 1.51fF
C348 SD2L.n81 SUB 1.51fF
C349 SD2L.n82 SUB 1.51fF
C350 SD2L.n83 SUB 1.51fF
C351 SD2L.n84 SUB 1.51fF
C352 SD2L.n85 SUB 1.34fF
C353 SD2L.n86 SUB 63.20fF
C354 SD2L.n87 SUB 10.27fF
C355 SD2L.n88 SUB 10.27fF
C356 SD2L.n89 SUB 10.27fF
C357 SD2L.n90 SUB 10.27fF
C358 SD2L.n91 SUB 10.27fF
C359 SD2L.n92 SUB 10.30fF
C360 SD2L.n93 SUB 10.27fF
C361 SD2L.n94 SUB 10.27fF
C362 SD2L.n95 SUB 10.27fF
C363 SD2L.n96 SUB 10.27fF
C364 SD2L.n97 SUB 10.27fF
C365 SD2L.n98 SUB 10.31fF
C366 SD2L.n99 SUB 3.09fF
C367 SD2L.n100 SUB 1.51fF
C368 SD2L.n101 SUB 1.51fF
C369 SD2L.n102 SUB 1.51fF
C370 SD2L.n103 SUB 10.28fF
C371 SD2L.n104 SUB 1.50fF
C372 SD2L.n105 SUB 1.51fF
C373 SD2L.n106 SUB 1.52fF
C374 SD2L.n107 SUB 1.51fF
C375 SD2L.n108 SUB 1.51fF
C376 SD2L.n109 SUB 1.51fF
C377 SD2L.n110 SUB 1.51fF
C378 SD2L.n111 SUB 1.22fF
C379 SD2L.n112 SUB 10.27fF
C380 SD2L.n113 SUB 10.31fF
C381 SD2L.n114 SUB 2.94fF
C382 SD2L.n115 SUB 79.17fF
C383 SD2L.n116 SUB 235.82fF
C384 SD2L.n117 SUB 137.14fF
C385 SD2L.n118 SUB 124.69fF
C386 SD1L.n0 SUB 78.95fF
C387 SD1L.n1 SUB 113.01fF
C388 SD1L.n2 SUB 10.89fF
C389 SD1L.n3 SUB 10.49fF
C390 SD1L.n4 SUB 10.60fF
C391 SD1L.n5 SUB 10.60fF
C392 SD1L.n6 SUB 10.60fF
C393 SD1L.n7 SUB 10.60fF
C394 SD1L.n8 SUB 10.60fF
C395 SD1L.n9 SUB 10.60fF
C396 SD1L.n10 SUB 10.60fF
C397 SD1L.t73 SUB 9.16fF $ **FLOATING
C398 SD1L.n11 SUB 5.46fF
C399 SD1L.n12 SUB 1.55fF
C400 SD1L.n13 SUB 1.55fF
C401 SD1L.n14 SUB 1.55fF
C402 SD1L.n15 SUB 1.55fF
C403 SD1L.n16 SUB 1.55fF
C404 SD1L.n17 SUB 1.44fF
C405 SD1L.n18 SUB 10.60fF
C406 SD1L.n19 SUB 10.60fF
C407 SD1L.n20 SUB 10.60fF
C408 SD1L.n21 SUB 10.60fF
C409 SD1L.n22 SUB 10.60fF
C410 SD1L.n23 SUB 10.60fF
C411 SD1L.n24 SUB 10.60fF
C412 SD1L.t35 SUB 9.16fF $ **FLOATING
C413 SD1L.n25 SUB 5.46fF
C414 SD1L.n26 SUB 1.55fF
C415 SD1L.n27 SUB 1.55fF
C416 SD1L.n28 SUB 1.55fF
C417 SD1L.n29 SUB 1.55fF
C418 SD1L.n30 SUB 1.55fF
C419 SD1L.n31 SUB 10.60fF
C420 SD1L.n32 SUB 10.60fF
C421 SD1L.n33 SUB 10.60fF
C422 SD1L.n34 SUB 10.60fF
C423 SD1L.n35 SUB 10.64fF
C424 SD1L.n36 SUB 3.19fF
C425 SD1L.n37 SUB 1.55fF
C426 SD1L.n38 SUB 1.55fF
C427 SD1L.n39 SUB 1.53fF
C428 SD1L.n40 SUB 10.60fF
C429 SD1L.n41 SUB 10.60fF
C430 SD1L.n42 SUB 10.63fF
C431 SD1L.n43 SUB 10.60fF
C432 SD1L.n44 SUB 10.60fF
C433 SD1L.n45 SUB 10.60fF
C434 SD1L.n46 SUB 10.60fF
C435 SD1L.n47 SUB 10.60fF
C436 SD1L.n48 SUB 10.60fF
C437 SD1L.n49 SUB 10.64fF
C438 SD1L.n50 SUB 3.19fF
C439 SD1L.n51 SUB 1.55fF
C440 SD1L.n52 SUB 1.55fF
C441 SD1L.n53 SUB 1.55fF
C442 SD1L.n54 SUB 1.55fF
C443 SD1L.n55 SUB 1.55fF
C444 SD1L.n56 SUB 1.56fF
C445 SD1L.n57 SUB 1.55fF
C446 SD1L.n58 SUB 10.60fF
C447 SD1L.n59 SUB 10.60fF
C448 SD1L.n60 SUB 10.60fF
C449 SD1L.n61 SUB 10.60fF
C450 SD1L.n62 SUB 10.60fF
C451 SD1L.n63 SUB 10.60fF
C452 SD1L.n64 SUB 10.60fF
C453 SD1L.t115 SUB 9.16fF $ **FLOATING
C454 SD1L.n65 SUB 5.46fF
C455 SD1L.n66 SUB 1.55fF
C456 SD1L.n67 SUB 1.55fF
C457 SD1L.n68 SUB 1.55fF
C458 SD1L.n69 SUB 1.55fF
C459 SD1L.n70 SUB 1.55fF
C460 SD1L.n71 SUB 1.44fF
C461 SD1L.n72 SUB 10.60fF
C462 SD1L.n73 SUB 10.60fF
C463 SD1L.n74 SUB 10.60fF
C464 SD1L.n75 SUB 10.60fF
C465 SD1L.n76 SUB 10.60fF
C466 SD1L.n77 SUB 10.60fF
C467 SD1L.n78 SUB 10.60fF
C468 SD1L.t98 SUB 9.16fF $ **FLOATING
C469 SD1L.n79 SUB 5.46fF
C470 SD1L.n80 SUB 1.55fF
C471 SD1L.n81 SUB 1.55fF
C472 SD1L.n82 SUB 1.55fF
C473 SD1L.n83 SUB 1.55fF
C474 SD1L.n84 SUB 1.55fF
C475 SD1L.n85 SUB 214.28fF
C476 SD1L.n86 SUB 153.28fF
C477 SD1L.n87 SUB 10.60fF
C478 SD1L.n88 SUB 10.60fF
C479 SD1L.n89 SUB 10.63fF
C480 SD1L.n90 SUB 10.60fF
C481 SD1L.n91 SUB 10.60fF
C482 SD1L.n92 SUB 10.60fF
C483 SD1L.n93 SUB 10.60fF
C484 SD1L.n94 SUB 10.60fF
C485 SD1L.n95 SUB 10.60fF
C486 SD1L.n96 SUB 10.64fF
C487 SD1L.n97 SUB 3.19fF
C488 SD1L.n98 SUB 1.55fF
C489 SD1L.n99 SUB 1.55fF
C490 SD1L.n100 SUB 1.55fF
C491 SD1L.n101 SUB 1.55fF
C492 SD1L.n102 SUB 1.55fF
C493 SD1L.n103 SUB 1.56fF
C494 SD1L.n104 SUB 1.55fF
C495 SD1L.n105 SUB 10.60fF
C496 SD1L.n106 SUB 10.60fF
C497 SD1L.n107 SUB 10.60fF
C498 SD1L.n108 SUB 10.64fF
C499 SD1L.n109 SUB 3.19fF
C500 SD1L.n110 SUB 10.60fF
C501 SD1L.n111 SUB 1.55fF
C502 SD1L.n112 SUB 1.55fF
C503 SD1L.n113 SUB 1.53fF
C504 SD1L.n114 SUB 116.77fF
.ends