magic
tech sky130A
timestamp 1659501813
<< metal3 >>
rect 5150 2850 6400 3000
rect 5150 2400 6150 2850
rect 6350 2550 6400 2850
rect 6350 2400 6450 2550
rect 6350 2250 6400 2400
rect 6150 2200 6400 2250
rect 5150 1250 6450 1850
<< via3 >>
rect 6150 2250 6350 2850
<< metal4 >>
rect 2500 4200 3600 4400
rect 4750 4250 5950 4300
rect 4750 3850 4800 4250
rect 5100 3850 5950 4250
rect 4750 3800 5150 3850
rect 6100 2850 6400 2900
rect 6100 2250 6150 2850
rect 6350 2250 6400 2850
rect 6100 2200 6400 2250
rect 4750 600 5900 650
rect 4750 200 4800 600
rect 5100 200 5900 600
rect 4750 150 5150 200
rect 2500 -100 3600 100
<< via4 >>
rect 4800 3850 5100 4250
rect 4800 200 5100 600
<< metal5 >>
rect 4750 4250 5150 4300
rect 4750 3850 4800 4250
rect 5100 3850 5150 4250
rect 4750 3800 5150 3850
rect 4750 600 5150 650
rect 4750 200 4800 600
rect 5100 200 5150 600
rect 4750 150 5150 200
use MIXER_5G_core  MIXER_5G_core_0
timestamp 1659323209
transform 1 0 580 0 1 2400
box -580 -2400 4940 1900
use OSC_5GHz_1  OSC_5GHz_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/OSC
timestamp 1659407314
transform 1 0 700 0 1 -1150
box 5000 -5450 28100 12050
use octal_ind_0p700n_5GHz  octal_ind_0p700n_5GHz_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1659405087
transform 0 -1 -8450 1 0 20200
box -16900 -16250 -4400 -3750
use octal_ind_0p700n_5GHz  octal_ind_0p700n_5GHz_1
timestamp 1659405087
transform 0 -1 -8450 -1 0 -15900
box -16900 -16250 -4400 -3750
<< end >>
