magic
tech sky130B
timestamp 1661649873
<< metal4 >>
rect 11000 5400 16000 5500
rect 10150 4700 10550 4750
rect 11000 4700 11100 5400
rect 10150 4100 11100 4700
rect 15900 4100 16000 5400
rect 11000 4000 16000 4100
rect 10150 2400 10550 2450
rect 11000 2400 16000 2500
rect 10150 1800 11100 2400
rect 11000 1100 11100 1800
rect 15900 1100 16000 2400
rect 11000 1000 16000 1100
<< via4 >>
rect 11100 4100 15900 5400
rect 11100 1100 15900 2400
<< metal5 >>
rect 13500 5500 16000 7500
rect 11000 5400 16000 5500
rect 11000 4100 11100 5400
rect 15900 4100 16000 5400
rect 11000 4000 16000 4100
rect 11000 2400 16000 2500
rect 11000 1100 11100 2400
rect 15900 1100 16000 2400
rect 11000 1000 16000 1100
rect 13500 -1000 16000 1000
use OSC_5GHz_wo_ind  OSC_5GHz_wo_ind_0
timestamp 1661123328
transform 1 0 7950 0 1 2500
box -2950 -1800 2600 3400
use octa_symm_thick_2t_275_200_flat  octa_symm_thick_2t_275_200_flat_0
timestamp 1661649517
transform 1 0 35161 0 1 13250
box -21661 -23750 -1150 3750
<< end >>
