magic
tech sky130B
magscale 1 2
timestamp 1660448881
<< error_p >>
rect -269 872 -211 878
rect -77 872 -19 878
rect 115 872 173 878
rect 307 872 365 878
rect -269 838 -257 872
rect -77 838 -65 872
rect 115 838 127 872
rect 307 838 319 872
rect -269 832 -211 838
rect -77 832 -19 838
rect 115 832 173 838
rect 307 832 365 838
rect -365 -838 -307 -832
rect -173 -838 -115 -832
rect 19 -838 77 -832
rect 211 -838 269 -832
rect -365 -872 -353 -838
rect -173 -872 -161 -838
rect 19 -872 31 -838
rect 211 -872 223 -838
rect -365 -878 -307 -872
rect -173 -878 -115 -872
rect 19 -878 77 -872
rect 211 -878 269 -872
<< pwell >>
rect -551 -1010 551 1010
<< nmos >>
rect -351 -800 -321 800
rect -255 -800 -225 800
rect -159 -800 -129 800
rect -63 -800 -33 800
rect 33 -800 63 800
rect 129 -800 159 800
rect 225 -800 255 800
rect 321 -800 351 800
<< ndiff >>
rect -413 788 -351 800
rect -413 -788 -401 788
rect -367 -788 -351 788
rect -413 -800 -351 -788
rect -321 788 -255 800
rect -321 -788 -305 788
rect -271 -788 -255 788
rect -321 -800 -255 -788
rect -225 788 -159 800
rect -225 -788 -209 788
rect -175 -788 -159 788
rect -225 -800 -159 -788
rect -129 788 -63 800
rect -129 -788 -113 788
rect -79 -788 -63 788
rect -129 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 129 800
rect 63 -788 79 788
rect 113 -788 129 788
rect 63 -800 129 -788
rect 159 788 225 800
rect 159 -788 175 788
rect 209 -788 225 788
rect 159 -800 225 -788
rect 255 788 321 800
rect 255 -788 271 788
rect 305 -788 321 788
rect 255 -800 321 -788
rect 351 788 413 800
rect 351 -788 367 788
rect 401 -788 413 788
rect 351 -800 413 -788
<< ndiffc >>
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
<< psubdiff >>
rect -515 940 -419 974
rect 419 940 515 974
rect -515 878 -481 940
rect 481 878 515 940
rect -515 -940 -481 -878
rect 481 -940 515 -878
rect -515 -974 -419 -940
rect 419 -974 515 -940
<< psubdiffcont >>
rect -419 940 419 974
rect -515 -878 -481 878
rect 481 -878 515 878
rect -419 -974 419 -940
<< poly >>
rect -273 872 -207 888
rect -273 838 -257 872
rect -223 838 -207 872
rect -351 800 -321 826
rect -273 822 -207 838
rect -81 872 -15 888
rect -81 838 -65 872
rect -31 838 -15 872
rect -255 800 -225 822
rect -159 800 -129 826
rect -81 822 -15 838
rect 111 872 177 888
rect 111 838 127 872
rect 161 838 177 872
rect -63 800 -33 822
rect 33 800 63 826
rect 111 822 177 838
rect 303 872 369 888
rect 303 838 319 872
rect 353 838 369 872
rect 129 800 159 822
rect 225 800 255 826
rect 303 822 369 838
rect 321 800 351 822
rect -351 -822 -321 -800
rect -369 -838 -303 -822
rect -255 -826 -225 -800
rect -159 -822 -129 -800
rect -369 -872 -353 -838
rect -319 -872 -303 -838
rect -369 -888 -303 -872
rect -177 -838 -111 -822
rect -63 -826 -33 -800
rect 33 -822 63 -800
rect -177 -872 -161 -838
rect -127 -872 -111 -838
rect -177 -888 -111 -872
rect 15 -838 81 -822
rect 129 -826 159 -800
rect 225 -822 255 -800
rect 15 -872 31 -838
rect 65 -872 81 -838
rect 15 -888 81 -872
rect 207 -838 273 -822
rect 321 -826 351 -800
rect 207 -872 223 -838
rect 257 -872 273 -838
rect 207 -888 273 -872
<< polycont >>
rect -257 838 -223 872
rect -65 838 -31 872
rect 127 838 161 872
rect 319 838 353 872
rect -353 -872 -319 -838
rect -161 -872 -127 -838
rect 31 -872 65 -838
rect 223 -872 257 -838
<< locali >>
rect -515 940 -419 974
rect 419 940 515 974
rect -515 878 -481 940
rect 481 878 515 940
rect -273 838 -257 872
rect -223 838 -207 872
rect -81 838 -65 872
rect -31 838 -15 872
rect 111 838 127 872
rect 161 838 177 872
rect 303 838 319 872
rect 353 838 369 872
rect -401 788 -367 804
rect -401 -804 -367 -788
rect -305 788 -271 804
rect -305 -804 -271 -788
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect 271 788 305 804
rect 271 -804 305 -788
rect 367 788 401 804
rect 367 -804 401 -788
rect -369 -872 -353 -838
rect -319 -872 -303 -838
rect -177 -872 -161 -838
rect -127 -872 -111 -838
rect 15 -872 31 -838
rect 65 -872 81 -838
rect 207 -872 223 -838
rect 257 -872 273 -838
rect -515 -940 -481 -878
rect 481 -940 515 -878
rect -515 -974 -419 -940
rect 419 -974 515 -940
<< viali >>
rect -257 838 -223 872
rect -65 838 -31 872
rect 127 838 161 872
rect 319 838 353 872
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect -353 -872 -319 -838
rect -161 -872 -127 -838
rect 31 -872 65 -838
rect 223 -872 257 -838
<< metal1 >>
rect -269 872 -211 878
rect -269 838 -257 872
rect -223 838 -211 872
rect -269 832 -211 838
rect -77 872 -19 878
rect -77 838 -65 872
rect -31 838 -19 872
rect -77 832 -19 838
rect 115 872 173 878
rect 115 838 127 872
rect 161 838 173 872
rect 115 832 173 838
rect 307 872 365 878
rect 307 838 319 872
rect 353 838 365 872
rect 307 832 365 838
rect -407 788 -361 800
rect -407 -788 -401 788
rect -367 -788 -361 788
rect -407 -800 -361 -788
rect -311 788 -265 800
rect -311 -788 -305 788
rect -271 -788 -265 788
rect -311 -800 -265 -788
rect -215 788 -169 800
rect -215 -788 -209 788
rect -175 -788 -169 788
rect -215 -800 -169 -788
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
rect 169 788 215 800
rect 169 -788 175 788
rect 209 -788 215 788
rect 169 -800 215 -788
rect 265 788 311 800
rect 265 -788 271 788
rect 305 -788 311 788
rect 265 -800 311 -788
rect 361 788 407 800
rect 361 -788 367 788
rect 401 -788 407 788
rect 361 -800 407 -788
rect -365 -838 -307 -832
rect -365 -872 -353 -838
rect -319 -872 -307 -838
rect -365 -878 -307 -872
rect -173 -838 -115 -832
rect -173 -872 -161 -838
rect -127 -872 -115 -838
rect -173 -878 -115 -872
rect 19 -838 77 -832
rect 19 -872 31 -838
rect 65 -872 77 -838
rect 19 -878 77 -872
rect 211 -838 269 -832
rect 211 -872 223 -838
rect 257 -872 269 -838
rect 211 -878 269 -872
<< properties >>
string FIXED_BBOX -498 -957 498 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
