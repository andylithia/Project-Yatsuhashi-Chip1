magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< nwell >>
rect -54 -54 204 1454
<< scpmos >>
rect 60 0 90 1400
<< pdiff >>
rect 0 0 60 1400
rect 90 0 150 1400
<< poly >>
rect 60 1400 90 1426
rect 60 -26 90 0
<< locali >>
rect 8 667 42 733
rect 108 667 142 733
use sky130_sram_1r1w_24x128_8_contact_11  sky130_sram_1r1w_24x128_8_contact_11_0
timestamp 1661296025
transform 1 0 100 0 1 667
box -59 -51 109 117
use sky130_sram_1r1w_24x128_8_contact_11  sky130_sram_1r1w_24x128_8_contact_11_1
timestamp 1661296025
transform 1 0 0 0 1 667
box -59 -51 109 117
<< labels >>
rlabel poly s 75 700 75 700 4 G
port 1 nsew
rlabel locali s 25 700 25 700 4 S
port 2 nsew
rlabel locali s 125 700 125 700 4 D
port 3 nsew
<< properties >>
string FIXED_BBOX -54 -54 204 1454
<< end >>
