magic
tech sky130B
magscale 1 2
timestamp 1662654558
<< metal1 >>
rect -83500 82880 100500 82900
rect -83500 82810 -83350 82880
rect -83150 82810 -82850 82880
rect -82650 82810 -82350 82880
rect -82150 82810 -81850 82880
rect -81650 82810 -81350 82880
rect -81150 82810 -80850 82880
rect -80650 82810 -80350 82880
rect -80150 82810 -79850 82880
rect -79650 82810 -79350 82880
rect -79150 82810 -78850 82880
rect -78650 82810 -78350 82880
rect -78150 82810 -77850 82880
rect -77650 82810 -77350 82880
rect -77150 82810 -76850 82880
rect -76650 82810 -76350 82880
rect -76150 82810 -75850 82880
rect -75650 82810 -75350 82880
rect -75150 82810 -74850 82880
rect -74650 82810 -74350 82880
rect -74150 82810 -73850 82880
rect -73650 82810 -73350 82880
rect -73150 82810 -72850 82880
rect -72650 82810 -72350 82880
rect -72150 82810 -71850 82880
rect -71650 82810 -71350 82880
rect -71150 82810 -70850 82880
rect -70650 82810 -70350 82880
rect -70150 82810 -69850 82880
rect -69650 82810 -69350 82880
rect -69150 82810 -68850 82880
rect -68650 82810 -68350 82880
rect -68150 82810 -67850 82880
rect -67650 82810 -67350 82880
rect -67150 82810 -66850 82880
rect -66650 82810 -66350 82880
rect -66150 82810 -65850 82880
rect -65650 82810 -65350 82880
rect -65150 82810 -64850 82880
rect -64650 82810 -64350 82880
rect -64150 82810 -63850 82880
rect -63650 82810 -63350 82880
rect -63150 82810 -62850 82880
rect -62650 82810 -62350 82880
rect -62150 82810 -61850 82880
rect -61650 82810 -61350 82880
rect -61150 82810 -60850 82880
rect -60650 82810 -60350 82880
rect -60150 82810 -59850 82880
rect -59650 82810 -59350 82880
rect -59150 82810 -58850 82880
rect -58650 82810 -58350 82880
rect -58150 82810 -57850 82880
rect -57650 82810 -57350 82880
rect -57150 82810 -56850 82880
rect -56650 82810 -56350 82880
rect -56150 82810 -55850 82880
rect -55650 82810 -55350 82880
rect -55150 82810 -54850 82880
rect -54650 82810 -54350 82880
rect -54150 82810 -53850 82880
rect -53650 82810 -53350 82880
rect -53150 82810 -52850 82880
rect -52650 82810 -52350 82880
rect -52150 82810 -51850 82880
rect -51650 82810 -51350 82880
rect -51150 82810 -50850 82880
rect -50650 82810 -50350 82880
rect -50150 82810 -49850 82880
rect -49650 82810 -49350 82880
rect -49150 82810 -48850 82880
rect -48650 82810 -48350 82880
rect -48150 82810 -47850 82880
rect -47650 82810 -47350 82880
rect -47150 82810 -46850 82880
rect -46650 82810 -46350 82880
rect -46150 82810 -45850 82880
rect -45650 82810 -45350 82880
rect -45150 82810 -44850 82880
rect -44650 82810 -44350 82880
rect -44150 82810 -43850 82880
rect -43650 82810 -43350 82880
rect -43150 82810 -42850 82880
rect -42650 82810 -42350 82880
rect -42150 82810 -41850 82880
rect -41650 82810 -41350 82880
rect -41150 82810 -40850 82880
rect -40650 82810 -40350 82880
rect -40150 82810 -39850 82880
rect -39650 82810 -39350 82880
rect -39150 82810 -38850 82880
rect -38650 82810 -38350 82880
rect -38150 82810 -37850 82880
rect -37650 82810 -37350 82880
rect -37150 82810 -36850 82880
rect -36650 82810 -36350 82880
rect -36150 82810 -35850 82880
rect -35650 82810 -35350 82880
rect -35150 82810 -34850 82880
rect -34650 82810 -34350 82880
rect -34150 82810 -33850 82880
rect -33650 82810 -33350 82880
rect -33150 82810 -32850 82880
rect -32650 82810 -32350 82880
rect -32150 82810 -31850 82880
rect -31650 82810 -31350 82880
rect -31150 82810 -30850 82880
rect -30650 82810 -30350 82880
rect -30150 82810 -29850 82880
rect -29650 82810 -29350 82880
rect -29150 82810 -28850 82880
rect -28650 82810 -28350 82880
rect -28150 82810 -27850 82880
rect -27650 82810 -27350 82880
rect -27150 82810 -26850 82880
rect -26650 82810 -26350 82880
rect -26150 82810 -25850 82880
rect -25650 82810 -25350 82880
rect -25150 82810 -24850 82880
rect -24650 82810 -24350 82880
rect -24150 82810 -23850 82880
rect -23650 82810 -23350 82880
rect -23150 82810 -22850 82880
rect -22650 82810 -22350 82880
rect -22150 82810 -21850 82880
rect -21650 82810 -21350 82880
rect -21150 82810 -20850 82880
rect -20650 82810 -20350 82880
rect -20150 82810 -19850 82880
rect -19650 82810 -19350 82880
rect -19150 82810 -18850 82880
rect -18650 82810 -18350 82880
rect -18150 82810 -17850 82880
rect -17650 82810 -17350 82880
rect -17150 82810 -16850 82880
rect -16650 82810 -16350 82880
rect -16150 82810 -15850 82880
rect -15650 82810 -15350 82880
rect -15150 82810 -14850 82880
rect -14650 82810 -14350 82880
rect -14150 82810 -13850 82880
rect -13650 82810 -13350 82880
rect -13150 82810 -12850 82880
rect -12650 82810 -12350 82880
rect -12150 82810 -11850 82880
rect -11650 82810 -11350 82880
rect -11150 82810 -10850 82880
rect -10650 82810 -10350 82880
rect -10150 82810 -9850 82880
rect -9650 82810 -9350 82880
rect -9150 82810 -8850 82880
rect -8650 82810 -8350 82880
rect -8150 82810 -7850 82880
rect -7650 82810 -7350 82880
rect -7150 82810 -6850 82880
rect -6650 82810 -6350 82880
rect -6150 82810 -5850 82880
rect -5650 82810 -5350 82880
rect -5150 82810 -4850 82880
rect -4650 82810 -4350 82880
rect -4150 82810 -3850 82880
rect -3650 82810 -3350 82880
rect -3150 82810 -2850 82880
rect -2650 82810 -2350 82880
rect -2150 82810 -1850 82880
rect -1650 82810 -1350 82880
rect -1150 82810 -850 82880
rect -650 82810 -350 82880
rect -150 82810 150 82880
rect 350 82810 650 82880
rect 850 82810 1150 82880
rect 1350 82810 1650 82880
rect 1850 82810 2150 82880
rect 2350 82810 2650 82880
rect 2850 82810 3150 82880
rect 3350 82810 3650 82880
rect 3850 82810 4150 82880
rect 4350 82810 4650 82880
rect 4850 82810 5150 82880
rect 5350 82810 5650 82880
rect 5850 82810 6150 82880
rect 6350 82810 6650 82880
rect 6850 82810 7150 82880
rect 7350 82810 7650 82880
rect 7850 82810 8150 82880
rect 8350 82810 8650 82880
rect 8850 82810 9150 82880
rect 9350 82810 9650 82880
rect 9850 82810 10150 82880
rect 10350 82810 10650 82880
rect 10850 82810 11150 82880
rect 11350 82810 11650 82880
rect 11850 82810 12150 82880
rect 12350 82810 12650 82880
rect 12850 82810 13150 82880
rect 13350 82810 13650 82880
rect 13850 82810 14150 82880
rect 14350 82810 14650 82880
rect 14850 82810 15150 82880
rect 15350 82810 15650 82880
rect 15850 82810 16150 82880
rect 16350 82810 16650 82880
rect 16850 82810 17150 82880
rect 17350 82810 17650 82880
rect 17850 82810 18150 82880
rect 18350 82810 18650 82880
rect 18850 82810 19150 82880
rect 19350 82810 19650 82880
rect 19850 82810 20150 82880
rect 20350 82810 20650 82880
rect 20850 82810 21150 82880
rect 21350 82810 21650 82880
rect 21850 82810 22150 82880
rect 22350 82810 22650 82880
rect 22850 82810 23150 82880
rect 23350 82810 23650 82880
rect 23850 82810 24150 82880
rect 24350 82810 24650 82880
rect 24850 82810 25150 82880
rect 25350 82810 25650 82880
rect 25850 82810 26150 82880
rect 26350 82810 26650 82880
rect 26850 82810 27150 82880
rect 27350 82810 27650 82880
rect 27850 82810 28150 82880
rect 28350 82810 28650 82880
rect 28850 82810 29150 82880
rect 29350 82810 29650 82880
rect 29850 82810 30150 82880
rect 30350 82810 30650 82880
rect 30850 82810 31150 82880
rect 31350 82810 31650 82880
rect 31850 82810 32150 82880
rect 32350 82810 32650 82880
rect 32850 82810 33150 82880
rect 33350 82810 33650 82880
rect 33850 82810 34150 82880
rect 34350 82810 34650 82880
rect 34850 82810 35150 82880
rect 35350 82810 35650 82880
rect 35850 82810 36150 82880
rect 36350 82810 36650 82880
rect 36850 82810 37150 82880
rect 37350 82810 37650 82880
rect 37850 82810 38150 82880
rect 38350 82810 38650 82880
rect 38850 82810 39150 82880
rect 39350 82810 39650 82880
rect 39850 82810 40150 82880
rect 40350 82810 40650 82880
rect 40850 82810 41150 82880
rect 41350 82810 41650 82880
rect 41850 82810 42150 82880
rect 42350 82810 42650 82880
rect 42850 82810 43150 82880
rect 43350 82810 43650 82880
rect 43850 82810 44150 82880
rect 44350 82810 44650 82880
rect 44850 82810 45150 82880
rect 45350 82810 45650 82880
rect 45850 82810 46150 82880
rect 46350 82810 46650 82880
rect 46850 82810 47150 82880
rect 47350 82810 47650 82880
rect 47850 82810 48150 82880
rect 48350 82810 48650 82880
rect 48850 82810 49150 82880
rect 49350 82810 49650 82880
rect 49850 82810 50150 82880
rect 50350 82810 50650 82880
rect 50850 82810 51150 82880
rect 51350 82810 51650 82880
rect 51850 82810 52150 82880
rect 52350 82810 52650 82880
rect 52850 82810 53150 82880
rect 53350 82810 53650 82880
rect 53850 82810 54150 82880
rect 54350 82810 54650 82880
rect 54850 82810 55150 82880
rect 55350 82810 55650 82880
rect 55850 82810 56150 82880
rect 56350 82810 56650 82880
rect 56850 82810 57150 82880
rect 57350 82810 57650 82880
rect 57850 82810 58150 82880
rect 58350 82810 58650 82880
rect 58850 82810 59150 82880
rect 59350 82810 59650 82880
rect 59850 82810 60150 82880
rect 60350 82810 60650 82880
rect 60850 82810 61150 82880
rect 61350 82810 61650 82880
rect 61850 82810 62150 82880
rect 62350 82810 62650 82880
rect 62850 82810 63150 82880
rect 63350 82810 63650 82880
rect 63850 82810 64150 82880
rect 64350 82810 64650 82880
rect 64850 82810 65150 82880
rect 65350 82810 65650 82880
rect 65850 82810 66150 82880
rect 66350 82810 66650 82880
rect 66850 82810 67150 82880
rect 67350 82810 67650 82880
rect 67850 82810 68150 82880
rect 68350 82810 68650 82880
rect 68850 82810 69150 82880
rect 69350 82810 69650 82880
rect 69850 82810 70150 82880
rect 70350 82810 70650 82880
rect 70850 82810 71150 82880
rect 71350 82810 71650 82880
rect 71850 82810 72150 82880
rect 72350 82810 72650 82880
rect 72850 82810 73150 82880
rect 73350 82810 73650 82880
rect 73850 82810 74150 82880
rect 74350 82810 74650 82880
rect 74850 82810 75150 82880
rect 75350 82810 75650 82880
rect 75850 82810 76150 82880
rect 76350 82810 76650 82880
rect 76850 82810 77150 82880
rect 77350 82810 77650 82880
rect 77850 82810 78150 82880
rect 78350 82810 78650 82880
rect 78850 82810 79150 82880
rect 79350 82810 79650 82880
rect 79850 82810 80150 82880
rect 80350 82810 80650 82880
rect 80850 82810 81150 82880
rect 81350 82810 81650 82880
rect 81850 82810 82150 82880
rect 82350 82810 82650 82880
rect 82850 82810 83150 82880
rect 83350 82810 83650 82880
rect 83850 82810 84150 82880
rect 84350 82810 84650 82880
rect 84850 82810 85150 82880
rect 85350 82810 85650 82880
rect 85850 82810 86150 82880
rect 86350 82810 86650 82880
rect 86850 82810 87150 82880
rect 87350 82810 87650 82880
rect 87850 82810 88150 82880
rect 88350 82810 88650 82880
rect 88850 82810 89150 82880
rect 89350 82810 89650 82880
rect 89850 82810 90150 82880
rect 90350 82810 90650 82880
rect 90850 82810 91150 82880
rect 91350 82810 91650 82880
rect 91850 82810 92150 82880
rect 92350 82810 92650 82880
rect 92850 82810 93150 82880
rect 93350 82810 93650 82880
rect 93850 82810 94150 82880
rect 94350 82810 94650 82880
rect 94850 82810 95150 82880
rect 95350 82810 95650 82880
rect 95850 82810 96150 82880
rect 96350 82810 96650 82880
rect 96850 82810 97150 82880
rect 97350 82810 97650 82880
rect 97850 82810 98150 82880
rect 98350 82810 98650 82880
rect 98850 82810 99150 82880
rect 99350 82810 99650 82880
rect 99850 82810 100150 82880
rect 100350 82810 100500 82880
rect -83500 82800 100500 82810
rect -83500 82780 -83380 82800
rect -83120 82780 -82880 82800
rect -82620 82780 -82380 82800
rect -82120 82780 -81880 82800
rect -81620 82780 -81380 82800
rect -81120 82780 -80880 82800
rect -80620 82780 -80380 82800
rect -80120 82780 -79880 82800
rect -79620 82780 -79380 82800
rect -79120 82780 -78880 82800
rect -78620 82780 -78380 82800
rect -78120 82780 -77880 82800
rect -77620 82780 -77380 82800
rect -77120 82780 -76880 82800
rect -76620 82780 -76380 82800
rect -76120 82780 -75880 82800
rect -75620 82780 -75380 82800
rect -75120 82780 -74880 82800
rect -74620 82780 -74380 82800
rect -74120 82780 -73880 82800
rect -73620 82780 -73380 82800
rect -73120 82780 -72880 82800
rect -72620 82780 -72380 82800
rect -72120 82780 -71880 82800
rect -71620 82780 -71380 82800
rect -71120 82780 -70880 82800
rect -70620 82780 -70380 82800
rect -70120 82780 -69880 82800
rect -69620 82780 -69380 82800
rect -69120 82780 -68880 82800
rect -68620 82780 -68380 82800
rect -68120 82780 -67880 82800
rect -67620 82780 -67380 82800
rect -67120 82780 -66880 82800
rect -66620 82780 -66380 82800
rect -66120 82780 -65880 82800
rect -65620 82780 -65380 82800
rect -65120 82780 -64880 82800
rect -64620 82780 -64380 82800
rect -64120 82780 -63880 82800
rect -63620 82780 -63380 82800
rect -63120 82780 -62880 82800
rect -62620 82780 -62380 82800
rect -62120 82780 -61880 82800
rect -61620 82780 -61380 82800
rect -61120 82780 -60880 82800
rect -60620 82780 -60380 82800
rect -60120 82780 -59880 82800
rect -59620 82780 -59380 82800
rect -59120 82780 -58880 82800
rect -58620 82780 -58380 82800
rect -58120 82780 -57880 82800
rect -57620 82780 -57380 82800
rect -57120 82780 -56880 82800
rect -56620 82780 -56380 82800
rect -56120 82780 -55880 82800
rect -55620 82780 -55380 82800
rect -55120 82780 -54880 82800
rect -54620 82780 -54380 82800
rect -54120 82780 -53880 82800
rect -53620 82780 -53380 82800
rect -53120 82780 -52880 82800
rect -52620 82780 -52380 82800
rect -52120 82780 -51880 82800
rect -51620 82780 -51380 82800
rect -51120 82780 -50880 82800
rect -50620 82780 -50380 82800
rect -50120 82780 -49880 82800
rect -49620 82780 -49380 82800
rect -49120 82780 -48880 82800
rect -48620 82780 -48380 82800
rect -48120 82780 -47880 82800
rect -47620 82780 -47380 82800
rect -47120 82780 -46880 82800
rect -46620 82780 -46380 82800
rect -46120 82780 -45880 82800
rect -45620 82780 -45380 82800
rect -45120 82780 -44880 82800
rect -44620 82780 -44380 82800
rect -44120 82780 -43880 82800
rect -43620 82780 -43380 82800
rect -43120 82780 -42880 82800
rect -42620 82780 -42380 82800
rect -42120 82780 -41880 82800
rect -41620 82780 -41380 82800
rect -41120 82780 -40880 82800
rect -40620 82780 -40380 82800
rect -40120 82780 -39880 82800
rect -39620 82780 -39380 82800
rect -39120 82780 -38880 82800
rect -38620 82780 -38380 82800
rect -38120 82780 -37880 82800
rect -37620 82780 -37380 82800
rect -37120 82780 -36880 82800
rect -36620 82780 -36380 82800
rect -36120 82780 -35880 82800
rect -35620 82780 -35380 82800
rect -35120 82780 -34880 82800
rect -34620 82780 -34380 82800
rect -34120 82780 -33880 82800
rect -33620 82780 -33380 82800
rect -33120 82780 -32880 82800
rect -32620 82780 -32380 82800
rect -32120 82780 -31880 82800
rect -31620 82780 -31380 82800
rect -31120 82780 -30880 82800
rect -30620 82780 -30380 82800
rect -30120 82780 -29880 82800
rect -29620 82780 -29380 82800
rect -29120 82780 -28880 82800
rect -28620 82780 -28380 82800
rect -28120 82780 -27880 82800
rect -27620 82780 -27380 82800
rect -27120 82780 -26880 82800
rect -26620 82780 -26380 82800
rect -26120 82780 -25880 82800
rect -25620 82780 -25380 82800
rect -25120 82780 -24880 82800
rect -24620 82780 -24380 82800
rect -24120 82780 -23880 82800
rect -23620 82780 -23380 82800
rect -23120 82780 -22880 82800
rect -22620 82780 -22380 82800
rect -22120 82780 -21880 82800
rect -21620 82780 -21380 82800
rect -21120 82780 -20880 82800
rect -20620 82780 -20380 82800
rect -20120 82780 -19880 82800
rect -19620 82780 -19380 82800
rect -19120 82780 -18880 82800
rect -18620 82780 -18380 82800
rect -18120 82780 -17880 82800
rect -17620 82780 -17380 82800
rect -17120 82780 -16880 82800
rect -16620 82780 -16380 82800
rect -16120 82780 -15880 82800
rect -15620 82780 -15380 82800
rect -15120 82780 -14880 82800
rect -14620 82780 -14380 82800
rect -14120 82780 -13880 82800
rect -13620 82780 -13380 82800
rect -13120 82780 -12880 82800
rect -12620 82780 -12380 82800
rect -12120 82780 -11880 82800
rect -11620 82780 -11380 82800
rect -11120 82780 -10880 82800
rect -10620 82780 -10380 82800
rect -10120 82780 -9880 82800
rect -9620 82780 -9380 82800
rect -9120 82780 -8880 82800
rect -8620 82780 -8380 82800
rect -8120 82780 -7880 82800
rect -7620 82780 -7380 82800
rect -7120 82780 -6880 82800
rect -6620 82780 -6380 82800
rect -6120 82780 -5880 82800
rect -5620 82780 -5380 82800
rect -5120 82780 -4880 82800
rect -4620 82780 -4380 82800
rect -4120 82780 -3880 82800
rect -3620 82780 -3380 82800
rect -3120 82780 -2880 82800
rect -2620 82780 -2380 82800
rect -2120 82780 -1880 82800
rect -1620 82780 -1380 82800
rect -1120 82780 -880 82800
rect -620 82780 -380 82800
rect -120 82780 120 82800
rect 380 82780 620 82800
rect 880 82780 1120 82800
rect 1380 82780 1620 82800
rect 1880 82780 2120 82800
rect 2380 82780 2620 82800
rect 2880 82780 3120 82800
rect 3380 82780 3620 82800
rect 3880 82780 4120 82800
rect 4380 82780 4620 82800
rect 4880 82780 5120 82800
rect 5380 82780 5620 82800
rect 5880 82780 6120 82800
rect 6380 82780 6620 82800
rect 6880 82780 7120 82800
rect 7380 82780 7620 82800
rect 7880 82780 8120 82800
rect 8380 82780 8620 82800
rect 8880 82780 9120 82800
rect 9380 82780 9620 82800
rect 9880 82780 10120 82800
rect 10380 82780 10620 82800
rect 10880 82780 11120 82800
rect 11380 82780 11620 82800
rect 11880 82780 12120 82800
rect 12380 82780 12620 82800
rect 12880 82780 13120 82800
rect 13380 82780 13620 82800
rect 13880 82780 14120 82800
rect 14380 82780 14620 82800
rect 14880 82780 15120 82800
rect 15380 82780 15620 82800
rect 15880 82780 16120 82800
rect 16380 82780 16620 82800
rect 16880 82780 17120 82800
rect 17380 82780 17620 82800
rect 17880 82780 18120 82800
rect 18380 82780 18620 82800
rect 18880 82780 19120 82800
rect 19380 82780 19620 82800
rect 19880 82780 20120 82800
rect 20380 82780 20620 82800
rect 20880 82780 21120 82800
rect 21380 82780 21620 82800
rect 21880 82780 22120 82800
rect 22380 82780 22620 82800
rect 22880 82780 23120 82800
rect 23380 82780 23620 82800
rect 23880 82780 24120 82800
rect 24380 82780 24620 82800
rect 24880 82780 25120 82800
rect 25380 82780 25620 82800
rect 25880 82780 26120 82800
rect 26380 82780 26620 82800
rect 26880 82780 27120 82800
rect 27380 82780 27620 82800
rect 27880 82780 28120 82800
rect 28380 82780 28620 82800
rect 28880 82780 29120 82800
rect 29380 82780 29620 82800
rect 29880 82780 30120 82800
rect 30380 82780 30620 82800
rect 30880 82780 31120 82800
rect 31380 82780 31620 82800
rect 31880 82780 32120 82800
rect 32380 82780 32620 82800
rect 32880 82780 33120 82800
rect 33380 82780 33620 82800
rect 33880 82780 34120 82800
rect 34380 82780 34620 82800
rect 34880 82780 35120 82800
rect 35380 82780 35620 82800
rect 35880 82780 36120 82800
rect 36380 82780 36620 82800
rect 36880 82780 37120 82800
rect 37380 82780 37620 82800
rect 37880 82780 38120 82800
rect 38380 82780 38620 82800
rect 38880 82780 39120 82800
rect 39380 82780 39620 82800
rect 39880 82780 40120 82800
rect 40380 82780 40620 82800
rect 40880 82780 41120 82800
rect 41380 82780 41620 82800
rect 41880 82780 42120 82800
rect 42380 82780 42620 82800
rect 42880 82780 43120 82800
rect 43380 82780 43620 82800
rect 43880 82780 44120 82800
rect 44380 82780 44620 82800
rect 44880 82780 45120 82800
rect 45380 82780 45620 82800
rect 45880 82780 46120 82800
rect 46380 82780 46620 82800
rect 46880 82780 47120 82800
rect 47380 82780 47620 82800
rect 47880 82780 48120 82800
rect 48380 82780 48620 82800
rect 48880 82780 49120 82800
rect 49380 82780 49620 82800
rect 49880 82780 50120 82800
rect 50380 82780 50620 82800
rect 50880 82780 51120 82800
rect 51380 82780 51620 82800
rect 51880 82780 52120 82800
rect 52380 82780 52620 82800
rect 52880 82780 53120 82800
rect 53380 82780 53620 82800
rect 53880 82780 54120 82800
rect 54380 82780 54620 82800
rect 54880 82780 55120 82800
rect 55380 82780 55620 82800
rect 55880 82780 56120 82800
rect 56380 82780 56620 82800
rect 56880 82780 57120 82800
rect 57380 82780 57620 82800
rect 57880 82780 58120 82800
rect 58380 82780 58620 82800
rect 58880 82780 59120 82800
rect 59380 82780 59620 82800
rect 59880 82780 60120 82800
rect 60380 82780 60620 82800
rect 60880 82780 61120 82800
rect 61380 82780 61620 82800
rect 61880 82780 62120 82800
rect 62380 82780 62620 82800
rect 62880 82780 63120 82800
rect 63380 82780 63620 82800
rect 63880 82780 64120 82800
rect 64380 82780 64620 82800
rect 64880 82780 65120 82800
rect 65380 82780 65620 82800
rect 65880 82780 66120 82800
rect 66380 82780 66620 82800
rect 66880 82780 67120 82800
rect 67380 82780 67620 82800
rect 67880 82780 68120 82800
rect 68380 82780 68620 82800
rect 68880 82780 69120 82800
rect 69380 82780 69620 82800
rect 69880 82780 70120 82800
rect 70380 82780 70620 82800
rect 70880 82780 71120 82800
rect 71380 82780 71620 82800
rect 71880 82780 72120 82800
rect 72380 82780 72620 82800
rect 72880 82780 73120 82800
rect 73380 82780 73620 82800
rect 73880 82780 74120 82800
rect 74380 82780 74620 82800
rect 74880 82780 75120 82800
rect 75380 82780 75620 82800
rect 75880 82780 76120 82800
rect 76380 82780 76620 82800
rect 76880 82780 77120 82800
rect 77380 82780 77620 82800
rect 77880 82780 78120 82800
rect 78380 82780 78620 82800
rect 78880 82780 79120 82800
rect 79380 82780 79620 82800
rect 79880 82780 80120 82800
rect 80380 82780 80620 82800
rect 80880 82780 81120 82800
rect 81380 82780 81620 82800
rect 81880 82780 82120 82800
rect 82380 82780 82620 82800
rect 82880 82780 83120 82800
rect 83380 82780 83620 82800
rect 83880 82780 84120 82800
rect 84380 82780 84620 82800
rect 84880 82780 85120 82800
rect 85380 82780 85620 82800
rect 85880 82780 86120 82800
rect 86380 82780 86620 82800
rect 86880 82780 87120 82800
rect 87380 82780 87620 82800
rect 87880 82780 88120 82800
rect 88380 82780 88620 82800
rect 88880 82780 89120 82800
rect 89380 82780 89620 82800
rect 89880 82780 90120 82800
rect 90380 82780 90620 82800
rect 90880 82780 91120 82800
rect 91380 82780 91620 82800
rect 91880 82780 92120 82800
rect 92380 82780 92620 82800
rect 92880 82780 93120 82800
rect 93380 82780 93620 82800
rect 93880 82780 94120 82800
rect 94380 82780 94620 82800
rect 94880 82780 95120 82800
rect 95380 82780 95620 82800
rect 95880 82780 96120 82800
rect 96380 82780 96620 82800
rect 96880 82780 97120 82800
rect 97380 82780 97620 82800
rect 97880 82780 98120 82800
rect 98380 82780 98620 82800
rect 98880 82780 99120 82800
rect 99380 82780 99620 82800
rect 99880 82780 100120 82800
rect 100380 82780 100500 82800
rect -83500 82750 -83400 82780
rect -83500 82550 -83480 82750
rect -83410 82550 -83400 82750
rect -83500 82520 -83400 82550
rect -83100 82750 -82900 82780
rect -83100 82550 -83090 82750
rect -83020 82550 -82980 82750
rect -82910 82550 -82900 82750
rect -83100 82520 -82900 82550
rect -82600 82750 -82400 82780
rect -82600 82550 -82590 82750
rect -82520 82550 -82480 82750
rect -82410 82550 -82400 82750
rect -82600 82520 -82400 82550
rect -82100 82750 -81900 82780
rect -82100 82550 -82090 82750
rect -82020 82550 -81980 82750
rect -81910 82550 -81900 82750
rect -82100 82520 -81900 82550
rect -81600 82750 -81400 82780
rect -81600 82550 -81590 82750
rect -81520 82550 -81480 82750
rect -81410 82550 -81400 82750
rect -81600 82520 -81400 82550
rect -81100 82750 -80900 82780
rect -81100 82550 -81090 82750
rect -81020 82550 -80980 82750
rect -80910 82550 -80900 82750
rect -81100 82520 -80900 82550
rect -80600 82750 -80400 82780
rect -80600 82550 -80590 82750
rect -80520 82550 -80480 82750
rect -80410 82550 -80400 82750
rect -80600 82520 -80400 82550
rect -80100 82750 -79900 82780
rect -80100 82550 -80090 82750
rect -80020 82550 -79980 82750
rect -79910 82550 -79900 82750
rect -80100 82520 -79900 82550
rect -79600 82750 -79400 82780
rect -79600 82550 -79590 82750
rect -79520 82550 -79480 82750
rect -79410 82550 -79400 82750
rect -79600 82520 -79400 82550
rect -79100 82750 -78900 82780
rect -79100 82550 -79090 82750
rect -79020 82550 -78980 82750
rect -78910 82550 -78900 82750
rect -79100 82520 -78900 82550
rect -78600 82750 -78400 82780
rect -78600 82550 -78590 82750
rect -78520 82550 -78480 82750
rect -78410 82550 -78400 82750
rect -78600 82520 -78400 82550
rect -78100 82750 -77900 82780
rect -78100 82550 -78090 82750
rect -78020 82550 -77980 82750
rect -77910 82550 -77900 82750
rect -78100 82520 -77900 82550
rect -77600 82750 -77400 82780
rect -77600 82550 -77590 82750
rect -77520 82550 -77480 82750
rect -77410 82550 -77400 82750
rect -77600 82520 -77400 82550
rect -77100 82750 -76900 82780
rect -77100 82550 -77090 82750
rect -77020 82550 -76980 82750
rect -76910 82550 -76900 82750
rect -77100 82520 -76900 82550
rect -76600 82750 -76400 82780
rect -76600 82550 -76590 82750
rect -76520 82550 -76480 82750
rect -76410 82550 -76400 82750
rect -76600 82520 -76400 82550
rect -76100 82750 -75900 82780
rect -76100 82550 -76090 82750
rect -76020 82550 -75980 82750
rect -75910 82550 -75900 82750
rect -76100 82520 -75900 82550
rect -75600 82750 -75400 82780
rect -75600 82550 -75590 82750
rect -75520 82550 -75480 82750
rect -75410 82550 -75400 82750
rect -75600 82520 -75400 82550
rect -75100 82750 -74900 82780
rect -75100 82550 -75090 82750
rect -75020 82550 -74980 82750
rect -74910 82550 -74900 82750
rect -75100 82520 -74900 82550
rect -74600 82750 -74400 82780
rect -74600 82550 -74590 82750
rect -74520 82550 -74480 82750
rect -74410 82550 -74400 82750
rect -74600 82520 -74400 82550
rect -74100 82750 -73900 82780
rect -74100 82550 -74090 82750
rect -74020 82550 -73980 82750
rect -73910 82550 -73900 82750
rect -74100 82520 -73900 82550
rect -73600 82750 -73400 82780
rect -73600 82550 -73590 82750
rect -73520 82550 -73480 82750
rect -73410 82550 -73400 82750
rect -73600 82520 -73400 82550
rect -73100 82750 -72900 82780
rect -73100 82550 -73090 82750
rect -73020 82550 -72980 82750
rect -72910 82550 -72900 82750
rect -73100 82520 -72900 82550
rect -72600 82750 -72400 82780
rect -72600 82550 -72590 82750
rect -72520 82550 -72480 82750
rect -72410 82550 -72400 82750
rect -72600 82520 -72400 82550
rect -72100 82750 -71900 82780
rect -72100 82550 -72090 82750
rect -72020 82550 -71980 82750
rect -71910 82550 -71900 82750
rect -72100 82520 -71900 82550
rect -71600 82750 -71400 82780
rect -71600 82550 -71590 82750
rect -71520 82550 -71480 82750
rect -71410 82550 -71400 82750
rect -71600 82520 -71400 82550
rect -71100 82750 -70900 82780
rect -71100 82550 -71090 82750
rect -71020 82550 -70980 82750
rect -70910 82550 -70900 82750
rect -71100 82520 -70900 82550
rect -70600 82750 -70400 82780
rect -70600 82550 -70590 82750
rect -70520 82550 -70480 82750
rect -70410 82550 -70400 82750
rect -70600 82520 -70400 82550
rect -70100 82750 -69900 82780
rect -70100 82550 -70090 82750
rect -70020 82550 -69980 82750
rect -69910 82550 -69900 82750
rect -70100 82520 -69900 82550
rect -69600 82750 -69400 82780
rect -69600 82550 -69590 82750
rect -69520 82550 -69480 82750
rect -69410 82550 -69400 82750
rect -69600 82520 -69400 82550
rect -69100 82750 -68900 82780
rect -69100 82550 -69090 82750
rect -69020 82550 -68980 82750
rect -68910 82550 -68900 82750
rect -69100 82520 -68900 82550
rect -68600 82750 -68400 82780
rect -68600 82550 -68590 82750
rect -68520 82550 -68480 82750
rect -68410 82550 -68400 82750
rect -68600 82520 -68400 82550
rect -68100 82750 -67900 82780
rect -68100 82550 -68090 82750
rect -68020 82550 -67980 82750
rect -67910 82550 -67900 82750
rect -68100 82520 -67900 82550
rect -67600 82750 -67400 82780
rect -67600 82550 -67590 82750
rect -67520 82550 -67480 82750
rect -67410 82550 -67400 82750
rect -67600 82520 -67400 82550
rect -67100 82750 -66900 82780
rect -67100 82550 -67090 82750
rect -67020 82550 -66980 82750
rect -66910 82550 -66900 82750
rect -67100 82520 -66900 82550
rect -66600 82750 -66400 82780
rect -66600 82550 -66590 82750
rect -66520 82550 -66480 82750
rect -66410 82550 -66400 82750
rect -66600 82520 -66400 82550
rect -66100 82750 -65900 82780
rect -66100 82550 -66090 82750
rect -66020 82550 -65980 82750
rect -65910 82550 -65900 82750
rect -66100 82520 -65900 82550
rect -65600 82750 -65400 82780
rect -65600 82550 -65590 82750
rect -65520 82550 -65480 82750
rect -65410 82550 -65400 82750
rect -65600 82520 -65400 82550
rect -65100 82750 -64900 82780
rect -65100 82550 -65090 82750
rect -65020 82550 -64980 82750
rect -64910 82550 -64900 82750
rect -65100 82520 -64900 82550
rect -64600 82750 -64400 82780
rect -64600 82550 -64590 82750
rect -64520 82550 -64480 82750
rect -64410 82550 -64400 82750
rect -64600 82520 -64400 82550
rect -64100 82750 -63900 82780
rect -64100 82550 -64090 82750
rect -64020 82550 -63980 82750
rect -63910 82550 -63900 82750
rect -64100 82520 -63900 82550
rect -63600 82750 -63400 82780
rect -63600 82550 -63590 82750
rect -63520 82550 -63480 82750
rect -63410 82550 -63400 82750
rect -63600 82520 -63400 82550
rect -63100 82750 -62900 82780
rect -63100 82550 -63090 82750
rect -63020 82550 -62980 82750
rect -62910 82550 -62900 82750
rect -63100 82520 -62900 82550
rect -62600 82750 -62400 82780
rect -62600 82550 -62590 82750
rect -62520 82550 -62480 82750
rect -62410 82550 -62400 82750
rect -62600 82520 -62400 82550
rect -62100 82750 -61900 82780
rect -62100 82550 -62090 82750
rect -62020 82550 -61980 82750
rect -61910 82550 -61900 82750
rect -62100 82520 -61900 82550
rect -61600 82750 -61400 82780
rect -61600 82550 -61590 82750
rect -61520 82550 -61480 82750
rect -61410 82550 -61400 82750
rect -61600 82520 -61400 82550
rect -61100 82750 -60900 82780
rect -61100 82550 -61090 82750
rect -61020 82550 -60980 82750
rect -60910 82550 -60900 82750
rect -61100 82520 -60900 82550
rect -60600 82750 -60400 82780
rect -60600 82550 -60590 82750
rect -60520 82550 -60480 82750
rect -60410 82550 -60400 82750
rect -60600 82520 -60400 82550
rect -60100 82750 -59900 82780
rect -60100 82550 -60090 82750
rect -60020 82550 -59980 82750
rect -59910 82550 -59900 82750
rect -60100 82520 -59900 82550
rect -59600 82750 -59400 82780
rect -59600 82550 -59590 82750
rect -59520 82550 -59480 82750
rect -59410 82550 -59400 82750
rect -59600 82520 -59400 82550
rect -59100 82750 -58900 82780
rect -59100 82550 -59090 82750
rect -59020 82550 -58980 82750
rect -58910 82550 -58900 82750
rect -59100 82520 -58900 82550
rect -58600 82750 -58400 82780
rect -58600 82550 -58590 82750
rect -58520 82550 -58480 82750
rect -58410 82550 -58400 82750
rect -58600 82520 -58400 82550
rect -58100 82750 -57900 82780
rect -58100 82550 -58090 82750
rect -58020 82550 -57980 82750
rect -57910 82550 -57900 82750
rect -58100 82520 -57900 82550
rect -57600 82750 -57400 82780
rect -57600 82550 -57590 82750
rect -57520 82550 -57480 82750
rect -57410 82550 -57400 82750
rect -57600 82520 -57400 82550
rect -57100 82750 -56900 82780
rect -57100 82550 -57090 82750
rect -57020 82550 -56980 82750
rect -56910 82550 -56900 82750
rect -57100 82520 -56900 82550
rect -56600 82750 -56400 82780
rect -56600 82550 -56590 82750
rect -56520 82550 -56480 82750
rect -56410 82550 -56400 82750
rect -56600 82520 -56400 82550
rect -56100 82750 -55900 82780
rect -56100 82550 -56090 82750
rect -56020 82550 -55980 82750
rect -55910 82550 -55900 82750
rect -56100 82520 -55900 82550
rect -55600 82750 -55400 82780
rect -55600 82550 -55590 82750
rect -55520 82550 -55480 82750
rect -55410 82550 -55400 82750
rect -55600 82520 -55400 82550
rect -55100 82750 -54900 82780
rect -55100 82550 -55090 82750
rect -55020 82550 -54980 82750
rect -54910 82550 -54900 82750
rect -55100 82520 -54900 82550
rect -54600 82750 -54400 82780
rect -54600 82550 -54590 82750
rect -54520 82550 -54480 82750
rect -54410 82550 -54400 82750
rect -54600 82520 -54400 82550
rect -54100 82750 -53900 82780
rect -54100 82550 -54090 82750
rect -54020 82550 -53980 82750
rect -53910 82550 -53900 82750
rect -54100 82520 -53900 82550
rect -53600 82750 -53400 82780
rect -53600 82550 -53590 82750
rect -53520 82550 -53480 82750
rect -53410 82550 -53400 82750
rect -53600 82520 -53400 82550
rect -53100 82750 -52900 82780
rect -53100 82550 -53090 82750
rect -53020 82550 -52980 82750
rect -52910 82550 -52900 82750
rect -53100 82520 -52900 82550
rect -52600 82750 -52400 82780
rect -52600 82550 -52590 82750
rect -52520 82550 -52480 82750
rect -52410 82550 -52400 82750
rect -52600 82520 -52400 82550
rect -52100 82750 -51900 82780
rect -52100 82550 -52090 82750
rect -52020 82550 -51980 82750
rect -51910 82550 -51900 82750
rect -52100 82520 -51900 82550
rect -51600 82750 -51400 82780
rect -51600 82550 -51590 82750
rect -51520 82550 -51480 82750
rect -51410 82550 -51400 82750
rect -51600 82520 -51400 82550
rect -51100 82750 -50900 82780
rect -51100 82550 -51090 82750
rect -51020 82550 -50980 82750
rect -50910 82550 -50900 82750
rect -51100 82520 -50900 82550
rect -50600 82750 -50400 82780
rect -50600 82550 -50590 82750
rect -50520 82550 -50480 82750
rect -50410 82550 -50400 82750
rect -50600 82520 -50400 82550
rect -50100 82750 -49900 82780
rect -50100 82550 -50090 82750
rect -50020 82550 -49980 82750
rect -49910 82550 -49900 82750
rect -50100 82520 -49900 82550
rect -49600 82750 -49400 82780
rect -49600 82550 -49590 82750
rect -49520 82550 -49480 82750
rect -49410 82550 -49400 82750
rect -49600 82520 -49400 82550
rect -49100 82750 -48900 82780
rect -49100 82550 -49090 82750
rect -49020 82550 -48980 82750
rect -48910 82550 -48900 82750
rect -49100 82520 -48900 82550
rect -48600 82750 -48400 82780
rect -48600 82550 -48590 82750
rect -48520 82550 -48480 82750
rect -48410 82550 -48400 82750
rect -48600 82520 -48400 82550
rect -48100 82750 -47900 82780
rect -48100 82550 -48090 82750
rect -48020 82550 -47980 82750
rect -47910 82550 -47900 82750
rect -48100 82520 -47900 82550
rect -47600 82750 -47400 82780
rect -47600 82550 -47590 82750
rect -47520 82550 -47480 82750
rect -47410 82550 -47400 82750
rect -47600 82520 -47400 82550
rect -47100 82750 -46900 82780
rect -47100 82550 -47090 82750
rect -47020 82550 -46980 82750
rect -46910 82550 -46900 82750
rect -47100 82520 -46900 82550
rect -46600 82750 -46400 82780
rect -46600 82550 -46590 82750
rect -46520 82550 -46480 82750
rect -46410 82550 -46400 82750
rect -46600 82520 -46400 82550
rect -46100 82750 -45900 82780
rect -46100 82550 -46090 82750
rect -46020 82550 -45980 82750
rect -45910 82550 -45900 82750
rect -46100 82520 -45900 82550
rect -45600 82750 -45400 82780
rect -45600 82550 -45590 82750
rect -45520 82550 -45480 82750
rect -45410 82550 -45400 82750
rect -45600 82520 -45400 82550
rect -45100 82750 -44900 82780
rect -45100 82550 -45090 82750
rect -45020 82550 -44980 82750
rect -44910 82550 -44900 82750
rect -45100 82520 -44900 82550
rect -44600 82750 -44400 82780
rect -44600 82550 -44590 82750
rect -44520 82550 -44480 82750
rect -44410 82550 -44400 82750
rect -44600 82520 -44400 82550
rect -44100 82750 -43900 82780
rect -44100 82550 -44090 82750
rect -44020 82550 -43980 82750
rect -43910 82550 -43900 82750
rect -44100 82520 -43900 82550
rect -43600 82750 -43400 82780
rect -43600 82550 -43590 82750
rect -43520 82550 -43480 82750
rect -43410 82550 -43400 82750
rect -43600 82520 -43400 82550
rect -43100 82750 -42900 82780
rect -43100 82550 -43090 82750
rect -43020 82550 -42980 82750
rect -42910 82550 -42900 82750
rect -43100 82520 -42900 82550
rect -42600 82750 -42400 82780
rect -42600 82550 -42590 82750
rect -42520 82550 -42480 82750
rect -42410 82550 -42400 82750
rect -42600 82520 -42400 82550
rect -42100 82750 -41900 82780
rect -42100 82550 -42090 82750
rect -42020 82550 -41980 82750
rect -41910 82550 -41900 82750
rect -42100 82520 -41900 82550
rect -41600 82750 -41400 82780
rect -41600 82550 -41590 82750
rect -41520 82550 -41480 82750
rect -41410 82550 -41400 82750
rect -41600 82520 -41400 82550
rect -41100 82750 -40900 82780
rect -41100 82550 -41090 82750
rect -41020 82550 -40980 82750
rect -40910 82550 -40900 82750
rect -41100 82520 -40900 82550
rect -40600 82750 -40400 82780
rect -40600 82550 -40590 82750
rect -40520 82550 -40480 82750
rect -40410 82550 -40400 82750
rect -40600 82520 -40400 82550
rect -40100 82750 -39900 82780
rect -40100 82550 -40090 82750
rect -40020 82550 -39980 82750
rect -39910 82550 -39900 82750
rect -40100 82520 -39900 82550
rect -39600 82750 -39400 82780
rect -39600 82550 -39590 82750
rect -39520 82550 -39480 82750
rect -39410 82550 -39400 82750
rect -39600 82520 -39400 82550
rect -39100 82750 -38900 82780
rect -39100 82550 -39090 82750
rect -39020 82550 -38980 82750
rect -38910 82550 -38900 82750
rect -39100 82520 -38900 82550
rect -38600 82750 -38400 82780
rect -38600 82550 -38590 82750
rect -38520 82550 -38480 82750
rect -38410 82550 -38400 82750
rect -38600 82520 -38400 82550
rect -38100 82750 -37900 82780
rect -38100 82550 -38090 82750
rect -38020 82550 -37980 82750
rect -37910 82550 -37900 82750
rect -38100 82520 -37900 82550
rect -37600 82750 -37400 82780
rect -37600 82550 -37590 82750
rect -37520 82550 -37480 82750
rect -37410 82550 -37400 82750
rect -37600 82520 -37400 82550
rect -37100 82750 -36900 82780
rect -37100 82550 -37090 82750
rect -37020 82550 -36980 82750
rect -36910 82550 -36900 82750
rect -37100 82520 -36900 82550
rect -36600 82750 -36400 82780
rect -36600 82550 -36590 82750
rect -36520 82550 -36480 82750
rect -36410 82550 -36400 82750
rect -36600 82520 -36400 82550
rect -36100 82750 -35900 82780
rect -36100 82550 -36090 82750
rect -36020 82550 -35980 82750
rect -35910 82550 -35900 82750
rect -36100 82520 -35900 82550
rect -35600 82750 -35400 82780
rect -35600 82550 -35590 82750
rect -35520 82550 -35480 82750
rect -35410 82550 -35400 82750
rect -35600 82520 -35400 82550
rect -35100 82750 -34900 82780
rect -35100 82550 -35090 82750
rect -35020 82550 -34980 82750
rect -34910 82550 -34900 82750
rect -35100 82520 -34900 82550
rect -34600 82750 -34400 82780
rect -34600 82550 -34590 82750
rect -34520 82550 -34480 82750
rect -34410 82550 -34400 82750
rect -34600 82520 -34400 82550
rect -34100 82750 -33900 82780
rect -34100 82550 -34090 82750
rect -34020 82550 -33980 82750
rect -33910 82550 -33900 82750
rect -34100 82520 -33900 82550
rect -33600 82750 -33400 82780
rect -33600 82550 -33590 82750
rect -33520 82550 -33480 82750
rect -33410 82550 -33400 82750
rect -33600 82520 -33400 82550
rect -33100 82750 -32900 82780
rect -33100 82550 -33090 82750
rect -33020 82550 -32980 82750
rect -32910 82550 -32900 82750
rect -33100 82520 -32900 82550
rect -32600 82750 -32400 82780
rect -32600 82550 -32590 82750
rect -32520 82550 -32480 82750
rect -32410 82550 -32400 82750
rect -32600 82520 -32400 82550
rect -32100 82750 -31900 82780
rect -32100 82550 -32090 82750
rect -32020 82550 -31980 82750
rect -31910 82550 -31900 82750
rect -32100 82520 -31900 82550
rect -31600 82750 -31400 82780
rect -31600 82550 -31590 82750
rect -31520 82550 -31480 82750
rect -31410 82550 -31400 82750
rect -31600 82520 -31400 82550
rect -31100 82750 -30900 82780
rect -31100 82550 -31090 82750
rect -31020 82550 -30980 82750
rect -30910 82550 -30900 82750
rect -31100 82520 -30900 82550
rect -30600 82750 -30400 82780
rect -30600 82550 -30590 82750
rect -30520 82550 -30480 82750
rect -30410 82550 -30400 82750
rect -30600 82520 -30400 82550
rect -30100 82750 -29900 82780
rect -30100 82550 -30090 82750
rect -30020 82550 -29980 82750
rect -29910 82550 -29900 82750
rect -30100 82520 -29900 82550
rect -29600 82750 -29400 82780
rect -29600 82550 -29590 82750
rect -29520 82550 -29480 82750
rect -29410 82550 -29400 82750
rect -29600 82520 -29400 82550
rect -29100 82750 -28900 82780
rect -29100 82550 -29090 82750
rect -29020 82550 -28980 82750
rect -28910 82550 -28900 82750
rect -29100 82520 -28900 82550
rect -28600 82750 -28400 82780
rect -28600 82550 -28590 82750
rect -28520 82550 -28480 82750
rect -28410 82550 -28400 82750
rect -28600 82520 -28400 82550
rect -28100 82750 -27900 82780
rect -28100 82550 -28090 82750
rect -28020 82550 -27980 82750
rect -27910 82550 -27900 82750
rect -28100 82520 -27900 82550
rect -27600 82750 -27400 82780
rect -27600 82550 -27590 82750
rect -27520 82550 -27480 82750
rect -27410 82550 -27400 82750
rect -27600 82520 -27400 82550
rect -27100 82750 -26900 82780
rect -27100 82550 -27090 82750
rect -27020 82550 -26980 82750
rect -26910 82550 -26900 82750
rect -27100 82520 -26900 82550
rect -26600 82750 -26400 82780
rect -26600 82550 -26590 82750
rect -26520 82550 -26480 82750
rect -26410 82550 -26400 82750
rect -26600 82520 -26400 82550
rect -26100 82750 -25900 82780
rect -26100 82550 -26090 82750
rect -26020 82550 -25980 82750
rect -25910 82550 -25900 82750
rect -26100 82520 -25900 82550
rect -25600 82750 -25400 82780
rect -25600 82550 -25590 82750
rect -25520 82550 -25480 82750
rect -25410 82550 -25400 82750
rect -25600 82520 -25400 82550
rect -25100 82750 -24900 82780
rect -25100 82550 -25090 82750
rect -25020 82550 -24980 82750
rect -24910 82550 -24900 82750
rect -25100 82520 -24900 82550
rect -24600 82750 -24400 82780
rect -24600 82550 -24590 82750
rect -24520 82550 -24480 82750
rect -24410 82550 -24400 82750
rect -24600 82520 -24400 82550
rect -24100 82750 -23900 82780
rect -24100 82550 -24090 82750
rect -24020 82550 -23980 82750
rect -23910 82550 -23900 82750
rect -24100 82520 -23900 82550
rect -23600 82750 -23400 82780
rect -23600 82550 -23590 82750
rect -23520 82550 -23480 82750
rect -23410 82550 -23400 82750
rect -23600 82520 -23400 82550
rect -23100 82750 -22900 82780
rect -23100 82550 -23090 82750
rect -23020 82550 -22980 82750
rect -22910 82550 -22900 82750
rect -23100 82520 -22900 82550
rect -22600 82750 -22400 82780
rect -22600 82550 -22590 82750
rect -22520 82550 -22480 82750
rect -22410 82550 -22400 82750
rect -22600 82520 -22400 82550
rect -22100 82750 -21900 82780
rect -22100 82550 -22090 82750
rect -22020 82550 -21980 82750
rect -21910 82550 -21900 82750
rect -22100 82520 -21900 82550
rect -21600 82750 -21400 82780
rect -21600 82550 -21590 82750
rect -21520 82550 -21480 82750
rect -21410 82550 -21400 82750
rect -21600 82520 -21400 82550
rect -21100 82750 -20900 82780
rect -21100 82550 -21090 82750
rect -21020 82550 -20980 82750
rect -20910 82550 -20900 82750
rect -21100 82520 -20900 82550
rect -20600 82750 -20400 82780
rect -20600 82550 -20590 82750
rect -20520 82550 -20480 82750
rect -20410 82550 -20400 82750
rect -20600 82520 -20400 82550
rect -20100 82750 -19900 82780
rect -20100 82550 -20090 82750
rect -20020 82550 -19980 82750
rect -19910 82550 -19900 82750
rect -20100 82520 -19900 82550
rect -19600 82750 -19400 82780
rect -19600 82550 -19590 82750
rect -19520 82550 -19480 82750
rect -19410 82550 -19400 82750
rect -19600 82520 -19400 82550
rect -19100 82750 -18900 82780
rect -19100 82550 -19090 82750
rect -19020 82550 -18980 82750
rect -18910 82550 -18900 82750
rect -19100 82520 -18900 82550
rect -18600 82750 -18400 82780
rect -18600 82550 -18590 82750
rect -18520 82550 -18480 82750
rect -18410 82550 -18400 82750
rect -18600 82520 -18400 82550
rect -18100 82750 -17900 82780
rect -18100 82550 -18090 82750
rect -18020 82550 -17980 82750
rect -17910 82550 -17900 82750
rect -18100 82520 -17900 82550
rect -17600 82750 -17400 82780
rect -17600 82550 -17590 82750
rect -17520 82550 -17480 82750
rect -17410 82550 -17400 82750
rect -17600 82520 -17400 82550
rect -17100 82750 -16900 82780
rect -17100 82550 -17090 82750
rect -17020 82550 -16980 82750
rect -16910 82550 -16900 82750
rect -17100 82520 -16900 82550
rect -16600 82750 -16400 82780
rect -16600 82550 -16590 82750
rect -16520 82550 -16480 82750
rect -16410 82550 -16400 82750
rect -16600 82520 -16400 82550
rect -16100 82750 -15900 82780
rect -16100 82550 -16090 82750
rect -16020 82550 -15980 82750
rect -15910 82550 -15900 82750
rect -16100 82520 -15900 82550
rect -15600 82750 -15400 82780
rect -15600 82550 -15590 82750
rect -15520 82550 -15480 82750
rect -15410 82550 -15400 82750
rect -15600 82520 -15400 82550
rect -15100 82750 -14900 82780
rect -15100 82550 -15090 82750
rect -15020 82550 -14980 82750
rect -14910 82550 -14900 82750
rect -15100 82520 -14900 82550
rect -14600 82750 -14400 82780
rect -14600 82550 -14590 82750
rect -14520 82550 -14480 82750
rect -14410 82550 -14400 82750
rect -14600 82520 -14400 82550
rect -14100 82750 -13900 82780
rect -14100 82550 -14090 82750
rect -14020 82550 -13980 82750
rect -13910 82550 -13900 82750
rect -14100 82520 -13900 82550
rect -13600 82750 -13400 82780
rect -13600 82550 -13590 82750
rect -13520 82550 -13480 82750
rect -13410 82550 -13400 82750
rect -13600 82520 -13400 82550
rect -13100 82750 -12900 82780
rect -13100 82550 -13090 82750
rect -13020 82550 -12980 82750
rect -12910 82550 -12900 82750
rect -13100 82520 -12900 82550
rect -12600 82750 -12400 82780
rect -12600 82550 -12590 82750
rect -12520 82550 -12480 82750
rect -12410 82550 -12400 82750
rect -12600 82520 -12400 82550
rect -12100 82750 -11900 82780
rect -12100 82550 -12090 82750
rect -12020 82550 -11980 82750
rect -11910 82550 -11900 82750
rect -12100 82520 -11900 82550
rect -11600 82750 -11400 82780
rect -11600 82550 -11590 82750
rect -11520 82550 -11480 82750
rect -11410 82550 -11400 82750
rect -11600 82520 -11400 82550
rect -11100 82750 -10900 82780
rect -11100 82550 -11090 82750
rect -11020 82550 -10980 82750
rect -10910 82550 -10900 82750
rect -11100 82520 -10900 82550
rect -10600 82750 -10400 82780
rect -10600 82550 -10590 82750
rect -10520 82550 -10480 82750
rect -10410 82550 -10400 82750
rect -10600 82520 -10400 82550
rect -10100 82750 -9900 82780
rect -10100 82550 -10090 82750
rect -10020 82550 -9980 82750
rect -9910 82550 -9900 82750
rect -10100 82520 -9900 82550
rect -9600 82750 -9400 82780
rect -9600 82550 -9590 82750
rect -9520 82550 -9480 82750
rect -9410 82550 -9400 82750
rect -9600 82520 -9400 82550
rect -9100 82750 -8900 82780
rect -9100 82550 -9090 82750
rect -9020 82550 -8980 82750
rect -8910 82550 -8900 82750
rect -9100 82520 -8900 82550
rect -8600 82750 -8400 82780
rect -8600 82550 -8590 82750
rect -8520 82550 -8480 82750
rect -8410 82550 -8400 82750
rect -8600 82520 -8400 82550
rect -8100 82750 -7900 82780
rect -8100 82550 -8090 82750
rect -8020 82550 -7980 82750
rect -7910 82550 -7900 82750
rect -8100 82520 -7900 82550
rect -7600 82750 -7400 82780
rect -7600 82550 -7590 82750
rect -7520 82550 -7480 82750
rect -7410 82550 -7400 82750
rect -7600 82520 -7400 82550
rect -7100 82750 -6900 82780
rect -7100 82550 -7090 82750
rect -7020 82550 -6980 82750
rect -6910 82550 -6900 82750
rect -7100 82520 -6900 82550
rect -6600 82750 -6400 82780
rect -6600 82550 -6590 82750
rect -6520 82550 -6480 82750
rect -6410 82550 -6400 82750
rect -6600 82520 -6400 82550
rect -6100 82750 -5900 82780
rect -6100 82550 -6090 82750
rect -6020 82550 -5980 82750
rect -5910 82550 -5900 82750
rect -6100 82520 -5900 82550
rect -5600 82750 -5400 82780
rect -5600 82550 -5590 82750
rect -5520 82550 -5480 82750
rect -5410 82550 -5400 82750
rect -5600 82520 -5400 82550
rect -5100 82750 -4900 82780
rect -5100 82550 -5090 82750
rect -5020 82550 -4980 82750
rect -4910 82550 -4900 82750
rect -5100 82520 -4900 82550
rect -4600 82750 -4400 82780
rect -4600 82550 -4590 82750
rect -4520 82550 -4480 82750
rect -4410 82550 -4400 82750
rect -4600 82520 -4400 82550
rect -4100 82750 -3900 82780
rect -4100 82550 -4090 82750
rect -4020 82550 -3980 82750
rect -3910 82550 -3900 82750
rect -4100 82520 -3900 82550
rect -3600 82750 -3400 82780
rect -3600 82550 -3590 82750
rect -3520 82550 -3480 82750
rect -3410 82550 -3400 82750
rect -3600 82520 -3400 82550
rect -3100 82750 -2900 82780
rect -3100 82550 -3090 82750
rect -3020 82550 -2980 82750
rect -2910 82550 -2900 82750
rect -3100 82520 -2900 82550
rect -2600 82750 -2400 82780
rect -2600 82550 -2590 82750
rect -2520 82550 -2480 82750
rect -2410 82550 -2400 82750
rect -2600 82520 -2400 82550
rect -2100 82750 -1900 82780
rect -2100 82550 -2090 82750
rect -2020 82550 -1980 82750
rect -1910 82550 -1900 82750
rect -2100 82520 -1900 82550
rect -1600 82750 -1400 82780
rect -1600 82550 -1590 82750
rect -1520 82550 -1480 82750
rect -1410 82550 -1400 82750
rect -1600 82520 -1400 82550
rect -1100 82750 -900 82780
rect -1100 82550 -1090 82750
rect -1020 82550 -980 82750
rect -910 82550 -900 82750
rect -1100 82520 -900 82550
rect -600 82750 -400 82780
rect -600 82550 -590 82750
rect -520 82550 -480 82750
rect -410 82550 -400 82750
rect -600 82520 -400 82550
rect -100 82750 100 82780
rect -100 82550 -90 82750
rect -20 82550 20 82750
rect 90 82550 100 82750
rect -100 82520 100 82550
rect 400 82750 600 82780
rect 400 82550 410 82750
rect 480 82550 520 82750
rect 590 82550 600 82750
rect 400 82520 600 82550
rect 900 82750 1100 82780
rect 900 82550 910 82750
rect 980 82550 1020 82750
rect 1090 82550 1100 82750
rect 900 82520 1100 82550
rect 1400 82750 1600 82780
rect 1400 82550 1410 82750
rect 1480 82550 1520 82750
rect 1590 82550 1600 82750
rect 1400 82520 1600 82550
rect 1900 82750 2100 82780
rect 1900 82550 1910 82750
rect 1980 82550 2020 82750
rect 2090 82550 2100 82750
rect 1900 82520 2100 82550
rect 2400 82750 2600 82780
rect 2400 82550 2410 82750
rect 2480 82550 2520 82750
rect 2590 82550 2600 82750
rect 2400 82520 2600 82550
rect 2900 82750 3100 82780
rect 2900 82550 2910 82750
rect 2980 82550 3020 82750
rect 3090 82550 3100 82750
rect 2900 82520 3100 82550
rect 3400 82750 3600 82780
rect 3400 82550 3410 82750
rect 3480 82550 3520 82750
rect 3590 82550 3600 82750
rect 3400 82520 3600 82550
rect 3900 82750 4100 82780
rect 3900 82550 3910 82750
rect 3980 82550 4020 82750
rect 4090 82550 4100 82750
rect 3900 82520 4100 82550
rect 4400 82750 4600 82780
rect 4400 82550 4410 82750
rect 4480 82550 4520 82750
rect 4590 82550 4600 82750
rect 4400 82520 4600 82550
rect 4900 82750 5100 82780
rect 4900 82550 4910 82750
rect 4980 82550 5020 82750
rect 5090 82550 5100 82750
rect 4900 82520 5100 82550
rect 5400 82750 5600 82780
rect 5400 82550 5410 82750
rect 5480 82550 5520 82750
rect 5590 82550 5600 82750
rect 5400 82520 5600 82550
rect 5900 82750 6100 82780
rect 5900 82550 5910 82750
rect 5980 82550 6020 82750
rect 6090 82550 6100 82750
rect 5900 82520 6100 82550
rect 6400 82750 6600 82780
rect 6400 82550 6410 82750
rect 6480 82550 6520 82750
rect 6590 82550 6600 82750
rect 6400 82520 6600 82550
rect 6900 82750 7100 82780
rect 6900 82550 6910 82750
rect 6980 82550 7020 82750
rect 7090 82550 7100 82750
rect 6900 82520 7100 82550
rect 7400 82750 7600 82780
rect 7400 82550 7410 82750
rect 7480 82550 7520 82750
rect 7590 82550 7600 82750
rect 7400 82520 7600 82550
rect 7900 82750 8100 82780
rect 7900 82550 7910 82750
rect 7980 82550 8020 82750
rect 8090 82550 8100 82750
rect 7900 82520 8100 82550
rect 8400 82750 8600 82780
rect 8400 82550 8410 82750
rect 8480 82550 8520 82750
rect 8590 82550 8600 82750
rect 8400 82520 8600 82550
rect 8900 82750 9100 82780
rect 8900 82550 8910 82750
rect 8980 82550 9020 82750
rect 9090 82550 9100 82750
rect 8900 82520 9100 82550
rect 9400 82750 9600 82780
rect 9400 82550 9410 82750
rect 9480 82550 9520 82750
rect 9590 82550 9600 82750
rect 9400 82520 9600 82550
rect 9900 82750 10100 82780
rect 9900 82550 9910 82750
rect 9980 82550 10020 82750
rect 10090 82550 10100 82750
rect 9900 82520 10100 82550
rect 10400 82750 10600 82780
rect 10400 82550 10410 82750
rect 10480 82550 10520 82750
rect 10590 82550 10600 82750
rect 10400 82520 10600 82550
rect 10900 82750 11100 82780
rect 10900 82550 10910 82750
rect 10980 82550 11020 82750
rect 11090 82550 11100 82750
rect 10900 82520 11100 82550
rect 11400 82750 11600 82780
rect 11400 82550 11410 82750
rect 11480 82550 11520 82750
rect 11590 82550 11600 82750
rect 11400 82520 11600 82550
rect 11900 82750 12100 82780
rect 11900 82550 11910 82750
rect 11980 82550 12020 82750
rect 12090 82550 12100 82750
rect 11900 82520 12100 82550
rect 12400 82750 12600 82780
rect 12400 82550 12410 82750
rect 12480 82550 12520 82750
rect 12590 82550 12600 82750
rect 12400 82520 12600 82550
rect 12900 82750 13100 82780
rect 12900 82550 12910 82750
rect 12980 82550 13020 82750
rect 13090 82550 13100 82750
rect 12900 82520 13100 82550
rect 13400 82750 13600 82780
rect 13400 82550 13410 82750
rect 13480 82550 13520 82750
rect 13590 82550 13600 82750
rect 13400 82520 13600 82550
rect 13900 82750 14100 82780
rect 13900 82550 13910 82750
rect 13980 82550 14020 82750
rect 14090 82550 14100 82750
rect 13900 82520 14100 82550
rect 14400 82750 14600 82780
rect 14400 82550 14410 82750
rect 14480 82550 14520 82750
rect 14590 82550 14600 82750
rect 14400 82520 14600 82550
rect 14900 82750 15100 82780
rect 14900 82550 14910 82750
rect 14980 82550 15020 82750
rect 15090 82550 15100 82750
rect 14900 82520 15100 82550
rect 15400 82750 15600 82780
rect 15400 82550 15410 82750
rect 15480 82550 15520 82750
rect 15590 82550 15600 82750
rect 15400 82520 15600 82550
rect 15900 82750 16100 82780
rect 15900 82550 15910 82750
rect 15980 82550 16020 82750
rect 16090 82550 16100 82750
rect 15900 82520 16100 82550
rect 16400 82750 16600 82780
rect 16400 82550 16410 82750
rect 16480 82550 16520 82750
rect 16590 82550 16600 82750
rect 16400 82520 16600 82550
rect 16900 82750 17100 82780
rect 16900 82550 16910 82750
rect 16980 82550 17020 82750
rect 17090 82550 17100 82750
rect 16900 82520 17100 82550
rect 17400 82750 17600 82780
rect 17400 82550 17410 82750
rect 17480 82550 17520 82750
rect 17590 82550 17600 82750
rect 17400 82520 17600 82550
rect 17900 82750 18100 82780
rect 17900 82550 17910 82750
rect 17980 82550 18020 82750
rect 18090 82550 18100 82750
rect 17900 82520 18100 82550
rect 18400 82750 18600 82780
rect 18400 82550 18410 82750
rect 18480 82550 18520 82750
rect 18590 82550 18600 82750
rect 18400 82520 18600 82550
rect 18900 82750 19100 82780
rect 18900 82550 18910 82750
rect 18980 82550 19020 82750
rect 19090 82550 19100 82750
rect 18900 82520 19100 82550
rect 19400 82750 19600 82780
rect 19400 82550 19410 82750
rect 19480 82550 19520 82750
rect 19590 82550 19600 82750
rect 19400 82520 19600 82550
rect 19900 82750 20100 82780
rect 19900 82550 19910 82750
rect 19980 82550 20020 82750
rect 20090 82550 20100 82750
rect 19900 82520 20100 82550
rect 20400 82750 20600 82780
rect 20400 82550 20410 82750
rect 20480 82550 20520 82750
rect 20590 82550 20600 82750
rect 20400 82520 20600 82550
rect 20900 82750 21100 82780
rect 20900 82550 20910 82750
rect 20980 82550 21020 82750
rect 21090 82550 21100 82750
rect 20900 82520 21100 82550
rect 21400 82750 21600 82780
rect 21400 82550 21410 82750
rect 21480 82550 21520 82750
rect 21590 82550 21600 82750
rect 21400 82520 21600 82550
rect 21900 82750 22100 82780
rect 21900 82550 21910 82750
rect 21980 82550 22020 82750
rect 22090 82550 22100 82750
rect 21900 82520 22100 82550
rect 22400 82750 22600 82780
rect 22400 82550 22410 82750
rect 22480 82550 22520 82750
rect 22590 82550 22600 82750
rect 22400 82520 22600 82550
rect 22900 82750 23100 82780
rect 22900 82550 22910 82750
rect 22980 82550 23020 82750
rect 23090 82550 23100 82750
rect 22900 82520 23100 82550
rect 23400 82750 23600 82780
rect 23400 82550 23410 82750
rect 23480 82550 23520 82750
rect 23590 82550 23600 82750
rect 23400 82520 23600 82550
rect 23900 82750 24100 82780
rect 23900 82550 23910 82750
rect 23980 82550 24020 82750
rect 24090 82550 24100 82750
rect 23900 82520 24100 82550
rect 24400 82750 24600 82780
rect 24400 82550 24410 82750
rect 24480 82550 24520 82750
rect 24590 82550 24600 82750
rect 24400 82520 24600 82550
rect 24900 82750 25100 82780
rect 24900 82550 24910 82750
rect 24980 82550 25020 82750
rect 25090 82550 25100 82750
rect 24900 82520 25100 82550
rect 25400 82750 25600 82780
rect 25400 82550 25410 82750
rect 25480 82550 25520 82750
rect 25590 82550 25600 82750
rect 25400 82520 25600 82550
rect 25900 82750 26100 82780
rect 25900 82550 25910 82750
rect 25980 82550 26020 82750
rect 26090 82550 26100 82750
rect 25900 82520 26100 82550
rect 26400 82750 26600 82780
rect 26400 82550 26410 82750
rect 26480 82550 26520 82750
rect 26590 82550 26600 82750
rect 26400 82520 26600 82550
rect 26900 82750 27100 82780
rect 26900 82550 26910 82750
rect 26980 82550 27020 82750
rect 27090 82550 27100 82750
rect 26900 82520 27100 82550
rect 27400 82750 27600 82780
rect 27400 82550 27410 82750
rect 27480 82550 27520 82750
rect 27590 82550 27600 82750
rect 27400 82520 27600 82550
rect 27900 82750 28100 82780
rect 27900 82550 27910 82750
rect 27980 82550 28020 82750
rect 28090 82550 28100 82750
rect 27900 82520 28100 82550
rect 28400 82750 28600 82780
rect 28400 82550 28410 82750
rect 28480 82550 28520 82750
rect 28590 82550 28600 82750
rect 28400 82520 28600 82550
rect 28900 82750 29100 82780
rect 28900 82550 28910 82750
rect 28980 82550 29020 82750
rect 29090 82550 29100 82750
rect 28900 82520 29100 82550
rect 29400 82750 29600 82780
rect 29400 82550 29410 82750
rect 29480 82550 29520 82750
rect 29590 82550 29600 82750
rect 29400 82520 29600 82550
rect 29900 82750 30100 82780
rect 29900 82550 29910 82750
rect 29980 82550 30020 82750
rect 30090 82550 30100 82750
rect 29900 82520 30100 82550
rect 30400 82750 30600 82780
rect 30400 82550 30410 82750
rect 30480 82550 30520 82750
rect 30590 82550 30600 82750
rect 30400 82520 30600 82550
rect 30900 82750 31100 82780
rect 30900 82550 30910 82750
rect 30980 82550 31020 82750
rect 31090 82550 31100 82750
rect 30900 82520 31100 82550
rect 31400 82750 31600 82780
rect 31400 82550 31410 82750
rect 31480 82550 31520 82750
rect 31590 82550 31600 82750
rect 31400 82520 31600 82550
rect 31900 82750 32100 82780
rect 31900 82550 31910 82750
rect 31980 82550 32020 82750
rect 32090 82550 32100 82750
rect 31900 82520 32100 82550
rect 32400 82750 32600 82780
rect 32400 82550 32410 82750
rect 32480 82550 32520 82750
rect 32590 82550 32600 82750
rect 32400 82520 32600 82550
rect 32900 82750 33100 82780
rect 32900 82550 32910 82750
rect 32980 82550 33020 82750
rect 33090 82550 33100 82750
rect 32900 82520 33100 82550
rect 33400 82750 33600 82780
rect 33400 82550 33410 82750
rect 33480 82550 33520 82750
rect 33590 82550 33600 82750
rect 33400 82520 33600 82550
rect 33900 82750 34100 82780
rect 33900 82550 33910 82750
rect 33980 82550 34020 82750
rect 34090 82550 34100 82750
rect 33900 82520 34100 82550
rect 34400 82750 34600 82780
rect 34400 82550 34410 82750
rect 34480 82550 34520 82750
rect 34590 82550 34600 82750
rect 34400 82520 34600 82550
rect 34900 82750 35100 82780
rect 34900 82550 34910 82750
rect 34980 82550 35020 82750
rect 35090 82550 35100 82750
rect 34900 82520 35100 82550
rect 35400 82750 35600 82780
rect 35400 82550 35410 82750
rect 35480 82550 35520 82750
rect 35590 82550 35600 82750
rect 35400 82520 35600 82550
rect 35900 82750 36100 82780
rect 35900 82550 35910 82750
rect 35980 82550 36020 82750
rect 36090 82550 36100 82750
rect 35900 82520 36100 82550
rect 36400 82750 36600 82780
rect 36400 82550 36410 82750
rect 36480 82550 36520 82750
rect 36590 82550 36600 82750
rect 36400 82520 36600 82550
rect 36900 82750 37100 82780
rect 36900 82550 36910 82750
rect 36980 82550 37020 82750
rect 37090 82550 37100 82750
rect 36900 82520 37100 82550
rect 37400 82750 37600 82780
rect 37400 82550 37410 82750
rect 37480 82550 37520 82750
rect 37590 82550 37600 82750
rect 37400 82520 37600 82550
rect 37900 82750 38100 82780
rect 37900 82550 37910 82750
rect 37980 82550 38020 82750
rect 38090 82550 38100 82750
rect 37900 82520 38100 82550
rect 38400 82750 38600 82780
rect 38400 82550 38410 82750
rect 38480 82550 38520 82750
rect 38590 82550 38600 82750
rect 38400 82520 38600 82550
rect 38900 82750 39100 82780
rect 38900 82550 38910 82750
rect 38980 82550 39020 82750
rect 39090 82550 39100 82750
rect 38900 82520 39100 82550
rect 39400 82750 39600 82780
rect 39400 82550 39410 82750
rect 39480 82550 39520 82750
rect 39590 82550 39600 82750
rect 39400 82520 39600 82550
rect 39900 82750 40100 82780
rect 39900 82550 39910 82750
rect 39980 82550 40020 82750
rect 40090 82550 40100 82750
rect 39900 82520 40100 82550
rect 40400 82750 40600 82780
rect 40400 82550 40410 82750
rect 40480 82550 40520 82750
rect 40590 82550 40600 82750
rect 40400 82520 40600 82550
rect 40900 82750 41100 82780
rect 40900 82550 40910 82750
rect 40980 82550 41020 82750
rect 41090 82550 41100 82750
rect 40900 82520 41100 82550
rect 41400 82750 41600 82780
rect 41400 82550 41410 82750
rect 41480 82550 41520 82750
rect 41590 82550 41600 82750
rect 41400 82520 41600 82550
rect 41900 82750 42100 82780
rect 41900 82550 41910 82750
rect 41980 82550 42020 82750
rect 42090 82550 42100 82750
rect 41900 82520 42100 82550
rect 42400 82750 42600 82780
rect 42400 82550 42410 82750
rect 42480 82550 42520 82750
rect 42590 82550 42600 82750
rect 42400 82520 42600 82550
rect 42900 82750 43100 82780
rect 42900 82550 42910 82750
rect 42980 82550 43020 82750
rect 43090 82550 43100 82750
rect 42900 82520 43100 82550
rect 43400 82750 43600 82780
rect 43400 82550 43410 82750
rect 43480 82550 43520 82750
rect 43590 82550 43600 82750
rect 43400 82520 43600 82550
rect 43900 82750 44100 82780
rect 43900 82550 43910 82750
rect 43980 82550 44020 82750
rect 44090 82550 44100 82750
rect 43900 82520 44100 82550
rect 44400 82750 44600 82780
rect 44400 82550 44410 82750
rect 44480 82550 44520 82750
rect 44590 82550 44600 82750
rect 44400 82520 44600 82550
rect 44900 82750 45100 82780
rect 44900 82550 44910 82750
rect 44980 82550 45020 82750
rect 45090 82550 45100 82750
rect 44900 82520 45100 82550
rect 45400 82750 45600 82780
rect 45400 82550 45410 82750
rect 45480 82550 45520 82750
rect 45590 82550 45600 82750
rect 45400 82520 45600 82550
rect 45900 82750 46100 82780
rect 45900 82550 45910 82750
rect 45980 82550 46020 82750
rect 46090 82550 46100 82750
rect 45900 82520 46100 82550
rect 46400 82750 46600 82780
rect 46400 82550 46410 82750
rect 46480 82550 46520 82750
rect 46590 82550 46600 82750
rect 46400 82520 46600 82550
rect 46900 82750 47100 82780
rect 46900 82550 46910 82750
rect 46980 82550 47020 82750
rect 47090 82550 47100 82750
rect 46900 82520 47100 82550
rect 47400 82750 47600 82780
rect 47400 82550 47410 82750
rect 47480 82550 47520 82750
rect 47590 82550 47600 82750
rect 47400 82520 47600 82550
rect 47900 82750 48100 82780
rect 47900 82550 47910 82750
rect 47980 82550 48020 82750
rect 48090 82550 48100 82750
rect 47900 82520 48100 82550
rect 48400 82750 48600 82780
rect 48400 82550 48410 82750
rect 48480 82550 48520 82750
rect 48590 82550 48600 82750
rect 48400 82520 48600 82550
rect 48900 82750 49100 82780
rect 48900 82550 48910 82750
rect 48980 82550 49020 82750
rect 49090 82550 49100 82750
rect 48900 82520 49100 82550
rect 49400 82750 49600 82780
rect 49400 82550 49410 82750
rect 49480 82550 49520 82750
rect 49590 82550 49600 82750
rect 49400 82520 49600 82550
rect 49900 82750 50100 82780
rect 49900 82550 49910 82750
rect 49980 82550 50020 82750
rect 50090 82550 50100 82750
rect 49900 82520 50100 82550
rect 50400 82750 50600 82780
rect 50400 82550 50410 82750
rect 50480 82550 50520 82750
rect 50590 82550 50600 82750
rect 50400 82520 50600 82550
rect 50900 82750 51100 82780
rect 50900 82550 50910 82750
rect 50980 82550 51020 82750
rect 51090 82550 51100 82750
rect 50900 82520 51100 82550
rect 51400 82750 51600 82780
rect 51400 82550 51410 82750
rect 51480 82550 51520 82750
rect 51590 82550 51600 82750
rect 51400 82520 51600 82550
rect 51900 82750 52100 82780
rect 51900 82550 51910 82750
rect 51980 82550 52020 82750
rect 52090 82550 52100 82750
rect 51900 82520 52100 82550
rect 52400 82750 52600 82780
rect 52400 82550 52410 82750
rect 52480 82550 52520 82750
rect 52590 82550 52600 82750
rect 52400 82520 52600 82550
rect 52900 82750 53100 82780
rect 52900 82550 52910 82750
rect 52980 82550 53020 82750
rect 53090 82550 53100 82750
rect 52900 82520 53100 82550
rect 53400 82750 53600 82780
rect 53400 82550 53410 82750
rect 53480 82550 53520 82750
rect 53590 82550 53600 82750
rect 53400 82520 53600 82550
rect 53900 82750 54100 82780
rect 53900 82550 53910 82750
rect 53980 82550 54020 82750
rect 54090 82550 54100 82750
rect 53900 82520 54100 82550
rect 54400 82750 54600 82780
rect 54400 82550 54410 82750
rect 54480 82550 54520 82750
rect 54590 82550 54600 82750
rect 54400 82520 54600 82550
rect 54900 82750 55100 82780
rect 54900 82550 54910 82750
rect 54980 82550 55020 82750
rect 55090 82550 55100 82750
rect 54900 82520 55100 82550
rect 55400 82750 55600 82780
rect 55400 82550 55410 82750
rect 55480 82550 55520 82750
rect 55590 82550 55600 82750
rect 55400 82520 55600 82550
rect 55900 82750 56100 82780
rect 55900 82550 55910 82750
rect 55980 82550 56020 82750
rect 56090 82550 56100 82750
rect 55900 82520 56100 82550
rect 56400 82750 56600 82780
rect 56400 82550 56410 82750
rect 56480 82550 56520 82750
rect 56590 82550 56600 82750
rect 56400 82520 56600 82550
rect 56900 82750 57100 82780
rect 56900 82550 56910 82750
rect 56980 82550 57020 82750
rect 57090 82550 57100 82750
rect 56900 82520 57100 82550
rect 57400 82750 57600 82780
rect 57400 82550 57410 82750
rect 57480 82550 57520 82750
rect 57590 82550 57600 82750
rect 57400 82520 57600 82550
rect 57900 82750 58100 82780
rect 57900 82550 57910 82750
rect 57980 82550 58020 82750
rect 58090 82550 58100 82750
rect 57900 82520 58100 82550
rect 58400 82750 58600 82780
rect 58400 82550 58410 82750
rect 58480 82550 58520 82750
rect 58590 82550 58600 82750
rect 58400 82520 58600 82550
rect 58900 82750 59100 82780
rect 58900 82550 58910 82750
rect 58980 82550 59020 82750
rect 59090 82550 59100 82750
rect 58900 82520 59100 82550
rect 59400 82750 59600 82780
rect 59400 82550 59410 82750
rect 59480 82550 59520 82750
rect 59590 82550 59600 82750
rect 59400 82520 59600 82550
rect 59900 82750 60100 82780
rect 59900 82550 59910 82750
rect 59980 82550 60020 82750
rect 60090 82550 60100 82750
rect 59900 82520 60100 82550
rect 60400 82750 60600 82780
rect 60400 82550 60410 82750
rect 60480 82550 60520 82750
rect 60590 82550 60600 82750
rect 60400 82520 60600 82550
rect 60900 82750 61100 82780
rect 60900 82550 60910 82750
rect 60980 82550 61020 82750
rect 61090 82550 61100 82750
rect 60900 82520 61100 82550
rect 61400 82750 61600 82780
rect 61400 82550 61410 82750
rect 61480 82550 61520 82750
rect 61590 82550 61600 82750
rect 61400 82520 61600 82550
rect 61900 82750 62100 82780
rect 61900 82550 61910 82750
rect 61980 82550 62020 82750
rect 62090 82550 62100 82750
rect 61900 82520 62100 82550
rect 62400 82750 62600 82780
rect 62400 82550 62410 82750
rect 62480 82550 62520 82750
rect 62590 82550 62600 82750
rect 62400 82520 62600 82550
rect 62900 82750 63100 82780
rect 62900 82550 62910 82750
rect 62980 82550 63020 82750
rect 63090 82550 63100 82750
rect 62900 82520 63100 82550
rect 63400 82750 63600 82780
rect 63400 82550 63410 82750
rect 63480 82550 63520 82750
rect 63590 82550 63600 82750
rect 63400 82520 63600 82550
rect 63900 82750 64100 82780
rect 63900 82550 63910 82750
rect 63980 82550 64020 82750
rect 64090 82550 64100 82750
rect 63900 82520 64100 82550
rect 64400 82750 64600 82780
rect 64400 82550 64410 82750
rect 64480 82550 64520 82750
rect 64590 82550 64600 82750
rect 64400 82520 64600 82550
rect 64900 82750 65100 82780
rect 64900 82550 64910 82750
rect 64980 82550 65020 82750
rect 65090 82550 65100 82750
rect 64900 82520 65100 82550
rect 65400 82750 65600 82780
rect 65400 82550 65410 82750
rect 65480 82550 65520 82750
rect 65590 82550 65600 82750
rect 65400 82520 65600 82550
rect 65900 82750 66100 82780
rect 65900 82550 65910 82750
rect 65980 82550 66020 82750
rect 66090 82550 66100 82750
rect 65900 82520 66100 82550
rect 66400 82750 66600 82780
rect 66400 82550 66410 82750
rect 66480 82550 66520 82750
rect 66590 82550 66600 82750
rect 66400 82520 66600 82550
rect 66900 82750 67100 82780
rect 66900 82550 66910 82750
rect 66980 82550 67020 82750
rect 67090 82550 67100 82750
rect 66900 82520 67100 82550
rect 67400 82750 67600 82780
rect 67400 82550 67410 82750
rect 67480 82550 67520 82750
rect 67590 82550 67600 82750
rect 67400 82520 67600 82550
rect 67900 82750 68100 82780
rect 67900 82550 67910 82750
rect 67980 82550 68020 82750
rect 68090 82550 68100 82750
rect 67900 82520 68100 82550
rect 68400 82750 68600 82780
rect 68400 82550 68410 82750
rect 68480 82550 68520 82750
rect 68590 82550 68600 82750
rect 68400 82520 68600 82550
rect 68900 82750 69100 82780
rect 68900 82550 68910 82750
rect 68980 82550 69020 82750
rect 69090 82550 69100 82750
rect 68900 82520 69100 82550
rect 69400 82750 69600 82780
rect 69400 82550 69410 82750
rect 69480 82550 69520 82750
rect 69590 82550 69600 82750
rect 69400 82520 69600 82550
rect 69900 82750 70100 82780
rect 69900 82550 69910 82750
rect 69980 82550 70020 82750
rect 70090 82550 70100 82750
rect 69900 82520 70100 82550
rect 70400 82750 70600 82780
rect 70400 82550 70410 82750
rect 70480 82550 70520 82750
rect 70590 82550 70600 82750
rect 70400 82520 70600 82550
rect 70900 82750 71100 82780
rect 70900 82550 70910 82750
rect 70980 82550 71020 82750
rect 71090 82550 71100 82750
rect 70900 82520 71100 82550
rect 71400 82750 71600 82780
rect 71400 82550 71410 82750
rect 71480 82550 71520 82750
rect 71590 82550 71600 82750
rect 71400 82520 71600 82550
rect 71900 82750 72100 82780
rect 71900 82550 71910 82750
rect 71980 82550 72020 82750
rect 72090 82550 72100 82750
rect 71900 82520 72100 82550
rect 72400 82750 72600 82780
rect 72400 82550 72410 82750
rect 72480 82550 72520 82750
rect 72590 82550 72600 82750
rect 72400 82520 72600 82550
rect 72900 82750 73100 82780
rect 72900 82550 72910 82750
rect 72980 82550 73020 82750
rect 73090 82550 73100 82750
rect 72900 82520 73100 82550
rect 73400 82750 73600 82780
rect 73400 82550 73410 82750
rect 73480 82550 73520 82750
rect 73590 82550 73600 82750
rect 73400 82520 73600 82550
rect 73900 82750 74100 82780
rect 73900 82550 73910 82750
rect 73980 82550 74020 82750
rect 74090 82550 74100 82750
rect 73900 82520 74100 82550
rect 74400 82750 74600 82780
rect 74400 82550 74410 82750
rect 74480 82550 74520 82750
rect 74590 82550 74600 82750
rect 74400 82520 74600 82550
rect 74900 82750 75100 82780
rect 74900 82550 74910 82750
rect 74980 82550 75020 82750
rect 75090 82550 75100 82750
rect 74900 82520 75100 82550
rect 75400 82750 75600 82780
rect 75400 82550 75410 82750
rect 75480 82550 75520 82750
rect 75590 82550 75600 82750
rect 75400 82520 75600 82550
rect 75900 82750 76100 82780
rect 75900 82550 75910 82750
rect 75980 82550 76020 82750
rect 76090 82550 76100 82750
rect 75900 82520 76100 82550
rect 76400 82750 76600 82780
rect 76400 82550 76410 82750
rect 76480 82550 76520 82750
rect 76590 82550 76600 82750
rect 76400 82520 76600 82550
rect 76900 82750 77100 82780
rect 76900 82550 76910 82750
rect 76980 82550 77020 82750
rect 77090 82550 77100 82750
rect 76900 82520 77100 82550
rect 77400 82750 77600 82780
rect 77400 82550 77410 82750
rect 77480 82550 77520 82750
rect 77590 82550 77600 82750
rect 77400 82520 77600 82550
rect 77900 82750 78100 82780
rect 77900 82550 77910 82750
rect 77980 82550 78020 82750
rect 78090 82550 78100 82750
rect 77900 82520 78100 82550
rect 78400 82750 78600 82780
rect 78400 82550 78410 82750
rect 78480 82550 78520 82750
rect 78590 82550 78600 82750
rect 78400 82520 78600 82550
rect 78900 82750 79100 82780
rect 78900 82550 78910 82750
rect 78980 82550 79020 82750
rect 79090 82550 79100 82750
rect 78900 82520 79100 82550
rect 79400 82750 79600 82780
rect 79400 82550 79410 82750
rect 79480 82550 79520 82750
rect 79590 82550 79600 82750
rect 79400 82520 79600 82550
rect 79900 82750 80100 82780
rect 79900 82550 79910 82750
rect 79980 82550 80020 82750
rect 80090 82550 80100 82750
rect 79900 82520 80100 82550
rect 80400 82750 80600 82780
rect 80400 82550 80410 82750
rect 80480 82550 80520 82750
rect 80590 82550 80600 82750
rect 80400 82520 80600 82550
rect 80900 82750 81100 82780
rect 80900 82550 80910 82750
rect 80980 82550 81020 82750
rect 81090 82550 81100 82750
rect 80900 82520 81100 82550
rect 81400 82750 81600 82780
rect 81400 82550 81410 82750
rect 81480 82550 81520 82750
rect 81590 82550 81600 82750
rect 81400 82520 81600 82550
rect 81900 82750 82100 82780
rect 81900 82550 81910 82750
rect 81980 82550 82020 82750
rect 82090 82550 82100 82750
rect 81900 82520 82100 82550
rect 82400 82750 82600 82780
rect 82400 82550 82410 82750
rect 82480 82550 82520 82750
rect 82590 82550 82600 82750
rect 82400 82520 82600 82550
rect 82900 82750 83100 82780
rect 82900 82550 82910 82750
rect 82980 82550 83020 82750
rect 83090 82550 83100 82750
rect 82900 82520 83100 82550
rect 83400 82750 83600 82780
rect 83400 82550 83410 82750
rect 83480 82550 83520 82750
rect 83590 82550 83600 82750
rect 83400 82520 83600 82550
rect 83900 82750 84100 82780
rect 83900 82550 83910 82750
rect 83980 82550 84020 82750
rect 84090 82550 84100 82750
rect 83900 82520 84100 82550
rect 84400 82750 84600 82780
rect 84400 82550 84410 82750
rect 84480 82550 84520 82750
rect 84590 82550 84600 82750
rect 84400 82520 84600 82550
rect 84900 82750 85100 82780
rect 84900 82550 84910 82750
rect 84980 82550 85020 82750
rect 85090 82550 85100 82750
rect 84900 82520 85100 82550
rect 85400 82750 85600 82780
rect 85400 82550 85410 82750
rect 85480 82550 85520 82750
rect 85590 82550 85600 82750
rect 85400 82520 85600 82550
rect 85900 82750 86100 82780
rect 85900 82550 85910 82750
rect 85980 82550 86020 82750
rect 86090 82550 86100 82750
rect 85900 82520 86100 82550
rect 86400 82750 86600 82780
rect 86400 82550 86410 82750
rect 86480 82550 86520 82750
rect 86590 82550 86600 82750
rect 86400 82520 86600 82550
rect 86900 82750 87100 82780
rect 86900 82550 86910 82750
rect 86980 82550 87020 82750
rect 87090 82550 87100 82750
rect 86900 82520 87100 82550
rect 87400 82750 87600 82780
rect 87400 82550 87410 82750
rect 87480 82550 87520 82750
rect 87590 82550 87600 82750
rect 87400 82520 87600 82550
rect 87900 82750 88100 82780
rect 87900 82550 87910 82750
rect 87980 82550 88020 82750
rect 88090 82550 88100 82750
rect 87900 82520 88100 82550
rect 88400 82750 88600 82780
rect 88400 82550 88410 82750
rect 88480 82550 88520 82750
rect 88590 82550 88600 82750
rect 88400 82520 88600 82550
rect 88900 82750 89100 82780
rect 88900 82550 88910 82750
rect 88980 82550 89020 82750
rect 89090 82550 89100 82750
rect 88900 82520 89100 82550
rect 89400 82750 89600 82780
rect 89400 82550 89410 82750
rect 89480 82550 89520 82750
rect 89590 82550 89600 82750
rect 89400 82520 89600 82550
rect 89900 82750 90100 82780
rect 89900 82550 89910 82750
rect 89980 82550 90020 82750
rect 90090 82550 90100 82750
rect 89900 82520 90100 82550
rect 90400 82750 90600 82780
rect 90400 82550 90410 82750
rect 90480 82550 90520 82750
rect 90590 82550 90600 82750
rect 90400 82520 90600 82550
rect 90900 82750 91100 82780
rect 90900 82550 90910 82750
rect 90980 82550 91020 82750
rect 91090 82550 91100 82750
rect 90900 82520 91100 82550
rect 91400 82750 91600 82780
rect 91400 82550 91410 82750
rect 91480 82550 91520 82750
rect 91590 82550 91600 82750
rect 91400 82520 91600 82550
rect 91900 82750 92100 82780
rect 91900 82550 91910 82750
rect 91980 82550 92020 82750
rect 92090 82550 92100 82750
rect 91900 82520 92100 82550
rect 92400 82750 92600 82780
rect 92400 82550 92410 82750
rect 92480 82550 92520 82750
rect 92590 82550 92600 82750
rect 92400 82520 92600 82550
rect 92900 82750 93100 82780
rect 92900 82550 92910 82750
rect 92980 82550 93020 82750
rect 93090 82550 93100 82750
rect 92900 82520 93100 82550
rect 93400 82750 93600 82780
rect 93400 82550 93410 82750
rect 93480 82550 93520 82750
rect 93590 82550 93600 82750
rect 93400 82520 93600 82550
rect 93900 82750 94100 82780
rect 93900 82550 93910 82750
rect 93980 82550 94020 82750
rect 94090 82550 94100 82750
rect 93900 82520 94100 82550
rect 94400 82750 94600 82780
rect 94400 82550 94410 82750
rect 94480 82550 94520 82750
rect 94590 82550 94600 82750
rect 94400 82520 94600 82550
rect 94900 82750 95100 82780
rect 94900 82550 94910 82750
rect 94980 82550 95020 82750
rect 95090 82550 95100 82750
rect 94900 82520 95100 82550
rect 95400 82750 95600 82780
rect 95400 82550 95410 82750
rect 95480 82550 95520 82750
rect 95590 82550 95600 82750
rect 95400 82520 95600 82550
rect 95900 82750 96100 82780
rect 95900 82550 95910 82750
rect 95980 82550 96020 82750
rect 96090 82550 96100 82750
rect 95900 82520 96100 82550
rect 96400 82750 96600 82780
rect 96400 82550 96410 82750
rect 96480 82550 96520 82750
rect 96590 82550 96600 82750
rect 96400 82520 96600 82550
rect 96900 82750 97100 82780
rect 96900 82550 96910 82750
rect 96980 82550 97020 82750
rect 97090 82550 97100 82750
rect 96900 82520 97100 82550
rect 97400 82750 97600 82780
rect 97400 82550 97410 82750
rect 97480 82550 97520 82750
rect 97590 82550 97600 82750
rect 97400 82520 97600 82550
rect 97900 82750 98100 82780
rect 97900 82550 97910 82750
rect 97980 82550 98020 82750
rect 98090 82550 98100 82750
rect 97900 82520 98100 82550
rect 98400 82750 98600 82780
rect 98400 82550 98410 82750
rect 98480 82550 98520 82750
rect 98590 82550 98600 82750
rect 98400 82520 98600 82550
rect 98900 82750 99100 82780
rect 98900 82550 98910 82750
rect 98980 82550 99020 82750
rect 99090 82550 99100 82750
rect 98900 82520 99100 82550
rect 99400 82750 99600 82780
rect 99400 82550 99410 82750
rect 99480 82550 99520 82750
rect 99590 82550 99600 82750
rect 99400 82520 99600 82550
rect 99900 82750 100100 82780
rect 99900 82550 99910 82750
rect 99980 82550 100020 82750
rect 100090 82550 100100 82750
rect 99900 82520 100100 82550
rect 100400 82750 100500 82780
rect 100400 82550 100410 82750
rect 100480 82550 100500 82750
rect 100400 82520 100500 82550
rect -83500 82500 -83380 82520
rect -83120 82500 -82880 82520
rect -82620 82500 -82380 82520
rect -82120 82500 -81880 82520
rect -81620 82500 -81380 82520
rect -81120 82500 -80880 82520
rect -80620 82500 -80380 82520
rect -80120 82500 -79880 82520
rect -79620 82500 -79380 82520
rect -79120 82500 -78880 82520
rect -78620 82500 -78380 82520
rect -78120 82500 -77880 82520
rect -77620 82500 -77380 82520
rect -77120 82500 -76880 82520
rect -76620 82500 -76380 82520
rect -76120 82500 -75880 82520
rect -75620 82500 -75380 82520
rect -75120 82500 -74880 82520
rect -74620 82500 -74380 82520
rect -74120 82500 -73880 82520
rect -73620 82500 -73380 82520
rect -73120 82500 -72880 82520
rect -72620 82500 -72380 82520
rect -72120 82500 -71880 82520
rect -71620 82500 -71380 82520
rect -71120 82500 -70880 82520
rect -70620 82500 -70380 82520
rect -70120 82500 -69880 82520
rect -69620 82500 -69380 82520
rect -69120 82500 -68880 82520
rect -68620 82500 -68380 82520
rect -68120 82500 -67880 82520
rect -67620 82500 -67380 82520
rect -67120 82500 -66880 82520
rect -66620 82500 -66380 82520
rect -66120 82500 -65880 82520
rect -65620 82500 -65380 82520
rect -65120 82500 -64880 82520
rect -64620 82500 -64380 82520
rect -64120 82500 -63880 82520
rect -63620 82500 -63380 82520
rect -63120 82500 -62880 82520
rect -62620 82500 -62380 82520
rect -62120 82500 -61880 82520
rect -61620 82500 -61380 82520
rect -61120 82500 -60880 82520
rect -60620 82500 -60380 82520
rect -60120 82500 -59880 82520
rect -59620 82500 -59380 82520
rect -59120 82500 -58880 82520
rect -58620 82500 -58380 82520
rect -58120 82500 -57880 82520
rect -57620 82500 -57380 82520
rect -57120 82500 -56880 82520
rect -56620 82500 -56380 82520
rect -56120 82500 -55880 82520
rect -55620 82500 -55380 82520
rect -55120 82500 -54880 82520
rect -54620 82500 -54380 82520
rect -54120 82500 -53880 82520
rect -53620 82500 -53380 82520
rect -53120 82500 -52880 82520
rect -52620 82500 -52380 82520
rect -52120 82500 -51880 82520
rect -51620 82500 -51380 82520
rect -51120 82500 -50880 82520
rect -50620 82500 -50380 82520
rect -50120 82500 -49880 82520
rect -49620 82500 -49380 82520
rect -49120 82500 -48880 82520
rect -48620 82500 -48380 82520
rect -48120 82500 -47880 82520
rect -47620 82500 -47380 82520
rect -47120 82500 -46880 82520
rect -46620 82500 -46380 82520
rect -46120 82500 -45880 82520
rect -45620 82500 -45380 82520
rect -45120 82500 -44880 82520
rect -44620 82500 -44380 82520
rect -44120 82500 -43880 82520
rect -43620 82500 -43380 82520
rect -43120 82500 -42880 82520
rect -42620 82500 -42380 82520
rect -42120 82500 -41880 82520
rect -41620 82500 -41380 82520
rect -41120 82500 -40880 82520
rect -40620 82500 -40380 82520
rect -40120 82500 -39880 82520
rect -39620 82500 -39380 82520
rect -39120 82500 -38880 82520
rect -38620 82500 -38380 82520
rect -38120 82500 -37880 82520
rect -37620 82500 -37380 82520
rect -37120 82500 -36880 82520
rect -36620 82500 -36380 82520
rect -36120 82500 -35880 82520
rect -35620 82500 -35380 82520
rect -35120 82500 -34880 82520
rect -34620 82500 -34380 82520
rect -34120 82500 -33880 82520
rect -33620 82500 -33380 82520
rect -33120 82500 -32880 82520
rect -32620 82500 -32380 82520
rect -32120 82500 -31880 82520
rect -31620 82500 -31380 82520
rect -31120 82500 -30880 82520
rect -30620 82500 -30380 82520
rect -30120 82500 -29880 82520
rect -29620 82500 -29380 82520
rect -29120 82500 -28880 82520
rect -28620 82500 -28380 82520
rect -28120 82500 -27880 82520
rect -27620 82500 -27380 82520
rect -27120 82500 -26880 82520
rect -26620 82500 -26380 82520
rect -26120 82500 -25880 82520
rect -25620 82500 -25380 82520
rect -25120 82500 -24880 82520
rect -24620 82500 -24380 82520
rect -24120 82500 -23880 82520
rect -23620 82500 -23380 82520
rect -23120 82500 -22880 82520
rect -22620 82500 -22380 82520
rect -22120 82500 -21880 82520
rect -21620 82500 -21380 82520
rect -21120 82500 -20880 82520
rect -20620 82500 -20380 82520
rect -20120 82500 -19880 82520
rect -19620 82500 -19380 82520
rect -19120 82500 -18880 82520
rect -18620 82500 -18380 82520
rect -18120 82500 -17880 82520
rect -17620 82500 -17380 82520
rect -17120 82500 -16880 82520
rect -16620 82500 -16380 82520
rect -16120 82500 -15880 82520
rect -15620 82500 -15380 82520
rect -15120 82500 -14880 82520
rect -14620 82500 -14380 82520
rect -14120 82500 -13880 82520
rect -13620 82500 -13380 82520
rect -13120 82500 -12880 82520
rect -12620 82500 -12380 82520
rect -12120 82500 -11880 82520
rect -11620 82500 -11380 82520
rect -11120 82500 -10880 82520
rect -10620 82500 -10380 82520
rect -10120 82500 -9880 82520
rect -9620 82500 -9380 82520
rect -9120 82500 -8880 82520
rect -8620 82500 -8380 82520
rect -8120 82500 -7880 82520
rect -7620 82500 -7380 82520
rect -7120 82500 -6880 82520
rect -6620 82500 -6380 82520
rect -6120 82500 -5880 82520
rect -5620 82500 -5380 82520
rect -5120 82500 -4880 82520
rect -4620 82500 -4380 82520
rect -4120 82500 -3880 82520
rect -3620 82500 -3380 82520
rect -3120 82500 -2880 82520
rect -2620 82500 -2380 82520
rect -2120 82500 -1880 82520
rect -1620 82500 -1380 82520
rect -1120 82500 -880 82520
rect -620 82500 -380 82520
rect -120 82500 120 82520
rect 380 82500 620 82520
rect 880 82500 1120 82520
rect 1380 82500 1620 82520
rect 1880 82500 2120 82520
rect 2380 82500 2620 82520
rect 2880 82500 3120 82520
rect 3380 82500 3620 82520
rect 3880 82500 4120 82520
rect 4380 82500 4620 82520
rect 4880 82500 5120 82520
rect 5380 82500 5620 82520
rect 5880 82500 6120 82520
rect 6380 82500 6620 82520
rect 6880 82500 7120 82520
rect 7380 82500 7620 82520
rect 7880 82500 8120 82520
rect 8380 82500 8620 82520
rect 8880 82500 9120 82520
rect 9380 82500 9620 82520
rect 9880 82500 10120 82520
rect 10380 82500 10620 82520
rect 10880 82500 11120 82520
rect 11380 82500 11620 82520
rect 11880 82500 12120 82520
rect 12380 82500 12620 82520
rect 12880 82500 13120 82520
rect 13380 82500 13620 82520
rect 13880 82500 14120 82520
rect 14380 82500 14620 82520
rect 14880 82500 15120 82520
rect 15380 82500 15620 82520
rect 15880 82500 16120 82520
rect 16380 82500 16620 82520
rect 16880 82500 17120 82520
rect 17380 82500 17620 82520
rect 17880 82500 18120 82520
rect 18380 82500 18620 82520
rect 18880 82500 19120 82520
rect 19380 82500 19620 82520
rect 19880 82500 20120 82520
rect 20380 82500 20620 82520
rect 20880 82500 21120 82520
rect 21380 82500 21620 82520
rect 21880 82500 22120 82520
rect 22380 82500 22620 82520
rect 22880 82500 23120 82520
rect 23380 82500 23620 82520
rect 23880 82500 24120 82520
rect 24380 82500 24620 82520
rect 24880 82500 25120 82520
rect 25380 82500 25620 82520
rect 25880 82500 26120 82520
rect 26380 82500 26620 82520
rect 26880 82500 27120 82520
rect 27380 82500 27620 82520
rect 27880 82500 28120 82520
rect 28380 82500 28620 82520
rect 28880 82500 29120 82520
rect 29380 82500 29620 82520
rect 29880 82500 30120 82520
rect 30380 82500 30620 82520
rect 30880 82500 31120 82520
rect 31380 82500 31620 82520
rect 31880 82500 32120 82520
rect 32380 82500 32620 82520
rect 32880 82500 33120 82520
rect 33380 82500 33620 82520
rect 33880 82500 34120 82520
rect 34380 82500 34620 82520
rect 34880 82500 35120 82520
rect 35380 82500 35620 82520
rect 35880 82500 36120 82520
rect 36380 82500 36620 82520
rect 36880 82500 37120 82520
rect 37380 82500 37620 82520
rect 37880 82500 38120 82520
rect 38380 82500 38620 82520
rect 38880 82500 39120 82520
rect 39380 82500 39620 82520
rect 39880 82500 40120 82520
rect 40380 82500 40620 82520
rect 40880 82500 41120 82520
rect 41380 82500 41620 82520
rect 41880 82500 42120 82520
rect 42380 82500 42620 82520
rect 42880 82500 43120 82520
rect 43380 82500 43620 82520
rect 43880 82500 44120 82520
rect 44380 82500 44620 82520
rect 44880 82500 45120 82520
rect 45380 82500 45620 82520
rect 45880 82500 46120 82520
rect 46380 82500 46620 82520
rect 46880 82500 47120 82520
rect 47380 82500 47620 82520
rect 47880 82500 48120 82520
rect 48380 82500 48620 82520
rect 48880 82500 49120 82520
rect 49380 82500 49620 82520
rect 49880 82500 50120 82520
rect 50380 82500 50620 82520
rect 50880 82500 51120 82520
rect 51380 82500 51620 82520
rect 51880 82500 52120 82520
rect 52380 82500 52620 82520
rect 52880 82500 53120 82520
rect 53380 82500 53620 82520
rect 53880 82500 54120 82520
rect 54380 82500 54620 82520
rect 54880 82500 55120 82520
rect 55380 82500 55620 82520
rect 55880 82500 56120 82520
rect 56380 82500 56620 82520
rect 56880 82500 57120 82520
rect 57380 82500 57620 82520
rect 57880 82500 58120 82520
rect 58380 82500 58620 82520
rect 58880 82500 59120 82520
rect 59380 82500 59620 82520
rect 59880 82500 60120 82520
rect 60380 82500 60620 82520
rect 60880 82500 61120 82520
rect 61380 82500 61620 82520
rect 61880 82500 62120 82520
rect 62380 82500 62620 82520
rect 62880 82500 63120 82520
rect 63380 82500 63620 82520
rect 63880 82500 64120 82520
rect 64380 82500 64620 82520
rect 64880 82500 65120 82520
rect 65380 82500 65620 82520
rect 65880 82500 66120 82520
rect 66380 82500 66620 82520
rect 66880 82500 67120 82520
rect 67380 82500 67620 82520
rect 67880 82500 68120 82520
rect 68380 82500 68620 82520
rect 68880 82500 69120 82520
rect 69380 82500 69620 82520
rect 69880 82500 70120 82520
rect 70380 82500 70620 82520
rect 70880 82500 71120 82520
rect 71380 82500 71620 82520
rect 71880 82500 72120 82520
rect 72380 82500 72620 82520
rect 72880 82500 73120 82520
rect 73380 82500 73620 82520
rect 73880 82500 74120 82520
rect 74380 82500 74620 82520
rect 74880 82500 75120 82520
rect 75380 82500 75620 82520
rect 75880 82500 76120 82520
rect 76380 82500 76620 82520
rect 76880 82500 77120 82520
rect 77380 82500 77620 82520
rect 77880 82500 78120 82520
rect 78380 82500 78620 82520
rect 78880 82500 79120 82520
rect 79380 82500 79620 82520
rect 79880 82500 80120 82520
rect 80380 82500 80620 82520
rect 80880 82500 81120 82520
rect 81380 82500 81620 82520
rect 81880 82500 82120 82520
rect 82380 82500 82620 82520
rect 82880 82500 83120 82520
rect 83380 82500 83620 82520
rect 83880 82500 84120 82520
rect 84380 82500 84620 82520
rect 84880 82500 85120 82520
rect 85380 82500 85620 82520
rect 85880 82500 86120 82520
rect 86380 82500 86620 82520
rect 86880 82500 87120 82520
rect 87380 82500 87620 82520
rect 87880 82500 88120 82520
rect 88380 82500 88620 82520
rect 88880 82500 89120 82520
rect 89380 82500 89620 82520
rect 89880 82500 90120 82520
rect 90380 82500 90620 82520
rect 90880 82500 91120 82520
rect 91380 82500 91620 82520
rect 91880 82500 92120 82520
rect 92380 82500 92620 82520
rect 92880 82500 93120 82520
rect 93380 82500 93620 82520
rect 93880 82500 94120 82520
rect 94380 82500 94620 82520
rect 94880 82500 95120 82520
rect 95380 82500 95620 82520
rect 95880 82500 96120 82520
rect 96380 82500 96620 82520
rect 96880 82500 97120 82520
rect 97380 82500 97620 82520
rect 97880 82500 98120 82520
rect 98380 82500 98620 82520
rect 98880 82500 99120 82520
rect 99380 82500 99620 82520
rect 99880 82500 100120 82520
rect 100380 82500 100500 82520
rect -83500 82490 100500 82500
rect -83500 82420 -83350 82490
rect -83150 82420 -82850 82490
rect -82650 82420 -82350 82490
rect -82150 82420 -81850 82490
rect -81650 82420 -81350 82490
rect -81150 82420 -80850 82490
rect -80650 82420 -80350 82490
rect -80150 82420 -79850 82490
rect -79650 82420 -79350 82490
rect -79150 82420 -78850 82490
rect -78650 82420 -78350 82490
rect -78150 82420 -77850 82490
rect -77650 82420 -77350 82490
rect -77150 82420 -76850 82490
rect -76650 82420 -76350 82490
rect -76150 82420 -75850 82490
rect -75650 82420 -75350 82490
rect -75150 82420 -74850 82490
rect -74650 82420 -74350 82490
rect -74150 82420 -73850 82490
rect -73650 82420 -73350 82490
rect -73150 82420 -72850 82490
rect -72650 82420 -72350 82490
rect -72150 82420 -71850 82490
rect -71650 82420 -71350 82490
rect -71150 82420 -70850 82490
rect -70650 82420 -70350 82490
rect -70150 82420 -69850 82490
rect -69650 82420 -69350 82490
rect -69150 82420 -68850 82490
rect -68650 82420 -68350 82490
rect -68150 82420 -67850 82490
rect -67650 82420 -67350 82490
rect -67150 82420 -66850 82490
rect -66650 82420 -66350 82490
rect -66150 82420 -65850 82490
rect -65650 82420 -65350 82490
rect -65150 82420 -64850 82490
rect -64650 82420 -64350 82490
rect -64150 82420 -63850 82490
rect -63650 82420 -63350 82490
rect -63150 82420 -62850 82490
rect -62650 82420 -62350 82490
rect -62150 82420 -61850 82490
rect -61650 82420 -61350 82490
rect -61150 82420 -60850 82490
rect -60650 82420 -60350 82490
rect -60150 82420 -59850 82490
rect -59650 82420 -59350 82490
rect -59150 82420 -58850 82490
rect -58650 82420 -58350 82490
rect -58150 82420 -57850 82490
rect -57650 82420 -57350 82490
rect -57150 82420 -56850 82490
rect -56650 82420 -56350 82490
rect -56150 82420 -55850 82490
rect -55650 82420 -55350 82490
rect -55150 82420 -54850 82490
rect -54650 82420 -54350 82490
rect -54150 82420 -53850 82490
rect -53650 82420 -53350 82490
rect -53150 82420 -52850 82490
rect -52650 82420 -52350 82490
rect -52150 82420 -51850 82490
rect -51650 82420 -51350 82490
rect -51150 82420 -50850 82490
rect -50650 82420 -50350 82490
rect -50150 82420 -49850 82490
rect -49650 82420 -49350 82490
rect -49150 82420 -48850 82490
rect -48650 82420 -48350 82490
rect -48150 82420 -47850 82490
rect -47650 82420 -47350 82490
rect -47150 82420 -46850 82490
rect -46650 82420 -46350 82490
rect -46150 82420 -45850 82490
rect -45650 82420 -45350 82490
rect -45150 82420 -44850 82490
rect -44650 82420 -44350 82490
rect -44150 82420 -43850 82490
rect -43650 82420 -43350 82490
rect -43150 82420 -42850 82490
rect -42650 82420 -42350 82490
rect -42150 82420 -41850 82490
rect -41650 82420 -41350 82490
rect -41150 82420 -40850 82490
rect -40650 82420 -40350 82490
rect -40150 82420 -39850 82490
rect -39650 82420 -39350 82490
rect -39150 82420 -38850 82490
rect -38650 82420 -38350 82490
rect -38150 82420 -37850 82490
rect -37650 82420 -37350 82490
rect -37150 82420 -36850 82490
rect -36650 82420 -36350 82490
rect -36150 82420 -35850 82490
rect -35650 82420 -35350 82490
rect -35150 82420 -34850 82490
rect -34650 82420 -34350 82490
rect -34150 82420 -33850 82490
rect -33650 82420 -33350 82490
rect -33150 82420 -32850 82490
rect -32650 82420 -32350 82490
rect -32150 82420 -31850 82490
rect -31650 82420 -31350 82490
rect -31150 82420 -30850 82490
rect -30650 82420 -30350 82490
rect -30150 82420 -29850 82490
rect -29650 82420 -29350 82490
rect -29150 82420 -28850 82490
rect -28650 82420 -28350 82490
rect -28150 82420 -27850 82490
rect -27650 82420 -27350 82490
rect -27150 82420 -26850 82490
rect -26650 82420 -26350 82490
rect -26150 82420 -25850 82490
rect -25650 82420 -25350 82490
rect -25150 82420 -24850 82490
rect -24650 82420 -24350 82490
rect -24150 82420 -23850 82490
rect -23650 82420 -23350 82490
rect -23150 82420 -22850 82490
rect -22650 82420 -22350 82490
rect -22150 82420 -21850 82490
rect -21650 82420 -21350 82490
rect -21150 82420 -20850 82490
rect -20650 82420 -20350 82490
rect -20150 82420 -19850 82490
rect -19650 82420 -19350 82490
rect -19150 82420 -18850 82490
rect -18650 82420 -18350 82490
rect -18150 82420 -17850 82490
rect -17650 82420 -17350 82490
rect -17150 82420 -16850 82490
rect -16650 82420 -16350 82490
rect -16150 82420 -15850 82490
rect -15650 82420 -15350 82490
rect -15150 82420 -14850 82490
rect -14650 82420 -14350 82490
rect -14150 82420 -13850 82490
rect -13650 82420 -13350 82490
rect -13150 82420 -12850 82490
rect -12650 82420 -12350 82490
rect -12150 82420 -11850 82490
rect -11650 82420 -11350 82490
rect -11150 82420 -10850 82490
rect -10650 82420 -10350 82490
rect -10150 82420 -9850 82490
rect -9650 82420 -9350 82490
rect -9150 82420 -8850 82490
rect -8650 82420 -8350 82490
rect -8150 82420 -7850 82490
rect -7650 82420 -7350 82490
rect -7150 82420 -6850 82490
rect -6650 82420 -6350 82490
rect -6150 82420 -5850 82490
rect -5650 82420 -5350 82490
rect -5150 82420 -4850 82490
rect -4650 82420 -4350 82490
rect -4150 82420 -3850 82490
rect -3650 82420 -3350 82490
rect -3150 82420 -2850 82490
rect -2650 82420 -2350 82490
rect -2150 82420 -1850 82490
rect -1650 82420 -1350 82490
rect -1150 82420 -850 82490
rect -650 82420 -350 82490
rect -150 82420 150 82490
rect 350 82420 650 82490
rect 850 82420 1150 82490
rect 1350 82420 1650 82490
rect 1850 82420 2150 82490
rect 2350 82420 2650 82490
rect 2850 82420 3150 82490
rect 3350 82420 3650 82490
rect 3850 82420 4150 82490
rect 4350 82420 4650 82490
rect 4850 82420 5150 82490
rect 5350 82420 5650 82490
rect 5850 82420 6150 82490
rect 6350 82420 6650 82490
rect 6850 82420 7150 82490
rect 7350 82420 7650 82490
rect 7850 82420 8150 82490
rect 8350 82420 8650 82490
rect 8850 82420 9150 82490
rect 9350 82420 9650 82490
rect 9850 82420 10150 82490
rect 10350 82420 10650 82490
rect 10850 82420 11150 82490
rect 11350 82420 11650 82490
rect 11850 82420 12150 82490
rect 12350 82420 12650 82490
rect 12850 82420 13150 82490
rect 13350 82420 13650 82490
rect 13850 82420 14150 82490
rect 14350 82420 14650 82490
rect 14850 82420 15150 82490
rect 15350 82420 15650 82490
rect 15850 82420 16150 82490
rect 16350 82420 16650 82490
rect 16850 82420 17150 82490
rect 17350 82420 17650 82490
rect 17850 82420 18150 82490
rect 18350 82420 18650 82490
rect 18850 82420 19150 82490
rect 19350 82420 19650 82490
rect 19850 82420 20150 82490
rect 20350 82420 20650 82490
rect 20850 82420 21150 82490
rect 21350 82420 21650 82490
rect 21850 82420 22150 82490
rect 22350 82420 22650 82490
rect 22850 82420 23150 82490
rect 23350 82420 23650 82490
rect 23850 82420 24150 82490
rect 24350 82420 24650 82490
rect 24850 82420 25150 82490
rect 25350 82420 25650 82490
rect 25850 82420 26150 82490
rect 26350 82420 26650 82490
rect 26850 82420 27150 82490
rect 27350 82420 27650 82490
rect 27850 82420 28150 82490
rect 28350 82420 28650 82490
rect 28850 82420 29150 82490
rect 29350 82420 29650 82490
rect 29850 82420 30150 82490
rect 30350 82420 30650 82490
rect 30850 82420 31150 82490
rect 31350 82420 31650 82490
rect 31850 82420 32150 82490
rect 32350 82420 32650 82490
rect 32850 82420 33150 82490
rect 33350 82420 33650 82490
rect 33850 82420 34150 82490
rect 34350 82420 34650 82490
rect 34850 82420 35150 82490
rect 35350 82420 35650 82490
rect 35850 82420 36150 82490
rect 36350 82420 36650 82490
rect 36850 82420 37150 82490
rect 37350 82420 37650 82490
rect 37850 82420 38150 82490
rect 38350 82420 38650 82490
rect 38850 82420 39150 82490
rect 39350 82420 39650 82490
rect 39850 82420 40150 82490
rect 40350 82420 40650 82490
rect 40850 82420 41150 82490
rect 41350 82420 41650 82490
rect 41850 82420 42150 82490
rect 42350 82420 42650 82490
rect 42850 82420 43150 82490
rect 43350 82420 43650 82490
rect 43850 82420 44150 82490
rect 44350 82420 44650 82490
rect 44850 82420 45150 82490
rect 45350 82420 45650 82490
rect 45850 82420 46150 82490
rect 46350 82420 46650 82490
rect 46850 82420 47150 82490
rect 47350 82420 47650 82490
rect 47850 82420 48150 82490
rect 48350 82420 48650 82490
rect 48850 82420 49150 82490
rect 49350 82420 49650 82490
rect 49850 82420 50150 82490
rect 50350 82420 50650 82490
rect 50850 82420 51150 82490
rect 51350 82420 51650 82490
rect 51850 82420 52150 82490
rect 52350 82420 52650 82490
rect 52850 82420 53150 82490
rect 53350 82420 53650 82490
rect 53850 82420 54150 82490
rect 54350 82420 54650 82490
rect 54850 82420 55150 82490
rect 55350 82420 55650 82490
rect 55850 82420 56150 82490
rect 56350 82420 56650 82490
rect 56850 82420 57150 82490
rect 57350 82420 57650 82490
rect 57850 82420 58150 82490
rect 58350 82420 58650 82490
rect 58850 82420 59150 82490
rect 59350 82420 59650 82490
rect 59850 82420 60150 82490
rect 60350 82420 60650 82490
rect 60850 82420 61150 82490
rect 61350 82420 61650 82490
rect 61850 82420 62150 82490
rect 62350 82420 62650 82490
rect 62850 82420 63150 82490
rect 63350 82420 63650 82490
rect 63850 82420 64150 82490
rect 64350 82420 64650 82490
rect 64850 82420 65150 82490
rect 65350 82420 65650 82490
rect 65850 82420 66150 82490
rect 66350 82420 66650 82490
rect 66850 82420 67150 82490
rect 67350 82420 67650 82490
rect 67850 82420 68150 82490
rect 68350 82420 68650 82490
rect 68850 82420 69150 82490
rect 69350 82420 69650 82490
rect 69850 82420 70150 82490
rect 70350 82420 70650 82490
rect 70850 82420 71150 82490
rect 71350 82420 71650 82490
rect 71850 82420 72150 82490
rect 72350 82420 72650 82490
rect 72850 82420 73150 82490
rect 73350 82420 73650 82490
rect 73850 82420 74150 82490
rect 74350 82420 74650 82490
rect 74850 82420 75150 82490
rect 75350 82420 75650 82490
rect 75850 82420 76150 82490
rect 76350 82420 76650 82490
rect 76850 82420 77150 82490
rect 77350 82420 77650 82490
rect 77850 82420 78150 82490
rect 78350 82420 78650 82490
rect 78850 82420 79150 82490
rect 79350 82420 79650 82490
rect 79850 82420 80150 82490
rect 80350 82420 80650 82490
rect 80850 82420 81150 82490
rect 81350 82420 81650 82490
rect 81850 82420 82150 82490
rect 82350 82420 82650 82490
rect 82850 82420 83150 82490
rect 83350 82420 83650 82490
rect 83850 82420 84150 82490
rect 84350 82420 84650 82490
rect 84850 82420 85150 82490
rect 85350 82420 85650 82490
rect 85850 82420 86150 82490
rect 86350 82420 86650 82490
rect 86850 82420 87150 82490
rect 87350 82420 87650 82490
rect 87850 82420 88150 82490
rect 88350 82420 88650 82490
rect 88850 82420 89150 82490
rect 89350 82420 89650 82490
rect 89850 82420 90150 82490
rect 90350 82420 90650 82490
rect 90850 82420 91150 82490
rect 91350 82420 91650 82490
rect 91850 82420 92150 82490
rect 92350 82420 92650 82490
rect 92850 82420 93150 82490
rect 93350 82420 93650 82490
rect 93850 82420 94150 82490
rect 94350 82420 94650 82490
rect 94850 82420 95150 82490
rect 95350 82420 95650 82490
rect 95850 82420 96150 82490
rect 96350 82420 96650 82490
rect 96850 82420 97150 82490
rect 97350 82420 97650 82490
rect 97850 82420 98150 82490
rect 98350 82420 98650 82490
rect 98850 82420 99150 82490
rect 99350 82420 99650 82490
rect 99850 82420 100150 82490
rect 100350 82420 100500 82490
rect -83500 82380 100500 82420
rect -83500 82310 -83350 82380
rect -83150 82310 -82850 82380
rect -82650 82310 -82350 82380
rect -82150 82310 -81850 82380
rect -81650 82310 -81350 82380
rect -81150 82310 -80850 82380
rect -80650 82310 -80350 82380
rect -80150 82310 -79850 82380
rect -79650 82310 -79350 82380
rect -79150 82310 -78850 82380
rect -78650 82310 -78350 82380
rect -78150 82310 -77850 82380
rect -77650 82310 -77350 82380
rect -77150 82310 -76850 82380
rect -76650 82310 -76350 82380
rect -76150 82310 -75850 82380
rect -75650 82310 -75350 82380
rect -75150 82310 -74850 82380
rect -74650 82310 -74350 82380
rect -74150 82310 -73850 82380
rect -73650 82310 -73350 82380
rect -73150 82310 -72850 82380
rect -72650 82310 -72350 82380
rect -72150 82310 -71850 82380
rect -71650 82310 -71350 82380
rect -71150 82310 -70850 82380
rect -70650 82310 -70350 82380
rect -70150 82310 -69850 82380
rect -69650 82310 -69350 82380
rect -69150 82310 -68850 82380
rect -68650 82310 -68350 82380
rect -68150 82310 -67850 82380
rect -67650 82310 -67350 82380
rect -67150 82310 -66850 82380
rect -66650 82310 -66350 82380
rect -66150 82310 -65850 82380
rect -65650 82310 -65350 82380
rect -65150 82310 -64850 82380
rect -64650 82310 -64350 82380
rect -64150 82310 -63850 82380
rect -63650 82310 -63350 82380
rect -63150 82310 -62850 82380
rect -62650 82310 -62350 82380
rect -62150 82310 -61850 82380
rect -61650 82310 -61350 82380
rect -61150 82310 -60850 82380
rect -60650 82310 -60350 82380
rect -60150 82310 -59850 82380
rect -59650 82310 -59350 82380
rect -59150 82310 -58850 82380
rect -58650 82310 -58350 82380
rect -58150 82310 -57850 82380
rect -57650 82310 -57350 82380
rect -57150 82310 -56850 82380
rect -56650 82310 -56350 82380
rect -56150 82310 -55850 82380
rect -55650 82310 -55350 82380
rect -55150 82310 -54850 82380
rect -54650 82310 -54350 82380
rect -54150 82310 -53850 82380
rect -53650 82310 -53350 82380
rect -53150 82310 -52850 82380
rect -52650 82310 -52350 82380
rect -52150 82310 -51850 82380
rect -51650 82310 -51350 82380
rect -51150 82310 -50850 82380
rect -50650 82310 -50350 82380
rect -50150 82310 -49850 82380
rect -49650 82310 -49350 82380
rect -49150 82310 -48850 82380
rect -48650 82310 -48350 82380
rect -48150 82310 -47850 82380
rect -47650 82310 -47350 82380
rect -47150 82310 -46850 82380
rect -46650 82310 -46350 82380
rect -46150 82310 -45850 82380
rect -45650 82310 -45350 82380
rect -45150 82310 -44850 82380
rect -44650 82310 -44350 82380
rect -44150 82310 -43850 82380
rect -43650 82310 -43350 82380
rect -43150 82310 -42850 82380
rect -42650 82310 -42350 82380
rect -42150 82310 -41850 82380
rect -41650 82310 -41350 82380
rect -41150 82310 -40850 82380
rect -40650 82310 -40350 82380
rect -40150 82310 -39850 82380
rect -39650 82310 -39350 82380
rect -39150 82310 -38850 82380
rect -38650 82310 -38350 82380
rect -38150 82310 -37850 82380
rect -37650 82310 -37350 82380
rect -37150 82310 -36850 82380
rect -36650 82310 -36350 82380
rect -36150 82310 -35850 82380
rect -35650 82310 -35350 82380
rect -35150 82310 -34850 82380
rect -34650 82310 -34350 82380
rect -34150 82310 -33850 82380
rect -33650 82310 -33350 82380
rect -33150 82310 -32850 82380
rect -32650 82310 -32350 82380
rect -32150 82310 -31850 82380
rect -31650 82310 -31350 82380
rect -31150 82310 -30850 82380
rect -30650 82310 -30350 82380
rect -30150 82310 -29850 82380
rect -29650 82310 -29350 82380
rect -29150 82310 -28850 82380
rect -28650 82310 -28350 82380
rect -28150 82310 -27850 82380
rect -27650 82310 -27350 82380
rect -27150 82310 -26850 82380
rect -26650 82310 -26350 82380
rect -26150 82310 -25850 82380
rect -25650 82310 -25350 82380
rect -25150 82310 -24850 82380
rect -24650 82310 -24350 82380
rect -24150 82310 -23850 82380
rect -23650 82310 -23350 82380
rect -23150 82310 -22850 82380
rect -22650 82310 -22350 82380
rect -22150 82310 -21850 82380
rect -21650 82310 -21350 82380
rect -21150 82310 -20850 82380
rect -20650 82310 -20350 82380
rect -20150 82310 -19850 82380
rect -19650 82310 -19350 82380
rect -19150 82310 -18850 82380
rect -18650 82310 -18350 82380
rect -18150 82310 -17850 82380
rect -17650 82310 -17350 82380
rect -17150 82310 -16850 82380
rect -16650 82310 -16350 82380
rect -16150 82310 -15850 82380
rect -15650 82310 -15350 82380
rect -15150 82310 -14850 82380
rect -14650 82310 -14350 82380
rect -14150 82310 -13850 82380
rect -13650 82310 -13350 82380
rect -13150 82310 -12850 82380
rect -12650 82310 -12350 82380
rect -12150 82310 -11850 82380
rect -11650 82310 -11350 82380
rect -11150 82310 -10850 82380
rect -10650 82310 -10350 82380
rect -10150 82310 -9850 82380
rect -9650 82310 -9350 82380
rect -9150 82310 -8850 82380
rect -8650 82310 -8350 82380
rect -8150 82310 -7850 82380
rect -7650 82310 -7350 82380
rect -7150 82310 -6850 82380
rect -6650 82310 -6350 82380
rect -6150 82310 -5850 82380
rect -5650 82310 -5350 82380
rect -5150 82310 -4850 82380
rect -4650 82310 -4350 82380
rect -4150 82310 -3850 82380
rect -3650 82310 -3350 82380
rect -3150 82310 -2850 82380
rect -2650 82310 -2350 82380
rect -2150 82310 -1850 82380
rect -1650 82310 -1350 82380
rect -1150 82310 -850 82380
rect -650 82310 -350 82380
rect -150 82310 150 82380
rect 350 82310 650 82380
rect 850 82310 1150 82380
rect 1350 82310 1650 82380
rect 1850 82310 2150 82380
rect 2350 82310 2650 82380
rect 2850 82310 3150 82380
rect 3350 82310 3650 82380
rect 3850 82310 4150 82380
rect 4350 82310 4650 82380
rect 4850 82310 5150 82380
rect 5350 82310 5650 82380
rect 5850 82310 6150 82380
rect 6350 82310 6650 82380
rect 6850 82310 7150 82380
rect 7350 82310 7650 82380
rect 7850 82310 8150 82380
rect 8350 82310 8650 82380
rect 8850 82310 9150 82380
rect 9350 82310 9650 82380
rect 9850 82310 10150 82380
rect 10350 82310 10650 82380
rect 10850 82310 11150 82380
rect 11350 82310 11650 82380
rect 11850 82310 12150 82380
rect 12350 82310 12650 82380
rect 12850 82310 13150 82380
rect 13350 82310 13650 82380
rect 13850 82310 14150 82380
rect 14350 82310 14650 82380
rect 14850 82310 15150 82380
rect 15350 82310 15650 82380
rect 15850 82310 16150 82380
rect 16350 82310 16650 82380
rect 16850 82310 17150 82380
rect 17350 82310 17650 82380
rect 17850 82310 18150 82380
rect 18350 82310 18650 82380
rect 18850 82310 19150 82380
rect 19350 82310 19650 82380
rect 19850 82310 20150 82380
rect 20350 82310 20650 82380
rect 20850 82310 21150 82380
rect 21350 82310 21650 82380
rect 21850 82310 22150 82380
rect 22350 82310 22650 82380
rect 22850 82310 23150 82380
rect 23350 82310 23650 82380
rect 23850 82310 24150 82380
rect 24350 82310 24650 82380
rect 24850 82310 25150 82380
rect 25350 82310 25650 82380
rect 25850 82310 26150 82380
rect 26350 82310 26650 82380
rect 26850 82310 27150 82380
rect 27350 82310 27650 82380
rect 27850 82310 28150 82380
rect 28350 82310 28650 82380
rect 28850 82310 29150 82380
rect 29350 82310 29650 82380
rect 29850 82310 30150 82380
rect 30350 82310 30650 82380
rect 30850 82310 31150 82380
rect 31350 82310 31650 82380
rect 31850 82310 32150 82380
rect 32350 82310 32650 82380
rect 32850 82310 33150 82380
rect 33350 82310 33650 82380
rect 33850 82310 34150 82380
rect 34350 82310 34650 82380
rect 34850 82310 35150 82380
rect 35350 82310 35650 82380
rect 35850 82310 36150 82380
rect 36350 82310 36650 82380
rect 36850 82310 37150 82380
rect 37350 82310 37650 82380
rect 37850 82310 38150 82380
rect 38350 82310 38650 82380
rect 38850 82310 39150 82380
rect 39350 82310 39650 82380
rect 39850 82310 40150 82380
rect 40350 82310 40650 82380
rect 40850 82310 41150 82380
rect 41350 82310 41650 82380
rect 41850 82310 42150 82380
rect 42350 82310 42650 82380
rect 42850 82310 43150 82380
rect 43350 82310 43650 82380
rect 43850 82310 44150 82380
rect 44350 82310 44650 82380
rect 44850 82310 45150 82380
rect 45350 82310 45650 82380
rect 45850 82310 46150 82380
rect 46350 82310 46650 82380
rect 46850 82310 47150 82380
rect 47350 82310 47650 82380
rect 47850 82310 48150 82380
rect 48350 82310 48650 82380
rect 48850 82310 49150 82380
rect 49350 82310 49650 82380
rect 49850 82310 50150 82380
rect 50350 82310 50650 82380
rect 50850 82310 51150 82380
rect 51350 82310 51650 82380
rect 51850 82310 52150 82380
rect 52350 82310 52650 82380
rect 52850 82310 53150 82380
rect 53350 82310 53650 82380
rect 53850 82310 54150 82380
rect 54350 82310 54650 82380
rect 54850 82310 55150 82380
rect 55350 82310 55650 82380
rect 55850 82310 56150 82380
rect 56350 82310 56650 82380
rect 56850 82310 57150 82380
rect 57350 82310 57650 82380
rect 57850 82310 58150 82380
rect 58350 82310 58650 82380
rect 58850 82310 59150 82380
rect 59350 82310 59650 82380
rect 59850 82310 60150 82380
rect 60350 82310 60650 82380
rect 60850 82310 61150 82380
rect 61350 82310 61650 82380
rect 61850 82310 62150 82380
rect 62350 82310 62650 82380
rect 62850 82310 63150 82380
rect 63350 82310 63650 82380
rect 63850 82310 64150 82380
rect 64350 82310 64650 82380
rect 64850 82310 65150 82380
rect 65350 82310 65650 82380
rect 65850 82310 66150 82380
rect 66350 82310 66650 82380
rect 66850 82310 67150 82380
rect 67350 82310 67650 82380
rect 67850 82310 68150 82380
rect 68350 82310 68650 82380
rect 68850 82310 69150 82380
rect 69350 82310 69650 82380
rect 69850 82310 70150 82380
rect 70350 82310 70650 82380
rect 70850 82310 71150 82380
rect 71350 82310 71650 82380
rect 71850 82310 72150 82380
rect 72350 82310 72650 82380
rect 72850 82310 73150 82380
rect 73350 82310 73650 82380
rect 73850 82310 74150 82380
rect 74350 82310 74650 82380
rect 74850 82310 75150 82380
rect 75350 82310 75650 82380
rect 75850 82310 76150 82380
rect 76350 82310 76650 82380
rect 76850 82310 77150 82380
rect 77350 82310 77650 82380
rect 77850 82310 78150 82380
rect 78350 82310 78650 82380
rect 78850 82310 79150 82380
rect 79350 82310 79650 82380
rect 79850 82310 80150 82380
rect 80350 82310 80650 82380
rect 80850 82310 81150 82380
rect 81350 82310 81650 82380
rect 81850 82310 82150 82380
rect 82350 82310 82650 82380
rect 82850 82310 83150 82380
rect 83350 82310 83650 82380
rect 83850 82310 84150 82380
rect 84350 82310 84650 82380
rect 84850 82310 85150 82380
rect 85350 82310 85650 82380
rect 85850 82310 86150 82380
rect 86350 82310 86650 82380
rect 86850 82310 87150 82380
rect 87350 82310 87650 82380
rect 87850 82310 88150 82380
rect 88350 82310 88650 82380
rect 88850 82310 89150 82380
rect 89350 82310 89650 82380
rect 89850 82310 90150 82380
rect 90350 82310 90650 82380
rect 90850 82310 91150 82380
rect 91350 82310 91650 82380
rect 91850 82310 92150 82380
rect 92350 82310 92650 82380
rect 92850 82310 93150 82380
rect 93350 82310 93650 82380
rect 93850 82310 94150 82380
rect 94350 82310 94650 82380
rect 94850 82310 95150 82380
rect 95350 82310 95650 82380
rect 95850 82310 96150 82380
rect 96350 82310 96650 82380
rect 96850 82310 97150 82380
rect 97350 82310 97650 82380
rect 97850 82310 98150 82380
rect 98350 82310 98650 82380
rect 98850 82310 99150 82380
rect 99350 82310 99650 82380
rect 99850 82310 100150 82380
rect 100350 82310 100500 82380
rect -83500 82300 100500 82310
rect -83500 82280 -83380 82300
rect -83120 82280 -82880 82300
rect -82620 82280 -82380 82300
rect -82120 82280 -81880 82300
rect -81620 82280 -81380 82300
rect -81120 82280 -80880 82300
rect -80620 82280 -80380 82300
rect -80120 82280 -79880 82300
rect -79620 82280 -79380 82300
rect -79120 82280 -78880 82300
rect -78620 82280 -78380 82300
rect -78120 82280 -77880 82300
rect -77620 82280 -77380 82300
rect -77120 82280 -76880 82300
rect -76620 82280 -76380 82300
rect -76120 82280 -75880 82300
rect -75620 82280 -75380 82300
rect -75120 82280 -74880 82300
rect -74620 82280 -74380 82300
rect -74120 82280 -73880 82300
rect -73620 82280 -73380 82300
rect -73120 82280 -72880 82300
rect -72620 82280 -72380 82300
rect -72120 82280 -71880 82300
rect -71620 82280 -71380 82300
rect -71120 82280 -70880 82300
rect -70620 82280 -70380 82300
rect -70120 82280 -69880 82300
rect -69620 82280 -69380 82300
rect -69120 82280 -68880 82300
rect -68620 82280 -68380 82300
rect -68120 82280 -67880 82300
rect -67620 82280 -67380 82300
rect -67120 82280 -66880 82300
rect -66620 82280 -66380 82300
rect -66120 82280 -65880 82300
rect -65620 82280 -65380 82300
rect -65120 82280 -64880 82300
rect -64620 82280 -64380 82300
rect -64120 82280 -63880 82300
rect -63620 82280 -63380 82300
rect -63120 82280 -62880 82300
rect -62620 82280 -62380 82300
rect -62120 82280 -61880 82300
rect -61620 82280 -61380 82300
rect -61120 82280 -60880 82300
rect -60620 82280 -60380 82300
rect -60120 82280 -59880 82300
rect -59620 82280 -59380 82300
rect -59120 82280 -58880 82300
rect -58620 82280 -58380 82300
rect -58120 82280 -57880 82300
rect -57620 82280 -57380 82300
rect -57120 82280 -56880 82300
rect -56620 82280 -56380 82300
rect -56120 82280 -55880 82300
rect -55620 82280 -55380 82300
rect -55120 82280 -54880 82300
rect -54620 82280 -54380 82300
rect -54120 82280 -53880 82300
rect -53620 82280 -53380 82300
rect -53120 82280 -52880 82300
rect -52620 82280 -52380 82300
rect -52120 82280 -51880 82300
rect -51620 82280 -51380 82300
rect -51120 82280 -50880 82300
rect -50620 82280 -50380 82300
rect -50120 82280 -49880 82300
rect -49620 82280 -49380 82300
rect -49120 82280 -48880 82300
rect -48620 82280 -48380 82300
rect -48120 82280 -47880 82300
rect -47620 82280 -47380 82300
rect -47120 82280 -46880 82300
rect -46620 82280 -46380 82300
rect -46120 82280 -45880 82300
rect -45620 82280 -45380 82300
rect -45120 82280 -44880 82300
rect -44620 82280 -44380 82300
rect -44120 82280 -43880 82300
rect -43620 82280 -43380 82300
rect -43120 82280 -42880 82300
rect -42620 82280 -42380 82300
rect -42120 82280 -41880 82300
rect -41620 82280 -41380 82300
rect -41120 82280 -40880 82300
rect -40620 82280 -40380 82300
rect -40120 82280 -39880 82300
rect -39620 82280 -39380 82300
rect -39120 82280 -38880 82300
rect -38620 82280 -38380 82300
rect -38120 82280 -37880 82300
rect -37620 82280 -37380 82300
rect -37120 82280 -36880 82300
rect -36620 82280 -36380 82300
rect -36120 82280 -35880 82300
rect -35620 82280 -35380 82300
rect -35120 82280 -34880 82300
rect -34620 82280 -34380 82300
rect -34120 82280 -33880 82300
rect -33620 82280 -33380 82300
rect -33120 82280 -32880 82300
rect -32620 82280 -32380 82300
rect -32120 82280 -31880 82300
rect -31620 82280 -31380 82300
rect -31120 82280 -30880 82300
rect -30620 82280 -30380 82300
rect -30120 82280 -29880 82300
rect -29620 82280 -29380 82300
rect -29120 82280 -28880 82300
rect -28620 82280 -28380 82300
rect -28120 82280 -27880 82300
rect -27620 82280 -27380 82300
rect -27120 82280 -26880 82300
rect -26620 82280 -26380 82300
rect -26120 82280 -25880 82300
rect -25620 82280 -25380 82300
rect -25120 82280 -24880 82300
rect -24620 82280 -24380 82300
rect -24120 82280 -23880 82300
rect -23620 82280 -23380 82300
rect -23120 82280 -22880 82300
rect -22620 82280 -22380 82300
rect -22120 82280 -21880 82300
rect -21620 82280 -21380 82300
rect -21120 82280 -20880 82300
rect -20620 82280 -20380 82300
rect -20120 82280 -19880 82300
rect -19620 82280 -19380 82300
rect -19120 82280 -18880 82300
rect -18620 82280 -18380 82300
rect -18120 82280 -17880 82300
rect -17620 82280 -17380 82300
rect -17120 82280 -16880 82300
rect -16620 82280 -16380 82300
rect -16120 82280 -15880 82300
rect -15620 82280 -15380 82300
rect -15120 82280 -14880 82300
rect -14620 82280 -14380 82300
rect -14120 82280 -13880 82300
rect -13620 82280 -13380 82300
rect -13120 82280 -12880 82300
rect -12620 82280 -12380 82300
rect -12120 82280 -11880 82300
rect -11620 82280 -11380 82300
rect -11120 82280 -10880 82300
rect -10620 82280 -10380 82300
rect -10120 82280 -9880 82300
rect -9620 82280 -9380 82300
rect -9120 82280 -8880 82300
rect -8620 82280 -8380 82300
rect -8120 82280 -7880 82300
rect -7620 82280 -7380 82300
rect -7120 82280 -6880 82300
rect -6620 82280 -6380 82300
rect -6120 82280 -5880 82300
rect -5620 82280 -5380 82300
rect -5120 82280 -4880 82300
rect -4620 82280 -4380 82300
rect -4120 82280 -3880 82300
rect -3620 82280 -3380 82300
rect -3120 82280 -2880 82300
rect -2620 82280 -2380 82300
rect -2120 82280 -1880 82300
rect -1620 82280 -1380 82300
rect -1120 82280 -880 82300
rect -620 82280 -380 82300
rect -120 82280 120 82300
rect 380 82280 620 82300
rect 880 82280 1120 82300
rect 1380 82280 1620 82300
rect 1880 82280 2120 82300
rect 2380 82280 2620 82300
rect 2880 82280 3120 82300
rect 3380 82280 3620 82300
rect 3880 82280 4120 82300
rect 4380 82280 4620 82300
rect 4880 82280 5120 82300
rect 5380 82280 5620 82300
rect 5880 82280 6120 82300
rect 6380 82280 6620 82300
rect 6880 82280 7120 82300
rect 7380 82280 7620 82300
rect 7880 82280 8120 82300
rect 8380 82280 8620 82300
rect 8880 82280 9120 82300
rect 9380 82280 9620 82300
rect 9880 82280 10120 82300
rect 10380 82280 10620 82300
rect 10880 82280 11120 82300
rect 11380 82280 11620 82300
rect 11880 82280 12120 82300
rect 12380 82280 12620 82300
rect 12880 82280 13120 82300
rect 13380 82280 13620 82300
rect 13880 82280 14120 82300
rect 14380 82280 14620 82300
rect 14880 82280 15120 82300
rect 15380 82280 15620 82300
rect 15880 82280 16120 82300
rect 16380 82280 16620 82300
rect 16880 82280 17120 82300
rect 17380 82280 17620 82300
rect 17880 82280 18120 82300
rect 18380 82280 18620 82300
rect 18880 82280 19120 82300
rect 19380 82280 19620 82300
rect 19880 82280 20120 82300
rect 20380 82280 20620 82300
rect 20880 82280 21120 82300
rect 21380 82280 21620 82300
rect 21880 82280 22120 82300
rect 22380 82280 22620 82300
rect 22880 82280 23120 82300
rect 23380 82280 23620 82300
rect 23880 82280 24120 82300
rect 24380 82280 24620 82300
rect 24880 82280 25120 82300
rect 25380 82280 25620 82300
rect 25880 82280 26120 82300
rect 26380 82280 26620 82300
rect 26880 82280 27120 82300
rect 27380 82280 27620 82300
rect 27880 82280 28120 82300
rect 28380 82280 28620 82300
rect 28880 82280 29120 82300
rect 29380 82280 29620 82300
rect 29880 82280 30120 82300
rect 30380 82280 30620 82300
rect 30880 82280 31120 82300
rect 31380 82280 31620 82300
rect 31880 82280 32120 82300
rect 32380 82280 32620 82300
rect 32880 82280 33120 82300
rect 33380 82280 33620 82300
rect 33880 82280 34120 82300
rect 34380 82280 34620 82300
rect 34880 82280 35120 82300
rect 35380 82280 35620 82300
rect 35880 82280 36120 82300
rect 36380 82280 36620 82300
rect 36880 82280 37120 82300
rect 37380 82280 37620 82300
rect 37880 82280 38120 82300
rect 38380 82280 38620 82300
rect 38880 82280 39120 82300
rect 39380 82280 39620 82300
rect 39880 82280 40120 82300
rect 40380 82280 40620 82300
rect 40880 82280 41120 82300
rect 41380 82280 41620 82300
rect 41880 82280 42120 82300
rect 42380 82280 42620 82300
rect 42880 82280 43120 82300
rect 43380 82280 43620 82300
rect 43880 82280 44120 82300
rect 44380 82280 44620 82300
rect 44880 82280 45120 82300
rect 45380 82280 45620 82300
rect 45880 82280 46120 82300
rect 46380 82280 46620 82300
rect 46880 82280 47120 82300
rect 47380 82280 47620 82300
rect 47880 82280 48120 82300
rect 48380 82280 48620 82300
rect 48880 82280 49120 82300
rect 49380 82280 49620 82300
rect 49880 82280 50120 82300
rect 50380 82280 50620 82300
rect 50880 82280 51120 82300
rect 51380 82280 51620 82300
rect 51880 82280 52120 82300
rect 52380 82280 52620 82300
rect 52880 82280 53120 82300
rect 53380 82280 53620 82300
rect 53880 82280 54120 82300
rect 54380 82280 54620 82300
rect 54880 82280 55120 82300
rect 55380 82280 55620 82300
rect 55880 82280 56120 82300
rect 56380 82280 56620 82300
rect 56880 82280 57120 82300
rect 57380 82280 57620 82300
rect 57880 82280 58120 82300
rect 58380 82280 58620 82300
rect 58880 82280 59120 82300
rect 59380 82280 59620 82300
rect 59880 82280 60120 82300
rect 60380 82280 60620 82300
rect 60880 82280 61120 82300
rect 61380 82280 61620 82300
rect 61880 82280 62120 82300
rect 62380 82280 62620 82300
rect 62880 82280 63120 82300
rect 63380 82280 63620 82300
rect 63880 82280 64120 82300
rect 64380 82280 64620 82300
rect 64880 82280 65120 82300
rect 65380 82280 65620 82300
rect 65880 82280 66120 82300
rect 66380 82280 66620 82300
rect 66880 82280 67120 82300
rect 67380 82280 67620 82300
rect 67880 82280 68120 82300
rect 68380 82280 68620 82300
rect 68880 82280 69120 82300
rect 69380 82280 69620 82300
rect 69880 82280 70120 82300
rect 70380 82280 70620 82300
rect 70880 82280 71120 82300
rect 71380 82280 71620 82300
rect 71880 82280 72120 82300
rect 72380 82280 72620 82300
rect 72880 82280 73120 82300
rect 73380 82280 73620 82300
rect 73880 82280 74120 82300
rect 74380 82280 74620 82300
rect 74880 82280 75120 82300
rect 75380 82280 75620 82300
rect 75880 82280 76120 82300
rect 76380 82280 76620 82300
rect 76880 82280 77120 82300
rect 77380 82280 77620 82300
rect 77880 82280 78120 82300
rect 78380 82280 78620 82300
rect 78880 82280 79120 82300
rect 79380 82280 79620 82300
rect 79880 82280 80120 82300
rect 80380 82280 80620 82300
rect 80880 82280 81120 82300
rect 81380 82280 81620 82300
rect 81880 82280 82120 82300
rect 82380 82280 82620 82300
rect 82880 82280 83120 82300
rect 83380 82280 83620 82300
rect 83880 82280 84120 82300
rect 84380 82280 84620 82300
rect 84880 82280 85120 82300
rect 85380 82280 85620 82300
rect 85880 82280 86120 82300
rect 86380 82280 86620 82300
rect 86880 82280 87120 82300
rect 87380 82280 87620 82300
rect 87880 82280 88120 82300
rect 88380 82280 88620 82300
rect 88880 82280 89120 82300
rect 89380 82280 89620 82300
rect 89880 82280 90120 82300
rect 90380 82280 90620 82300
rect 90880 82280 91120 82300
rect 91380 82280 91620 82300
rect 91880 82280 92120 82300
rect 92380 82280 92620 82300
rect 92880 82280 93120 82300
rect 93380 82280 93620 82300
rect 93880 82280 94120 82300
rect 94380 82280 94620 82300
rect 94880 82280 95120 82300
rect 95380 82280 95620 82300
rect 95880 82280 96120 82300
rect 96380 82280 96620 82300
rect 96880 82280 97120 82300
rect 97380 82280 97620 82300
rect 97880 82280 98120 82300
rect 98380 82280 98620 82300
rect 98880 82280 99120 82300
rect 99380 82280 99620 82300
rect 99880 82280 100120 82300
rect 100380 82280 100500 82300
rect -83500 82250 -83400 82280
rect -83500 82050 -83480 82250
rect -83410 82050 -83400 82250
rect -83500 82020 -83400 82050
rect -83100 82250 -82900 82280
rect -83100 82050 -83090 82250
rect -83020 82050 -82980 82250
rect -82910 82050 -82900 82250
rect -83100 82020 -82900 82050
rect -82600 82250 -82400 82280
rect -82600 82050 -82590 82250
rect -82520 82050 -82480 82250
rect -82410 82050 -82400 82250
rect -82600 82020 -82400 82050
rect -82100 82250 -81900 82280
rect -82100 82050 -82090 82250
rect -82020 82050 -81980 82250
rect -81910 82050 -81900 82250
rect -82100 82020 -81900 82050
rect -81600 82250 -81400 82280
rect -81600 82050 -81590 82250
rect -81520 82050 -81480 82250
rect -81410 82050 -81400 82250
rect -81600 82020 -81400 82050
rect -81100 82250 -80900 82280
rect -81100 82050 -81090 82250
rect -81020 82050 -80980 82250
rect -80910 82050 -80900 82250
rect -81100 82020 -80900 82050
rect -80600 82250 -80400 82280
rect -80600 82050 -80590 82250
rect -80520 82050 -80480 82250
rect -80410 82050 -80400 82250
rect -80600 82020 -80400 82050
rect -80100 82250 -79900 82280
rect -80100 82050 -80090 82250
rect -80020 82050 -79980 82250
rect -79910 82050 -79900 82250
rect -80100 82020 -79900 82050
rect -79600 82250 -79400 82280
rect -79600 82050 -79590 82250
rect -79520 82050 -79480 82250
rect -79410 82050 -79400 82250
rect -79600 82020 -79400 82050
rect -79100 82250 -78900 82280
rect -79100 82050 -79090 82250
rect -79020 82050 -78980 82250
rect -78910 82050 -78900 82250
rect -79100 82020 -78900 82050
rect -78600 82250 -78400 82280
rect -78600 82050 -78590 82250
rect -78520 82050 -78480 82250
rect -78410 82050 -78400 82250
rect -78600 82020 -78400 82050
rect -78100 82250 -77900 82280
rect -78100 82050 -78090 82250
rect -78020 82050 -77980 82250
rect -77910 82050 -77900 82250
rect -78100 82020 -77900 82050
rect -77600 82250 -77400 82280
rect -77600 82050 -77590 82250
rect -77520 82050 -77480 82250
rect -77410 82050 -77400 82250
rect -77600 82020 -77400 82050
rect -77100 82250 -76900 82280
rect -77100 82050 -77090 82250
rect -77020 82050 -76980 82250
rect -76910 82050 -76900 82250
rect -77100 82020 -76900 82050
rect -76600 82250 -76400 82280
rect -76600 82050 -76590 82250
rect -76520 82050 -76480 82250
rect -76410 82050 -76400 82250
rect -76600 82020 -76400 82050
rect -76100 82250 -75900 82280
rect -76100 82050 -76090 82250
rect -76020 82050 -75980 82250
rect -75910 82050 -75900 82250
rect -76100 82020 -75900 82050
rect -75600 82250 -75400 82280
rect -75600 82050 -75590 82250
rect -75520 82050 -75480 82250
rect -75410 82050 -75400 82250
rect -75600 82020 -75400 82050
rect -75100 82250 -74900 82280
rect -75100 82050 -75090 82250
rect -75020 82050 -74980 82250
rect -74910 82050 -74900 82250
rect -75100 82020 -74900 82050
rect -74600 82250 -74400 82280
rect -74600 82050 -74590 82250
rect -74520 82050 -74480 82250
rect -74410 82050 -74400 82250
rect -74600 82020 -74400 82050
rect -74100 82250 -73900 82280
rect -74100 82050 -74090 82250
rect -74020 82050 -73980 82250
rect -73910 82050 -73900 82250
rect -74100 82020 -73900 82050
rect -73600 82250 -73400 82280
rect -73600 82050 -73590 82250
rect -73520 82050 -73480 82250
rect -73410 82050 -73400 82250
rect -73600 82020 -73400 82050
rect -73100 82250 -72900 82280
rect -73100 82050 -73090 82250
rect -73020 82050 -72980 82250
rect -72910 82050 -72900 82250
rect -73100 82020 -72900 82050
rect -72600 82250 -72400 82280
rect -72600 82050 -72590 82250
rect -72520 82050 -72480 82250
rect -72410 82050 -72400 82250
rect -72600 82020 -72400 82050
rect -72100 82250 -71900 82280
rect -72100 82050 -72090 82250
rect -72020 82050 -71980 82250
rect -71910 82050 -71900 82250
rect -72100 82020 -71900 82050
rect -71600 82250 -71400 82280
rect -71600 82050 -71590 82250
rect -71520 82050 -71480 82250
rect -71410 82050 -71400 82250
rect -71600 82020 -71400 82050
rect -71100 82250 -70900 82280
rect -71100 82050 -71090 82250
rect -71020 82050 -70980 82250
rect -70910 82050 -70900 82250
rect -71100 82020 -70900 82050
rect -70600 82250 -70400 82280
rect -70600 82050 -70590 82250
rect -70520 82050 -70480 82250
rect -70410 82050 -70400 82250
rect -70600 82020 -70400 82050
rect -70100 82250 -69900 82280
rect -70100 82050 -70090 82250
rect -70020 82050 -69980 82250
rect -69910 82050 -69900 82250
rect -70100 82020 -69900 82050
rect -69600 82250 -69400 82280
rect -69600 82050 -69590 82250
rect -69520 82050 -69480 82250
rect -69410 82050 -69400 82250
rect -69600 82020 -69400 82050
rect -69100 82250 -68900 82280
rect -69100 82050 -69090 82250
rect -69020 82050 -68980 82250
rect -68910 82050 -68900 82250
rect -69100 82020 -68900 82050
rect -68600 82250 -68400 82280
rect -68600 82050 -68590 82250
rect -68520 82050 -68480 82250
rect -68410 82050 -68400 82250
rect -68600 82020 -68400 82050
rect -68100 82250 -67900 82280
rect -68100 82050 -68090 82250
rect -68020 82050 -67980 82250
rect -67910 82050 -67900 82250
rect -68100 82020 -67900 82050
rect -67600 82250 -67400 82280
rect -67600 82050 -67590 82250
rect -67520 82050 -67480 82250
rect -67410 82050 -67400 82250
rect -67600 82020 -67400 82050
rect -67100 82250 -66900 82280
rect -67100 82050 -67090 82250
rect -67020 82050 -66980 82250
rect -66910 82050 -66900 82250
rect -67100 82020 -66900 82050
rect -66600 82250 -66400 82280
rect -66600 82050 -66590 82250
rect -66520 82050 -66480 82250
rect -66410 82050 -66400 82250
rect -66600 82020 -66400 82050
rect -66100 82250 -65900 82280
rect -66100 82050 -66090 82250
rect -66020 82050 -65980 82250
rect -65910 82050 -65900 82250
rect -66100 82020 -65900 82050
rect -65600 82250 -65400 82280
rect -65600 82050 -65590 82250
rect -65520 82050 -65480 82250
rect -65410 82050 -65400 82250
rect -65600 82020 -65400 82050
rect -65100 82250 -64900 82280
rect -65100 82050 -65090 82250
rect -65020 82050 -64980 82250
rect -64910 82050 -64900 82250
rect -65100 82020 -64900 82050
rect -64600 82250 -64400 82280
rect -64600 82050 -64590 82250
rect -64520 82050 -64480 82250
rect -64410 82050 -64400 82250
rect -64600 82020 -64400 82050
rect -64100 82250 -63900 82280
rect -64100 82050 -64090 82250
rect -64020 82050 -63980 82250
rect -63910 82050 -63900 82250
rect -64100 82020 -63900 82050
rect -63600 82250 -63400 82280
rect -63600 82050 -63590 82250
rect -63520 82050 -63480 82250
rect -63410 82050 -63400 82250
rect -63600 82020 -63400 82050
rect -63100 82250 -62900 82280
rect -63100 82050 -63090 82250
rect -63020 82050 -62980 82250
rect -62910 82050 -62900 82250
rect -63100 82020 -62900 82050
rect -62600 82250 -62400 82280
rect -62600 82050 -62590 82250
rect -62520 82050 -62480 82250
rect -62410 82050 -62400 82250
rect -62600 82020 -62400 82050
rect -62100 82250 -61900 82280
rect -62100 82050 -62090 82250
rect -62020 82050 -61980 82250
rect -61910 82050 -61900 82250
rect -62100 82020 -61900 82050
rect -61600 82250 -61400 82280
rect -61600 82050 -61590 82250
rect -61520 82050 -61480 82250
rect -61410 82050 -61400 82250
rect -61600 82020 -61400 82050
rect -61100 82250 -60900 82280
rect -61100 82050 -61090 82250
rect -61020 82050 -60980 82250
rect -60910 82050 -60900 82250
rect -61100 82020 -60900 82050
rect -60600 82250 -60400 82280
rect -60600 82050 -60590 82250
rect -60520 82050 -60480 82250
rect -60410 82050 -60400 82250
rect -60600 82020 -60400 82050
rect -60100 82250 -59900 82280
rect -60100 82050 -60090 82250
rect -60020 82050 -59980 82250
rect -59910 82050 -59900 82250
rect -60100 82020 -59900 82050
rect -59600 82250 -59400 82280
rect -59600 82050 -59590 82250
rect -59520 82050 -59480 82250
rect -59410 82050 -59400 82250
rect -59600 82020 -59400 82050
rect -59100 82250 -58900 82280
rect -59100 82050 -59090 82250
rect -59020 82050 -58980 82250
rect -58910 82050 -58900 82250
rect -59100 82020 -58900 82050
rect -58600 82250 -58400 82280
rect -58600 82050 -58590 82250
rect -58520 82050 -58480 82250
rect -58410 82050 -58400 82250
rect -58600 82020 -58400 82050
rect -58100 82250 -57900 82280
rect -58100 82050 -58090 82250
rect -58020 82050 -57980 82250
rect -57910 82050 -57900 82250
rect -58100 82020 -57900 82050
rect -57600 82250 -57400 82280
rect -57600 82050 -57590 82250
rect -57520 82050 -57480 82250
rect -57410 82050 -57400 82250
rect -57600 82020 -57400 82050
rect -57100 82250 -56900 82280
rect -57100 82050 -57090 82250
rect -57020 82050 -56980 82250
rect -56910 82050 -56900 82250
rect -57100 82020 -56900 82050
rect -56600 82250 -56400 82280
rect -56600 82050 -56590 82250
rect -56520 82050 -56480 82250
rect -56410 82050 -56400 82250
rect -56600 82020 -56400 82050
rect -56100 82250 -55900 82280
rect -56100 82050 -56090 82250
rect -56020 82050 -55980 82250
rect -55910 82050 -55900 82250
rect -56100 82020 -55900 82050
rect -55600 82250 -55400 82280
rect -55600 82050 -55590 82250
rect -55520 82050 -55480 82250
rect -55410 82050 -55400 82250
rect -55600 82020 -55400 82050
rect -55100 82250 -54900 82280
rect -55100 82050 -55090 82250
rect -55020 82050 -54980 82250
rect -54910 82050 -54900 82250
rect -55100 82020 -54900 82050
rect -54600 82250 -54400 82280
rect -54600 82050 -54590 82250
rect -54520 82050 -54480 82250
rect -54410 82050 -54400 82250
rect -54600 82020 -54400 82050
rect -54100 82250 -53900 82280
rect -54100 82050 -54090 82250
rect -54020 82050 -53980 82250
rect -53910 82050 -53900 82250
rect -54100 82020 -53900 82050
rect -53600 82250 -53400 82280
rect -53600 82050 -53590 82250
rect -53520 82050 -53480 82250
rect -53410 82050 -53400 82250
rect -53600 82020 -53400 82050
rect -53100 82250 -52900 82280
rect -53100 82050 -53090 82250
rect -53020 82050 -52980 82250
rect -52910 82050 -52900 82250
rect -53100 82020 -52900 82050
rect -52600 82250 -52400 82280
rect -52600 82050 -52590 82250
rect -52520 82050 -52480 82250
rect -52410 82050 -52400 82250
rect -52600 82020 -52400 82050
rect -52100 82250 -51900 82280
rect -52100 82050 -52090 82250
rect -52020 82050 -51980 82250
rect -51910 82050 -51900 82250
rect -52100 82020 -51900 82050
rect -51600 82250 -51400 82280
rect -51600 82050 -51590 82250
rect -51520 82050 -51480 82250
rect -51410 82050 -51400 82250
rect -51600 82020 -51400 82050
rect -51100 82250 -50900 82280
rect -51100 82050 -51090 82250
rect -51020 82050 -50980 82250
rect -50910 82050 -50900 82250
rect -51100 82020 -50900 82050
rect -50600 82250 -50400 82280
rect -50600 82050 -50590 82250
rect -50520 82050 -50480 82250
rect -50410 82050 -50400 82250
rect -50600 82020 -50400 82050
rect -50100 82250 -49900 82280
rect -50100 82050 -50090 82250
rect -50020 82050 -49980 82250
rect -49910 82050 -49900 82250
rect -50100 82020 -49900 82050
rect -49600 82250 -49400 82280
rect -49600 82050 -49590 82250
rect -49520 82050 -49480 82250
rect -49410 82050 -49400 82250
rect -49600 82020 -49400 82050
rect -49100 82250 -48900 82280
rect -49100 82050 -49090 82250
rect -49020 82050 -48980 82250
rect -48910 82050 -48900 82250
rect -49100 82020 -48900 82050
rect -48600 82250 -48400 82280
rect -48600 82050 -48590 82250
rect -48520 82050 -48480 82250
rect -48410 82050 -48400 82250
rect -48600 82020 -48400 82050
rect -48100 82250 -47900 82280
rect -48100 82050 -48090 82250
rect -48020 82050 -47980 82250
rect -47910 82050 -47900 82250
rect -48100 82020 -47900 82050
rect -47600 82250 -47400 82280
rect -47600 82050 -47590 82250
rect -47520 82050 -47480 82250
rect -47410 82050 -47400 82250
rect -47600 82020 -47400 82050
rect -47100 82250 -46900 82280
rect -47100 82050 -47090 82250
rect -47020 82050 -46980 82250
rect -46910 82050 -46900 82250
rect -47100 82020 -46900 82050
rect -46600 82250 -46400 82280
rect -46600 82050 -46590 82250
rect -46520 82050 -46480 82250
rect -46410 82050 -46400 82250
rect -46600 82020 -46400 82050
rect -46100 82250 -45900 82280
rect -46100 82050 -46090 82250
rect -46020 82050 -45980 82250
rect -45910 82050 -45900 82250
rect -46100 82020 -45900 82050
rect -45600 82250 -45400 82280
rect -45600 82050 -45590 82250
rect -45520 82050 -45480 82250
rect -45410 82050 -45400 82250
rect -45600 82020 -45400 82050
rect -45100 82250 -44900 82280
rect -45100 82050 -45090 82250
rect -45020 82050 -44980 82250
rect -44910 82050 -44900 82250
rect -45100 82020 -44900 82050
rect -44600 82250 -44400 82280
rect -44600 82050 -44590 82250
rect -44520 82050 -44480 82250
rect -44410 82050 -44400 82250
rect -44600 82020 -44400 82050
rect -44100 82250 -43900 82280
rect -44100 82050 -44090 82250
rect -44020 82050 -43980 82250
rect -43910 82050 -43900 82250
rect -44100 82020 -43900 82050
rect -43600 82250 -43400 82280
rect -43600 82050 -43590 82250
rect -43520 82050 -43480 82250
rect -43410 82050 -43400 82250
rect -43600 82020 -43400 82050
rect -43100 82250 -42900 82280
rect -43100 82050 -43090 82250
rect -43020 82050 -42980 82250
rect -42910 82050 -42900 82250
rect -43100 82020 -42900 82050
rect -42600 82250 -42400 82280
rect -42600 82050 -42590 82250
rect -42520 82050 -42480 82250
rect -42410 82050 -42400 82250
rect -42600 82020 -42400 82050
rect -42100 82250 -41900 82280
rect -42100 82050 -42090 82250
rect -42020 82050 -41980 82250
rect -41910 82050 -41900 82250
rect -42100 82020 -41900 82050
rect -41600 82250 -41400 82280
rect -41600 82050 -41590 82250
rect -41520 82050 -41480 82250
rect -41410 82050 -41400 82250
rect -41600 82020 -41400 82050
rect -41100 82250 -40900 82280
rect -41100 82050 -41090 82250
rect -41020 82050 -40980 82250
rect -40910 82050 -40900 82250
rect -41100 82020 -40900 82050
rect -40600 82250 -40400 82280
rect -40600 82050 -40590 82250
rect -40520 82050 -40480 82250
rect -40410 82050 -40400 82250
rect -40600 82020 -40400 82050
rect -40100 82250 -39900 82280
rect -40100 82050 -40090 82250
rect -40020 82050 -39980 82250
rect -39910 82050 -39900 82250
rect -40100 82020 -39900 82050
rect -39600 82250 -39400 82280
rect -39600 82050 -39590 82250
rect -39520 82050 -39480 82250
rect -39410 82050 -39400 82250
rect -39600 82020 -39400 82050
rect -39100 82250 -38900 82280
rect -39100 82050 -39090 82250
rect -39020 82050 -38980 82250
rect -38910 82050 -38900 82250
rect -39100 82020 -38900 82050
rect -38600 82250 -38400 82280
rect -38600 82050 -38590 82250
rect -38520 82050 -38480 82250
rect -38410 82050 -38400 82250
rect -38600 82020 -38400 82050
rect -38100 82250 -37900 82280
rect -38100 82050 -38090 82250
rect -38020 82050 -37980 82250
rect -37910 82050 -37900 82250
rect -38100 82020 -37900 82050
rect -37600 82250 -37400 82280
rect -37600 82050 -37590 82250
rect -37520 82050 -37480 82250
rect -37410 82050 -37400 82250
rect -37600 82020 -37400 82050
rect -37100 82250 -36900 82280
rect -37100 82050 -37090 82250
rect -37020 82050 -36980 82250
rect -36910 82050 -36900 82250
rect -37100 82020 -36900 82050
rect -36600 82250 -36400 82280
rect -36600 82050 -36590 82250
rect -36520 82050 -36480 82250
rect -36410 82050 -36400 82250
rect -36600 82020 -36400 82050
rect -36100 82250 -35900 82280
rect -36100 82050 -36090 82250
rect -36020 82050 -35980 82250
rect -35910 82050 -35900 82250
rect -36100 82020 -35900 82050
rect -35600 82250 -35400 82280
rect -35600 82050 -35590 82250
rect -35520 82050 -35480 82250
rect -35410 82050 -35400 82250
rect -35600 82020 -35400 82050
rect -35100 82250 -34900 82280
rect -35100 82050 -35090 82250
rect -35020 82050 -34980 82250
rect -34910 82050 -34900 82250
rect -35100 82020 -34900 82050
rect -34600 82250 -34400 82280
rect -34600 82050 -34590 82250
rect -34520 82050 -34480 82250
rect -34410 82050 -34400 82250
rect -34600 82020 -34400 82050
rect -34100 82250 -33900 82280
rect -34100 82050 -34090 82250
rect -34020 82050 -33980 82250
rect -33910 82050 -33900 82250
rect -34100 82020 -33900 82050
rect -33600 82250 -33400 82280
rect -33600 82050 -33590 82250
rect -33520 82050 -33480 82250
rect -33410 82050 -33400 82250
rect -33600 82020 -33400 82050
rect -33100 82250 -32900 82280
rect -33100 82050 -33090 82250
rect -33020 82050 -32980 82250
rect -32910 82050 -32900 82250
rect -33100 82020 -32900 82050
rect -32600 82250 -32400 82280
rect -32600 82050 -32590 82250
rect -32520 82050 -32480 82250
rect -32410 82050 -32400 82250
rect -32600 82020 -32400 82050
rect -32100 82250 -31900 82280
rect -32100 82050 -32090 82250
rect -32020 82050 -31980 82250
rect -31910 82050 -31900 82250
rect -32100 82020 -31900 82050
rect -31600 82250 -31400 82280
rect -31600 82050 -31590 82250
rect -31520 82050 -31480 82250
rect -31410 82050 -31400 82250
rect -31600 82020 -31400 82050
rect -31100 82250 -30900 82280
rect -31100 82050 -31090 82250
rect -31020 82050 -30980 82250
rect -30910 82050 -30900 82250
rect -31100 82020 -30900 82050
rect -30600 82250 -30400 82280
rect -30600 82050 -30590 82250
rect -30520 82050 -30480 82250
rect -30410 82050 -30400 82250
rect -30600 82020 -30400 82050
rect -30100 82250 -29900 82280
rect -30100 82050 -30090 82250
rect -30020 82050 -29980 82250
rect -29910 82050 -29900 82250
rect -30100 82020 -29900 82050
rect -29600 82250 -29400 82280
rect -29600 82050 -29590 82250
rect -29520 82050 -29480 82250
rect -29410 82050 -29400 82250
rect -29600 82020 -29400 82050
rect -29100 82250 -28900 82280
rect -29100 82050 -29090 82250
rect -29020 82050 -28980 82250
rect -28910 82050 -28900 82250
rect -29100 82020 -28900 82050
rect -28600 82250 -28400 82280
rect -28600 82050 -28590 82250
rect -28520 82050 -28480 82250
rect -28410 82050 -28400 82250
rect -28600 82020 -28400 82050
rect -28100 82250 -27900 82280
rect -28100 82050 -28090 82250
rect -28020 82050 -27980 82250
rect -27910 82050 -27900 82250
rect -28100 82020 -27900 82050
rect -27600 82250 -27400 82280
rect -27600 82050 -27590 82250
rect -27520 82050 -27480 82250
rect -27410 82050 -27400 82250
rect -27600 82020 -27400 82050
rect -27100 82250 -26900 82280
rect -27100 82050 -27090 82250
rect -27020 82050 -26980 82250
rect -26910 82050 -26900 82250
rect -27100 82020 -26900 82050
rect -26600 82250 -26400 82280
rect -26600 82050 -26590 82250
rect -26520 82050 -26480 82250
rect -26410 82050 -26400 82250
rect -26600 82020 -26400 82050
rect -26100 82250 -25900 82280
rect -26100 82050 -26090 82250
rect -26020 82050 -25980 82250
rect -25910 82050 -25900 82250
rect -26100 82020 -25900 82050
rect -25600 82250 -25400 82280
rect -25600 82050 -25590 82250
rect -25520 82050 -25480 82250
rect -25410 82050 -25400 82250
rect -25600 82020 -25400 82050
rect -25100 82250 -24900 82280
rect -25100 82050 -25090 82250
rect -25020 82050 -24980 82250
rect -24910 82050 -24900 82250
rect -25100 82020 -24900 82050
rect -24600 82250 -24400 82280
rect -24600 82050 -24590 82250
rect -24520 82050 -24480 82250
rect -24410 82050 -24400 82250
rect -24600 82020 -24400 82050
rect -24100 82250 -23900 82280
rect -24100 82050 -24090 82250
rect -24020 82050 -23980 82250
rect -23910 82050 -23900 82250
rect -24100 82020 -23900 82050
rect -23600 82250 -23400 82280
rect -23600 82050 -23590 82250
rect -23520 82050 -23480 82250
rect -23410 82050 -23400 82250
rect -23600 82020 -23400 82050
rect -23100 82250 -22900 82280
rect -23100 82050 -23090 82250
rect -23020 82050 -22980 82250
rect -22910 82050 -22900 82250
rect -23100 82020 -22900 82050
rect -22600 82250 -22400 82280
rect -22600 82050 -22590 82250
rect -22520 82050 -22480 82250
rect -22410 82050 -22400 82250
rect -22600 82020 -22400 82050
rect -22100 82250 -21900 82280
rect -22100 82050 -22090 82250
rect -22020 82050 -21980 82250
rect -21910 82050 -21900 82250
rect -22100 82020 -21900 82050
rect -21600 82250 -21400 82280
rect -21600 82050 -21590 82250
rect -21520 82050 -21480 82250
rect -21410 82050 -21400 82250
rect -21600 82020 -21400 82050
rect -21100 82250 -20900 82280
rect -21100 82050 -21090 82250
rect -21020 82050 -20980 82250
rect -20910 82050 -20900 82250
rect -21100 82020 -20900 82050
rect -20600 82250 -20400 82280
rect -20600 82050 -20590 82250
rect -20520 82050 -20480 82250
rect -20410 82050 -20400 82250
rect -20600 82020 -20400 82050
rect -20100 82250 -19900 82280
rect -20100 82050 -20090 82250
rect -20020 82050 -19980 82250
rect -19910 82050 -19900 82250
rect -20100 82020 -19900 82050
rect -19600 82250 -19400 82280
rect -19600 82050 -19590 82250
rect -19520 82050 -19480 82250
rect -19410 82050 -19400 82250
rect -19600 82020 -19400 82050
rect -19100 82250 -18900 82280
rect -19100 82050 -19090 82250
rect -19020 82050 -18980 82250
rect -18910 82050 -18900 82250
rect -19100 82020 -18900 82050
rect -18600 82250 -18400 82280
rect -18600 82050 -18590 82250
rect -18520 82050 -18480 82250
rect -18410 82050 -18400 82250
rect -18600 82020 -18400 82050
rect -18100 82250 -17900 82280
rect -18100 82050 -18090 82250
rect -18020 82050 -17980 82250
rect -17910 82050 -17900 82250
rect -18100 82020 -17900 82050
rect -17600 82250 -17400 82280
rect -17600 82050 -17590 82250
rect -17520 82050 -17480 82250
rect -17410 82050 -17400 82250
rect -17600 82020 -17400 82050
rect -17100 82250 -16900 82280
rect -17100 82050 -17090 82250
rect -17020 82050 -16980 82250
rect -16910 82050 -16900 82250
rect -17100 82020 -16900 82050
rect -16600 82250 -16400 82280
rect -16600 82050 -16590 82250
rect -16520 82050 -16480 82250
rect -16410 82050 -16400 82250
rect -16600 82020 -16400 82050
rect -16100 82250 -15900 82280
rect -16100 82050 -16090 82250
rect -16020 82050 -15980 82250
rect -15910 82050 -15900 82250
rect -16100 82020 -15900 82050
rect -15600 82250 -15400 82280
rect -15600 82050 -15590 82250
rect -15520 82050 -15480 82250
rect -15410 82050 -15400 82250
rect -15600 82020 -15400 82050
rect -15100 82250 -14900 82280
rect -15100 82050 -15090 82250
rect -15020 82050 -14980 82250
rect -14910 82050 -14900 82250
rect -15100 82020 -14900 82050
rect -14600 82250 -14400 82280
rect -14600 82050 -14590 82250
rect -14520 82050 -14480 82250
rect -14410 82050 -14400 82250
rect -14600 82020 -14400 82050
rect -14100 82250 -13900 82280
rect -14100 82050 -14090 82250
rect -14020 82050 -13980 82250
rect -13910 82050 -13900 82250
rect -14100 82020 -13900 82050
rect -13600 82250 -13400 82280
rect -13600 82050 -13590 82250
rect -13520 82050 -13480 82250
rect -13410 82050 -13400 82250
rect -13600 82020 -13400 82050
rect -13100 82250 -12900 82280
rect -13100 82050 -13090 82250
rect -13020 82050 -12980 82250
rect -12910 82050 -12900 82250
rect -13100 82020 -12900 82050
rect -12600 82250 -12400 82280
rect -12600 82050 -12590 82250
rect -12520 82050 -12480 82250
rect -12410 82050 -12400 82250
rect -12600 82020 -12400 82050
rect -12100 82250 -11900 82280
rect -12100 82050 -12090 82250
rect -12020 82050 -11980 82250
rect -11910 82050 -11900 82250
rect -12100 82020 -11900 82050
rect -11600 82250 -11400 82280
rect -11600 82050 -11590 82250
rect -11520 82050 -11480 82250
rect -11410 82050 -11400 82250
rect -11600 82020 -11400 82050
rect -11100 82250 -10900 82280
rect -11100 82050 -11090 82250
rect -11020 82050 -10980 82250
rect -10910 82050 -10900 82250
rect -11100 82020 -10900 82050
rect -10600 82250 -10400 82280
rect -10600 82050 -10590 82250
rect -10520 82050 -10480 82250
rect -10410 82050 -10400 82250
rect -10600 82020 -10400 82050
rect -10100 82250 -9900 82280
rect -10100 82050 -10090 82250
rect -10020 82050 -9980 82250
rect -9910 82050 -9900 82250
rect -10100 82020 -9900 82050
rect -9600 82250 -9400 82280
rect -9600 82050 -9590 82250
rect -9520 82050 -9480 82250
rect -9410 82050 -9400 82250
rect -9600 82020 -9400 82050
rect -9100 82250 -8900 82280
rect -9100 82050 -9090 82250
rect -9020 82050 -8980 82250
rect -8910 82050 -8900 82250
rect -9100 82020 -8900 82050
rect -8600 82250 -8400 82280
rect -8600 82050 -8590 82250
rect -8520 82050 -8480 82250
rect -8410 82050 -8400 82250
rect -8600 82020 -8400 82050
rect -8100 82250 -7900 82280
rect -8100 82050 -8090 82250
rect -8020 82050 -7980 82250
rect -7910 82050 -7900 82250
rect -8100 82020 -7900 82050
rect -7600 82250 -7400 82280
rect -7600 82050 -7590 82250
rect -7520 82050 -7480 82250
rect -7410 82050 -7400 82250
rect -7600 82020 -7400 82050
rect -7100 82250 -6900 82280
rect -7100 82050 -7090 82250
rect -7020 82050 -6980 82250
rect -6910 82050 -6900 82250
rect -7100 82020 -6900 82050
rect -6600 82250 -6400 82280
rect -6600 82050 -6590 82250
rect -6520 82050 -6480 82250
rect -6410 82050 -6400 82250
rect -6600 82020 -6400 82050
rect -6100 82250 -5900 82280
rect -6100 82050 -6090 82250
rect -6020 82050 -5980 82250
rect -5910 82050 -5900 82250
rect -6100 82020 -5900 82050
rect -5600 82250 -5400 82280
rect -5600 82050 -5590 82250
rect -5520 82050 -5480 82250
rect -5410 82050 -5400 82250
rect -5600 82020 -5400 82050
rect -5100 82250 -4900 82280
rect -5100 82050 -5090 82250
rect -5020 82050 -4980 82250
rect -4910 82050 -4900 82250
rect -5100 82020 -4900 82050
rect -4600 82250 -4400 82280
rect -4600 82050 -4590 82250
rect -4520 82050 -4480 82250
rect -4410 82050 -4400 82250
rect -4600 82020 -4400 82050
rect -4100 82250 -3900 82280
rect -4100 82050 -4090 82250
rect -4020 82050 -3980 82250
rect -3910 82050 -3900 82250
rect -4100 82020 -3900 82050
rect -3600 82250 -3400 82280
rect -3600 82050 -3590 82250
rect -3520 82050 -3480 82250
rect -3410 82050 -3400 82250
rect -3600 82020 -3400 82050
rect -3100 82250 -2900 82280
rect -3100 82050 -3090 82250
rect -3020 82050 -2980 82250
rect -2910 82050 -2900 82250
rect -3100 82020 -2900 82050
rect -2600 82250 -2400 82280
rect -2600 82050 -2590 82250
rect -2520 82050 -2480 82250
rect -2410 82050 -2400 82250
rect -2600 82020 -2400 82050
rect -2100 82250 -1900 82280
rect -2100 82050 -2090 82250
rect -2020 82050 -1980 82250
rect -1910 82050 -1900 82250
rect -2100 82020 -1900 82050
rect -1600 82250 -1400 82280
rect -1600 82050 -1590 82250
rect -1520 82050 -1480 82250
rect -1410 82050 -1400 82250
rect -1600 82020 -1400 82050
rect -1100 82250 -900 82280
rect -1100 82050 -1090 82250
rect -1020 82050 -980 82250
rect -910 82050 -900 82250
rect -1100 82020 -900 82050
rect -600 82250 -400 82280
rect -600 82050 -590 82250
rect -520 82050 -480 82250
rect -410 82050 -400 82250
rect -600 82020 -400 82050
rect -100 82250 100 82280
rect -100 82050 -90 82250
rect -20 82050 20 82250
rect 90 82050 100 82250
rect -100 82020 100 82050
rect 400 82250 600 82280
rect 400 82050 410 82250
rect 480 82050 520 82250
rect 590 82050 600 82250
rect 400 82020 600 82050
rect 900 82250 1100 82280
rect 900 82050 910 82250
rect 980 82050 1020 82250
rect 1090 82050 1100 82250
rect 900 82020 1100 82050
rect 1400 82250 1600 82280
rect 1400 82050 1410 82250
rect 1480 82050 1520 82250
rect 1590 82050 1600 82250
rect 1400 82020 1600 82050
rect 1900 82250 2100 82280
rect 1900 82050 1910 82250
rect 1980 82050 2020 82250
rect 2090 82050 2100 82250
rect 1900 82020 2100 82050
rect 2400 82250 2600 82280
rect 2400 82050 2410 82250
rect 2480 82050 2520 82250
rect 2590 82050 2600 82250
rect 2400 82020 2600 82050
rect 2900 82250 3100 82280
rect 2900 82050 2910 82250
rect 2980 82050 3020 82250
rect 3090 82050 3100 82250
rect 2900 82020 3100 82050
rect 3400 82250 3600 82280
rect 3400 82050 3410 82250
rect 3480 82050 3520 82250
rect 3590 82050 3600 82250
rect 3400 82020 3600 82050
rect 3900 82250 4100 82280
rect 3900 82050 3910 82250
rect 3980 82050 4020 82250
rect 4090 82050 4100 82250
rect 3900 82020 4100 82050
rect 4400 82250 4600 82280
rect 4400 82050 4410 82250
rect 4480 82050 4520 82250
rect 4590 82050 4600 82250
rect 4400 82020 4600 82050
rect 4900 82250 5100 82280
rect 4900 82050 4910 82250
rect 4980 82050 5020 82250
rect 5090 82050 5100 82250
rect 4900 82020 5100 82050
rect 5400 82250 5600 82280
rect 5400 82050 5410 82250
rect 5480 82050 5520 82250
rect 5590 82050 5600 82250
rect 5400 82020 5600 82050
rect 5900 82250 6100 82280
rect 5900 82050 5910 82250
rect 5980 82050 6020 82250
rect 6090 82050 6100 82250
rect 5900 82020 6100 82050
rect 6400 82250 6600 82280
rect 6400 82050 6410 82250
rect 6480 82050 6520 82250
rect 6590 82050 6600 82250
rect 6400 82020 6600 82050
rect 6900 82250 7100 82280
rect 6900 82050 6910 82250
rect 6980 82050 7020 82250
rect 7090 82050 7100 82250
rect 6900 82020 7100 82050
rect 7400 82250 7600 82280
rect 7400 82050 7410 82250
rect 7480 82050 7520 82250
rect 7590 82050 7600 82250
rect 7400 82020 7600 82050
rect 7900 82250 8100 82280
rect 7900 82050 7910 82250
rect 7980 82050 8020 82250
rect 8090 82050 8100 82250
rect 7900 82020 8100 82050
rect 8400 82250 8600 82280
rect 8400 82050 8410 82250
rect 8480 82050 8520 82250
rect 8590 82050 8600 82250
rect 8400 82020 8600 82050
rect 8900 82250 9100 82280
rect 8900 82050 8910 82250
rect 8980 82050 9020 82250
rect 9090 82050 9100 82250
rect 8900 82020 9100 82050
rect 9400 82250 9600 82280
rect 9400 82050 9410 82250
rect 9480 82050 9520 82250
rect 9590 82050 9600 82250
rect 9400 82020 9600 82050
rect 9900 82250 10100 82280
rect 9900 82050 9910 82250
rect 9980 82050 10020 82250
rect 10090 82050 10100 82250
rect 9900 82020 10100 82050
rect 10400 82250 10600 82280
rect 10400 82050 10410 82250
rect 10480 82050 10520 82250
rect 10590 82050 10600 82250
rect 10400 82020 10600 82050
rect 10900 82250 11100 82280
rect 10900 82050 10910 82250
rect 10980 82050 11020 82250
rect 11090 82050 11100 82250
rect 10900 82020 11100 82050
rect 11400 82250 11600 82280
rect 11400 82050 11410 82250
rect 11480 82050 11520 82250
rect 11590 82050 11600 82250
rect 11400 82020 11600 82050
rect 11900 82250 12100 82280
rect 11900 82050 11910 82250
rect 11980 82050 12020 82250
rect 12090 82050 12100 82250
rect 11900 82020 12100 82050
rect 12400 82250 12600 82280
rect 12400 82050 12410 82250
rect 12480 82050 12520 82250
rect 12590 82050 12600 82250
rect 12400 82020 12600 82050
rect 12900 82250 13100 82280
rect 12900 82050 12910 82250
rect 12980 82050 13020 82250
rect 13090 82050 13100 82250
rect 12900 82020 13100 82050
rect 13400 82250 13600 82280
rect 13400 82050 13410 82250
rect 13480 82050 13520 82250
rect 13590 82050 13600 82250
rect 13400 82020 13600 82050
rect 13900 82250 14100 82280
rect 13900 82050 13910 82250
rect 13980 82050 14020 82250
rect 14090 82050 14100 82250
rect 13900 82020 14100 82050
rect 14400 82250 14600 82280
rect 14400 82050 14410 82250
rect 14480 82050 14520 82250
rect 14590 82050 14600 82250
rect 14400 82020 14600 82050
rect 14900 82250 15100 82280
rect 14900 82050 14910 82250
rect 14980 82050 15020 82250
rect 15090 82050 15100 82250
rect 14900 82020 15100 82050
rect 15400 82250 15600 82280
rect 15400 82050 15410 82250
rect 15480 82050 15520 82250
rect 15590 82050 15600 82250
rect 15400 82020 15600 82050
rect 15900 82250 16100 82280
rect 15900 82050 15910 82250
rect 15980 82050 16020 82250
rect 16090 82050 16100 82250
rect 15900 82020 16100 82050
rect 16400 82250 16600 82280
rect 16400 82050 16410 82250
rect 16480 82050 16520 82250
rect 16590 82050 16600 82250
rect 16400 82020 16600 82050
rect 16900 82250 17100 82280
rect 16900 82050 16910 82250
rect 16980 82050 17020 82250
rect 17090 82050 17100 82250
rect 16900 82020 17100 82050
rect 17400 82250 17600 82280
rect 17400 82050 17410 82250
rect 17480 82050 17520 82250
rect 17590 82050 17600 82250
rect 17400 82020 17600 82050
rect 17900 82250 18100 82280
rect 17900 82050 17910 82250
rect 17980 82050 18020 82250
rect 18090 82050 18100 82250
rect 17900 82020 18100 82050
rect 18400 82250 18600 82280
rect 18400 82050 18410 82250
rect 18480 82050 18520 82250
rect 18590 82050 18600 82250
rect 18400 82020 18600 82050
rect 18900 82250 19100 82280
rect 18900 82050 18910 82250
rect 18980 82050 19020 82250
rect 19090 82050 19100 82250
rect 18900 82020 19100 82050
rect 19400 82250 19600 82280
rect 19400 82050 19410 82250
rect 19480 82050 19520 82250
rect 19590 82050 19600 82250
rect 19400 82020 19600 82050
rect 19900 82250 20100 82280
rect 19900 82050 19910 82250
rect 19980 82050 20020 82250
rect 20090 82050 20100 82250
rect 19900 82020 20100 82050
rect 20400 82250 20600 82280
rect 20400 82050 20410 82250
rect 20480 82050 20520 82250
rect 20590 82050 20600 82250
rect 20400 82020 20600 82050
rect 20900 82250 21100 82280
rect 20900 82050 20910 82250
rect 20980 82050 21020 82250
rect 21090 82050 21100 82250
rect 20900 82020 21100 82050
rect 21400 82250 21600 82280
rect 21400 82050 21410 82250
rect 21480 82050 21520 82250
rect 21590 82050 21600 82250
rect 21400 82020 21600 82050
rect 21900 82250 22100 82280
rect 21900 82050 21910 82250
rect 21980 82050 22020 82250
rect 22090 82050 22100 82250
rect 21900 82020 22100 82050
rect 22400 82250 22600 82280
rect 22400 82050 22410 82250
rect 22480 82050 22520 82250
rect 22590 82050 22600 82250
rect 22400 82020 22600 82050
rect 22900 82250 23100 82280
rect 22900 82050 22910 82250
rect 22980 82050 23020 82250
rect 23090 82050 23100 82250
rect 22900 82020 23100 82050
rect 23400 82250 23600 82280
rect 23400 82050 23410 82250
rect 23480 82050 23520 82250
rect 23590 82050 23600 82250
rect 23400 82020 23600 82050
rect 23900 82250 24100 82280
rect 23900 82050 23910 82250
rect 23980 82050 24020 82250
rect 24090 82050 24100 82250
rect 23900 82020 24100 82050
rect 24400 82250 24600 82280
rect 24400 82050 24410 82250
rect 24480 82050 24520 82250
rect 24590 82050 24600 82250
rect 24400 82020 24600 82050
rect 24900 82250 25100 82280
rect 24900 82050 24910 82250
rect 24980 82050 25020 82250
rect 25090 82050 25100 82250
rect 24900 82020 25100 82050
rect 25400 82250 25600 82280
rect 25400 82050 25410 82250
rect 25480 82050 25520 82250
rect 25590 82050 25600 82250
rect 25400 82020 25600 82050
rect 25900 82250 26100 82280
rect 25900 82050 25910 82250
rect 25980 82050 26020 82250
rect 26090 82050 26100 82250
rect 25900 82020 26100 82050
rect 26400 82250 26600 82280
rect 26400 82050 26410 82250
rect 26480 82050 26520 82250
rect 26590 82050 26600 82250
rect 26400 82020 26600 82050
rect 26900 82250 27100 82280
rect 26900 82050 26910 82250
rect 26980 82050 27020 82250
rect 27090 82050 27100 82250
rect 26900 82020 27100 82050
rect 27400 82250 27600 82280
rect 27400 82050 27410 82250
rect 27480 82050 27520 82250
rect 27590 82050 27600 82250
rect 27400 82020 27600 82050
rect 27900 82250 28100 82280
rect 27900 82050 27910 82250
rect 27980 82050 28020 82250
rect 28090 82050 28100 82250
rect 27900 82020 28100 82050
rect 28400 82250 28600 82280
rect 28400 82050 28410 82250
rect 28480 82050 28520 82250
rect 28590 82050 28600 82250
rect 28400 82020 28600 82050
rect 28900 82250 29100 82280
rect 28900 82050 28910 82250
rect 28980 82050 29020 82250
rect 29090 82050 29100 82250
rect 28900 82020 29100 82050
rect 29400 82250 29600 82280
rect 29400 82050 29410 82250
rect 29480 82050 29520 82250
rect 29590 82050 29600 82250
rect 29400 82020 29600 82050
rect 29900 82250 30100 82280
rect 29900 82050 29910 82250
rect 29980 82050 30020 82250
rect 30090 82050 30100 82250
rect 29900 82020 30100 82050
rect 30400 82250 30600 82280
rect 30400 82050 30410 82250
rect 30480 82050 30520 82250
rect 30590 82050 30600 82250
rect 30400 82020 30600 82050
rect 30900 82250 31100 82280
rect 30900 82050 30910 82250
rect 30980 82050 31020 82250
rect 31090 82050 31100 82250
rect 30900 82020 31100 82050
rect 31400 82250 31600 82280
rect 31400 82050 31410 82250
rect 31480 82050 31520 82250
rect 31590 82050 31600 82250
rect 31400 82020 31600 82050
rect 31900 82250 32100 82280
rect 31900 82050 31910 82250
rect 31980 82050 32020 82250
rect 32090 82050 32100 82250
rect 31900 82020 32100 82050
rect 32400 82250 32600 82280
rect 32400 82050 32410 82250
rect 32480 82050 32520 82250
rect 32590 82050 32600 82250
rect 32400 82020 32600 82050
rect 32900 82250 33100 82280
rect 32900 82050 32910 82250
rect 32980 82050 33020 82250
rect 33090 82050 33100 82250
rect 32900 82020 33100 82050
rect 33400 82250 33600 82280
rect 33400 82050 33410 82250
rect 33480 82050 33520 82250
rect 33590 82050 33600 82250
rect 33400 82020 33600 82050
rect 33900 82250 34100 82280
rect 33900 82050 33910 82250
rect 33980 82050 34020 82250
rect 34090 82050 34100 82250
rect 33900 82020 34100 82050
rect 34400 82250 34600 82280
rect 34400 82050 34410 82250
rect 34480 82050 34520 82250
rect 34590 82050 34600 82250
rect 34400 82020 34600 82050
rect 34900 82250 35100 82280
rect 34900 82050 34910 82250
rect 34980 82050 35020 82250
rect 35090 82050 35100 82250
rect 34900 82020 35100 82050
rect 35400 82250 35600 82280
rect 35400 82050 35410 82250
rect 35480 82050 35520 82250
rect 35590 82050 35600 82250
rect 35400 82020 35600 82050
rect 35900 82250 36100 82280
rect 35900 82050 35910 82250
rect 35980 82050 36020 82250
rect 36090 82050 36100 82250
rect 35900 82020 36100 82050
rect 36400 82250 36600 82280
rect 36400 82050 36410 82250
rect 36480 82050 36520 82250
rect 36590 82050 36600 82250
rect 36400 82020 36600 82050
rect 36900 82250 37100 82280
rect 36900 82050 36910 82250
rect 36980 82050 37020 82250
rect 37090 82050 37100 82250
rect 36900 82020 37100 82050
rect 37400 82250 37600 82280
rect 37400 82050 37410 82250
rect 37480 82050 37520 82250
rect 37590 82050 37600 82250
rect 37400 82020 37600 82050
rect 37900 82250 38100 82280
rect 37900 82050 37910 82250
rect 37980 82050 38020 82250
rect 38090 82050 38100 82250
rect 37900 82020 38100 82050
rect 38400 82250 38600 82280
rect 38400 82050 38410 82250
rect 38480 82050 38520 82250
rect 38590 82050 38600 82250
rect 38400 82020 38600 82050
rect 38900 82250 39100 82280
rect 38900 82050 38910 82250
rect 38980 82050 39020 82250
rect 39090 82050 39100 82250
rect 38900 82020 39100 82050
rect 39400 82250 39600 82280
rect 39400 82050 39410 82250
rect 39480 82050 39520 82250
rect 39590 82050 39600 82250
rect 39400 82020 39600 82050
rect 39900 82250 40100 82280
rect 39900 82050 39910 82250
rect 39980 82050 40020 82250
rect 40090 82050 40100 82250
rect 39900 82020 40100 82050
rect 40400 82250 40600 82280
rect 40400 82050 40410 82250
rect 40480 82050 40520 82250
rect 40590 82050 40600 82250
rect 40400 82020 40600 82050
rect 40900 82250 41100 82280
rect 40900 82050 40910 82250
rect 40980 82050 41020 82250
rect 41090 82050 41100 82250
rect 40900 82020 41100 82050
rect 41400 82250 41600 82280
rect 41400 82050 41410 82250
rect 41480 82050 41520 82250
rect 41590 82050 41600 82250
rect 41400 82020 41600 82050
rect 41900 82250 42100 82280
rect 41900 82050 41910 82250
rect 41980 82050 42020 82250
rect 42090 82050 42100 82250
rect 41900 82020 42100 82050
rect 42400 82250 42600 82280
rect 42400 82050 42410 82250
rect 42480 82050 42520 82250
rect 42590 82050 42600 82250
rect 42400 82020 42600 82050
rect 42900 82250 43100 82280
rect 42900 82050 42910 82250
rect 42980 82050 43020 82250
rect 43090 82050 43100 82250
rect 42900 82020 43100 82050
rect 43400 82250 43600 82280
rect 43400 82050 43410 82250
rect 43480 82050 43520 82250
rect 43590 82050 43600 82250
rect 43400 82020 43600 82050
rect 43900 82250 44100 82280
rect 43900 82050 43910 82250
rect 43980 82050 44020 82250
rect 44090 82050 44100 82250
rect 43900 82020 44100 82050
rect 44400 82250 44600 82280
rect 44400 82050 44410 82250
rect 44480 82050 44520 82250
rect 44590 82050 44600 82250
rect 44400 82020 44600 82050
rect 44900 82250 45100 82280
rect 44900 82050 44910 82250
rect 44980 82050 45020 82250
rect 45090 82050 45100 82250
rect 44900 82020 45100 82050
rect 45400 82250 45600 82280
rect 45400 82050 45410 82250
rect 45480 82050 45520 82250
rect 45590 82050 45600 82250
rect 45400 82020 45600 82050
rect 45900 82250 46100 82280
rect 45900 82050 45910 82250
rect 45980 82050 46020 82250
rect 46090 82050 46100 82250
rect 45900 82020 46100 82050
rect 46400 82250 46600 82280
rect 46400 82050 46410 82250
rect 46480 82050 46520 82250
rect 46590 82050 46600 82250
rect 46400 82020 46600 82050
rect 46900 82250 47100 82280
rect 46900 82050 46910 82250
rect 46980 82050 47020 82250
rect 47090 82050 47100 82250
rect 46900 82020 47100 82050
rect 47400 82250 47600 82280
rect 47400 82050 47410 82250
rect 47480 82050 47520 82250
rect 47590 82050 47600 82250
rect 47400 82020 47600 82050
rect 47900 82250 48100 82280
rect 47900 82050 47910 82250
rect 47980 82050 48020 82250
rect 48090 82050 48100 82250
rect 47900 82020 48100 82050
rect 48400 82250 48600 82280
rect 48400 82050 48410 82250
rect 48480 82050 48520 82250
rect 48590 82050 48600 82250
rect 48400 82020 48600 82050
rect 48900 82250 49100 82280
rect 48900 82050 48910 82250
rect 48980 82050 49020 82250
rect 49090 82050 49100 82250
rect 48900 82020 49100 82050
rect 49400 82250 49600 82280
rect 49400 82050 49410 82250
rect 49480 82050 49520 82250
rect 49590 82050 49600 82250
rect 49400 82020 49600 82050
rect 49900 82250 50100 82280
rect 49900 82050 49910 82250
rect 49980 82050 50020 82250
rect 50090 82050 50100 82250
rect 49900 82020 50100 82050
rect 50400 82250 50600 82280
rect 50400 82050 50410 82250
rect 50480 82050 50520 82250
rect 50590 82050 50600 82250
rect 50400 82020 50600 82050
rect 50900 82250 51100 82280
rect 50900 82050 50910 82250
rect 50980 82050 51020 82250
rect 51090 82050 51100 82250
rect 50900 82020 51100 82050
rect 51400 82250 51600 82280
rect 51400 82050 51410 82250
rect 51480 82050 51520 82250
rect 51590 82050 51600 82250
rect 51400 82020 51600 82050
rect 51900 82250 52100 82280
rect 51900 82050 51910 82250
rect 51980 82050 52020 82250
rect 52090 82050 52100 82250
rect 51900 82020 52100 82050
rect 52400 82250 52600 82280
rect 52400 82050 52410 82250
rect 52480 82050 52520 82250
rect 52590 82050 52600 82250
rect 52400 82020 52600 82050
rect 52900 82250 53100 82280
rect 52900 82050 52910 82250
rect 52980 82050 53020 82250
rect 53090 82050 53100 82250
rect 52900 82020 53100 82050
rect 53400 82250 53600 82280
rect 53400 82050 53410 82250
rect 53480 82050 53520 82250
rect 53590 82050 53600 82250
rect 53400 82020 53600 82050
rect 53900 82250 54100 82280
rect 53900 82050 53910 82250
rect 53980 82050 54020 82250
rect 54090 82050 54100 82250
rect 53900 82020 54100 82050
rect 54400 82250 54600 82280
rect 54400 82050 54410 82250
rect 54480 82050 54520 82250
rect 54590 82050 54600 82250
rect 54400 82020 54600 82050
rect 54900 82250 55100 82280
rect 54900 82050 54910 82250
rect 54980 82050 55020 82250
rect 55090 82050 55100 82250
rect 54900 82020 55100 82050
rect 55400 82250 55600 82280
rect 55400 82050 55410 82250
rect 55480 82050 55520 82250
rect 55590 82050 55600 82250
rect 55400 82020 55600 82050
rect 55900 82250 56100 82280
rect 55900 82050 55910 82250
rect 55980 82050 56020 82250
rect 56090 82050 56100 82250
rect 55900 82020 56100 82050
rect 56400 82250 56600 82280
rect 56400 82050 56410 82250
rect 56480 82050 56520 82250
rect 56590 82050 56600 82250
rect 56400 82020 56600 82050
rect 56900 82250 57100 82280
rect 56900 82050 56910 82250
rect 56980 82050 57020 82250
rect 57090 82050 57100 82250
rect 56900 82020 57100 82050
rect 57400 82250 57600 82280
rect 57400 82050 57410 82250
rect 57480 82050 57520 82250
rect 57590 82050 57600 82250
rect 57400 82020 57600 82050
rect 57900 82250 58100 82280
rect 57900 82050 57910 82250
rect 57980 82050 58020 82250
rect 58090 82050 58100 82250
rect 57900 82020 58100 82050
rect 58400 82250 58600 82280
rect 58400 82050 58410 82250
rect 58480 82050 58520 82250
rect 58590 82050 58600 82250
rect 58400 82020 58600 82050
rect 58900 82250 59100 82280
rect 58900 82050 58910 82250
rect 58980 82050 59020 82250
rect 59090 82050 59100 82250
rect 58900 82020 59100 82050
rect 59400 82250 59600 82280
rect 59400 82050 59410 82250
rect 59480 82050 59520 82250
rect 59590 82050 59600 82250
rect 59400 82020 59600 82050
rect 59900 82250 60100 82280
rect 59900 82050 59910 82250
rect 59980 82050 60020 82250
rect 60090 82050 60100 82250
rect 59900 82020 60100 82050
rect 60400 82250 60600 82280
rect 60400 82050 60410 82250
rect 60480 82050 60520 82250
rect 60590 82050 60600 82250
rect 60400 82020 60600 82050
rect 60900 82250 61100 82280
rect 60900 82050 60910 82250
rect 60980 82050 61020 82250
rect 61090 82050 61100 82250
rect 60900 82020 61100 82050
rect 61400 82250 61600 82280
rect 61400 82050 61410 82250
rect 61480 82050 61520 82250
rect 61590 82050 61600 82250
rect 61400 82020 61600 82050
rect 61900 82250 62100 82280
rect 61900 82050 61910 82250
rect 61980 82050 62020 82250
rect 62090 82050 62100 82250
rect 61900 82020 62100 82050
rect 62400 82250 62600 82280
rect 62400 82050 62410 82250
rect 62480 82050 62520 82250
rect 62590 82050 62600 82250
rect 62400 82020 62600 82050
rect 62900 82250 63100 82280
rect 62900 82050 62910 82250
rect 62980 82050 63020 82250
rect 63090 82050 63100 82250
rect 62900 82020 63100 82050
rect 63400 82250 63600 82280
rect 63400 82050 63410 82250
rect 63480 82050 63520 82250
rect 63590 82050 63600 82250
rect 63400 82020 63600 82050
rect 63900 82250 64100 82280
rect 63900 82050 63910 82250
rect 63980 82050 64020 82250
rect 64090 82050 64100 82250
rect 63900 82020 64100 82050
rect 64400 82250 64600 82280
rect 64400 82050 64410 82250
rect 64480 82050 64520 82250
rect 64590 82050 64600 82250
rect 64400 82020 64600 82050
rect 64900 82250 65100 82280
rect 64900 82050 64910 82250
rect 64980 82050 65020 82250
rect 65090 82050 65100 82250
rect 64900 82020 65100 82050
rect 65400 82250 65600 82280
rect 65400 82050 65410 82250
rect 65480 82050 65520 82250
rect 65590 82050 65600 82250
rect 65400 82020 65600 82050
rect 65900 82250 66100 82280
rect 65900 82050 65910 82250
rect 65980 82050 66020 82250
rect 66090 82050 66100 82250
rect 65900 82020 66100 82050
rect 66400 82250 66600 82280
rect 66400 82050 66410 82250
rect 66480 82050 66520 82250
rect 66590 82050 66600 82250
rect 66400 82020 66600 82050
rect 66900 82250 67100 82280
rect 66900 82050 66910 82250
rect 66980 82050 67020 82250
rect 67090 82050 67100 82250
rect 66900 82020 67100 82050
rect 67400 82250 67600 82280
rect 67400 82050 67410 82250
rect 67480 82050 67520 82250
rect 67590 82050 67600 82250
rect 67400 82020 67600 82050
rect 67900 82250 68100 82280
rect 67900 82050 67910 82250
rect 67980 82050 68020 82250
rect 68090 82050 68100 82250
rect 67900 82020 68100 82050
rect 68400 82250 68600 82280
rect 68400 82050 68410 82250
rect 68480 82050 68520 82250
rect 68590 82050 68600 82250
rect 68400 82020 68600 82050
rect 68900 82250 69100 82280
rect 68900 82050 68910 82250
rect 68980 82050 69020 82250
rect 69090 82050 69100 82250
rect 68900 82020 69100 82050
rect 69400 82250 69600 82280
rect 69400 82050 69410 82250
rect 69480 82050 69520 82250
rect 69590 82050 69600 82250
rect 69400 82020 69600 82050
rect 69900 82250 70100 82280
rect 69900 82050 69910 82250
rect 69980 82050 70020 82250
rect 70090 82050 70100 82250
rect 69900 82020 70100 82050
rect 70400 82250 70600 82280
rect 70400 82050 70410 82250
rect 70480 82050 70520 82250
rect 70590 82050 70600 82250
rect 70400 82020 70600 82050
rect 70900 82250 71100 82280
rect 70900 82050 70910 82250
rect 70980 82050 71020 82250
rect 71090 82050 71100 82250
rect 70900 82020 71100 82050
rect 71400 82250 71600 82280
rect 71400 82050 71410 82250
rect 71480 82050 71520 82250
rect 71590 82050 71600 82250
rect 71400 82020 71600 82050
rect 71900 82250 72100 82280
rect 71900 82050 71910 82250
rect 71980 82050 72020 82250
rect 72090 82050 72100 82250
rect 71900 82020 72100 82050
rect 72400 82250 72600 82280
rect 72400 82050 72410 82250
rect 72480 82050 72520 82250
rect 72590 82050 72600 82250
rect 72400 82020 72600 82050
rect 72900 82250 73100 82280
rect 72900 82050 72910 82250
rect 72980 82050 73020 82250
rect 73090 82050 73100 82250
rect 72900 82020 73100 82050
rect 73400 82250 73600 82280
rect 73400 82050 73410 82250
rect 73480 82050 73520 82250
rect 73590 82050 73600 82250
rect 73400 82020 73600 82050
rect 73900 82250 74100 82280
rect 73900 82050 73910 82250
rect 73980 82050 74020 82250
rect 74090 82050 74100 82250
rect 73900 82020 74100 82050
rect 74400 82250 74600 82280
rect 74400 82050 74410 82250
rect 74480 82050 74520 82250
rect 74590 82050 74600 82250
rect 74400 82020 74600 82050
rect 74900 82250 75100 82280
rect 74900 82050 74910 82250
rect 74980 82050 75020 82250
rect 75090 82050 75100 82250
rect 74900 82020 75100 82050
rect 75400 82250 75600 82280
rect 75400 82050 75410 82250
rect 75480 82050 75520 82250
rect 75590 82050 75600 82250
rect 75400 82020 75600 82050
rect 75900 82250 76100 82280
rect 75900 82050 75910 82250
rect 75980 82050 76020 82250
rect 76090 82050 76100 82250
rect 75900 82020 76100 82050
rect 76400 82250 76600 82280
rect 76400 82050 76410 82250
rect 76480 82050 76520 82250
rect 76590 82050 76600 82250
rect 76400 82020 76600 82050
rect 76900 82250 77100 82280
rect 76900 82050 76910 82250
rect 76980 82050 77020 82250
rect 77090 82050 77100 82250
rect 76900 82020 77100 82050
rect 77400 82250 77600 82280
rect 77400 82050 77410 82250
rect 77480 82050 77520 82250
rect 77590 82050 77600 82250
rect 77400 82020 77600 82050
rect 77900 82250 78100 82280
rect 77900 82050 77910 82250
rect 77980 82050 78020 82250
rect 78090 82050 78100 82250
rect 77900 82020 78100 82050
rect 78400 82250 78600 82280
rect 78400 82050 78410 82250
rect 78480 82050 78520 82250
rect 78590 82050 78600 82250
rect 78400 82020 78600 82050
rect 78900 82250 79100 82280
rect 78900 82050 78910 82250
rect 78980 82050 79020 82250
rect 79090 82050 79100 82250
rect 78900 82020 79100 82050
rect 79400 82250 79600 82280
rect 79400 82050 79410 82250
rect 79480 82050 79520 82250
rect 79590 82050 79600 82250
rect 79400 82020 79600 82050
rect 79900 82250 80100 82280
rect 79900 82050 79910 82250
rect 79980 82050 80020 82250
rect 80090 82050 80100 82250
rect 79900 82020 80100 82050
rect 80400 82250 80600 82280
rect 80400 82050 80410 82250
rect 80480 82050 80520 82250
rect 80590 82050 80600 82250
rect 80400 82020 80600 82050
rect 80900 82250 81100 82280
rect 80900 82050 80910 82250
rect 80980 82050 81020 82250
rect 81090 82050 81100 82250
rect 80900 82020 81100 82050
rect 81400 82250 81600 82280
rect 81400 82050 81410 82250
rect 81480 82050 81520 82250
rect 81590 82050 81600 82250
rect 81400 82020 81600 82050
rect 81900 82250 82100 82280
rect 81900 82050 81910 82250
rect 81980 82050 82020 82250
rect 82090 82050 82100 82250
rect 81900 82020 82100 82050
rect 82400 82250 82600 82280
rect 82400 82050 82410 82250
rect 82480 82050 82520 82250
rect 82590 82050 82600 82250
rect 82400 82020 82600 82050
rect 82900 82250 83100 82280
rect 82900 82050 82910 82250
rect 82980 82050 83020 82250
rect 83090 82050 83100 82250
rect 82900 82020 83100 82050
rect 83400 82250 83600 82280
rect 83400 82050 83410 82250
rect 83480 82050 83520 82250
rect 83590 82050 83600 82250
rect 83400 82020 83600 82050
rect 83900 82250 84100 82280
rect 83900 82050 83910 82250
rect 83980 82050 84020 82250
rect 84090 82050 84100 82250
rect 83900 82020 84100 82050
rect 84400 82250 84600 82280
rect 84400 82050 84410 82250
rect 84480 82050 84520 82250
rect 84590 82050 84600 82250
rect 84400 82020 84600 82050
rect 84900 82250 85100 82280
rect 84900 82050 84910 82250
rect 84980 82050 85020 82250
rect 85090 82050 85100 82250
rect 84900 82020 85100 82050
rect 85400 82250 85600 82280
rect 85400 82050 85410 82250
rect 85480 82050 85520 82250
rect 85590 82050 85600 82250
rect 85400 82020 85600 82050
rect 85900 82250 86100 82280
rect 85900 82050 85910 82250
rect 85980 82050 86020 82250
rect 86090 82050 86100 82250
rect 85900 82020 86100 82050
rect 86400 82250 86600 82280
rect 86400 82050 86410 82250
rect 86480 82050 86520 82250
rect 86590 82050 86600 82250
rect 86400 82020 86600 82050
rect 86900 82250 87100 82280
rect 86900 82050 86910 82250
rect 86980 82050 87020 82250
rect 87090 82050 87100 82250
rect 86900 82020 87100 82050
rect 87400 82250 87600 82280
rect 87400 82050 87410 82250
rect 87480 82050 87520 82250
rect 87590 82050 87600 82250
rect 87400 82020 87600 82050
rect 87900 82250 88100 82280
rect 87900 82050 87910 82250
rect 87980 82050 88020 82250
rect 88090 82050 88100 82250
rect 87900 82020 88100 82050
rect 88400 82250 88600 82280
rect 88400 82050 88410 82250
rect 88480 82050 88520 82250
rect 88590 82050 88600 82250
rect 88400 82020 88600 82050
rect 88900 82250 89100 82280
rect 88900 82050 88910 82250
rect 88980 82050 89020 82250
rect 89090 82050 89100 82250
rect 88900 82020 89100 82050
rect 89400 82250 89600 82280
rect 89400 82050 89410 82250
rect 89480 82050 89520 82250
rect 89590 82050 89600 82250
rect 89400 82020 89600 82050
rect 89900 82250 90100 82280
rect 89900 82050 89910 82250
rect 89980 82050 90020 82250
rect 90090 82050 90100 82250
rect 89900 82020 90100 82050
rect 90400 82250 90600 82280
rect 90400 82050 90410 82250
rect 90480 82050 90520 82250
rect 90590 82050 90600 82250
rect 90400 82020 90600 82050
rect 90900 82250 91100 82280
rect 90900 82050 90910 82250
rect 90980 82050 91020 82250
rect 91090 82050 91100 82250
rect 90900 82020 91100 82050
rect 91400 82250 91600 82280
rect 91400 82050 91410 82250
rect 91480 82050 91520 82250
rect 91590 82050 91600 82250
rect 91400 82020 91600 82050
rect 91900 82250 92100 82280
rect 91900 82050 91910 82250
rect 91980 82050 92020 82250
rect 92090 82050 92100 82250
rect 91900 82020 92100 82050
rect 92400 82250 92600 82280
rect 92400 82050 92410 82250
rect 92480 82050 92520 82250
rect 92590 82050 92600 82250
rect 92400 82020 92600 82050
rect 92900 82250 93100 82280
rect 92900 82050 92910 82250
rect 92980 82050 93020 82250
rect 93090 82050 93100 82250
rect 92900 82020 93100 82050
rect 93400 82250 93600 82280
rect 93400 82050 93410 82250
rect 93480 82050 93520 82250
rect 93590 82050 93600 82250
rect 93400 82020 93600 82050
rect 93900 82250 94100 82280
rect 93900 82050 93910 82250
rect 93980 82050 94020 82250
rect 94090 82050 94100 82250
rect 93900 82020 94100 82050
rect 94400 82250 94600 82280
rect 94400 82050 94410 82250
rect 94480 82050 94520 82250
rect 94590 82050 94600 82250
rect 94400 82020 94600 82050
rect 94900 82250 95100 82280
rect 94900 82050 94910 82250
rect 94980 82050 95020 82250
rect 95090 82050 95100 82250
rect 94900 82020 95100 82050
rect 95400 82250 95600 82280
rect 95400 82050 95410 82250
rect 95480 82050 95520 82250
rect 95590 82050 95600 82250
rect 95400 82020 95600 82050
rect 95900 82250 96100 82280
rect 95900 82050 95910 82250
rect 95980 82050 96020 82250
rect 96090 82050 96100 82250
rect 95900 82020 96100 82050
rect 96400 82250 96600 82280
rect 96400 82050 96410 82250
rect 96480 82050 96520 82250
rect 96590 82050 96600 82250
rect 96400 82020 96600 82050
rect 96900 82250 97100 82280
rect 96900 82050 96910 82250
rect 96980 82050 97020 82250
rect 97090 82050 97100 82250
rect 96900 82020 97100 82050
rect 97400 82250 97600 82280
rect 97400 82050 97410 82250
rect 97480 82050 97520 82250
rect 97590 82050 97600 82250
rect 97400 82020 97600 82050
rect 97900 82250 98100 82280
rect 97900 82050 97910 82250
rect 97980 82050 98020 82250
rect 98090 82050 98100 82250
rect 97900 82020 98100 82050
rect 98400 82250 98600 82280
rect 98400 82050 98410 82250
rect 98480 82050 98520 82250
rect 98590 82050 98600 82250
rect 98400 82020 98600 82050
rect 98900 82250 99100 82280
rect 98900 82050 98910 82250
rect 98980 82050 99020 82250
rect 99090 82050 99100 82250
rect 98900 82020 99100 82050
rect 99400 82250 99600 82280
rect 99400 82050 99410 82250
rect 99480 82050 99520 82250
rect 99590 82050 99600 82250
rect 99400 82020 99600 82050
rect 99900 82250 100100 82280
rect 99900 82050 99910 82250
rect 99980 82050 100020 82250
rect 100090 82050 100100 82250
rect 99900 82020 100100 82050
rect 100400 82250 100500 82280
rect 100400 82050 100410 82250
rect 100480 82050 100500 82250
rect 100400 82020 100500 82050
rect -83500 82000 -83380 82020
rect -83120 82000 -82880 82020
rect -82620 82000 -82380 82020
rect -82120 82000 -81880 82020
rect -81620 82000 -81380 82020
rect -81120 82000 -80880 82020
rect -80620 82000 -80380 82020
rect -80120 82000 -79880 82020
rect -79620 82000 -79380 82020
rect -79120 82000 -78880 82020
rect -78620 82000 -78380 82020
rect -78120 82000 -77880 82020
rect -77620 82000 -77380 82020
rect -77120 82000 -76880 82020
rect -76620 82000 -76380 82020
rect -76120 82000 -75880 82020
rect -75620 82000 -75380 82020
rect -75120 82000 -74880 82020
rect -74620 82000 -74380 82020
rect -74120 82000 -73880 82020
rect -73620 82000 -73380 82020
rect -73120 82000 -72880 82020
rect -72620 82000 -72380 82020
rect -72120 82000 -71880 82020
rect -71620 82000 -71380 82020
rect -71120 82000 -70880 82020
rect -70620 82000 -70380 82020
rect -70120 82000 -69880 82020
rect -69620 82000 -69380 82020
rect -69120 82000 -68880 82020
rect -68620 82000 -68380 82020
rect -68120 82000 -67880 82020
rect -67620 82000 -67380 82020
rect -67120 82000 -66880 82020
rect -66620 82000 -66380 82020
rect -66120 82000 -65880 82020
rect -65620 82000 -65380 82020
rect -65120 82000 -64880 82020
rect -64620 82000 -64380 82020
rect -64120 82000 -63880 82020
rect -63620 82000 -63380 82020
rect -63120 82000 -62880 82020
rect -62620 82000 -62380 82020
rect -62120 82000 -61880 82020
rect -61620 82000 -61380 82020
rect -61120 82000 -60880 82020
rect -60620 82000 -60380 82020
rect -60120 82000 -59880 82020
rect -59620 82000 -59380 82020
rect -59120 82000 -58880 82020
rect -58620 82000 -58380 82020
rect -58120 82000 -57880 82020
rect -57620 82000 -57380 82020
rect -57120 82000 -56880 82020
rect -56620 82000 -56380 82020
rect -56120 82000 -55880 82020
rect -55620 82000 -55380 82020
rect -55120 82000 -54880 82020
rect -54620 82000 -54380 82020
rect -54120 82000 -53880 82020
rect -53620 82000 -53380 82020
rect -53120 82000 -52880 82020
rect -52620 82000 -52380 82020
rect -52120 82000 -51880 82020
rect -51620 82000 -51380 82020
rect -51120 82000 -50880 82020
rect -50620 82000 -50380 82020
rect -50120 82000 -49880 82020
rect -49620 82000 -49380 82020
rect -49120 82000 -48880 82020
rect -48620 82000 -48380 82020
rect -48120 82000 -47880 82020
rect -47620 82000 -47380 82020
rect -47120 82000 -46880 82020
rect -46620 82000 -46380 82020
rect -46120 82000 -45880 82020
rect -45620 82000 -45380 82020
rect -45120 82000 -44880 82020
rect -44620 82000 -44380 82020
rect -44120 82000 -43880 82020
rect -43620 82000 -43380 82020
rect -43120 82000 -42880 82020
rect -42620 82000 -42380 82020
rect -42120 82000 -41880 82020
rect -41620 82000 -41380 82020
rect -41120 82000 -40880 82020
rect -40620 82000 -40380 82020
rect -40120 82000 -39880 82020
rect -39620 82000 -39380 82020
rect -39120 82000 -38880 82020
rect -38620 82000 -38380 82020
rect -38120 82000 -37880 82020
rect -37620 82000 -37380 82020
rect -37120 82000 -36880 82020
rect -36620 82000 -36380 82020
rect -36120 82000 -35880 82020
rect -35620 82000 -35380 82020
rect -35120 82000 -34880 82020
rect -34620 82000 -34380 82020
rect -34120 82000 -33880 82020
rect -33620 82000 -33380 82020
rect -33120 82000 -32880 82020
rect -32620 82000 -32380 82020
rect -32120 82000 -31880 82020
rect -31620 82000 -31380 82020
rect -31120 82000 -30880 82020
rect -30620 82000 -30380 82020
rect -30120 82000 -29880 82020
rect -29620 82000 -29380 82020
rect -29120 82000 -28880 82020
rect -28620 82000 -28380 82020
rect -28120 82000 -27880 82020
rect -27620 82000 -27380 82020
rect -27120 82000 -26880 82020
rect -26620 82000 -26380 82020
rect -26120 82000 -25880 82020
rect -25620 82000 -25380 82020
rect -25120 82000 -24880 82020
rect -24620 82000 -24380 82020
rect -24120 82000 -23880 82020
rect -23620 82000 -23380 82020
rect -23120 82000 -22880 82020
rect -22620 82000 -22380 82020
rect -22120 82000 -21880 82020
rect -21620 82000 -21380 82020
rect -21120 82000 -20880 82020
rect -20620 82000 -20380 82020
rect -20120 82000 -19880 82020
rect -19620 82000 -19380 82020
rect -19120 82000 -18880 82020
rect -18620 82000 -18380 82020
rect -18120 82000 -17880 82020
rect -17620 82000 -17380 82020
rect -17120 82000 -16880 82020
rect -16620 82000 -16380 82020
rect -16120 82000 -15880 82020
rect -15620 82000 -15380 82020
rect -15120 82000 -14880 82020
rect -14620 82000 -14380 82020
rect -14120 82000 -13880 82020
rect -13620 82000 -13380 82020
rect -13120 82000 -12880 82020
rect -12620 82000 -12380 82020
rect -12120 82000 -11880 82020
rect -11620 82000 -11380 82020
rect -11120 82000 -10880 82020
rect -10620 82000 -10380 82020
rect -10120 82000 -9880 82020
rect -9620 82000 -9380 82020
rect -9120 82000 -8880 82020
rect -8620 82000 -8380 82020
rect -8120 82000 -7880 82020
rect -7620 82000 -7380 82020
rect -7120 82000 -6880 82020
rect -6620 82000 -6380 82020
rect -6120 82000 -5880 82020
rect -5620 82000 -5380 82020
rect -5120 82000 -4880 82020
rect -4620 82000 -4380 82020
rect -4120 82000 -3880 82020
rect -3620 82000 -3380 82020
rect -3120 82000 -2880 82020
rect -2620 82000 -2380 82020
rect -2120 82000 -1880 82020
rect -1620 82000 -1380 82020
rect -1120 82000 -880 82020
rect -620 82000 -380 82020
rect -120 82000 120 82020
rect 380 82000 620 82020
rect 880 82000 1120 82020
rect 1380 82000 1620 82020
rect 1880 82000 2120 82020
rect 2380 82000 2620 82020
rect 2880 82000 3120 82020
rect 3380 82000 3620 82020
rect 3880 82000 4120 82020
rect 4380 82000 4620 82020
rect 4880 82000 5120 82020
rect 5380 82000 5620 82020
rect 5880 82000 6120 82020
rect 6380 82000 6620 82020
rect 6880 82000 7120 82020
rect 7380 82000 7620 82020
rect 7880 82000 8120 82020
rect 8380 82000 8620 82020
rect 8880 82000 9120 82020
rect 9380 82000 9620 82020
rect 9880 82000 10120 82020
rect 10380 82000 10620 82020
rect 10880 82000 11120 82020
rect 11380 82000 11620 82020
rect 11880 82000 12120 82020
rect 12380 82000 12620 82020
rect 12880 82000 13120 82020
rect 13380 82000 13620 82020
rect 13880 82000 14120 82020
rect 14380 82000 14620 82020
rect 14880 82000 15120 82020
rect 15380 82000 15620 82020
rect 15880 82000 16120 82020
rect 16380 82000 16620 82020
rect 16880 82000 17120 82020
rect 17380 82000 17620 82020
rect 17880 82000 18120 82020
rect 18380 82000 18620 82020
rect 18880 82000 19120 82020
rect 19380 82000 19620 82020
rect 19880 82000 20120 82020
rect 20380 82000 20620 82020
rect 20880 82000 21120 82020
rect 21380 82000 21620 82020
rect 21880 82000 22120 82020
rect 22380 82000 22620 82020
rect 22880 82000 23120 82020
rect 23380 82000 23620 82020
rect 23880 82000 24120 82020
rect 24380 82000 24620 82020
rect 24880 82000 25120 82020
rect 25380 82000 25620 82020
rect 25880 82000 26120 82020
rect 26380 82000 26620 82020
rect 26880 82000 27120 82020
rect 27380 82000 27620 82020
rect 27880 82000 28120 82020
rect 28380 82000 28620 82020
rect 28880 82000 29120 82020
rect 29380 82000 29620 82020
rect 29880 82000 30120 82020
rect 30380 82000 30620 82020
rect 30880 82000 31120 82020
rect 31380 82000 31620 82020
rect 31880 82000 32120 82020
rect 32380 82000 32620 82020
rect 32880 82000 33120 82020
rect 33380 82000 33620 82020
rect 33880 82000 34120 82020
rect 34380 82000 34620 82020
rect 34880 82000 35120 82020
rect 35380 82000 35620 82020
rect 35880 82000 36120 82020
rect 36380 82000 36620 82020
rect 36880 82000 37120 82020
rect 37380 82000 37620 82020
rect 37880 82000 38120 82020
rect 38380 82000 38620 82020
rect 38880 82000 39120 82020
rect 39380 82000 39620 82020
rect 39880 82000 40120 82020
rect 40380 82000 40620 82020
rect 40880 82000 41120 82020
rect 41380 82000 41620 82020
rect 41880 82000 42120 82020
rect 42380 82000 42620 82020
rect 42880 82000 43120 82020
rect 43380 82000 43620 82020
rect 43880 82000 44120 82020
rect 44380 82000 44620 82020
rect 44880 82000 45120 82020
rect 45380 82000 45620 82020
rect 45880 82000 46120 82020
rect 46380 82000 46620 82020
rect 46880 82000 47120 82020
rect 47380 82000 47620 82020
rect 47880 82000 48120 82020
rect 48380 82000 48620 82020
rect 48880 82000 49120 82020
rect 49380 82000 49620 82020
rect 49880 82000 50120 82020
rect 50380 82000 50620 82020
rect 50880 82000 51120 82020
rect 51380 82000 51620 82020
rect 51880 82000 52120 82020
rect 52380 82000 52620 82020
rect 52880 82000 53120 82020
rect 53380 82000 53620 82020
rect 53880 82000 54120 82020
rect 54380 82000 54620 82020
rect 54880 82000 55120 82020
rect 55380 82000 55620 82020
rect 55880 82000 56120 82020
rect 56380 82000 56620 82020
rect 56880 82000 57120 82020
rect 57380 82000 57620 82020
rect 57880 82000 58120 82020
rect 58380 82000 58620 82020
rect 58880 82000 59120 82020
rect 59380 82000 59620 82020
rect 59880 82000 60120 82020
rect 60380 82000 60620 82020
rect 60880 82000 61120 82020
rect 61380 82000 61620 82020
rect 61880 82000 62120 82020
rect 62380 82000 62620 82020
rect 62880 82000 63120 82020
rect 63380 82000 63620 82020
rect 63880 82000 64120 82020
rect 64380 82000 64620 82020
rect 64880 82000 65120 82020
rect 65380 82000 65620 82020
rect 65880 82000 66120 82020
rect 66380 82000 66620 82020
rect 66880 82000 67120 82020
rect 67380 82000 67620 82020
rect 67880 82000 68120 82020
rect 68380 82000 68620 82020
rect 68880 82000 69120 82020
rect 69380 82000 69620 82020
rect 69880 82000 70120 82020
rect 70380 82000 70620 82020
rect 70880 82000 71120 82020
rect 71380 82000 71620 82020
rect 71880 82000 72120 82020
rect 72380 82000 72620 82020
rect 72880 82000 73120 82020
rect 73380 82000 73620 82020
rect 73880 82000 74120 82020
rect 74380 82000 74620 82020
rect 74880 82000 75120 82020
rect 75380 82000 75620 82020
rect 75880 82000 76120 82020
rect 76380 82000 76620 82020
rect 76880 82000 77120 82020
rect 77380 82000 77620 82020
rect 77880 82000 78120 82020
rect 78380 82000 78620 82020
rect 78880 82000 79120 82020
rect 79380 82000 79620 82020
rect 79880 82000 80120 82020
rect 80380 82000 80620 82020
rect 80880 82000 81120 82020
rect 81380 82000 81620 82020
rect 81880 82000 82120 82020
rect 82380 82000 82620 82020
rect 82880 82000 83120 82020
rect 83380 82000 83620 82020
rect 83880 82000 84120 82020
rect 84380 82000 84620 82020
rect 84880 82000 85120 82020
rect 85380 82000 85620 82020
rect 85880 82000 86120 82020
rect 86380 82000 86620 82020
rect 86880 82000 87120 82020
rect 87380 82000 87620 82020
rect 87880 82000 88120 82020
rect 88380 82000 88620 82020
rect 88880 82000 89120 82020
rect 89380 82000 89620 82020
rect 89880 82000 90120 82020
rect 90380 82000 90620 82020
rect 90880 82000 91120 82020
rect 91380 82000 91620 82020
rect 91880 82000 92120 82020
rect 92380 82000 92620 82020
rect 92880 82000 93120 82020
rect 93380 82000 93620 82020
rect 93880 82000 94120 82020
rect 94380 82000 94620 82020
rect 94880 82000 95120 82020
rect 95380 82000 95620 82020
rect 95880 82000 96120 82020
rect 96380 82000 96620 82020
rect 96880 82000 97120 82020
rect 97380 82000 97620 82020
rect 97880 82000 98120 82020
rect 98380 82000 98620 82020
rect 98880 82000 99120 82020
rect 99380 82000 99620 82020
rect 99880 82000 100120 82020
rect 100380 82000 100500 82020
rect -83500 81990 100500 82000
rect -83500 81920 -83350 81990
rect -83150 81920 -82850 81990
rect -82650 81920 -82350 81990
rect -82150 81920 -81850 81990
rect -81650 81920 -81350 81990
rect -81150 81920 -80850 81990
rect -80650 81920 -80350 81990
rect -80150 81920 -79850 81990
rect -79650 81920 -79350 81990
rect -79150 81920 -78850 81990
rect -78650 81920 -78350 81990
rect -78150 81920 -77850 81990
rect -77650 81920 -77350 81990
rect -77150 81920 -76850 81990
rect -76650 81920 -76350 81990
rect -76150 81920 -75850 81990
rect -75650 81920 -75350 81990
rect -75150 81920 -74850 81990
rect -74650 81920 -74350 81990
rect -74150 81920 -73850 81990
rect -73650 81920 -73350 81990
rect -73150 81920 -72850 81990
rect -72650 81920 -72350 81990
rect -72150 81920 -71850 81990
rect -71650 81920 -71350 81990
rect -71150 81920 -70850 81990
rect -70650 81920 -70350 81990
rect -70150 81920 -69850 81990
rect -69650 81920 -69350 81990
rect -69150 81920 -68850 81990
rect -68650 81920 -68350 81990
rect -68150 81920 -67850 81990
rect -67650 81920 -67350 81990
rect -67150 81920 -66850 81990
rect -66650 81920 -66350 81990
rect -66150 81920 -65850 81990
rect -65650 81920 -65350 81990
rect -65150 81920 -64850 81990
rect -64650 81920 -64350 81990
rect -64150 81920 -63850 81990
rect -63650 81920 -63350 81990
rect -63150 81920 -62850 81990
rect -62650 81920 -62350 81990
rect -62150 81920 -61850 81990
rect -61650 81920 -61350 81990
rect -61150 81920 -60850 81990
rect -60650 81920 -60350 81990
rect -60150 81920 -59850 81990
rect -59650 81920 -59350 81990
rect -59150 81920 -58850 81990
rect -58650 81920 -58350 81990
rect -58150 81920 -57850 81990
rect -57650 81920 -57350 81990
rect -57150 81920 -56850 81990
rect -56650 81920 -56350 81990
rect -56150 81920 -55850 81990
rect -55650 81920 -55350 81990
rect -55150 81920 -54850 81990
rect -54650 81920 -54350 81990
rect -54150 81920 -53850 81990
rect -53650 81920 -53350 81990
rect -53150 81920 -52850 81990
rect -52650 81920 -52350 81990
rect -52150 81920 -51850 81990
rect -51650 81920 -51350 81990
rect -51150 81920 -50850 81990
rect -50650 81920 -50350 81990
rect -50150 81920 -49850 81990
rect -49650 81920 -49350 81990
rect -49150 81920 -48850 81990
rect -48650 81920 -48350 81990
rect -48150 81920 -47850 81990
rect -47650 81920 -47350 81990
rect -47150 81920 -46850 81990
rect -46650 81920 -46350 81990
rect -46150 81920 -45850 81990
rect -45650 81920 -45350 81990
rect -45150 81920 -44850 81990
rect -44650 81920 -44350 81990
rect -44150 81920 -43850 81990
rect -43650 81920 -43350 81990
rect -43150 81920 -42850 81990
rect -42650 81920 -42350 81990
rect -42150 81920 -41850 81990
rect -41650 81920 -41350 81990
rect -41150 81920 -40850 81990
rect -40650 81920 -40350 81990
rect -40150 81920 -39850 81990
rect -39650 81920 -39350 81990
rect -39150 81920 -38850 81990
rect -38650 81920 -38350 81990
rect -38150 81920 -37850 81990
rect -37650 81920 -37350 81990
rect -37150 81920 -36850 81990
rect -36650 81920 -36350 81990
rect -36150 81920 -35850 81990
rect -35650 81920 -35350 81990
rect -35150 81920 -34850 81990
rect -34650 81920 -34350 81990
rect -34150 81920 -33850 81990
rect -33650 81920 -33350 81990
rect -33150 81920 -32850 81990
rect -32650 81920 -32350 81990
rect -32150 81920 -31850 81990
rect -31650 81920 -31350 81990
rect -31150 81920 -30850 81990
rect -30650 81920 -30350 81990
rect -30150 81920 -29850 81990
rect -29650 81920 -29350 81990
rect -29150 81920 -28850 81990
rect -28650 81920 -28350 81990
rect -28150 81920 -27850 81990
rect -27650 81920 -27350 81990
rect -27150 81920 -26850 81990
rect -26650 81920 -26350 81990
rect -26150 81920 -25850 81990
rect -25650 81920 -25350 81990
rect -25150 81920 -24850 81990
rect -24650 81920 -24350 81990
rect -24150 81920 -23850 81990
rect -23650 81920 -23350 81990
rect -23150 81920 -22850 81990
rect -22650 81920 -22350 81990
rect -22150 81920 -21850 81990
rect -21650 81920 -21350 81990
rect -21150 81920 -20850 81990
rect -20650 81920 -20350 81990
rect -20150 81920 -19850 81990
rect -19650 81920 -19350 81990
rect -19150 81920 -18850 81990
rect -18650 81920 -18350 81990
rect -18150 81920 -17850 81990
rect -17650 81920 -17350 81990
rect -17150 81920 -16850 81990
rect -16650 81920 -16350 81990
rect -16150 81920 -15850 81990
rect -15650 81920 -15350 81990
rect -15150 81920 -14850 81990
rect -14650 81920 -14350 81990
rect -14150 81920 -13850 81990
rect -13650 81920 -13350 81990
rect -13150 81920 -12850 81990
rect -12650 81920 -12350 81990
rect -12150 81920 -11850 81990
rect -11650 81920 -11350 81990
rect -11150 81920 -10850 81990
rect -10650 81920 -10350 81990
rect -10150 81920 -9850 81990
rect -9650 81920 -9350 81990
rect -9150 81920 -8850 81990
rect -8650 81920 -8350 81990
rect -8150 81920 -7850 81990
rect -7650 81920 -7350 81990
rect -7150 81920 -6850 81990
rect -6650 81920 -6350 81990
rect -6150 81920 -5850 81990
rect -5650 81920 -5350 81990
rect -5150 81920 -4850 81990
rect -4650 81920 -4350 81990
rect -4150 81920 -3850 81990
rect -3650 81920 -3350 81990
rect -3150 81920 -2850 81990
rect -2650 81920 -2350 81990
rect -2150 81920 -1850 81990
rect -1650 81920 -1350 81990
rect -1150 81920 -850 81990
rect -650 81920 -350 81990
rect -150 81920 150 81990
rect 350 81920 650 81990
rect 850 81920 1150 81990
rect 1350 81920 1650 81990
rect 1850 81920 2150 81990
rect 2350 81920 2650 81990
rect 2850 81920 3150 81990
rect 3350 81920 3650 81990
rect 3850 81920 4150 81990
rect 4350 81920 4650 81990
rect 4850 81920 5150 81990
rect 5350 81920 5650 81990
rect 5850 81920 6150 81990
rect 6350 81920 6650 81990
rect 6850 81920 7150 81990
rect 7350 81920 7650 81990
rect 7850 81920 8150 81990
rect 8350 81920 8650 81990
rect 8850 81920 9150 81990
rect 9350 81920 9650 81990
rect 9850 81920 10150 81990
rect 10350 81920 10650 81990
rect 10850 81920 11150 81990
rect 11350 81920 11650 81990
rect 11850 81920 12150 81990
rect 12350 81920 12650 81990
rect 12850 81920 13150 81990
rect 13350 81920 13650 81990
rect 13850 81920 14150 81990
rect 14350 81920 14650 81990
rect 14850 81920 15150 81990
rect 15350 81920 15650 81990
rect 15850 81920 16150 81990
rect 16350 81920 16650 81990
rect 16850 81920 17150 81990
rect 17350 81920 17650 81990
rect 17850 81920 18150 81990
rect 18350 81920 18650 81990
rect 18850 81920 19150 81990
rect 19350 81920 19650 81990
rect 19850 81920 20150 81990
rect 20350 81920 20650 81990
rect 20850 81920 21150 81990
rect 21350 81920 21650 81990
rect 21850 81920 22150 81990
rect 22350 81920 22650 81990
rect 22850 81920 23150 81990
rect 23350 81920 23650 81990
rect 23850 81920 24150 81990
rect 24350 81920 24650 81990
rect 24850 81920 25150 81990
rect 25350 81920 25650 81990
rect 25850 81920 26150 81990
rect 26350 81920 26650 81990
rect 26850 81920 27150 81990
rect 27350 81920 27650 81990
rect 27850 81920 28150 81990
rect 28350 81920 28650 81990
rect 28850 81920 29150 81990
rect 29350 81920 29650 81990
rect 29850 81920 30150 81990
rect 30350 81920 30650 81990
rect 30850 81920 31150 81990
rect 31350 81920 31650 81990
rect 31850 81920 32150 81990
rect 32350 81920 32650 81990
rect 32850 81920 33150 81990
rect 33350 81920 33650 81990
rect 33850 81920 34150 81990
rect 34350 81920 34650 81990
rect 34850 81920 35150 81990
rect 35350 81920 35650 81990
rect 35850 81920 36150 81990
rect 36350 81920 36650 81990
rect 36850 81920 37150 81990
rect 37350 81920 37650 81990
rect 37850 81920 38150 81990
rect 38350 81920 38650 81990
rect 38850 81920 39150 81990
rect 39350 81920 39650 81990
rect 39850 81920 40150 81990
rect 40350 81920 40650 81990
rect 40850 81920 41150 81990
rect 41350 81920 41650 81990
rect 41850 81920 42150 81990
rect 42350 81920 42650 81990
rect 42850 81920 43150 81990
rect 43350 81920 43650 81990
rect 43850 81920 44150 81990
rect 44350 81920 44650 81990
rect 44850 81920 45150 81990
rect 45350 81920 45650 81990
rect 45850 81920 46150 81990
rect 46350 81920 46650 81990
rect 46850 81920 47150 81990
rect 47350 81920 47650 81990
rect 47850 81920 48150 81990
rect 48350 81920 48650 81990
rect 48850 81920 49150 81990
rect 49350 81920 49650 81990
rect 49850 81920 50150 81990
rect 50350 81920 50650 81990
rect 50850 81920 51150 81990
rect 51350 81920 51650 81990
rect 51850 81920 52150 81990
rect 52350 81920 52650 81990
rect 52850 81920 53150 81990
rect 53350 81920 53650 81990
rect 53850 81920 54150 81990
rect 54350 81920 54650 81990
rect 54850 81920 55150 81990
rect 55350 81920 55650 81990
rect 55850 81920 56150 81990
rect 56350 81920 56650 81990
rect 56850 81920 57150 81990
rect 57350 81920 57650 81990
rect 57850 81920 58150 81990
rect 58350 81920 58650 81990
rect 58850 81920 59150 81990
rect 59350 81920 59650 81990
rect 59850 81920 60150 81990
rect 60350 81920 60650 81990
rect 60850 81920 61150 81990
rect 61350 81920 61650 81990
rect 61850 81920 62150 81990
rect 62350 81920 62650 81990
rect 62850 81920 63150 81990
rect 63350 81920 63650 81990
rect 63850 81920 64150 81990
rect 64350 81920 64650 81990
rect 64850 81920 65150 81990
rect 65350 81920 65650 81990
rect 65850 81920 66150 81990
rect 66350 81920 66650 81990
rect 66850 81920 67150 81990
rect 67350 81920 67650 81990
rect 67850 81920 68150 81990
rect 68350 81920 68650 81990
rect 68850 81920 69150 81990
rect 69350 81920 69650 81990
rect 69850 81920 70150 81990
rect 70350 81920 70650 81990
rect 70850 81920 71150 81990
rect 71350 81920 71650 81990
rect 71850 81920 72150 81990
rect 72350 81920 72650 81990
rect 72850 81920 73150 81990
rect 73350 81920 73650 81990
rect 73850 81920 74150 81990
rect 74350 81920 74650 81990
rect 74850 81920 75150 81990
rect 75350 81920 75650 81990
rect 75850 81920 76150 81990
rect 76350 81920 76650 81990
rect 76850 81920 77150 81990
rect 77350 81920 77650 81990
rect 77850 81920 78150 81990
rect 78350 81920 78650 81990
rect 78850 81920 79150 81990
rect 79350 81920 79650 81990
rect 79850 81920 80150 81990
rect 80350 81920 80650 81990
rect 80850 81920 81150 81990
rect 81350 81920 81650 81990
rect 81850 81920 82150 81990
rect 82350 81920 82650 81990
rect 82850 81920 83150 81990
rect 83350 81920 83650 81990
rect 83850 81920 84150 81990
rect 84350 81920 84650 81990
rect 84850 81920 85150 81990
rect 85350 81920 85650 81990
rect 85850 81920 86150 81990
rect 86350 81920 86650 81990
rect 86850 81920 87150 81990
rect 87350 81920 87650 81990
rect 87850 81920 88150 81990
rect 88350 81920 88650 81990
rect 88850 81920 89150 81990
rect 89350 81920 89650 81990
rect 89850 81920 90150 81990
rect 90350 81920 90650 81990
rect 90850 81920 91150 81990
rect 91350 81920 91650 81990
rect 91850 81920 92150 81990
rect 92350 81920 92650 81990
rect 92850 81920 93150 81990
rect 93350 81920 93650 81990
rect 93850 81920 94150 81990
rect 94350 81920 94650 81990
rect 94850 81920 95150 81990
rect 95350 81920 95650 81990
rect 95850 81920 96150 81990
rect 96350 81920 96650 81990
rect 96850 81920 97150 81990
rect 97350 81920 97650 81990
rect 97850 81920 98150 81990
rect 98350 81920 98650 81990
rect 98850 81920 99150 81990
rect 99350 81920 99650 81990
rect 99850 81920 100150 81990
rect 100350 81920 100500 81990
rect -83500 81880 100500 81920
rect -83500 81810 -83350 81880
rect -83150 81810 -82850 81880
rect -82650 81810 -82350 81880
rect -82150 81810 -81850 81880
rect -81650 81810 -81350 81880
rect -81150 81810 -80850 81880
rect -80650 81810 -80350 81880
rect -80150 81810 -79850 81880
rect -79650 81810 -79350 81880
rect -79150 81810 -78850 81880
rect -78650 81810 -78350 81880
rect -78150 81810 -77850 81880
rect -77650 81810 -77350 81880
rect -77150 81810 -76850 81880
rect -76650 81810 -76350 81880
rect -76150 81810 -75850 81880
rect -75650 81810 -75350 81880
rect -75150 81810 -74850 81880
rect -74650 81810 -74350 81880
rect -74150 81810 -73850 81880
rect -73650 81810 -73350 81880
rect -73150 81810 -72850 81880
rect -72650 81810 -72350 81880
rect -72150 81810 -71850 81880
rect -71650 81810 -71350 81880
rect -71150 81810 -70850 81880
rect -70650 81810 -70350 81880
rect -70150 81810 -69850 81880
rect -69650 81810 -69350 81880
rect -69150 81810 -68850 81880
rect -68650 81810 -68350 81880
rect -68150 81810 -67850 81880
rect -67650 81810 -67350 81880
rect -67150 81810 -66850 81880
rect -66650 81810 -66350 81880
rect -66150 81810 -65850 81880
rect -65650 81810 -65350 81880
rect -65150 81810 -64850 81880
rect -64650 81810 -64350 81880
rect -64150 81810 -63850 81880
rect -63650 81810 -63350 81880
rect -63150 81810 -62850 81880
rect -62650 81810 -62350 81880
rect -62150 81810 -61850 81880
rect -61650 81810 -61350 81880
rect -61150 81810 -60850 81880
rect -60650 81810 -60350 81880
rect -60150 81810 -59850 81880
rect -59650 81810 -59350 81880
rect -59150 81810 -58850 81880
rect -58650 81810 -58350 81880
rect -58150 81810 -57850 81880
rect -57650 81810 -57350 81880
rect -57150 81810 -56850 81880
rect -56650 81810 -56350 81880
rect -56150 81810 -55850 81880
rect -55650 81810 -55350 81880
rect -55150 81810 -54850 81880
rect -54650 81810 -54350 81880
rect -54150 81810 -53850 81880
rect -53650 81810 -53350 81880
rect -53150 81810 -52850 81880
rect -52650 81810 -52350 81880
rect -52150 81810 -51850 81880
rect -51650 81810 -51350 81880
rect -51150 81810 -50850 81880
rect -50650 81810 -50350 81880
rect -50150 81810 -49850 81880
rect -49650 81810 -49350 81880
rect -49150 81810 -48850 81880
rect -48650 81810 -48350 81880
rect -48150 81810 -47850 81880
rect -47650 81810 -47350 81880
rect -47150 81810 -46850 81880
rect -46650 81810 -46350 81880
rect -46150 81810 -45850 81880
rect -45650 81810 -45350 81880
rect -45150 81810 -44850 81880
rect -44650 81810 -44350 81880
rect -44150 81810 -43850 81880
rect -43650 81810 -43350 81880
rect -43150 81810 -42850 81880
rect -42650 81810 -42350 81880
rect -42150 81810 -41850 81880
rect -41650 81810 -41350 81880
rect -41150 81810 -40850 81880
rect -40650 81810 -40350 81880
rect -40150 81810 -39850 81880
rect -39650 81810 -39350 81880
rect -39150 81810 -38850 81880
rect -38650 81810 -38350 81880
rect -38150 81810 -37850 81880
rect -37650 81810 -37350 81880
rect -37150 81810 -36850 81880
rect -36650 81810 -36350 81880
rect -36150 81810 -35850 81880
rect -35650 81810 -35350 81880
rect -35150 81810 -34850 81880
rect -34650 81810 -34350 81880
rect -34150 81810 -33850 81880
rect -33650 81810 -33350 81880
rect -33150 81810 -32850 81880
rect -32650 81810 -32350 81880
rect -32150 81810 -31850 81880
rect -31650 81810 -31350 81880
rect -31150 81810 -30850 81880
rect -30650 81810 -30350 81880
rect -30150 81810 -29850 81880
rect -29650 81810 -29350 81880
rect -29150 81810 -28850 81880
rect -28650 81810 -28350 81880
rect -28150 81810 -27850 81880
rect -27650 81810 -27350 81880
rect -27150 81810 -26850 81880
rect -26650 81810 -26350 81880
rect -26150 81810 -25850 81880
rect -25650 81810 -25350 81880
rect -25150 81810 -24850 81880
rect -24650 81810 -24350 81880
rect -24150 81810 -23850 81880
rect -23650 81810 -23350 81880
rect -23150 81810 -22850 81880
rect -22650 81810 -22350 81880
rect -22150 81810 -21850 81880
rect -21650 81810 -21350 81880
rect -21150 81810 -20850 81880
rect -20650 81810 -20350 81880
rect -20150 81810 -19850 81880
rect -19650 81810 -19350 81880
rect -19150 81810 -18850 81880
rect -18650 81810 -18350 81880
rect -18150 81810 -17850 81880
rect -17650 81810 -17350 81880
rect -17150 81810 -16850 81880
rect -16650 81810 -16350 81880
rect -16150 81810 -15850 81880
rect -15650 81810 -15350 81880
rect -15150 81810 -14850 81880
rect -14650 81810 -14350 81880
rect -14150 81810 -13850 81880
rect -13650 81810 -13350 81880
rect -13150 81810 -12850 81880
rect -12650 81810 -12350 81880
rect -12150 81810 -11850 81880
rect -11650 81810 -11350 81880
rect -11150 81810 -10850 81880
rect -10650 81810 -10350 81880
rect -10150 81810 -9850 81880
rect -9650 81810 -9350 81880
rect -9150 81810 -8850 81880
rect -8650 81810 -8350 81880
rect -8150 81810 -7850 81880
rect -7650 81810 -7350 81880
rect -7150 81810 -6850 81880
rect -6650 81810 -6350 81880
rect -6150 81810 -5850 81880
rect -5650 81810 -5350 81880
rect -5150 81810 -4850 81880
rect -4650 81810 -4350 81880
rect -4150 81810 -3850 81880
rect -3650 81810 -3350 81880
rect -3150 81810 -2850 81880
rect -2650 81810 -2350 81880
rect -2150 81810 -1850 81880
rect -1650 81810 -1350 81880
rect -1150 81810 -850 81880
rect -650 81810 -350 81880
rect -150 81810 150 81880
rect 350 81810 650 81880
rect 850 81810 1150 81880
rect 1350 81810 1650 81880
rect 1850 81810 2150 81880
rect 2350 81810 2650 81880
rect 2850 81810 3150 81880
rect 3350 81810 3650 81880
rect 3850 81810 4150 81880
rect 4350 81810 4650 81880
rect 4850 81810 5150 81880
rect 5350 81810 5650 81880
rect 5850 81810 6150 81880
rect 6350 81810 6650 81880
rect 6850 81810 7150 81880
rect 7350 81810 7650 81880
rect 7850 81810 8150 81880
rect 8350 81810 8650 81880
rect 8850 81810 9150 81880
rect 9350 81810 9650 81880
rect 9850 81810 10150 81880
rect 10350 81810 10650 81880
rect 10850 81810 11150 81880
rect 11350 81810 11650 81880
rect 11850 81810 12150 81880
rect 12350 81810 12650 81880
rect 12850 81810 13150 81880
rect 13350 81810 13650 81880
rect 13850 81810 14150 81880
rect 14350 81810 14650 81880
rect 14850 81810 15150 81880
rect 15350 81810 15650 81880
rect 15850 81810 16150 81880
rect 16350 81810 16650 81880
rect 16850 81810 17150 81880
rect 17350 81810 17650 81880
rect 17850 81810 18150 81880
rect 18350 81810 18650 81880
rect 18850 81810 19150 81880
rect 19350 81810 19650 81880
rect 19850 81810 20150 81880
rect 20350 81810 20650 81880
rect 20850 81810 21150 81880
rect 21350 81810 21650 81880
rect 21850 81810 22150 81880
rect 22350 81810 22650 81880
rect 22850 81810 23150 81880
rect 23350 81810 23650 81880
rect 23850 81810 24150 81880
rect 24350 81810 24650 81880
rect 24850 81810 25150 81880
rect 25350 81810 25650 81880
rect 25850 81810 26150 81880
rect 26350 81810 26650 81880
rect 26850 81810 27150 81880
rect 27350 81810 27650 81880
rect 27850 81810 28150 81880
rect 28350 81810 28650 81880
rect 28850 81810 29150 81880
rect 29350 81810 29650 81880
rect 29850 81810 30150 81880
rect 30350 81810 30650 81880
rect 30850 81810 31150 81880
rect 31350 81810 31650 81880
rect 31850 81810 32150 81880
rect 32350 81810 32650 81880
rect 32850 81810 33150 81880
rect 33350 81810 33650 81880
rect 33850 81810 34150 81880
rect 34350 81810 34650 81880
rect 34850 81810 35150 81880
rect 35350 81810 35650 81880
rect 35850 81810 36150 81880
rect 36350 81810 36650 81880
rect 36850 81810 37150 81880
rect 37350 81810 37650 81880
rect 37850 81810 38150 81880
rect 38350 81810 38650 81880
rect 38850 81810 39150 81880
rect 39350 81810 39650 81880
rect 39850 81810 40150 81880
rect 40350 81810 40650 81880
rect 40850 81810 41150 81880
rect 41350 81810 41650 81880
rect 41850 81810 42150 81880
rect 42350 81810 42650 81880
rect 42850 81810 43150 81880
rect 43350 81810 43650 81880
rect 43850 81810 44150 81880
rect 44350 81810 44650 81880
rect 44850 81810 45150 81880
rect 45350 81810 45650 81880
rect 45850 81810 46150 81880
rect 46350 81810 46650 81880
rect 46850 81810 47150 81880
rect 47350 81810 47650 81880
rect 47850 81810 48150 81880
rect 48350 81810 48650 81880
rect 48850 81810 49150 81880
rect 49350 81810 49650 81880
rect 49850 81810 50150 81880
rect 50350 81810 50650 81880
rect 50850 81810 51150 81880
rect 51350 81810 51650 81880
rect 51850 81810 52150 81880
rect 52350 81810 52650 81880
rect 52850 81810 53150 81880
rect 53350 81810 53650 81880
rect 53850 81810 54150 81880
rect 54350 81810 54650 81880
rect 54850 81810 55150 81880
rect 55350 81810 55650 81880
rect 55850 81810 56150 81880
rect 56350 81810 56650 81880
rect 56850 81810 57150 81880
rect 57350 81810 57650 81880
rect 57850 81810 58150 81880
rect 58350 81810 58650 81880
rect 58850 81810 59150 81880
rect 59350 81810 59650 81880
rect 59850 81810 60150 81880
rect 60350 81810 60650 81880
rect 60850 81810 61150 81880
rect 61350 81810 61650 81880
rect 61850 81810 62150 81880
rect 62350 81810 62650 81880
rect 62850 81810 63150 81880
rect 63350 81810 63650 81880
rect 63850 81810 64150 81880
rect 64350 81810 64650 81880
rect 64850 81810 65150 81880
rect 65350 81810 65650 81880
rect 65850 81810 66150 81880
rect 66350 81810 66650 81880
rect 66850 81810 67150 81880
rect 67350 81810 67650 81880
rect 67850 81810 68150 81880
rect 68350 81810 68650 81880
rect 68850 81810 69150 81880
rect 69350 81810 69650 81880
rect 69850 81810 70150 81880
rect 70350 81810 70650 81880
rect 70850 81810 71150 81880
rect 71350 81810 71650 81880
rect 71850 81810 72150 81880
rect 72350 81810 72650 81880
rect 72850 81810 73150 81880
rect 73350 81810 73650 81880
rect 73850 81810 74150 81880
rect 74350 81810 74650 81880
rect 74850 81810 75150 81880
rect 75350 81810 75650 81880
rect 75850 81810 76150 81880
rect 76350 81810 76650 81880
rect 76850 81810 77150 81880
rect 77350 81810 77650 81880
rect 77850 81810 78150 81880
rect 78350 81810 78650 81880
rect 78850 81810 79150 81880
rect 79350 81810 79650 81880
rect 79850 81810 80150 81880
rect 80350 81810 80650 81880
rect 80850 81810 81150 81880
rect 81350 81810 81650 81880
rect 81850 81810 82150 81880
rect 82350 81810 82650 81880
rect 82850 81810 83150 81880
rect 83350 81810 83650 81880
rect 83850 81810 84150 81880
rect 84350 81810 84650 81880
rect 84850 81810 85150 81880
rect 85350 81810 85650 81880
rect 85850 81810 86150 81880
rect 86350 81810 86650 81880
rect 86850 81810 87150 81880
rect 87350 81810 87650 81880
rect 87850 81810 88150 81880
rect 88350 81810 88650 81880
rect 88850 81810 89150 81880
rect 89350 81810 89650 81880
rect 89850 81810 90150 81880
rect 90350 81810 90650 81880
rect 90850 81810 91150 81880
rect 91350 81810 91650 81880
rect 91850 81810 92150 81880
rect 92350 81810 92650 81880
rect 92850 81810 93150 81880
rect 93350 81810 93650 81880
rect 93850 81810 94150 81880
rect 94350 81810 94650 81880
rect 94850 81810 95150 81880
rect 95350 81810 95650 81880
rect 95850 81810 96150 81880
rect 96350 81810 96650 81880
rect 96850 81810 97150 81880
rect 97350 81810 97650 81880
rect 97850 81810 98150 81880
rect 98350 81810 98650 81880
rect 98850 81810 99150 81880
rect 99350 81810 99650 81880
rect 99850 81810 100150 81880
rect 100350 81810 100500 81880
rect -83500 81800 100500 81810
rect -83500 81780 -83380 81800
rect -83120 81780 -82880 81800
rect -82620 81780 -82380 81800
rect -82120 81780 -81880 81800
rect -81620 81780 -81380 81800
rect -81120 81780 -80880 81800
rect -80620 81780 -80380 81800
rect -80120 81780 -79880 81800
rect -79620 81780 -79380 81800
rect -79120 81780 -78880 81800
rect -78620 81780 -78380 81800
rect -78120 81780 -77880 81800
rect -77620 81780 -77380 81800
rect -77120 81780 -76880 81800
rect -76620 81780 -76380 81800
rect -76120 81780 -75880 81800
rect -75620 81780 -75380 81800
rect -75120 81780 -74880 81800
rect -74620 81780 -74380 81800
rect -74120 81780 -73880 81800
rect -73620 81780 -73380 81800
rect -73120 81780 -72880 81800
rect -72620 81780 -72380 81800
rect -72120 81780 -71880 81800
rect -71620 81780 -71380 81800
rect -71120 81780 -70880 81800
rect -70620 81780 -70380 81800
rect -70120 81780 -69880 81800
rect -69620 81780 -69380 81800
rect -69120 81780 -68880 81800
rect -68620 81780 -68380 81800
rect -68120 81780 -67880 81800
rect -67620 81780 -67380 81800
rect -67120 81780 -66880 81800
rect -66620 81780 -66380 81800
rect -66120 81780 -65880 81800
rect -65620 81780 -65380 81800
rect -65120 81780 -64880 81800
rect -64620 81780 -64380 81800
rect -64120 81780 -63880 81800
rect -63620 81780 -63380 81800
rect -63120 81780 -62880 81800
rect -62620 81780 -62380 81800
rect -62120 81780 -61880 81800
rect -61620 81780 -61380 81800
rect -61120 81780 -60880 81800
rect -60620 81780 -60380 81800
rect -60120 81780 -59880 81800
rect -59620 81780 -59380 81800
rect -59120 81780 -58880 81800
rect -58620 81780 -58380 81800
rect -58120 81780 -57880 81800
rect -57620 81780 -57380 81800
rect -57120 81780 -56880 81800
rect -56620 81780 -56380 81800
rect -56120 81780 -55880 81800
rect -55620 81780 -55380 81800
rect -55120 81780 -54880 81800
rect -54620 81780 -54380 81800
rect -54120 81780 -53880 81800
rect -53620 81780 -53380 81800
rect -53120 81780 -52880 81800
rect -52620 81780 -52380 81800
rect -52120 81780 -51880 81800
rect -51620 81780 -51380 81800
rect -51120 81780 -50880 81800
rect -50620 81780 -50380 81800
rect -50120 81780 -49880 81800
rect -49620 81780 -49380 81800
rect -49120 81780 -48880 81800
rect -48620 81780 -48380 81800
rect -48120 81780 -47880 81800
rect -47620 81780 -47380 81800
rect -47120 81780 -46880 81800
rect -46620 81780 -46380 81800
rect -46120 81780 -45880 81800
rect -45620 81780 -45380 81800
rect -45120 81780 -44880 81800
rect -44620 81780 -44380 81800
rect -44120 81780 -43880 81800
rect -43620 81780 -43380 81800
rect -43120 81780 -42880 81800
rect -42620 81780 -42380 81800
rect -42120 81780 -41880 81800
rect -41620 81780 -41380 81800
rect -41120 81780 -40880 81800
rect -40620 81780 -40380 81800
rect -40120 81780 -39880 81800
rect -39620 81780 -39380 81800
rect -39120 81780 -38880 81800
rect -38620 81780 -38380 81800
rect -38120 81780 -37880 81800
rect -37620 81780 -37380 81800
rect -37120 81780 -36880 81800
rect -36620 81780 -36380 81800
rect -36120 81780 -35880 81800
rect -35620 81780 -35380 81800
rect -35120 81780 -34880 81800
rect -34620 81780 -34380 81800
rect -34120 81780 -33880 81800
rect -33620 81780 -33380 81800
rect -33120 81780 -32880 81800
rect -32620 81780 -32380 81800
rect -32120 81780 -31880 81800
rect -31620 81780 -31380 81800
rect -31120 81780 -30880 81800
rect -30620 81780 -30380 81800
rect -30120 81780 -29880 81800
rect -29620 81780 -29380 81800
rect -29120 81780 -28880 81800
rect -28620 81780 -28380 81800
rect -28120 81780 -27880 81800
rect -27620 81780 -27380 81800
rect -27120 81780 -26880 81800
rect -26620 81780 -26380 81800
rect -26120 81780 -25880 81800
rect -25620 81780 -25380 81800
rect -25120 81780 -24880 81800
rect -24620 81780 -24380 81800
rect -24120 81780 -23880 81800
rect -23620 81780 -23380 81800
rect -23120 81780 -22880 81800
rect -22620 81780 -22380 81800
rect -22120 81780 -21880 81800
rect -21620 81780 -21380 81800
rect -21120 81780 -20880 81800
rect -20620 81780 -20380 81800
rect -20120 81780 -19880 81800
rect -19620 81780 -19380 81800
rect -19120 81780 -18880 81800
rect -18620 81780 -18380 81800
rect -18120 81780 -17880 81800
rect -17620 81780 -17380 81800
rect -17120 81780 -16880 81800
rect -16620 81780 -16380 81800
rect -16120 81780 -15880 81800
rect -15620 81780 -15380 81800
rect -15120 81780 -14880 81800
rect -14620 81780 -14380 81800
rect -14120 81780 -13880 81800
rect -13620 81780 -13380 81800
rect -13120 81780 -12880 81800
rect -12620 81780 -12380 81800
rect -12120 81780 -11880 81800
rect -11620 81780 -11380 81800
rect -11120 81780 -10880 81800
rect -10620 81780 -10380 81800
rect -10120 81780 -9880 81800
rect -9620 81780 -9380 81800
rect -9120 81780 -8880 81800
rect -8620 81780 -8380 81800
rect -8120 81780 -7880 81800
rect -7620 81780 -7380 81800
rect -7120 81780 -6880 81800
rect -6620 81780 -6380 81800
rect -6120 81780 -5880 81800
rect -5620 81780 -5380 81800
rect -5120 81780 -4880 81800
rect -4620 81780 -4380 81800
rect -4120 81780 -3880 81800
rect -3620 81780 -3380 81800
rect -3120 81780 -2880 81800
rect -2620 81780 -2380 81800
rect -2120 81780 -1880 81800
rect -1620 81780 -1380 81800
rect -1120 81780 -880 81800
rect -620 81780 -380 81800
rect -120 81780 120 81800
rect 380 81780 620 81800
rect 880 81780 1120 81800
rect 1380 81780 1620 81800
rect 1880 81780 2120 81800
rect 2380 81780 2620 81800
rect 2880 81780 3120 81800
rect 3380 81780 3620 81800
rect 3880 81780 4120 81800
rect 4380 81780 4620 81800
rect 4880 81780 5120 81800
rect 5380 81780 5620 81800
rect 5880 81780 6120 81800
rect 6380 81780 6620 81800
rect 6880 81780 7120 81800
rect 7380 81780 7620 81800
rect 7880 81780 8120 81800
rect 8380 81780 8620 81800
rect 8880 81780 9120 81800
rect 9380 81780 9620 81800
rect 9880 81780 10120 81800
rect 10380 81780 10620 81800
rect 10880 81780 11120 81800
rect 11380 81780 11620 81800
rect 11880 81780 12120 81800
rect 12380 81780 12620 81800
rect 12880 81780 13120 81800
rect 13380 81780 13620 81800
rect 13880 81780 14120 81800
rect 14380 81780 14620 81800
rect 14880 81780 15120 81800
rect 15380 81780 15620 81800
rect 15880 81780 16120 81800
rect 16380 81780 16620 81800
rect 16880 81780 17120 81800
rect 17380 81780 17620 81800
rect 17880 81780 18120 81800
rect 18380 81780 18620 81800
rect 18880 81780 19120 81800
rect 19380 81780 19620 81800
rect 19880 81780 20120 81800
rect 20380 81780 20620 81800
rect 20880 81780 21120 81800
rect 21380 81780 21620 81800
rect 21880 81780 22120 81800
rect 22380 81780 22620 81800
rect 22880 81780 23120 81800
rect 23380 81780 23620 81800
rect 23880 81780 24120 81800
rect 24380 81780 24620 81800
rect 24880 81780 25120 81800
rect 25380 81780 25620 81800
rect 25880 81780 26120 81800
rect 26380 81780 26620 81800
rect 26880 81780 27120 81800
rect 27380 81780 27620 81800
rect 27880 81780 28120 81800
rect 28380 81780 28620 81800
rect 28880 81780 29120 81800
rect 29380 81780 29620 81800
rect 29880 81780 30120 81800
rect 30380 81780 30620 81800
rect 30880 81780 31120 81800
rect 31380 81780 31620 81800
rect 31880 81780 32120 81800
rect 32380 81780 32620 81800
rect 32880 81780 33120 81800
rect 33380 81780 33620 81800
rect 33880 81780 34120 81800
rect 34380 81780 34620 81800
rect 34880 81780 35120 81800
rect 35380 81780 35620 81800
rect 35880 81780 36120 81800
rect 36380 81780 36620 81800
rect 36880 81780 37120 81800
rect 37380 81780 37620 81800
rect 37880 81780 38120 81800
rect 38380 81780 38620 81800
rect 38880 81780 39120 81800
rect 39380 81780 39620 81800
rect 39880 81780 40120 81800
rect 40380 81780 40620 81800
rect 40880 81780 41120 81800
rect 41380 81780 41620 81800
rect 41880 81780 42120 81800
rect 42380 81780 42620 81800
rect 42880 81780 43120 81800
rect 43380 81780 43620 81800
rect 43880 81780 44120 81800
rect 44380 81780 44620 81800
rect 44880 81780 45120 81800
rect 45380 81780 45620 81800
rect 45880 81780 46120 81800
rect 46380 81780 46620 81800
rect 46880 81780 47120 81800
rect 47380 81780 47620 81800
rect 47880 81780 48120 81800
rect 48380 81780 48620 81800
rect 48880 81780 49120 81800
rect 49380 81780 49620 81800
rect 49880 81780 50120 81800
rect 50380 81780 50620 81800
rect 50880 81780 51120 81800
rect 51380 81780 51620 81800
rect 51880 81780 52120 81800
rect 52380 81780 52620 81800
rect 52880 81780 53120 81800
rect 53380 81780 53620 81800
rect 53880 81780 54120 81800
rect 54380 81780 54620 81800
rect 54880 81780 55120 81800
rect 55380 81780 55620 81800
rect 55880 81780 56120 81800
rect 56380 81780 56620 81800
rect 56880 81780 57120 81800
rect 57380 81780 57620 81800
rect 57880 81780 58120 81800
rect 58380 81780 58620 81800
rect 58880 81780 59120 81800
rect 59380 81780 59620 81800
rect 59880 81780 60120 81800
rect 60380 81780 60620 81800
rect 60880 81780 61120 81800
rect 61380 81780 61620 81800
rect 61880 81780 62120 81800
rect 62380 81780 62620 81800
rect 62880 81780 63120 81800
rect 63380 81780 63620 81800
rect 63880 81780 64120 81800
rect 64380 81780 64620 81800
rect 64880 81780 65120 81800
rect 65380 81780 65620 81800
rect 65880 81780 66120 81800
rect 66380 81780 66620 81800
rect 66880 81780 67120 81800
rect 67380 81780 67620 81800
rect 67880 81780 68120 81800
rect 68380 81780 68620 81800
rect 68880 81780 69120 81800
rect 69380 81780 69620 81800
rect 69880 81780 70120 81800
rect 70380 81780 70620 81800
rect 70880 81780 71120 81800
rect 71380 81780 71620 81800
rect 71880 81780 72120 81800
rect 72380 81780 72620 81800
rect 72880 81780 73120 81800
rect 73380 81780 73620 81800
rect 73880 81780 74120 81800
rect 74380 81780 74620 81800
rect 74880 81780 75120 81800
rect 75380 81780 75620 81800
rect 75880 81780 76120 81800
rect 76380 81780 76620 81800
rect 76880 81780 77120 81800
rect 77380 81780 77620 81800
rect 77880 81780 78120 81800
rect 78380 81780 78620 81800
rect 78880 81780 79120 81800
rect 79380 81780 79620 81800
rect 79880 81780 80120 81800
rect 80380 81780 80620 81800
rect 80880 81780 81120 81800
rect 81380 81780 81620 81800
rect 81880 81780 82120 81800
rect 82380 81780 82620 81800
rect 82880 81780 83120 81800
rect 83380 81780 83620 81800
rect 83880 81780 84120 81800
rect 84380 81780 84620 81800
rect 84880 81780 85120 81800
rect 85380 81780 85620 81800
rect 85880 81780 86120 81800
rect 86380 81780 86620 81800
rect 86880 81780 87120 81800
rect 87380 81780 87620 81800
rect 87880 81780 88120 81800
rect 88380 81780 88620 81800
rect 88880 81780 89120 81800
rect 89380 81780 89620 81800
rect 89880 81780 90120 81800
rect 90380 81780 90620 81800
rect 90880 81780 91120 81800
rect 91380 81780 91620 81800
rect 91880 81780 92120 81800
rect 92380 81780 92620 81800
rect 92880 81780 93120 81800
rect 93380 81780 93620 81800
rect 93880 81780 94120 81800
rect 94380 81780 94620 81800
rect 94880 81780 95120 81800
rect 95380 81780 95620 81800
rect 95880 81780 96120 81800
rect 96380 81780 96620 81800
rect 96880 81780 97120 81800
rect 97380 81780 97620 81800
rect 97880 81780 98120 81800
rect 98380 81780 98620 81800
rect 98880 81780 99120 81800
rect 99380 81780 99620 81800
rect 99880 81780 100120 81800
rect 100380 81780 100500 81800
rect -83500 81750 -83400 81780
rect -83500 81550 -83480 81750
rect -83410 81550 -83400 81750
rect -83500 81520 -83400 81550
rect -83100 81750 -82900 81780
rect -83100 81550 -83090 81750
rect -83020 81550 -82980 81750
rect -82910 81550 -82900 81750
rect -83100 81520 -82900 81550
rect -82600 81750 -82400 81780
rect -82600 81550 -82590 81750
rect -82520 81550 -82480 81750
rect -82410 81550 -82400 81750
rect -82600 81520 -82400 81550
rect -82100 81750 -81900 81780
rect -82100 81550 -82090 81750
rect -82020 81550 -81980 81750
rect -81910 81550 -81900 81750
rect -82100 81520 -81900 81550
rect -81600 81750 -81400 81780
rect -81600 81550 -81590 81750
rect -81520 81550 -81480 81750
rect -81410 81550 -81400 81750
rect -81600 81520 -81400 81550
rect -81100 81750 -80900 81780
rect -81100 81550 -81090 81750
rect -81020 81550 -80980 81750
rect -80910 81550 -80900 81750
rect -81100 81520 -80900 81550
rect -80600 81750 -80400 81780
rect -80600 81550 -80590 81750
rect -80520 81550 -80480 81750
rect -80410 81550 -80400 81750
rect -80600 81520 -80400 81550
rect -80100 81750 -79900 81780
rect -80100 81550 -80090 81750
rect -80020 81550 -79980 81750
rect -79910 81550 -79900 81750
rect -80100 81520 -79900 81550
rect -79600 81750 -79400 81780
rect -79600 81550 -79590 81750
rect -79520 81550 -79480 81750
rect -79410 81550 -79400 81750
rect -79600 81520 -79400 81550
rect -79100 81750 -78900 81780
rect -79100 81550 -79090 81750
rect -79020 81550 -78980 81750
rect -78910 81550 -78900 81750
rect -79100 81520 -78900 81550
rect -78600 81750 -78400 81780
rect -78600 81550 -78590 81750
rect -78520 81550 -78480 81750
rect -78410 81550 -78400 81750
rect -78600 81520 -78400 81550
rect -78100 81750 -77900 81780
rect -78100 81550 -78090 81750
rect -78020 81550 -77980 81750
rect -77910 81550 -77900 81750
rect -78100 81520 -77900 81550
rect -77600 81750 -77400 81780
rect -77600 81550 -77590 81750
rect -77520 81550 -77480 81750
rect -77410 81550 -77400 81750
rect -77600 81520 -77400 81550
rect -77100 81750 -76900 81780
rect -77100 81550 -77090 81750
rect -77020 81550 -76980 81750
rect -76910 81550 -76900 81750
rect -77100 81520 -76900 81550
rect -76600 81750 -76400 81780
rect -76600 81550 -76590 81750
rect -76520 81550 -76480 81750
rect -76410 81550 -76400 81750
rect -76600 81520 -76400 81550
rect -76100 81750 -75900 81780
rect -76100 81550 -76090 81750
rect -76020 81550 -75980 81750
rect -75910 81550 -75900 81750
rect -76100 81520 -75900 81550
rect -75600 81750 -75400 81780
rect -75600 81550 -75590 81750
rect -75520 81550 -75480 81750
rect -75410 81550 -75400 81750
rect -75600 81520 -75400 81550
rect -75100 81750 -74900 81780
rect -75100 81550 -75090 81750
rect -75020 81550 -74980 81750
rect -74910 81550 -74900 81750
rect -75100 81520 -74900 81550
rect -74600 81750 -74400 81780
rect -74600 81550 -74590 81750
rect -74520 81550 -74480 81750
rect -74410 81550 -74400 81750
rect -74600 81520 -74400 81550
rect -74100 81750 -73900 81780
rect -74100 81550 -74090 81750
rect -74020 81550 -73980 81750
rect -73910 81550 -73900 81750
rect -74100 81520 -73900 81550
rect -73600 81750 -73400 81780
rect -73600 81550 -73590 81750
rect -73520 81550 -73480 81750
rect -73410 81550 -73400 81750
rect -73600 81520 -73400 81550
rect -73100 81750 -72900 81780
rect -73100 81550 -73090 81750
rect -73020 81550 -72980 81750
rect -72910 81550 -72900 81750
rect -73100 81520 -72900 81550
rect -72600 81750 -72400 81780
rect -72600 81550 -72590 81750
rect -72520 81550 -72480 81750
rect -72410 81550 -72400 81750
rect -72600 81520 -72400 81550
rect -72100 81750 -71900 81780
rect -72100 81550 -72090 81750
rect -72020 81550 -71980 81750
rect -71910 81550 -71900 81750
rect -72100 81520 -71900 81550
rect -71600 81750 -71400 81780
rect -71600 81550 -71590 81750
rect -71520 81550 -71480 81750
rect -71410 81550 -71400 81750
rect -71600 81520 -71400 81550
rect -71100 81750 -70900 81780
rect -71100 81550 -71090 81750
rect -71020 81550 -70980 81750
rect -70910 81550 -70900 81750
rect -71100 81520 -70900 81550
rect -70600 81750 -70400 81780
rect -70600 81550 -70590 81750
rect -70520 81550 -70480 81750
rect -70410 81550 -70400 81750
rect -70600 81520 -70400 81550
rect -70100 81750 -69900 81780
rect -70100 81550 -70090 81750
rect -70020 81550 -69980 81750
rect -69910 81550 -69900 81750
rect -70100 81520 -69900 81550
rect -69600 81750 -69400 81780
rect -69600 81550 -69590 81750
rect -69520 81550 -69480 81750
rect -69410 81550 -69400 81750
rect -69600 81520 -69400 81550
rect -69100 81750 -68900 81780
rect -69100 81550 -69090 81750
rect -69020 81550 -68980 81750
rect -68910 81550 -68900 81750
rect -69100 81520 -68900 81550
rect -68600 81750 -68400 81780
rect -68600 81550 -68590 81750
rect -68520 81550 -68480 81750
rect -68410 81550 -68400 81750
rect -68600 81520 -68400 81550
rect -68100 81750 -67900 81780
rect -68100 81550 -68090 81750
rect -68020 81550 -67980 81750
rect -67910 81550 -67900 81750
rect -68100 81520 -67900 81550
rect -67600 81750 -67400 81780
rect -67600 81550 -67590 81750
rect -67520 81550 -67480 81750
rect -67410 81550 -67400 81750
rect -67600 81520 -67400 81550
rect -67100 81750 -66900 81780
rect -67100 81550 -67090 81750
rect -67020 81550 -66980 81750
rect -66910 81550 -66900 81750
rect -67100 81520 -66900 81550
rect -66600 81750 -66400 81780
rect -66600 81550 -66590 81750
rect -66520 81550 -66480 81750
rect -66410 81550 -66400 81750
rect -66600 81520 -66400 81550
rect -66100 81750 -65900 81780
rect -66100 81550 -66090 81750
rect -66020 81550 -65980 81750
rect -65910 81550 -65900 81750
rect -66100 81520 -65900 81550
rect -65600 81750 -65400 81780
rect -65600 81550 -65590 81750
rect -65520 81550 -65480 81750
rect -65410 81550 -65400 81750
rect -65600 81520 -65400 81550
rect -65100 81750 -64900 81780
rect -65100 81550 -65090 81750
rect -65020 81550 -64980 81750
rect -64910 81550 -64900 81750
rect -65100 81520 -64900 81550
rect -64600 81750 -64400 81780
rect -64600 81550 -64590 81750
rect -64520 81550 -64480 81750
rect -64410 81550 -64400 81750
rect -64600 81520 -64400 81550
rect -64100 81750 -63900 81780
rect -64100 81550 -64090 81750
rect -64020 81550 -63980 81750
rect -63910 81550 -63900 81750
rect -64100 81520 -63900 81550
rect -63600 81750 -63400 81780
rect -63600 81550 -63590 81750
rect -63520 81550 -63480 81750
rect -63410 81550 -63400 81750
rect -63600 81520 -63400 81550
rect -63100 81750 -62900 81780
rect -63100 81550 -63090 81750
rect -63020 81550 -62980 81750
rect -62910 81550 -62900 81750
rect -63100 81520 -62900 81550
rect -62600 81750 -62400 81780
rect -62600 81550 -62590 81750
rect -62520 81550 -62480 81750
rect -62410 81550 -62400 81750
rect -62600 81520 -62400 81550
rect -62100 81750 -61900 81780
rect -62100 81550 -62090 81750
rect -62020 81550 -61980 81750
rect -61910 81550 -61900 81750
rect -62100 81520 -61900 81550
rect -61600 81750 -61400 81780
rect -61600 81550 -61590 81750
rect -61520 81550 -61480 81750
rect -61410 81550 -61400 81750
rect -61600 81520 -61400 81550
rect -61100 81750 -60900 81780
rect -61100 81550 -61090 81750
rect -61020 81550 -60980 81750
rect -60910 81550 -60900 81750
rect -61100 81520 -60900 81550
rect -60600 81750 -60400 81780
rect -60600 81550 -60590 81750
rect -60520 81550 -60480 81750
rect -60410 81550 -60400 81750
rect -60600 81520 -60400 81550
rect -60100 81750 -59900 81780
rect -60100 81550 -60090 81750
rect -60020 81550 -59980 81750
rect -59910 81550 -59900 81750
rect -60100 81520 -59900 81550
rect -59600 81750 -59400 81780
rect -59600 81550 -59590 81750
rect -59520 81550 -59480 81750
rect -59410 81550 -59400 81750
rect -59600 81520 -59400 81550
rect -59100 81750 -58900 81780
rect -59100 81550 -59090 81750
rect -59020 81550 -58980 81750
rect -58910 81550 -58900 81750
rect -59100 81520 -58900 81550
rect -58600 81750 -58400 81780
rect -58600 81550 -58590 81750
rect -58520 81550 -58480 81750
rect -58410 81550 -58400 81750
rect -58600 81520 -58400 81550
rect -58100 81750 -57900 81780
rect -58100 81550 -58090 81750
rect -58020 81550 -57980 81750
rect -57910 81550 -57900 81750
rect -58100 81520 -57900 81550
rect -57600 81750 -57400 81780
rect -57600 81550 -57590 81750
rect -57520 81550 -57480 81750
rect -57410 81550 -57400 81750
rect -57600 81520 -57400 81550
rect -57100 81750 -56900 81780
rect -57100 81550 -57090 81750
rect -57020 81550 -56980 81750
rect -56910 81550 -56900 81750
rect -57100 81520 -56900 81550
rect -56600 81750 -56400 81780
rect -56600 81550 -56590 81750
rect -56520 81550 -56480 81750
rect -56410 81550 -56400 81750
rect -56600 81520 -56400 81550
rect -56100 81750 -55900 81780
rect -56100 81550 -56090 81750
rect -56020 81550 -55980 81750
rect -55910 81550 -55900 81750
rect -56100 81520 -55900 81550
rect -55600 81750 -55400 81780
rect -55600 81550 -55590 81750
rect -55520 81550 -55480 81750
rect -55410 81550 -55400 81750
rect -55600 81520 -55400 81550
rect -55100 81750 -54900 81780
rect -55100 81550 -55090 81750
rect -55020 81550 -54980 81750
rect -54910 81550 -54900 81750
rect -55100 81520 -54900 81550
rect -54600 81750 -54400 81780
rect -54600 81550 -54590 81750
rect -54520 81550 -54480 81750
rect -54410 81550 -54400 81750
rect -54600 81520 -54400 81550
rect -54100 81750 -53900 81780
rect -54100 81550 -54090 81750
rect -54020 81550 -53980 81750
rect -53910 81550 -53900 81750
rect -54100 81520 -53900 81550
rect -53600 81750 -53400 81780
rect -53600 81550 -53590 81750
rect -53520 81550 -53480 81750
rect -53410 81550 -53400 81750
rect -53600 81520 -53400 81550
rect -53100 81750 -52900 81780
rect -53100 81550 -53090 81750
rect -53020 81550 -52980 81750
rect -52910 81550 -52900 81750
rect -53100 81520 -52900 81550
rect -52600 81750 -52400 81780
rect -52600 81550 -52590 81750
rect -52520 81550 -52480 81750
rect -52410 81550 -52400 81750
rect -52600 81520 -52400 81550
rect -52100 81750 -51900 81780
rect -52100 81550 -52090 81750
rect -52020 81550 -51980 81750
rect -51910 81550 -51900 81750
rect -52100 81520 -51900 81550
rect -51600 81750 -51400 81780
rect -51600 81550 -51590 81750
rect -51520 81550 -51480 81750
rect -51410 81550 -51400 81750
rect -51600 81520 -51400 81550
rect -51100 81750 -50900 81780
rect -51100 81550 -51090 81750
rect -51020 81550 -50980 81750
rect -50910 81550 -50900 81750
rect -51100 81520 -50900 81550
rect -50600 81750 -50400 81780
rect -50600 81550 -50590 81750
rect -50520 81550 -50480 81750
rect -50410 81550 -50400 81750
rect -50600 81520 -50400 81550
rect -50100 81750 -49900 81780
rect -50100 81550 -50090 81750
rect -50020 81550 -49980 81750
rect -49910 81550 -49900 81750
rect -50100 81520 -49900 81550
rect -49600 81750 -49400 81780
rect -49600 81550 -49590 81750
rect -49520 81550 -49480 81750
rect -49410 81550 -49400 81750
rect -49600 81520 -49400 81550
rect -49100 81750 -48900 81780
rect -49100 81550 -49090 81750
rect -49020 81550 -48980 81750
rect -48910 81550 -48900 81750
rect -49100 81520 -48900 81550
rect -48600 81750 -48400 81780
rect -48600 81550 -48590 81750
rect -48520 81550 -48480 81750
rect -48410 81550 -48400 81750
rect -48600 81520 -48400 81550
rect -48100 81750 -47900 81780
rect -48100 81550 -48090 81750
rect -48020 81550 -47980 81750
rect -47910 81550 -47900 81750
rect -48100 81520 -47900 81550
rect -47600 81750 -47400 81780
rect -47600 81550 -47590 81750
rect -47520 81550 -47480 81750
rect -47410 81550 -47400 81750
rect -47600 81520 -47400 81550
rect -47100 81750 -46900 81780
rect -47100 81550 -47090 81750
rect -47020 81550 -46980 81750
rect -46910 81550 -46900 81750
rect -47100 81520 -46900 81550
rect -46600 81750 -46400 81780
rect -46600 81550 -46590 81750
rect -46520 81550 -46480 81750
rect -46410 81550 -46400 81750
rect -46600 81520 -46400 81550
rect -46100 81750 -45900 81780
rect -46100 81550 -46090 81750
rect -46020 81550 -45980 81750
rect -45910 81550 -45900 81750
rect -46100 81520 -45900 81550
rect -45600 81750 -45400 81780
rect -45600 81550 -45590 81750
rect -45520 81550 -45480 81750
rect -45410 81550 -45400 81750
rect -45600 81520 -45400 81550
rect -45100 81750 -44900 81780
rect -45100 81550 -45090 81750
rect -45020 81550 -44980 81750
rect -44910 81550 -44900 81750
rect -45100 81520 -44900 81550
rect -44600 81750 -44400 81780
rect -44600 81550 -44590 81750
rect -44520 81550 -44480 81750
rect -44410 81550 -44400 81750
rect -44600 81520 -44400 81550
rect -44100 81750 -43900 81780
rect -44100 81550 -44090 81750
rect -44020 81550 -43980 81750
rect -43910 81550 -43900 81750
rect -44100 81520 -43900 81550
rect -43600 81750 -43400 81780
rect -43600 81550 -43590 81750
rect -43520 81550 -43480 81750
rect -43410 81550 -43400 81750
rect -43600 81520 -43400 81550
rect -43100 81750 -42900 81780
rect -43100 81550 -43090 81750
rect -43020 81550 -42980 81750
rect -42910 81550 -42900 81750
rect -43100 81520 -42900 81550
rect -42600 81750 -42400 81780
rect -42600 81550 -42590 81750
rect -42520 81550 -42480 81750
rect -42410 81550 -42400 81750
rect -42600 81520 -42400 81550
rect -42100 81750 -41900 81780
rect -42100 81550 -42090 81750
rect -42020 81550 -41980 81750
rect -41910 81550 -41900 81750
rect -42100 81520 -41900 81550
rect -41600 81750 -41400 81780
rect -41600 81550 -41590 81750
rect -41520 81550 -41480 81750
rect -41410 81550 -41400 81750
rect -41600 81520 -41400 81550
rect -41100 81750 -40900 81780
rect -41100 81550 -41090 81750
rect -41020 81550 -40980 81750
rect -40910 81550 -40900 81750
rect -41100 81520 -40900 81550
rect -40600 81750 -40400 81780
rect -40600 81550 -40590 81750
rect -40520 81550 -40480 81750
rect -40410 81550 -40400 81750
rect -40600 81520 -40400 81550
rect -40100 81750 -39900 81780
rect -40100 81550 -40090 81750
rect -40020 81550 -39980 81750
rect -39910 81550 -39900 81750
rect -40100 81520 -39900 81550
rect -39600 81750 -39400 81780
rect -39600 81550 -39590 81750
rect -39520 81550 -39480 81750
rect -39410 81550 -39400 81750
rect -39600 81520 -39400 81550
rect -39100 81750 -38900 81780
rect -39100 81550 -39090 81750
rect -39020 81550 -38980 81750
rect -38910 81550 -38900 81750
rect -39100 81520 -38900 81550
rect -38600 81750 -38400 81780
rect -38600 81550 -38590 81750
rect -38520 81550 -38480 81750
rect -38410 81550 -38400 81750
rect -38600 81520 -38400 81550
rect -38100 81750 -37900 81780
rect -38100 81550 -38090 81750
rect -38020 81550 -37980 81750
rect -37910 81550 -37900 81750
rect -38100 81520 -37900 81550
rect -37600 81750 -37400 81780
rect -37600 81550 -37590 81750
rect -37520 81550 -37480 81750
rect -37410 81550 -37400 81750
rect -37600 81520 -37400 81550
rect -37100 81750 -36900 81780
rect -37100 81550 -37090 81750
rect -37020 81550 -36980 81750
rect -36910 81550 -36900 81750
rect -37100 81520 -36900 81550
rect -36600 81750 -36400 81780
rect -36600 81550 -36590 81750
rect -36520 81550 -36480 81750
rect -36410 81550 -36400 81750
rect -36600 81520 -36400 81550
rect -36100 81750 -35900 81780
rect -36100 81550 -36090 81750
rect -36020 81550 -35980 81750
rect -35910 81550 -35900 81750
rect -36100 81520 -35900 81550
rect -35600 81750 -35400 81780
rect -35600 81550 -35590 81750
rect -35520 81550 -35480 81750
rect -35410 81550 -35400 81750
rect -35600 81520 -35400 81550
rect -35100 81750 -34900 81780
rect -35100 81550 -35090 81750
rect -35020 81550 -34980 81750
rect -34910 81550 -34900 81750
rect -35100 81520 -34900 81550
rect -34600 81750 -34400 81780
rect -34600 81550 -34590 81750
rect -34520 81550 -34480 81750
rect -34410 81550 -34400 81750
rect -34600 81520 -34400 81550
rect -34100 81750 -33900 81780
rect -34100 81550 -34090 81750
rect -34020 81550 -33980 81750
rect -33910 81550 -33900 81750
rect -34100 81520 -33900 81550
rect -33600 81750 -33400 81780
rect -33600 81550 -33590 81750
rect -33520 81550 -33480 81750
rect -33410 81550 -33400 81750
rect -33600 81520 -33400 81550
rect -33100 81750 -32900 81780
rect -33100 81550 -33090 81750
rect -33020 81550 -32980 81750
rect -32910 81550 -32900 81750
rect -33100 81520 -32900 81550
rect -32600 81750 -32400 81780
rect -32600 81550 -32590 81750
rect -32520 81550 -32480 81750
rect -32410 81550 -32400 81750
rect -32600 81520 -32400 81550
rect -32100 81750 -31900 81780
rect -32100 81550 -32090 81750
rect -32020 81550 -31980 81750
rect -31910 81550 -31900 81750
rect -32100 81520 -31900 81550
rect -31600 81750 -31400 81780
rect -31600 81550 -31590 81750
rect -31520 81550 -31480 81750
rect -31410 81550 -31400 81750
rect -31600 81520 -31400 81550
rect -31100 81750 -30900 81780
rect -31100 81550 -31090 81750
rect -31020 81550 -30980 81750
rect -30910 81550 -30900 81750
rect -31100 81520 -30900 81550
rect -30600 81750 -30400 81780
rect -30600 81550 -30590 81750
rect -30520 81550 -30480 81750
rect -30410 81550 -30400 81750
rect -30600 81520 -30400 81550
rect -30100 81750 -29900 81780
rect -30100 81550 -30090 81750
rect -30020 81550 -29980 81750
rect -29910 81550 -29900 81750
rect -30100 81520 -29900 81550
rect -29600 81750 -29400 81780
rect -29600 81550 -29590 81750
rect -29520 81550 -29480 81750
rect -29410 81550 -29400 81750
rect -29600 81520 -29400 81550
rect -29100 81750 -28900 81780
rect -29100 81550 -29090 81750
rect -29020 81550 -28980 81750
rect -28910 81550 -28900 81750
rect -29100 81520 -28900 81550
rect -28600 81750 -28400 81780
rect -28600 81550 -28590 81750
rect -28520 81550 -28480 81750
rect -28410 81550 -28400 81750
rect -28600 81520 -28400 81550
rect -28100 81750 -27900 81780
rect -28100 81550 -28090 81750
rect -28020 81550 -27980 81750
rect -27910 81550 -27900 81750
rect -28100 81520 -27900 81550
rect -27600 81750 -27400 81780
rect -27600 81550 -27590 81750
rect -27520 81550 -27480 81750
rect -27410 81550 -27400 81750
rect -27600 81520 -27400 81550
rect -27100 81750 -26900 81780
rect -27100 81550 -27090 81750
rect -27020 81550 -26980 81750
rect -26910 81550 -26900 81750
rect -27100 81520 -26900 81550
rect -26600 81750 -26400 81780
rect -26600 81550 -26590 81750
rect -26520 81550 -26480 81750
rect -26410 81550 -26400 81750
rect -26600 81520 -26400 81550
rect -26100 81750 -25900 81780
rect -26100 81550 -26090 81750
rect -26020 81550 -25980 81750
rect -25910 81550 -25900 81750
rect -26100 81520 -25900 81550
rect -25600 81750 -25400 81780
rect -25600 81550 -25590 81750
rect -25520 81550 -25480 81750
rect -25410 81550 -25400 81750
rect -25600 81520 -25400 81550
rect -25100 81750 -24900 81780
rect -25100 81550 -25090 81750
rect -25020 81550 -24980 81750
rect -24910 81550 -24900 81750
rect -25100 81520 -24900 81550
rect -24600 81750 -24400 81780
rect -24600 81550 -24590 81750
rect -24520 81550 -24480 81750
rect -24410 81550 -24400 81750
rect -24600 81520 -24400 81550
rect -24100 81750 -23900 81780
rect -24100 81550 -24090 81750
rect -24020 81550 -23980 81750
rect -23910 81550 -23900 81750
rect -24100 81520 -23900 81550
rect -23600 81750 -23400 81780
rect -23600 81550 -23590 81750
rect -23520 81550 -23480 81750
rect -23410 81550 -23400 81750
rect -23600 81520 -23400 81550
rect -23100 81750 -22900 81780
rect -23100 81550 -23090 81750
rect -23020 81550 -22980 81750
rect -22910 81550 -22900 81750
rect -23100 81520 -22900 81550
rect -22600 81750 -22400 81780
rect -22600 81550 -22590 81750
rect -22520 81550 -22480 81750
rect -22410 81550 -22400 81750
rect -22600 81520 -22400 81550
rect -22100 81750 -21900 81780
rect -22100 81550 -22090 81750
rect -22020 81550 -21980 81750
rect -21910 81550 -21900 81750
rect -22100 81520 -21900 81550
rect -21600 81750 -21400 81780
rect -21600 81550 -21590 81750
rect -21520 81550 -21480 81750
rect -21410 81550 -21400 81750
rect -21600 81520 -21400 81550
rect -21100 81750 -20900 81780
rect -21100 81550 -21090 81750
rect -21020 81550 -20980 81750
rect -20910 81550 -20900 81750
rect -21100 81520 -20900 81550
rect -20600 81750 -20400 81780
rect -20600 81550 -20590 81750
rect -20520 81550 -20480 81750
rect -20410 81550 -20400 81750
rect -20600 81520 -20400 81550
rect -20100 81750 -19900 81780
rect -20100 81550 -20090 81750
rect -20020 81550 -19980 81750
rect -19910 81550 -19900 81750
rect -20100 81520 -19900 81550
rect -19600 81750 -19400 81780
rect -19600 81550 -19590 81750
rect -19520 81550 -19480 81750
rect -19410 81550 -19400 81750
rect -19600 81520 -19400 81550
rect -19100 81750 -18900 81780
rect -19100 81550 -19090 81750
rect -19020 81550 -18980 81750
rect -18910 81550 -18900 81750
rect -19100 81520 -18900 81550
rect -18600 81750 -18400 81780
rect -18600 81550 -18590 81750
rect -18520 81550 -18480 81750
rect -18410 81550 -18400 81750
rect -18600 81520 -18400 81550
rect -18100 81750 -17900 81780
rect -18100 81550 -18090 81750
rect -18020 81550 -17980 81750
rect -17910 81550 -17900 81750
rect -18100 81520 -17900 81550
rect -17600 81750 -17400 81780
rect -17600 81550 -17590 81750
rect -17520 81550 -17480 81750
rect -17410 81550 -17400 81750
rect -17600 81520 -17400 81550
rect -17100 81750 -16900 81780
rect -17100 81550 -17090 81750
rect -17020 81550 -16980 81750
rect -16910 81550 -16900 81750
rect -17100 81520 -16900 81550
rect -16600 81750 -16400 81780
rect -16600 81550 -16590 81750
rect -16520 81550 -16480 81750
rect -16410 81550 -16400 81750
rect -16600 81520 -16400 81550
rect -16100 81750 -15900 81780
rect -16100 81550 -16090 81750
rect -16020 81550 -15980 81750
rect -15910 81550 -15900 81750
rect -16100 81520 -15900 81550
rect -15600 81750 -15400 81780
rect -15600 81550 -15590 81750
rect -15520 81550 -15480 81750
rect -15410 81550 -15400 81750
rect -15600 81520 -15400 81550
rect -15100 81750 -14900 81780
rect -15100 81550 -15090 81750
rect -15020 81550 -14980 81750
rect -14910 81550 -14900 81750
rect -15100 81520 -14900 81550
rect -14600 81750 -14400 81780
rect -14600 81550 -14590 81750
rect -14520 81550 -14480 81750
rect -14410 81550 -14400 81750
rect -14600 81520 -14400 81550
rect -14100 81750 -13900 81780
rect -14100 81550 -14090 81750
rect -14020 81550 -13980 81750
rect -13910 81550 -13900 81750
rect -14100 81520 -13900 81550
rect -13600 81750 -13400 81780
rect -13600 81550 -13590 81750
rect -13520 81550 -13480 81750
rect -13410 81550 -13400 81750
rect -13600 81520 -13400 81550
rect -13100 81750 -12900 81780
rect -13100 81550 -13090 81750
rect -13020 81550 -12980 81750
rect -12910 81550 -12900 81750
rect -13100 81520 -12900 81550
rect -12600 81750 -12400 81780
rect -12600 81550 -12590 81750
rect -12520 81550 -12480 81750
rect -12410 81550 -12400 81750
rect -12600 81520 -12400 81550
rect -12100 81750 -11900 81780
rect -12100 81550 -12090 81750
rect -12020 81550 -11980 81750
rect -11910 81550 -11900 81750
rect -12100 81520 -11900 81550
rect -11600 81750 -11400 81780
rect -11600 81550 -11590 81750
rect -11520 81550 -11480 81750
rect -11410 81550 -11400 81750
rect -11600 81520 -11400 81550
rect -11100 81750 -10900 81780
rect -11100 81550 -11090 81750
rect -11020 81550 -10980 81750
rect -10910 81550 -10900 81750
rect -11100 81520 -10900 81550
rect -10600 81750 -10400 81780
rect -10600 81550 -10590 81750
rect -10520 81550 -10480 81750
rect -10410 81550 -10400 81750
rect -10600 81520 -10400 81550
rect -10100 81750 -9900 81780
rect -10100 81550 -10090 81750
rect -10020 81550 -9980 81750
rect -9910 81550 -9900 81750
rect -10100 81520 -9900 81550
rect -9600 81750 -9400 81780
rect -9600 81550 -9590 81750
rect -9520 81550 -9480 81750
rect -9410 81550 -9400 81750
rect -9600 81520 -9400 81550
rect -9100 81750 -8900 81780
rect -9100 81550 -9090 81750
rect -9020 81550 -8980 81750
rect -8910 81550 -8900 81750
rect -9100 81520 -8900 81550
rect -8600 81750 -8400 81780
rect -8600 81550 -8590 81750
rect -8520 81550 -8480 81750
rect -8410 81550 -8400 81750
rect -8600 81520 -8400 81550
rect -8100 81750 -7900 81780
rect -8100 81550 -8090 81750
rect -8020 81550 -7980 81750
rect -7910 81550 -7900 81750
rect -8100 81520 -7900 81550
rect -7600 81750 -7400 81780
rect -7600 81550 -7590 81750
rect -7520 81550 -7480 81750
rect -7410 81550 -7400 81750
rect -7600 81520 -7400 81550
rect -7100 81750 -6900 81780
rect -7100 81550 -7090 81750
rect -7020 81550 -6980 81750
rect -6910 81550 -6900 81750
rect -7100 81520 -6900 81550
rect -6600 81750 -6400 81780
rect -6600 81550 -6590 81750
rect -6520 81550 -6480 81750
rect -6410 81550 -6400 81750
rect -6600 81520 -6400 81550
rect -6100 81750 -5900 81780
rect -6100 81550 -6090 81750
rect -6020 81550 -5980 81750
rect -5910 81550 -5900 81750
rect -6100 81520 -5900 81550
rect -5600 81750 -5400 81780
rect -5600 81550 -5590 81750
rect -5520 81550 -5480 81750
rect -5410 81550 -5400 81750
rect -5600 81520 -5400 81550
rect -5100 81750 -4900 81780
rect -5100 81550 -5090 81750
rect -5020 81550 -4980 81750
rect -4910 81550 -4900 81750
rect -5100 81520 -4900 81550
rect -4600 81750 -4400 81780
rect -4600 81550 -4590 81750
rect -4520 81550 -4480 81750
rect -4410 81550 -4400 81750
rect -4600 81520 -4400 81550
rect -4100 81750 -3900 81780
rect -4100 81550 -4090 81750
rect -4020 81550 -3980 81750
rect -3910 81550 -3900 81750
rect -4100 81520 -3900 81550
rect -3600 81750 -3400 81780
rect -3600 81550 -3590 81750
rect -3520 81550 -3480 81750
rect -3410 81550 -3400 81750
rect -3600 81520 -3400 81550
rect -3100 81750 -2900 81780
rect -3100 81550 -3090 81750
rect -3020 81550 -2980 81750
rect -2910 81550 -2900 81750
rect -3100 81520 -2900 81550
rect -2600 81750 -2400 81780
rect -2600 81550 -2590 81750
rect -2520 81550 -2480 81750
rect -2410 81550 -2400 81750
rect -2600 81520 -2400 81550
rect -2100 81750 -1900 81780
rect -2100 81550 -2090 81750
rect -2020 81550 -1980 81750
rect -1910 81550 -1900 81750
rect -2100 81520 -1900 81550
rect -1600 81750 -1400 81780
rect -1600 81550 -1590 81750
rect -1520 81550 -1480 81750
rect -1410 81550 -1400 81750
rect -1600 81520 -1400 81550
rect -1100 81750 -900 81780
rect -1100 81550 -1090 81750
rect -1020 81550 -980 81750
rect -910 81550 -900 81750
rect -1100 81520 -900 81550
rect -600 81750 -400 81780
rect -600 81550 -590 81750
rect -520 81550 -480 81750
rect -410 81550 -400 81750
rect -600 81520 -400 81550
rect -100 81750 100 81780
rect -100 81550 -90 81750
rect -20 81550 20 81750
rect 90 81550 100 81750
rect -100 81520 100 81550
rect 400 81750 600 81780
rect 400 81550 410 81750
rect 480 81550 520 81750
rect 590 81550 600 81750
rect 400 81520 600 81550
rect 900 81750 1100 81780
rect 900 81550 910 81750
rect 980 81550 1020 81750
rect 1090 81550 1100 81750
rect 900 81520 1100 81550
rect 1400 81750 1600 81780
rect 1400 81550 1410 81750
rect 1480 81550 1520 81750
rect 1590 81550 1600 81750
rect 1400 81520 1600 81550
rect 1900 81750 2100 81780
rect 1900 81550 1910 81750
rect 1980 81550 2020 81750
rect 2090 81550 2100 81750
rect 1900 81520 2100 81550
rect 2400 81750 2600 81780
rect 2400 81550 2410 81750
rect 2480 81550 2520 81750
rect 2590 81550 2600 81750
rect 2400 81520 2600 81550
rect 2900 81750 3100 81780
rect 2900 81550 2910 81750
rect 2980 81550 3020 81750
rect 3090 81550 3100 81750
rect 2900 81520 3100 81550
rect 3400 81750 3600 81780
rect 3400 81550 3410 81750
rect 3480 81550 3520 81750
rect 3590 81550 3600 81750
rect 3400 81520 3600 81550
rect 3900 81750 4100 81780
rect 3900 81550 3910 81750
rect 3980 81550 4020 81750
rect 4090 81550 4100 81750
rect 3900 81520 4100 81550
rect 4400 81750 4600 81780
rect 4400 81550 4410 81750
rect 4480 81550 4520 81750
rect 4590 81550 4600 81750
rect 4400 81520 4600 81550
rect 4900 81750 5100 81780
rect 4900 81550 4910 81750
rect 4980 81550 5020 81750
rect 5090 81550 5100 81750
rect 4900 81520 5100 81550
rect 5400 81750 5600 81780
rect 5400 81550 5410 81750
rect 5480 81550 5520 81750
rect 5590 81550 5600 81750
rect 5400 81520 5600 81550
rect 5900 81750 6100 81780
rect 5900 81550 5910 81750
rect 5980 81550 6020 81750
rect 6090 81550 6100 81750
rect 5900 81520 6100 81550
rect 6400 81750 6600 81780
rect 6400 81550 6410 81750
rect 6480 81550 6520 81750
rect 6590 81550 6600 81750
rect 6400 81520 6600 81550
rect 6900 81750 7100 81780
rect 6900 81550 6910 81750
rect 6980 81550 7020 81750
rect 7090 81550 7100 81750
rect 6900 81520 7100 81550
rect 7400 81750 7600 81780
rect 7400 81550 7410 81750
rect 7480 81550 7520 81750
rect 7590 81550 7600 81750
rect 7400 81520 7600 81550
rect 7900 81750 8100 81780
rect 7900 81550 7910 81750
rect 7980 81550 8020 81750
rect 8090 81550 8100 81750
rect 7900 81520 8100 81550
rect 8400 81750 8600 81780
rect 8400 81550 8410 81750
rect 8480 81550 8520 81750
rect 8590 81550 8600 81750
rect 8400 81520 8600 81550
rect 8900 81750 9100 81780
rect 8900 81550 8910 81750
rect 8980 81550 9020 81750
rect 9090 81550 9100 81750
rect 8900 81520 9100 81550
rect 9400 81750 9600 81780
rect 9400 81550 9410 81750
rect 9480 81550 9520 81750
rect 9590 81550 9600 81750
rect 9400 81520 9600 81550
rect 9900 81750 10100 81780
rect 9900 81550 9910 81750
rect 9980 81550 10020 81750
rect 10090 81550 10100 81750
rect 9900 81520 10100 81550
rect 10400 81750 10600 81780
rect 10400 81550 10410 81750
rect 10480 81550 10520 81750
rect 10590 81550 10600 81750
rect 10400 81520 10600 81550
rect 10900 81750 11100 81780
rect 10900 81550 10910 81750
rect 10980 81550 11020 81750
rect 11090 81550 11100 81750
rect 10900 81520 11100 81550
rect 11400 81750 11600 81780
rect 11400 81550 11410 81750
rect 11480 81550 11520 81750
rect 11590 81550 11600 81750
rect 11400 81520 11600 81550
rect 11900 81750 12100 81780
rect 11900 81550 11910 81750
rect 11980 81550 12020 81750
rect 12090 81550 12100 81750
rect 11900 81520 12100 81550
rect 12400 81750 12600 81780
rect 12400 81550 12410 81750
rect 12480 81550 12520 81750
rect 12590 81550 12600 81750
rect 12400 81520 12600 81550
rect 12900 81750 13100 81780
rect 12900 81550 12910 81750
rect 12980 81550 13020 81750
rect 13090 81550 13100 81750
rect 12900 81520 13100 81550
rect 13400 81750 13600 81780
rect 13400 81550 13410 81750
rect 13480 81550 13520 81750
rect 13590 81550 13600 81750
rect 13400 81520 13600 81550
rect 13900 81750 14100 81780
rect 13900 81550 13910 81750
rect 13980 81550 14020 81750
rect 14090 81550 14100 81750
rect 13900 81520 14100 81550
rect 14400 81750 14600 81780
rect 14400 81550 14410 81750
rect 14480 81550 14520 81750
rect 14590 81550 14600 81750
rect 14400 81520 14600 81550
rect 14900 81750 15100 81780
rect 14900 81550 14910 81750
rect 14980 81550 15020 81750
rect 15090 81550 15100 81750
rect 14900 81520 15100 81550
rect 15400 81750 15600 81780
rect 15400 81550 15410 81750
rect 15480 81550 15520 81750
rect 15590 81550 15600 81750
rect 15400 81520 15600 81550
rect 15900 81750 16100 81780
rect 15900 81550 15910 81750
rect 15980 81550 16020 81750
rect 16090 81550 16100 81750
rect 15900 81520 16100 81550
rect 16400 81750 16600 81780
rect 16400 81550 16410 81750
rect 16480 81550 16520 81750
rect 16590 81550 16600 81750
rect 16400 81520 16600 81550
rect 16900 81750 17100 81780
rect 16900 81550 16910 81750
rect 16980 81550 17020 81750
rect 17090 81550 17100 81750
rect 16900 81520 17100 81550
rect 17400 81750 17600 81780
rect 17400 81550 17410 81750
rect 17480 81550 17520 81750
rect 17590 81550 17600 81750
rect 17400 81520 17600 81550
rect 17900 81750 18100 81780
rect 17900 81550 17910 81750
rect 17980 81550 18020 81750
rect 18090 81550 18100 81750
rect 17900 81520 18100 81550
rect 18400 81750 18600 81780
rect 18400 81550 18410 81750
rect 18480 81550 18520 81750
rect 18590 81550 18600 81750
rect 18400 81520 18600 81550
rect 18900 81750 19100 81780
rect 18900 81550 18910 81750
rect 18980 81550 19020 81750
rect 19090 81550 19100 81750
rect 18900 81520 19100 81550
rect 19400 81750 19600 81780
rect 19400 81550 19410 81750
rect 19480 81550 19520 81750
rect 19590 81550 19600 81750
rect 19400 81520 19600 81550
rect 19900 81750 20100 81780
rect 19900 81550 19910 81750
rect 19980 81550 20020 81750
rect 20090 81550 20100 81750
rect 19900 81520 20100 81550
rect 20400 81750 20600 81780
rect 20400 81550 20410 81750
rect 20480 81550 20520 81750
rect 20590 81550 20600 81750
rect 20400 81520 20600 81550
rect 20900 81750 21100 81780
rect 20900 81550 20910 81750
rect 20980 81550 21020 81750
rect 21090 81550 21100 81750
rect 20900 81520 21100 81550
rect 21400 81750 21600 81780
rect 21400 81550 21410 81750
rect 21480 81550 21520 81750
rect 21590 81550 21600 81750
rect 21400 81520 21600 81550
rect 21900 81750 22100 81780
rect 21900 81550 21910 81750
rect 21980 81550 22020 81750
rect 22090 81550 22100 81750
rect 21900 81520 22100 81550
rect 22400 81750 22600 81780
rect 22400 81550 22410 81750
rect 22480 81550 22520 81750
rect 22590 81550 22600 81750
rect 22400 81520 22600 81550
rect 22900 81750 23100 81780
rect 22900 81550 22910 81750
rect 22980 81550 23020 81750
rect 23090 81550 23100 81750
rect 22900 81520 23100 81550
rect 23400 81750 23600 81780
rect 23400 81550 23410 81750
rect 23480 81550 23520 81750
rect 23590 81550 23600 81750
rect 23400 81520 23600 81550
rect 23900 81750 24100 81780
rect 23900 81550 23910 81750
rect 23980 81550 24020 81750
rect 24090 81550 24100 81750
rect 23900 81520 24100 81550
rect 24400 81750 24600 81780
rect 24400 81550 24410 81750
rect 24480 81550 24520 81750
rect 24590 81550 24600 81750
rect 24400 81520 24600 81550
rect 24900 81750 25100 81780
rect 24900 81550 24910 81750
rect 24980 81550 25020 81750
rect 25090 81550 25100 81750
rect 24900 81520 25100 81550
rect 25400 81750 25600 81780
rect 25400 81550 25410 81750
rect 25480 81550 25520 81750
rect 25590 81550 25600 81750
rect 25400 81520 25600 81550
rect 25900 81750 26100 81780
rect 25900 81550 25910 81750
rect 25980 81550 26020 81750
rect 26090 81550 26100 81750
rect 25900 81520 26100 81550
rect 26400 81750 26600 81780
rect 26400 81550 26410 81750
rect 26480 81550 26520 81750
rect 26590 81550 26600 81750
rect 26400 81520 26600 81550
rect 26900 81750 27100 81780
rect 26900 81550 26910 81750
rect 26980 81550 27020 81750
rect 27090 81550 27100 81750
rect 26900 81520 27100 81550
rect 27400 81750 27600 81780
rect 27400 81550 27410 81750
rect 27480 81550 27520 81750
rect 27590 81550 27600 81750
rect 27400 81520 27600 81550
rect 27900 81750 28100 81780
rect 27900 81550 27910 81750
rect 27980 81550 28020 81750
rect 28090 81550 28100 81750
rect 27900 81520 28100 81550
rect 28400 81750 28600 81780
rect 28400 81550 28410 81750
rect 28480 81550 28520 81750
rect 28590 81550 28600 81750
rect 28400 81520 28600 81550
rect 28900 81750 29100 81780
rect 28900 81550 28910 81750
rect 28980 81550 29020 81750
rect 29090 81550 29100 81750
rect 28900 81520 29100 81550
rect 29400 81750 29600 81780
rect 29400 81550 29410 81750
rect 29480 81550 29520 81750
rect 29590 81550 29600 81750
rect 29400 81520 29600 81550
rect 29900 81750 30100 81780
rect 29900 81550 29910 81750
rect 29980 81550 30020 81750
rect 30090 81550 30100 81750
rect 29900 81520 30100 81550
rect 30400 81750 30600 81780
rect 30400 81550 30410 81750
rect 30480 81550 30520 81750
rect 30590 81550 30600 81750
rect 30400 81520 30600 81550
rect 30900 81750 31100 81780
rect 30900 81550 30910 81750
rect 30980 81550 31020 81750
rect 31090 81550 31100 81750
rect 30900 81520 31100 81550
rect 31400 81750 31600 81780
rect 31400 81550 31410 81750
rect 31480 81550 31520 81750
rect 31590 81550 31600 81750
rect 31400 81520 31600 81550
rect 31900 81750 32100 81780
rect 31900 81550 31910 81750
rect 31980 81550 32020 81750
rect 32090 81550 32100 81750
rect 31900 81520 32100 81550
rect 32400 81750 32600 81780
rect 32400 81550 32410 81750
rect 32480 81550 32520 81750
rect 32590 81550 32600 81750
rect 32400 81520 32600 81550
rect 32900 81750 33100 81780
rect 32900 81550 32910 81750
rect 32980 81550 33020 81750
rect 33090 81550 33100 81750
rect 32900 81520 33100 81550
rect 33400 81750 33600 81780
rect 33400 81550 33410 81750
rect 33480 81550 33520 81750
rect 33590 81550 33600 81750
rect 33400 81520 33600 81550
rect 33900 81750 34100 81780
rect 33900 81550 33910 81750
rect 33980 81550 34020 81750
rect 34090 81550 34100 81750
rect 33900 81520 34100 81550
rect 34400 81750 34600 81780
rect 34400 81550 34410 81750
rect 34480 81550 34520 81750
rect 34590 81550 34600 81750
rect 34400 81520 34600 81550
rect 34900 81750 35100 81780
rect 34900 81550 34910 81750
rect 34980 81550 35020 81750
rect 35090 81550 35100 81750
rect 34900 81520 35100 81550
rect 35400 81750 35600 81780
rect 35400 81550 35410 81750
rect 35480 81550 35520 81750
rect 35590 81550 35600 81750
rect 35400 81520 35600 81550
rect 35900 81750 36100 81780
rect 35900 81550 35910 81750
rect 35980 81550 36020 81750
rect 36090 81550 36100 81750
rect 35900 81520 36100 81550
rect 36400 81750 36600 81780
rect 36400 81550 36410 81750
rect 36480 81550 36520 81750
rect 36590 81550 36600 81750
rect 36400 81520 36600 81550
rect 36900 81750 37100 81780
rect 36900 81550 36910 81750
rect 36980 81550 37020 81750
rect 37090 81550 37100 81750
rect 36900 81520 37100 81550
rect 37400 81750 37600 81780
rect 37400 81550 37410 81750
rect 37480 81550 37520 81750
rect 37590 81550 37600 81750
rect 37400 81520 37600 81550
rect 37900 81750 38100 81780
rect 37900 81550 37910 81750
rect 37980 81550 38020 81750
rect 38090 81550 38100 81750
rect 37900 81520 38100 81550
rect 38400 81750 38600 81780
rect 38400 81550 38410 81750
rect 38480 81550 38520 81750
rect 38590 81550 38600 81750
rect 38400 81520 38600 81550
rect 38900 81750 39100 81780
rect 38900 81550 38910 81750
rect 38980 81550 39020 81750
rect 39090 81550 39100 81750
rect 38900 81520 39100 81550
rect 39400 81750 39600 81780
rect 39400 81550 39410 81750
rect 39480 81550 39520 81750
rect 39590 81550 39600 81750
rect 39400 81520 39600 81550
rect 39900 81750 40100 81780
rect 39900 81550 39910 81750
rect 39980 81550 40020 81750
rect 40090 81550 40100 81750
rect 39900 81520 40100 81550
rect 40400 81750 40600 81780
rect 40400 81550 40410 81750
rect 40480 81550 40520 81750
rect 40590 81550 40600 81750
rect 40400 81520 40600 81550
rect 40900 81750 41100 81780
rect 40900 81550 40910 81750
rect 40980 81550 41020 81750
rect 41090 81550 41100 81750
rect 40900 81520 41100 81550
rect 41400 81750 41600 81780
rect 41400 81550 41410 81750
rect 41480 81550 41520 81750
rect 41590 81550 41600 81750
rect 41400 81520 41600 81550
rect 41900 81750 42100 81780
rect 41900 81550 41910 81750
rect 41980 81550 42020 81750
rect 42090 81550 42100 81750
rect 41900 81520 42100 81550
rect 42400 81750 42600 81780
rect 42400 81550 42410 81750
rect 42480 81550 42520 81750
rect 42590 81550 42600 81750
rect 42400 81520 42600 81550
rect 42900 81750 43100 81780
rect 42900 81550 42910 81750
rect 42980 81550 43020 81750
rect 43090 81550 43100 81750
rect 42900 81520 43100 81550
rect 43400 81750 43600 81780
rect 43400 81550 43410 81750
rect 43480 81550 43520 81750
rect 43590 81550 43600 81750
rect 43400 81520 43600 81550
rect 43900 81750 44100 81780
rect 43900 81550 43910 81750
rect 43980 81550 44020 81750
rect 44090 81550 44100 81750
rect 43900 81520 44100 81550
rect 44400 81750 44600 81780
rect 44400 81550 44410 81750
rect 44480 81550 44520 81750
rect 44590 81550 44600 81750
rect 44400 81520 44600 81550
rect 44900 81750 45100 81780
rect 44900 81550 44910 81750
rect 44980 81550 45020 81750
rect 45090 81550 45100 81750
rect 44900 81520 45100 81550
rect 45400 81750 45600 81780
rect 45400 81550 45410 81750
rect 45480 81550 45520 81750
rect 45590 81550 45600 81750
rect 45400 81520 45600 81550
rect 45900 81750 46100 81780
rect 45900 81550 45910 81750
rect 45980 81550 46020 81750
rect 46090 81550 46100 81750
rect 45900 81520 46100 81550
rect 46400 81750 46600 81780
rect 46400 81550 46410 81750
rect 46480 81550 46520 81750
rect 46590 81550 46600 81750
rect 46400 81520 46600 81550
rect 46900 81750 47100 81780
rect 46900 81550 46910 81750
rect 46980 81550 47020 81750
rect 47090 81550 47100 81750
rect 46900 81520 47100 81550
rect 47400 81750 47600 81780
rect 47400 81550 47410 81750
rect 47480 81550 47520 81750
rect 47590 81550 47600 81750
rect 47400 81520 47600 81550
rect 47900 81750 48100 81780
rect 47900 81550 47910 81750
rect 47980 81550 48020 81750
rect 48090 81550 48100 81750
rect 47900 81520 48100 81550
rect 48400 81750 48600 81780
rect 48400 81550 48410 81750
rect 48480 81550 48520 81750
rect 48590 81550 48600 81750
rect 48400 81520 48600 81550
rect 48900 81750 49100 81780
rect 48900 81550 48910 81750
rect 48980 81550 49020 81750
rect 49090 81550 49100 81750
rect 48900 81520 49100 81550
rect 49400 81750 49600 81780
rect 49400 81550 49410 81750
rect 49480 81550 49520 81750
rect 49590 81550 49600 81750
rect 49400 81520 49600 81550
rect 49900 81750 50100 81780
rect 49900 81550 49910 81750
rect 49980 81550 50020 81750
rect 50090 81550 50100 81750
rect 49900 81520 50100 81550
rect 50400 81750 50600 81780
rect 50400 81550 50410 81750
rect 50480 81550 50520 81750
rect 50590 81550 50600 81750
rect 50400 81520 50600 81550
rect 50900 81750 51100 81780
rect 50900 81550 50910 81750
rect 50980 81550 51020 81750
rect 51090 81550 51100 81750
rect 50900 81520 51100 81550
rect 51400 81750 51600 81780
rect 51400 81550 51410 81750
rect 51480 81550 51520 81750
rect 51590 81550 51600 81750
rect 51400 81520 51600 81550
rect 51900 81750 52100 81780
rect 51900 81550 51910 81750
rect 51980 81550 52020 81750
rect 52090 81550 52100 81750
rect 51900 81520 52100 81550
rect 52400 81750 52600 81780
rect 52400 81550 52410 81750
rect 52480 81550 52520 81750
rect 52590 81550 52600 81750
rect 52400 81520 52600 81550
rect 52900 81750 53100 81780
rect 52900 81550 52910 81750
rect 52980 81550 53020 81750
rect 53090 81550 53100 81750
rect 52900 81520 53100 81550
rect 53400 81750 53600 81780
rect 53400 81550 53410 81750
rect 53480 81550 53520 81750
rect 53590 81550 53600 81750
rect 53400 81520 53600 81550
rect 53900 81750 54100 81780
rect 53900 81550 53910 81750
rect 53980 81550 54020 81750
rect 54090 81550 54100 81750
rect 53900 81520 54100 81550
rect 54400 81750 54600 81780
rect 54400 81550 54410 81750
rect 54480 81550 54520 81750
rect 54590 81550 54600 81750
rect 54400 81520 54600 81550
rect 54900 81750 55100 81780
rect 54900 81550 54910 81750
rect 54980 81550 55020 81750
rect 55090 81550 55100 81750
rect 54900 81520 55100 81550
rect 55400 81750 55600 81780
rect 55400 81550 55410 81750
rect 55480 81550 55520 81750
rect 55590 81550 55600 81750
rect 55400 81520 55600 81550
rect 55900 81750 56100 81780
rect 55900 81550 55910 81750
rect 55980 81550 56020 81750
rect 56090 81550 56100 81750
rect 55900 81520 56100 81550
rect 56400 81750 56600 81780
rect 56400 81550 56410 81750
rect 56480 81550 56520 81750
rect 56590 81550 56600 81750
rect 56400 81520 56600 81550
rect 56900 81750 57100 81780
rect 56900 81550 56910 81750
rect 56980 81550 57020 81750
rect 57090 81550 57100 81750
rect 56900 81520 57100 81550
rect 57400 81750 57600 81780
rect 57400 81550 57410 81750
rect 57480 81550 57520 81750
rect 57590 81550 57600 81750
rect 57400 81520 57600 81550
rect 57900 81750 58100 81780
rect 57900 81550 57910 81750
rect 57980 81550 58020 81750
rect 58090 81550 58100 81750
rect 57900 81520 58100 81550
rect 58400 81750 58600 81780
rect 58400 81550 58410 81750
rect 58480 81550 58520 81750
rect 58590 81550 58600 81750
rect 58400 81520 58600 81550
rect 58900 81750 59100 81780
rect 58900 81550 58910 81750
rect 58980 81550 59020 81750
rect 59090 81550 59100 81750
rect 58900 81520 59100 81550
rect 59400 81750 59600 81780
rect 59400 81550 59410 81750
rect 59480 81550 59520 81750
rect 59590 81550 59600 81750
rect 59400 81520 59600 81550
rect 59900 81750 60100 81780
rect 59900 81550 59910 81750
rect 59980 81550 60020 81750
rect 60090 81550 60100 81750
rect 59900 81520 60100 81550
rect 60400 81750 60600 81780
rect 60400 81550 60410 81750
rect 60480 81550 60520 81750
rect 60590 81550 60600 81750
rect 60400 81520 60600 81550
rect 60900 81750 61100 81780
rect 60900 81550 60910 81750
rect 60980 81550 61020 81750
rect 61090 81550 61100 81750
rect 60900 81520 61100 81550
rect 61400 81750 61600 81780
rect 61400 81550 61410 81750
rect 61480 81550 61520 81750
rect 61590 81550 61600 81750
rect 61400 81520 61600 81550
rect 61900 81750 62100 81780
rect 61900 81550 61910 81750
rect 61980 81550 62020 81750
rect 62090 81550 62100 81750
rect 61900 81520 62100 81550
rect 62400 81750 62600 81780
rect 62400 81550 62410 81750
rect 62480 81550 62520 81750
rect 62590 81550 62600 81750
rect 62400 81520 62600 81550
rect 62900 81750 63100 81780
rect 62900 81550 62910 81750
rect 62980 81550 63020 81750
rect 63090 81550 63100 81750
rect 62900 81520 63100 81550
rect 63400 81750 63600 81780
rect 63400 81550 63410 81750
rect 63480 81550 63520 81750
rect 63590 81550 63600 81750
rect 63400 81520 63600 81550
rect 63900 81750 64100 81780
rect 63900 81550 63910 81750
rect 63980 81550 64020 81750
rect 64090 81550 64100 81750
rect 63900 81520 64100 81550
rect 64400 81750 64600 81780
rect 64400 81550 64410 81750
rect 64480 81550 64520 81750
rect 64590 81550 64600 81750
rect 64400 81520 64600 81550
rect 64900 81750 65100 81780
rect 64900 81550 64910 81750
rect 64980 81550 65020 81750
rect 65090 81550 65100 81750
rect 64900 81520 65100 81550
rect 65400 81750 65600 81780
rect 65400 81550 65410 81750
rect 65480 81550 65520 81750
rect 65590 81550 65600 81750
rect 65400 81520 65600 81550
rect 65900 81750 66100 81780
rect 65900 81550 65910 81750
rect 65980 81550 66020 81750
rect 66090 81550 66100 81750
rect 65900 81520 66100 81550
rect 66400 81750 66600 81780
rect 66400 81550 66410 81750
rect 66480 81550 66520 81750
rect 66590 81550 66600 81750
rect 66400 81520 66600 81550
rect 66900 81750 67100 81780
rect 66900 81550 66910 81750
rect 66980 81550 67020 81750
rect 67090 81550 67100 81750
rect 66900 81520 67100 81550
rect 67400 81750 67600 81780
rect 67400 81550 67410 81750
rect 67480 81550 67520 81750
rect 67590 81550 67600 81750
rect 67400 81520 67600 81550
rect 67900 81750 68100 81780
rect 67900 81550 67910 81750
rect 67980 81550 68020 81750
rect 68090 81550 68100 81750
rect 67900 81520 68100 81550
rect 68400 81750 68600 81780
rect 68400 81550 68410 81750
rect 68480 81550 68520 81750
rect 68590 81550 68600 81750
rect 68400 81520 68600 81550
rect 68900 81750 69100 81780
rect 68900 81550 68910 81750
rect 68980 81550 69020 81750
rect 69090 81550 69100 81750
rect 68900 81520 69100 81550
rect 69400 81750 69600 81780
rect 69400 81550 69410 81750
rect 69480 81550 69520 81750
rect 69590 81550 69600 81750
rect 69400 81520 69600 81550
rect 69900 81750 70100 81780
rect 69900 81550 69910 81750
rect 69980 81550 70020 81750
rect 70090 81550 70100 81750
rect 69900 81520 70100 81550
rect 70400 81750 70600 81780
rect 70400 81550 70410 81750
rect 70480 81550 70520 81750
rect 70590 81550 70600 81750
rect 70400 81520 70600 81550
rect 70900 81750 71100 81780
rect 70900 81550 70910 81750
rect 70980 81550 71020 81750
rect 71090 81550 71100 81750
rect 70900 81520 71100 81550
rect 71400 81750 71600 81780
rect 71400 81550 71410 81750
rect 71480 81550 71520 81750
rect 71590 81550 71600 81750
rect 71400 81520 71600 81550
rect 71900 81750 72100 81780
rect 71900 81550 71910 81750
rect 71980 81550 72020 81750
rect 72090 81550 72100 81750
rect 71900 81520 72100 81550
rect 72400 81750 72600 81780
rect 72400 81550 72410 81750
rect 72480 81550 72520 81750
rect 72590 81550 72600 81750
rect 72400 81520 72600 81550
rect 72900 81750 73100 81780
rect 72900 81550 72910 81750
rect 72980 81550 73020 81750
rect 73090 81550 73100 81750
rect 72900 81520 73100 81550
rect 73400 81750 73600 81780
rect 73400 81550 73410 81750
rect 73480 81550 73520 81750
rect 73590 81550 73600 81750
rect 73400 81520 73600 81550
rect 73900 81750 74100 81780
rect 73900 81550 73910 81750
rect 73980 81550 74020 81750
rect 74090 81550 74100 81750
rect 73900 81520 74100 81550
rect 74400 81750 74600 81780
rect 74400 81550 74410 81750
rect 74480 81550 74520 81750
rect 74590 81550 74600 81750
rect 74400 81520 74600 81550
rect 74900 81750 75100 81780
rect 74900 81550 74910 81750
rect 74980 81550 75020 81750
rect 75090 81550 75100 81750
rect 74900 81520 75100 81550
rect 75400 81750 75600 81780
rect 75400 81550 75410 81750
rect 75480 81550 75520 81750
rect 75590 81550 75600 81750
rect 75400 81520 75600 81550
rect 75900 81750 76100 81780
rect 75900 81550 75910 81750
rect 75980 81550 76020 81750
rect 76090 81550 76100 81750
rect 75900 81520 76100 81550
rect 76400 81750 76600 81780
rect 76400 81550 76410 81750
rect 76480 81550 76520 81750
rect 76590 81550 76600 81750
rect 76400 81520 76600 81550
rect 76900 81750 77100 81780
rect 76900 81550 76910 81750
rect 76980 81550 77020 81750
rect 77090 81550 77100 81750
rect 76900 81520 77100 81550
rect 77400 81750 77600 81780
rect 77400 81550 77410 81750
rect 77480 81550 77520 81750
rect 77590 81550 77600 81750
rect 77400 81520 77600 81550
rect 77900 81750 78100 81780
rect 77900 81550 77910 81750
rect 77980 81550 78020 81750
rect 78090 81550 78100 81750
rect 77900 81520 78100 81550
rect 78400 81750 78600 81780
rect 78400 81550 78410 81750
rect 78480 81550 78520 81750
rect 78590 81550 78600 81750
rect 78400 81520 78600 81550
rect 78900 81750 79100 81780
rect 78900 81550 78910 81750
rect 78980 81550 79020 81750
rect 79090 81550 79100 81750
rect 78900 81520 79100 81550
rect 79400 81750 79600 81780
rect 79400 81550 79410 81750
rect 79480 81550 79520 81750
rect 79590 81550 79600 81750
rect 79400 81520 79600 81550
rect 79900 81750 80100 81780
rect 79900 81550 79910 81750
rect 79980 81550 80020 81750
rect 80090 81550 80100 81750
rect 79900 81520 80100 81550
rect 80400 81750 80600 81780
rect 80400 81550 80410 81750
rect 80480 81550 80520 81750
rect 80590 81550 80600 81750
rect 80400 81520 80600 81550
rect 80900 81750 81100 81780
rect 80900 81550 80910 81750
rect 80980 81550 81020 81750
rect 81090 81550 81100 81750
rect 80900 81520 81100 81550
rect 81400 81750 81600 81780
rect 81400 81550 81410 81750
rect 81480 81550 81520 81750
rect 81590 81550 81600 81750
rect 81400 81520 81600 81550
rect 81900 81750 82100 81780
rect 81900 81550 81910 81750
rect 81980 81550 82020 81750
rect 82090 81550 82100 81750
rect 81900 81520 82100 81550
rect 82400 81750 82600 81780
rect 82400 81550 82410 81750
rect 82480 81550 82520 81750
rect 82590 81550 82600 81750
rect 82400 81520 82600 81550
rect 82900 81750 83100 81780
rect 82900 81550 82910 81750
rect 82980 81550 83020 81750
rect 83090 81550 83100 81750
rect 82900 81520 83100 81550
rect 83400 81750 83600 81780
rect 83400 81550 83410 81750
rect 83480 81550 83520 81750
rect 83590 81550 83600 81750
rect 83400 81520 83600 81550
rect 83900 81750 84100 81780
rect 83900 81550 83910 81750
rect 83980 81550 84020 81750
rect 84090 81550 84100 81750
rect 83900 81520 84100 81550
rect 84400 81750 84600 81780
rect 84400 81550 84410 81750
rect 84480 81550 84520 81750
rect 84590 81550 84600 81750
rect 84400 81520 84600 81550
rect 84900 81750 85100 81780
rect 84900 81550 84910 81750
rect 84980 81550 85020 81750
rect 85090 81550 85100 81750
rect 84900 81520 85100 81550
rect 85400 81750 85600 81780
rect 85400 81550 85410 81750
rect 85480 81550 85520 81750
rect 85590 81550 85600 81750
rect 85400 81520 85600 81550
rect 85900 81750 86100 81780
rect 85900 81550 85910 81750
rect 85980 81550 86020 81750
rect 86090 81550 86100 81750
rect 85900 81520 86100 81550
rect 86400 81750 86600 81780
rect 86400 81550 86410 81750
rect 86480 81550 86520 81750
rect 86590 81550 86600 81750
rect 86400 81520 86600 81550
rect 86900 81750 87100 81780
rect 86900 81550 86910 81750
rect 86980 81550 87020 81750
rect 87090 81550 87100 81750
rect 86900 81520 87100 81550
rect 87400 81750 87600 81780
rect 87400 81550 87410 81750
rect 87480 81550 87520 81750
rect 87590 81550 87600 81750
rect 87400 81520 87600 81550
rect 87900 81750 88100 81780
rect 87900 81550 87910 81750
rect 87980 81550 88020 81750
rect 88090 81550 88100 81750
rect 87900 81520 88100 81550
rect 88400 81750 88600 81780
rect 88400 81550 88410 81750
rect 88480 81550 88520 81750
rect 88590 81550 88600 81750
rect 88400 81520 88600 81550
rect 88900 81750 89100 81780
rect 88900 81550 88910 81750
rect 88980 81550 89020 81750
rect 89090 81550 89100 81750
rect 88900 81520 89100 81550
rect 89400 81750 89600 81780
rect 89400 81550 89410 81750
rect 89480 81550 89520 81750
rect 89590 81550 89600 81750
rect 89400 81520 89600 81550
rect 89900 81750 90100 81780
rect 89900 81550 89910 81750
rect 89980 81550 90020 81750
rect 90090 81550 90100 81750
rect 89900 81520 90100 81550
rect 90400 81750 90600 81780
rect 90400 81550 90410 81750
rect 90480 81550 90520 81750
rect 90590 81550 90600 81750
rect 90400 81520 90600 81550
rect 90900 81750 91100 81780
rect 90900 81550 90910 81750
rect 90980 81550 91020 81750
rect 91090 81550 91100 81750
rect 90900 81520 91100 81550
rect 91400 81750 91600 81780
rect 91400 81550 91410 81750
rect 91480 81550 91520 81750
rect 91590 81550 91600 81750
rect 91400 81520 91600 81550
rect 91900 81750 92100 81780
rect 91900 81550 91910 81750
rect 91980 81550 92020 81750
rect 92090 81550 92100 81750
rect 91900 81520 92100 81550
rect 92400 81750 92600 81780
rect 92400 81550 92410 81750
rect 92480 81550 92520 81750
rect 92590 81550 92600 81750
rect 92400 81520 92600 81550
rect 92900 81750 93100 81780
rect 92900 81550 92910 81750
rect 92980 81550 93020 81750
rect 93090 81550 93100 81750
rect 92900 81520 93100 81550
rect 93400 81750 93600 81780
rect 93400 81550 93410 81750
rect 93480 81550 93520 81750
rect 93590 81550 93600 81750
rect 93400 81520 93600 81550
rect 93900 81750 94100 81780
rect 93900 81550 93910 81750
rect 93980 81550 94020 81750
rect 94090 81550 94100 81750
rect 93900 81520 94100 81550
rect 94400 81750 94600 81780
rect 94400 81550 94410 81750
rect 94480 81550 94520 81750
rect 94590 81550 94600 81750
rect 94400 81520 94600 81550
rect 94900 81750 95100 81780
rect 94900 81550 94910 81750
rect 94980 81550 95020 81750
rect 95090 81550 95100 81750
rect 94900 81520 95100 81550
rect 95400 81750 95600 81780
rect 95400 81550 95410 81750
rect 95480 81550 95520 81750
rect 95590 81550 95600 81750
rect 95400 81520 95600 81550
rect 95900 81750 96100 81780
rect 95900 81550 95910 81750
rect 95980 81550 96020 81750
rect 96090 81550 96100 81750
rect 95900 81520 96100 81550
rect 96400 81750 96600 81780
rect 96400 81550 96410 81750
rect 96480 81550 96520 81750
rect 96590 81550 96600 81750
rect 96400 81520 96600 81550
rect 96900 81750 97100 81780
rect 96900 81550 96910 81750
rect 96980 81550 97020 81750
rect 97090 81550 97100 81750
rect 96900 81520 97100 81550
rect 97400 81750 97600 81780
rect 97400 81550 97410 81750
rect 97480 81550 97520 81750
rect 97590 81550 97600 81750
rect 97400 81520 97600 81550
rect 97900 81750 98100 81780
rect 97900 81550 97910 81750
rect 97980 81550 98020 81750
rect 98090 81550 98100 81750
rect 97900 81520 98100 81550
rect 98400 81750 98600 81780
rect 98400 81550 98410 81750
rect 98480 81550 98520 81750
rect 98590 81550 98600 81750
rect 98400 81520 98600 81550
rect 98900 81750 99100 81780
rect 98900 81550 98910 81750
rect 98980 81550 99020 81750
rect 99090 81550 99100 81750
rect 98900 81520 99100 81550
rect 99400 81750 99600 81780
rect 99400 81550 99410 81750
rect 99480 81550 99520 81750
rect 99590 81550 99600 81750
rect 99400 81520 99600 81550
rect 99900 81750 100100 81780
rect 99900 81550 99910 81750
rect 99980 81550 100020 81750
rect 100090 81550 100100 81750
rect 99900 81520 100100 81550
rect 100400 81750 100500 81780
rect 100400 81550 100410 81750
rect 100480 81550 100500 81750
rect 100400 81520 100500 81550
rect -83500 81500 -83380 81520
rect -83120 81500 -82880 81520
rect -82620 81500 -82380 81520
rect -82120 81500 -81880 81520
rect -81620 81500 -81380 81520
rect -81120 81500 -80880 81520
rect -80620 81500 -80380 81520
rect -80120 81500 -79880 81520
rect -79620 81500 -79380 81520
rect -79120 81500 -78880 81520
rect -78620 81500 -78380 81520
rect -78120 81500 -77880 81520
rect -77620 81500 -77380 81520
rect -77120 81500 -76880 81520
rect -76620 81500 -76380 81520
rect -76120 81500 -75880 81520
rect -75620 81500 -75380 81520
rect -75120 81500 -74880 81520
rect -74620 81500 -74380 81520
rect -74120 81500 -73880 81520
rect -73620 81500 -73380 81520
rect -73120 81500 -72880 81520
rect -72620 81500 -72380 81520
rect -72120 81500 -71880 81520
rect -71620 81500 -71380 81520
rect -71120 81500 -70880 81520
rect -70620 81500 -70380 81520
rect -70120 81500 -69880 81520
rect -69620 81500 -69380 81520
rect -69120 81500 -68880 81520
rect -68620 81500 -68380 81520
rect -68120 81500 -67880 81520
rect -67620 81500 -67380 81520
rect -67120 81500 -66880 81520
rect -66620 81500 -66380 81520
rect -66120 81500 -65880 81520
rect -65620 81500 -65380 81520
rect -65120 81500 -64880 81520
rect -64620 81500 -64380 81520
rect -64120 81500 -63880 81520
rect -63620 81500 -63380 81520
rect -63120 81500 -62880 81520
rect -62620 81500 -62380 81520
rect -62120 81500 -61880 81520
rect -61620 81500 -61380 81520
rect -61120 81500 -60880 81520
rect -60620 81500 -60380 81520
rect -60120 81500 -59880 81520
rect -59620 81500 -59380 81520
rect -59120 81500 -58880 81520
rect -58620 81500 -58380 81520
rect -58120 81500 -57880 81520
rect -57620 81500 -57380 81520
rect -57120 81500 -56880 81520
rect -56620 81500 -56380 81520
rect -56120 81500 -55880 81520
rect -55620 81500 -55380 81520
rect -55120 81500 -54880 81520
rect -54620 81500 -54380 81520
rect -54120 81500 -53880 81520
rect -53620 81500 -53380 81520
rect -53120 81500 -52880 81520
rect -52620 81500 -52380 81520
rect -52120 81500 -51880 81520
rect -51620 81500 -51380 81520
rect -51120 81500 -50880 81520
rect -50620 81500 -50380 81520
rect -50120 81500 -49880 81520
rect -49620 81500 -49380 81520
rect -49120 81500 -48880 81520
rect -48620 81500 -48380 81520
rect -48120 81500 -47880 81520
rect -47620 81500 -47380 81520
rect -47120 81500 -46880 81520
rect -46620 81500 -46380 81520
rect -46120 81500 -45880 81520
rect -45620 81500 -45380 81520
rect -45120 81500 -44880 81520
rect -44620 81500 -44380 81520
rect -44120 81500 -43880 81520
rect -43620 81500 -43380 81520
rect -43120 81500 -42880 81520
rect -42620 81500 -42380 81520
rect -42120 81500 -41880 81520
rect -41620 81500 -41380 81520
rect -41120 81500 -40880 81520
rect -40620 81500 -40380 81520
rect -40120 81500 -39880 81520
rect -39620 81500 -39380 81520
rect -39120 81500 -38880 81520
rect -38620 81500 -38380 81520
rect -38120 81500 -37880 81520
rect -37620 81500 -37380 81520
rect -37120 81500 -36880 81520
rect -36620 81500 -36380 81520
rect -36120 81500 -35880 81520
rect -35620 81500 -35380 81520
rect -35120 81500 -34880 81520
rect -34620 81500 -34380 81520
rect -34120 81500 -33880 81520
rect -33620 81500 -33380 81520
rect -33120 81500 -32880 81520
rect -32620 81500 -32380 81520
rect -32120 81500 -31880 81520
rect -31620 81500 -31380 81520
rect -31120 81500 -30880 81520
rect -30620 81500 -30380 81520
rect -30120 81500 -29880 81520
rect -29620 81500 -29380 81520
rect -29120 81500 -28880 81520
rect -28620 81500 -28380 81520
rect -28120 81500 -27880 81520
rect -27620 81500 -27380 81520
rect -27120 81500 -26880 81520
rect -26620 81500 -26380 81520
rect -26120 81500 -25880 81520
rect -25620 81500 -25380 81520
rect -25120 81500 -24880 81520
rect -24620 81500 -24380 81520
rect -24120 81500 -23880 81520
rect -23620 81500 -23380 81520
rect -23120 81500 -22880 81520
rect -22620 81500 -22380 81520
rect -22120 81500 -21880 81520
rect -21620 81500 -21380 81520
rect -21120 81500 -20880 81520
rect -20620 81500 -20380 81520
rect -20120 81500 -19880 81520
rect -19620 81500 -19380 81520
rect -19120 81500 -18880 81520
rect -18620 81500 -18380 81520
rect -18120 81500 -17880 81520
rect -17620 81500 -17380 81520
rect -17120 81500 -16880 81520
rect -16620 81500 -16380 81520
rect -16120 81500 -15880 81520
rect -15620 81500 -15380 81520
rect -15120 81500 -14880 81520
rect -14620 81500 -14380 81520
rect -14120 81500 -13880 81520
rect -13620 81500 -13380 81520
rect -13120 81500 -12880 81520
rect -12620 81500 -12380 81520
rect -12120 81500 -11880 81520
rect -11620 81500 -11380 81520
rect -11120 81500 -10880 81520
rect -10620 81500 -10380 81520
rect -10120 81500 -9880 81520
rect -9620 81500 -9380 81520
rect -9120 81500 -8880 81520
rect -8620 81500 -8380 81520
rect -8120 81500 -7880 81520
rect -7620 81500 -7380 81520
rect -7120 81500 -6880 81520
rect -6620 81500 -6380 81520
rect -6120 81500 -5880 81520
rect -5620 81500 -5380 81520
rect -5120 81500 -4880 81520
rect -4620 81500 -4380 81520
rect -4120 81500 -3880 81520
rect -3620 81500 -3380 81520
rect -3120 81500 -2880 81520
rect -2620 81500 -2380 81520
rect -2120 81500 -1880 81520
rect -1620 81500 -1380 81520
rect -1120 81500 -880 81520
rect -620 81500 -380 81520
rect -120 81500 120 81520
rect 380 81500 620 81520
rect 880 81500 1120 81520
rect 1380 81500 1620 81520
rect 1880 81500 2120 81520
rect 2380 81500 2620 81520
rect 2880 81500 3120 81520
rect 3380 81500 3620 81520
rect 3880 81500 4120 81520
rect 4380 81500 4620 81520
rect 4880 81500 5120 81520
rect 5380 81500 5620 81520
rect 5880 81500 6120 81520
rect 6380 81500 6620 81520
rect 6880 81500 7120 81520
rect 7380 81500 7620 81520
rect 7880 81500 8120 81520
rect 8380 81500 8620 81520
rect 8880 81500 9120 81520
rect 9380 81500 9620 81520
rect 9880 81500 10120 81520
rect 10380 81500 10620 81520
rect 10880 81500 11120 81520
rect 11380 81500 11620 81520
rect 11880 81500 12120 81520
rect 12380 81500 12620 81520
rect 12880 81500 13120 81520
rect 13380 81500 13620 81520
rect 13880 81500 14120 81520
rect 14380 81500 14620 81520
rect 14880 81500 15120 81520
rect 15380 81500 15620 81520
rect 15880 81500 16120 81520
rect 16380 81500 16620 81520
rect 16880 81500 17120 81520
rect 17380 81500 17620 81520
rect 17880 81500 18120 81520
rect 18380 81500 18620 81520
rect 18880 81500 19120 81520
rect 19380 81500 19620 81520
rect 19880 81500 20120 81520
rect 20380 81500 20620 81520
rect 20880 81500 21120 81520
rect 21380 81500 21620 81520
rect 21880 81500 22120 81520
rect 22380 81500 22620 81520
rect 22880 81500 23120 81520
rect 23380 81500 23620 81520
rect 23880 81500 24120 81520
rect 24380 81500 24620 81520
rect 24880 81500 25120 81520
rect 25380 81500 25620 81520
rect 25880 81500 26120 81520
rect 26380 81500 26620 81520
rect 26880 81500 27120 81520
rect 27380 81500 27620 81520
rect 27880 81500 28120 81520
rect 28380 81500 28620 81520
rect 28880 81500 29120 81520
rect 29380 81500 29620 81520
rect 29880 81500 30120 81520
rect 30380 81500 30620 81520
rect 30880 81500 31120 81520
rect 31380 81500 31620 81520
rect 31880 81500 32120 81520
rect 32380 81500 32620 81520
rect 32880 81500 33120 81520
rect 33380 81500 33620 81520
rect 33880 81500 34120 81520
rect 34380 81500 34620 81520
rect 34880 81500 35120 81520
rect 35380 81500 35620 81520
rect 35880 81500 36120 81520
rect 36380 81500 36620 81520
rect 36880 81500 37120 81520
rect 37380 81500 37620 81520
rect 37880 81500 38120 81520
rect 38380 81500 38620 81520
rect 38880 81500 39120 81520
rect 39380 81500 39620 81520
rect 39880 81500 40120 81520
rect 40380 81500 40620 81520
rect 40880 81500 41120 81520
rect 41380 81500 41620 81520
rect 41880 81500 42120 81520
rect 42380 81500 42620 81520
rect 42880 81500 43120 81520
rect 43380 81500 43620 81520
rect 43880 81500 44120 81520
rect 44380 81500 44620 81520
rect 44880 81500 45120 81520
rect 45380 81500 45620 81520
rect 45880 81500 46120 81520
rect 46380 81500 46620 81520
rect 46880 81500 47120 81520
rect 47380 81500 47620 81520
rect 47880 81500 48120 81520
rect 48380 81500 48620 81520
rect 48880 81500 49120 81520
rect 49380 81500 49620 81520
rect 49880 81500 50120 81520
rect 50380 81500 50620 81520
rect 50880 81500 51120 81520
rect 51380 81500 51620 81520
rect 51880 81500 52120 81520
rect 52380 81500 52620 81520
rect 52880 81500 53120 81520
rect 53380 81500 53620 81520
rect 53880 81500 54120 81520
rect 54380 81500 54620 81520
rect 54880 81500 55120 81520
rect 55380 81500 55620 81520
rect 55880 81500 56120 81520
rect 56380 81500 56620 81520
rect 56880 81500 57120 81520
rect 57380 81500 57620 81520
rect 57880 81500 58120 81520
rect 58380 81500 58620 81520
rect 58880 81500 59120 81520
rect 59380 81500 59620 81520
rect 59880 81500 60120 81520
rect 60380 81500 60620 81520
rect 60880 81500 61120 81520
rect 61380 81500 61620 81520
rect 61880 81500 62120 81520
rect 62380 81500 62620 81520
rect 62880 81500 63120 81520
rect 63380 81500 63620 81520
rect 63880 81500 64120 81520
rect 64380 81500 64620 81520
rect 64880 81500 65120 81520
rect 65380 81500 65620 81520
rect 65880 81500 66120 81520
rect 66380 81500 66620 81520
rect 66880 81500 67120 81520
rect 67380 81500 67620 81520
rect 67880 81500 68120 81520
rect 68380 81500 68620 81520
rect 68880 81500 69120 81520
rect 69380 81500 69620 81520
rect 69880 81500 70120 81520
rect 70380 81500 70620 81520
rect 70880 81500 71120 81520
rect 71380 81500 71620 81520
rect 71880 81500 72120 81520
rect 72380 81500 72620 81520
rect 72880 81500 73120 81520
rect 73380 81500 73620 81520
rect 73880 81500 74120 81520
rect 74380 81500 74620 81520
rect 74880 81500 75120 81520
rect 75380 81500 75620 81520
rect 75880 81500 76120 81520
rect 76380 81500 76620 81520
rect 76880 81500 77120 81520
rect 77380 81500 77620 81520
rect 77880 81500 78120 81520
rect 78380 81500 78620 81520
rect 78880 81500 79120 81520
rect 79380 81500 79620 81520
rect 79880 81500 80120 81520
rect 80380 81500 80620 81520
rect 80880 81500 81120 81520
rect 81380 81500 81620 81520
rect 81880 81500 82120 81520
rect 82380 81500 82620 81520
rect 82880 81500 83120 81520
rect 83380 81500 83620 81520
rect 83880 81500 84120 81520
rect 84380 81500 84620 81520
rect 84880 81500 85120 81520
rect 85380 81500 85620 81520
rect 85880 81500 86120 81520
rect 86380 81500 86620 81520
rect 86880 81500 87120 81520
rect 87380 81500 87620 81520
rect 87880 81500 88120 81520
rect 88380 81500 88620 81520
rect 88880 81500 89120 81520
rect 89380 81500 89620 81520
rect 89880 81500 90120 81520
rect 90380 81500 90620 81520
rect 90880 81500 91120 81520
rect 91380 81500 91620 81520
rect 91880 81500 92120 81520
rect 92380 81500 92620 81520
rect 92880 81500 93120 81520
rect 93380 81500 93620 81520
rect 93880 81500 94120 81520
rect 94380 81500 94620 81520
rect 94880 81500 95120 81520
rect 95380 81500 95620 81520
rect 95880 81500 96120 81520
rect 96380 81500 96620 81520
rect 96880 81500 97120 81520
rect 97380 81500 97620 81520
rect 97880 81500 98120 81520
rect 98380 81500 98620 81520
rect 98880 81500 99120 81520
rect 99380 81500 99620 81520
rect 99880 81500 100120 81520
rect 100380 81500 100500 81520
rect -83500 81490 100500 81500
rect -83500 81420 -83350 81490
rect -83150 81420 -82850 81490
rect -82650 81420 -82350 81490
rect -82150 81420 -81850 81490
rect -81650 81420 -81350 81490
rect -81150 81420 -80850 81490
rect -80650 81420 -80350 81490
rect -80150 81420 -79850 81490
rect -79650 81420 -79350 81490
rect -79150 81420 -78850 81490
rect -78650 81420 -78350 81490
rect -78150 81420 -77850 81490
rect -77650 81420 -77350 81490
rect -77150 81420 -76850 81490
rect -76650 81420 -76350 81490
rect -76150 81420 -75850 81490
rect -75650 81420 -75350 81490
rect -75150 81420 -74850 81490
rect -74650 81420 -74350 81490
rect -74150 81420 -73850 81490
rect -73650 81420 -73350 81490
rect -73150 81420 -72850 81490
rect -72650 81420 -72350 81490
rect -72150 81420 -71850 81490
rect -71650 81420 -71350 81490
rect -71150 81420 -70850 81490
rect -70650 81420 -70350 81490
rect -70150 81420 -69850 81490
rect -69650 81420 -69350 81490
rect -69150 81420 -68850 81490
rect -68650 81420 -68350 81490
rect -68150 81420 -67850 81490
rect -67650 81420 -67350 81490
rect -67150 81420 -66850 81490
rect -66650 81420 -66350 81490
rect -66150 81420 -65850 81490
rect -65650 81420 -65350 81490
rect -65150 81420 -64850 81490
rect -64650 81420 -64350 81490
rect -64150 81420 -63850 81490
rect -63650 81420 -63350 81490
rect -63150 81420 -62850 81490
rect -62650 81420 -62350 81490
rect -62150 81420 -61850 81490
rect -61650 81420 -61350 81490
rect -61150 81420 -60850 81490
rect -60650 81420 -60350 81490
rect -60150 81420 -59850 81490
rect -59650 81420 -59350 81490
rect -59150 81420 -58850 81490
rect -58650 81420 -58350 81490
rect -58150 81420 -57850 81490
rect -57650 81420 -57350 81490
rect -57150 81420 -56850 81490
rect -56650 81420 -56350 81490
rect -56150 81420 -55850 81490
rect -55650 81420 -55350 81490
rect -55150 81420 -54850 81490
rect -54650 81420 -54350 81490
rect -54150 81420 -53850 81490
rect -53650 81420 -53350 81490
rect -53150 81420 -52850 81490
rect -52650 81420 -52350 81490
rect -52150 81420 -51850 81490
rect -51650 81420 -51350 81490
rect -51150 81420 -50850 81490
rect -50650 81420 -50350 81490
rect -50150 81420 -49850 81490
rect -49650 81420 -49350 81490
rect -49150 81420 -48850 81490
rect -48650 81420 -48350 81490
rect -48150 81420 -47850 81490
rect -47650 81420 -47350 81490
rect -47150 81420 -46850 81490
rect -46650 81420 -46350 81490
rect -46150 81420 -45850 81490
rect -45650 81420 -45350 81490
rect -45150 81420 -44850 81490
rect -44650 81420 -44350 81490
rect -44150 81420 -43850 81490
rect -43650 81420 -43350 81490
rect -43150 81420 -42850 81490
rect -42650 81420 -42350 81490
rect -42150 81420 -41850 81490
rect -41650 81420 -41350 81490
rect -41150 81420 -40850 81490
rect -40650 81420 -40350 81490
rect -40150 81420 -39850 81490
rect -39650 81420 -39350 81490
rect -39150 81420 -38850 81490
rect -38650 81420 -38350 81490
rect -38150 81420 -37850 81490
rect -37650 81420 -37350 81490
rect -37150 81420 -36850 81490
rect -36650 81420 -36350 81490
rect -36150 81420 -35850 81490
rect -35650 81420 -35350 81490
rect -35150 81420 -34850 81490
rect -34650 81420 -34350 81490
rect -34150 81420 -33850 81490
rect -33650 81420 -33350 81490
rect -33150 81420 -32850 81490
rect -32650 81420 -32350 81490
rect -32150 81420 -31850 81490
rect -31650 81420 -31350 81490
rect -31150 81420 -30850 81490
rect -30650 81420 -30350 81490
rect -30150 81420 -29850 81490
rect -29650 81420 -29350 81490
rect -29150 81420 -28850 81490
rect -28650 81420 -28350 81490
rect -28150 81420 -27850 81490
rect -27650 81420 -27350 81490
rect -27150 81420 -26850 81490
rect -26650 81420 -26350 81490
rect -26150 81420 -25850 81490
rect -25650 81420 -25350 81490
rect -25150 81420 -24850 81490
rect -24650 81420 -24350 81490
rect -24150 81420 -23850 81490
rect -23650 81420 -23350 81490
rect -23150 81420 -22850 81490
rect -22650 81420 -22350 81490
rect -22150 81420 -21850 81490
rect -21650 81420 -21350 81490
rect -21150 81420 -20850 81490
rect -20650 81420 -20350 81490
rect -20150 81420 -19850 81490
rect -19650 81420 -19350 81490
rect -19150 81420 -18850 81490
rect -18650 81420 -18350 81490
rect -18150 81420 -17850 81490
rect -17650 81420 -17350 81490
rect -17150 81420 -16850 81490
rect -16650 81420 -16350 81490
rect -16150 81420 -15850 81490
rect -15650 81420 -15350 81490
rect -15150 81420 -14850 81490
rect -14650 81420 -14350 81490
rect -14150 81420 -13850 81490
rect -13650 81420 -13350 81490
rect -13150 81420 -12850 81490
rect -12650 81420 -12350 81490
rect -12150 81420 -11850 81490
rect -11650 81420 -11350 81490
rect -11150 81420 -10850 81490
rect -10650 81420 -10350 81490
rect -10150 81420 -9850 81490
rect -9650 81420 -9350 81490
rect -9150 81420 -8850 81490
rect -8650 81420 -8350 81490
rect -8150 81420 -7850 81490
rect -7650 81420 -7350 81490
rect -7150 81420 -6850 81490
rect -6650 81420 -6350 81490
rect -6150 81420 -5850 81490
rect -5650 81420 -5350 81490
rect -5150 81420 -4850 81490
rect -4650 81420 -4350 81490
rect -4150 81420 -3850 81490
rect -3650 81420 -3350 81490
rect -3150 81420 -2850 81490
rect -2650 81420 -2350 81490
rect -2150 81420 -1850 81490
rect -1650 81420 -1350 81490
rect -1150 81420 -850 81490
rect -650 81420 -350 81490
rect -150 81420 150 81490
rect 350 81420 650 81490
rect 850 81420 1150 81490
rect 1350 81420 1650 81490
rect 1850 81420 2150 81490
rect 2350 81420 2650 81490
rect 2850 81420 3150 81490
rect 3350 81420 3650 81490
rect 3850 81420 4150 81490
rect 4350 81420 4650 81490
rect 4850 81420 5150 81490
rect 5350 81420 5650 81490
rect 5850 81420 6150 81490
rect 6350 81420 6650 81490
rect 6850 81420 7150 81490
rect 7350 81420 7650 81490
rect 7850 81420 8150 81490
rect 8350 81420 8650 81490
rect 8850 81420 9150 81490
rect 9350 81420 9650 81490
rect 9850 81420 10150 81490
rect 10350 81420 10650 81490
rect 10850 81420 11150 81490
rect 11350 81420 11650 81490
rect 11850 81420 12150 81490
rect 12350 81420 12650 81490
rect 12850 81420 13150 81490
rect 13350 81420 13650 81490
rect 13850 81420 14150 81490
rect 14350 81420 14650 81490
rect 14850 81420 15150 81490
rect 15350 81420 15650 81490
rect 15850 81420 16150 81490
rect 16350 81420 16650 81490
rect 16850 81420 17150 81490
rect 17350 81420 17650 81490
rect 17850 81420 18150 81490
rect 18350 81420 18650 81490
rect 18850 81420 19150 81490
rect 19350 81420 19650 81490
rect 19850 81420 20150 81490
rect 20350 81420 20650 81490
rect 20850 81420 21150 81490
rect 21350 81420 21650 81490
rect 21850 81420 22150 81490
rect 22350 81420 22650 81490
rect 22850 81420 23150 81490
rect 23350 81420 23650 81490
rect 23850 81420 24150 81490
rect 24350 81420 24650 81490
rect 24850 81420 25150 81490
rect 25350 81420 25650 81490
rect 25850 81420 26150 81490
rect 26350 81420 26650 81490
rect 26850 81420 27150 81490
rect 27350 81420 27650 81490
rect 27850 81420 28150 81490
rect 28350 81420 28650 81490
rect 28850 81420 29150 81490
rect 29350 81420 29650 81490
rect 29850 81420 30150 81490
rect 30350 81420 30650 81490
rect 30850 81420 31150 81490
rect 31350 81420 31650 81490
rect 31850 81420 32150 81490
rect 32350 81420 32650 81490
rect 32850 81420 33150 81490
rect 33350 81420 33650 81490
rect 33850 81420 34150 81490
rect 34350 81420 34650 81490
rect 34850 81420 35150 81490
rect 35350 81420 35650 81490
rect 35850 81420 36150 81490
rect 36350 81420 36650 81490
rect 36850 81420 37150 81490
rect 37350 81420 37650 81490
rect 37850 81420 38150 81490
rect 38350 81420 38650 81490
rect 38850 81420 39150 81490
rect 39350 81420 39650 81490
rect 39850 81420 40150 81490
rect 40350 81420 40650 81490
rect 40850 81420 41150 81490
rect 41350 81420 41650 81490
rect 41850 81420 42150 81490
rect 42350 81420 42650 81490
rect 42850 81420 43150 81490
rect 43350 81420 43650 81490
rect 43850 81420 44150 81490
rect 44350 81420 44650 81490
rect 44850 81420 45150 81490
rect 45350 81420 45650 81490
rect 45850 81420 46150 81490
rect 46350 81420 46650 81490
rect 46850 81420 47150 81490
rect 47350 81420 47650 81490
rect 47850 81420 48150 81490
rect 48350 81420 48650 81490
rect 48850 81420 49150 81490
rect 49350 81420 49650 81490
rect 49850 81420 50150 81490
rect 50350 81420 50650 81490
rect 50850 81420 51150 81490
rect 51350 81420 51650 81490
rect 51850 81420 52150 81490
rect 52350 81420 52650 81490
rect 52850 81420 53150 81490
rect 53350 81420 53650 81490
rect 53850 81420 54150 81490
rect 54350 81420 54650 81490
rect 54850 81420 55150 81490
rect 55350 81420 55650 81490
rect 55850 81420 56150 81490
rect 56350 81420 56650 81490
rect 56850 81420 57150 81490
rect 57350 81420 57650 81490
rect 57850 81420 58150 81490
rect 58350 81420 58650 81490
rect 58850 81420 59150 81490
rect 59350 81420 59650 81490
rect 59850 81420 60150 81490
rect 60350 81420 60650 81490
rect 60850 81420 61150 81490
rect 61350 81420 61650 81490
rect 61850 81420 62150 81490
rect 62350 81420 62650 81490
rect 62850 81420 63150 81490
rect 63350 81420 63650 81490
rect 63850 81420 64150 81490
rect 64350 81420 64650 81490
rect 64850 81420 65150 81490
rect 65350 81420 65650 81490
rect 65850 81420 66150 81490
rect 66350 81420 66650 81490
rect 66850 81420 67150 81490
rect 67350 81420 67650 81490
rect 67850 81420 68150 81490
rect 68350 81420 68650 81490
rect 68850 81420 69150 81490
rect 69350 81420 69650 81490
rect 69850 81420 70150 81490
rect 70350 81420 70650 81490
rect 70850 81420 71150 81490
rect 71350 81420 71650 81490
rect 71850 81420 72150 81490
rect 72350 81420 72650 81490
rect 72850 81420 73150 81490
rect 73350 81420 73650 81490
rect 73850 81420 74150 81490
rect 74350 81420 74650 81490
rect 74850 81420 75150 81490
rect 75350 81420 75650 81490
rect 75850 81420 76150 81490
rect 76350 81420 76650 81490
rect 76850 81420 77150 81490
rect 77350 81420 77650 81490
rect 77850 81420 78150 81490
rect 78350 81420 78650 81490
rect 78850 81420 79150 81490
rect 79350 81420 79650 81490
rect 79850 81420 80150 81490
rect 80350 81420 80650 81490
rect 80850 81420 81150 81490
rect 81350 81420 81650 81490
rect 81850 81420 82150 81490
rect 82350 81420 82650 81490
rect 82850 81420 83150 81490
rect 83350 81420 83650 81490
rect 83850 81420 84150 81490
rect 84350 81420 84650 81490
rect 84850 81420 85150 81490
rect 85350 81420 85650 81490
rect 85850 81420 86150 81490
rect 86350 81420 86650 81490
rect 86850 81420 87150 81490
rect 87350 81420 87650 81490
rect 87850 81420 88150 81490
rect 88350 81420 88650 81490
rect 88850 81420 89150 81490
rect 89350 81420 89650 81490
rect 89850 81420 90150 81490
rect 90350 81420 90650 81490
rect 90850 81420 91150 81490
rect 91350 81420 91650 81490
rect 91850 81420 92150 81490
rect 92350 81420 92650 81490
rect 92850 81420 93150 81490
rect 93350 81420 93650 81490
rect 93850 81420 94150 81490
rect 94350 81420 94650 81490
rect 94850 81420 95150 81490
rect 95350 81420 95650 81490
rect 95850 81420 96150 81490
rect 96350 81420 96650 81490
rect 96850 81420 97150 81490
rect 97350 81420 97650 81490
rect 97850 81420 98150 81490
rect 98350 81420 98650 81490
rect 98850 81420 99150 81490
rect 99350 81420 99650 81490
rect 99850 81420 100150 81490
rect 100350 81420 100500 81490
rect -83500 81380 100500 81420
rect -83500 81310 -83350 81380
rect -83150 81310 -82850 81380
rect -82650 81310 -82350 81380
rect -82150 81310 -81850 81380
rect -81650 81310 -81350 81380
rect -81150 81310 -80850 81380
rect -80650 81310 -80350 81380
rect -80150 81310 -79850 81380
rect -79650 81310 -79350 81380
rect -79150 81310 -78850 81380
rect -78650 81310 -78350 81380
rect -78150 81310 -77850 81380
rect -77650 81310 -77350 81380
rect -77150 81310 -76850 81380
rect -76650 81310 -76350 81380
rect -76150 81310 -75850 81380
rect -75650 81310 -75350 81380
rect -75150 81310 -74850 81380
rect -74650 81310 -74350 81380
rect -74150 81310 -73850 81380
rect -73650 81310 -73350 81380
rect -73150 81310 -72850 81380
rect -72650 81310 -72350 81380
rect -72150 81310 -71850 81380
rect -71650 81310 -71350 81380
rect -71150 81310 -70850 81380
rect -70650 81310 -70350 81380
rect -70150 81310 -69850 81380
rect -69650 81310 -69350 81380
rect -69150 81310 -68850 81380
rect -68650 81310 -68350 81380
rect -68150 81310 -67850 81380
rect -67650 81310 -67350 81380
rect -67150 81310 -66850 81380
rect -66650 81310 -66350 81380
rect -66150 81310 -65850 81380
rect -65650 81310 -65350 81380
rect -65150 81310 -64850 81380
rect -64650 81310 -64350 81380
rect -64150 81310 -63850 81380
rect -63650 81310 -63350 81380
rect -63150 81310 -62850 81380
rect -62650 81310 -62350 81380
rect -62150 81310 -61850 81380
rect -61650 81310 -61350 81380
rect -61150 81310 -60850 81380
rect -60650 81310 -60350 81380
rect -60150 81310 -59850 81380
rect -59650 81310 -59350 81380
rect -59150 81310 -58850 81380
rect -58650 81310 -58350 81380
rect -58150 81310 -57850 81380
rect -57650 81310 -57350 81380
rect -57150 81310 -56850 81380
rect -56650 81310 -56350 81380
rect -56150 81310 -55850 81380
rect -55650 81310 -55350 81380
rect -55150 81310 -54850 81380
rect -54650 81310 -54350 81380
rect -54150 81310 -53850 81380
rect -53650 81310 -53350 81380
rect -53150 81310 -52850 81380
rect -52650 81310 -52350 81380
rect -52150 81310 -51850 81380
rect -51650 81310 -51350 81380
rect -51150 81310 -50850 81380
rect -50650 81310 -50350 81380
rect -50150 81310 -49850 81380
rect -49650 81310 -49350 81380
rect -49150 81310 -48850 81380
rect -48650 81310 -48350 81380
rect -48150 81310 -47850 81380
rect -47650 81310 -47350 81380
rect -47150 81310 -46850 81380
rect -46650 81310 -46350 81380
rect -46150 81310 -45850 81380
rect -45650 81310 -45350 81380
rect -45150 81310 -44850 81380
rect -44650 81310 -44350 81380
rect -44150 81310 -43850 81380
rect -43650 81310 -43350 81380
rect -43150 81310 -42850 81380
rect -42650 81310 -42350 81380
rect -42150 81310 -41850 81380
rect -41650 81310 -41350 81380
rect -41150 81310 -40850 81380
rect -40650 81310 -40350 81380
rect -40150 81310 -39850 81380
rect -39650 81310 -39350 81380
rect -39150 81310 -38850 81380
rect -38650 81310 -38350 81380
rect -38150 81310 -37850 81380
rect -37650 81310 -37350 81380
rect -37150 81310 -36850 81380
rect -36650 81310 -36350 81380
rect -36150 81310 -35850 81380
rect -35650 81310 -35350 81380
rect -35150 81310 -34850 81380
rect -34650 81310 -34350 81380
rect -34150 81310 -33850 81380
rect -33650 81310 -33350 81380
rect -33150 81310 -32850 81380
rect -32650 81310 -32350 81380
rect -32150 81310 -31850 81380
rect -31650 81310 -31350 81380
rect -31150 81310 -30850 81380
rect -30650 81310 -30350 81380
rect -30150 81310 -29850 81380
rect -29650 81310 -29350 81380
rect -29150 81310 -28850 81380
rect -28650 81310 -28350 81380
rect -28150 81310 -27850 81380
rect -27650 81310 -27350 81380
rect -27150 81310 -26850 81380
rect -26650 81310 -26350 81380
rect -26150 81310 -25850 81380
rect -25650 81310 -25350 81380
rect -25150 81310 -24850 81380
rect -24650 81310 -24350 81380
rect -24150 81310 -23850 81380
rect -23650 81310 -23350 81380
rect -23150 81310 -22850 81380
rect -22650 81310 -22350 81380
rect -22150 81310 -21850 81380
rect -21650 81310 -21350 81380
rect -21150 81310 -20850 81380
rect -20650 81310 -20350 81380
rect -20150 81310 -19850 81380
rect -19650 81310 -19350 81380
rect -19150 81310 -18850 81380
rect -18650 81310 -18350 81380
rect -18150 81310 -17850 81380
rect -17650 81310 -17350 81380
rect -17150 81310 -16850 81380
rect -16650 81310 -16350 81380
rect -16150 81310 -15850 81380
rect -15650 81310 -15350 81380
rect -15150 81310 -14850 81380
rect -14650 81310 -14350 81380
rect -14150 81310 -13850 81380
rect -13650 81310 -13350 81380
rect -13150 81310 -12850 81380
rect -12650 81310 -12350 81380
rect -12150 81310 -11850 81380
rect -11650 81310 -11350 81380
rect -11150 81310 -10850 81380
rect -10650 81310 -10350 81380
rect -10150 81310 -9850 81380
rect -9650 81310 -9350 81380
rect -9150 81310 -8850 81380
rect -8650 81310 -8350 81380
rect -8150 81310 -7850 81380
rect -7650 81310 -7350 81380
rect -7150 81310 -6850 81380
rect -6650 81310 -6350 81380
rect -6150 81310 -5850 81380
rect -5650 81310 -5350 81380
rect -5150 81310 -4850 81380
rect -4650 81310 -4350 81380
rect -4150 81310 -3850 81380
rect -3650 81310 -3350 81380
rect -3150 81310 -2850 81380
rect -2650 81310 -2350 81380
rect -2150 81310 -1850 81380
rect -1650 81310 -1350 81380
rect -1150 81310 -850 81380
rect -650 81310 -350 81380
rect -150 81310 150 81380
rect 350 81310 650 81380
rect 850 81310 1150 81380
rect 1350 81310 1650 81380
rect 1850 81310 2150 81380
rect 2350 81310 2650 81380
rect 2850 81310 3150 81380
rect 3350 81310 3650 81380
rect 3850 81310 4150 81380
rect 4350 81310 4650 81380
rect 4850 81310 5150 81380
rect 5350 81310 5650 81380
rect 5850 81310 6150 81380
rect 6350 81310 6650 81380
rect 6850 81310 7150 81380
rect 7350 81310 7650 81380
rect 7850 81310 8150 81380
rect 8350 81310 8650 81380
rect 8850 81310 9150 81380
rect 9350 81310 9650 81380
rect 9850 81310 10150 81380
rect 10350 81310 10650 81380
rect 10850 81310 11150 81380
rect 11350 81310 11650 81380
rect 11850 81310 12150 81380
rect 12350 81310 12650 81380
rect 12850 81310 13150 81380
rect 13350 81310 13650 81380
rect 13850 81310 14150 81380
rect 14350 81310 14650 81380
rect 14850 81310 15150 81380
rect 15350 81310 15650 81380
rect 15850 81310 16150 81380
rect 16350 81310 16650 81380
rect 16850 81310 17150 81380
rect 17350 81310 17650 81380
rect 17850 81310 18150 81380
rect 18350 81310 18650 81380
rect 18850 81310 19150 81380
rect 19350 81310 19650 81380
rect 19850 81310 20150 81380
rect 20350 81310 20650 81380
rect 20850 81310 21150 81380
rect 21350 81310 21650 81380
rect 21850 81310 22150 81380
rect 22350 81310 22650 81380
rect 22850 81310 23150 81380
rect 23350 81310 23650 81380
rect 23850 81310 24150 81380
rect 24350 81310 24650 81380
rect 24850 81310 25150 81380
rect 25350 81310 25650 81380
rect 25850 81310 26150 81380
rect 26350 81310 26650 81380
rect 26850 81310 27150 81380
rect 27350 81310 27650 81380
rect 27850 81310 28150 81380
rect 28350 81310 28650 81380
rect 28850 81310 29150 81380
rect 29350 81310 29650 81380
rect 29850 81310 30150 81380
rect 30350 81310 30650 81380
rect 30850 81310 31150 81380
rect 31350 81310 31650 81380
rect 31850 81310 32150 81380
rect 32350 81310 32650 81380
rect 32850 81310 33150 81380
rect 33350 81310 33650 81380
rect 33850 81310 34150 81380
rect 34350 81310 34650 81380
rect 34850 81310 35150 81380
rect 35350 81310 35650 81380
rect 35850 81310 36150 81380
rect 36350 81310 36650 81380
rect 36850 81310 37150 81380
rect 37350 81310 37650 81380
rect 37850 81310 38150 81380
rect 38350 81310 38650 81380
rect 38850 81310 39150 81380
rect 39350 81310 39650 81380
rect 39850 81310 40150 81380
rect 40350 81310 40650 81380
rect 40850 81310 41150 81380
rect 41350 81310 41650 81380
rect 41850 81310 42150 81380
rect 42350 81310 42650 81380
rect 42850 81310 43150 81380
rect 43350 81310 43650 81380
rect 43850 81310 44150 81380
rect 44350 81310 44650 81380
rect 44850 81310 45150 81380
rect 45350 81310 45650 81380
rect 45850 81310 46150 81380
rect 46350 81310 46650 81380
rect 46850 81310 47150 81380
rect 47350 81310 47650 81380
rect 47850 81310 48150 81380
rect 48350 81310 48650 81380
rect 48850 81310 49150 81380
rect 49350 81310 49650 81380
rect 49850 81310 50150 81380
rect 50350 81310 50650 81380
rect 50850 81310 51150 81380
rect 51350 81310 51650 81380
rect 51850 81310 52150 81380
rect 52350 81310 52650 81380
rect 52850 81310 53150 81380
rect 53350 81310 53650 81380
rect 53850 81310 54150 81380
rect 54350 81310 54650 81380
rect 54850 81310 55150 81380
rect 55350 81310 55650 81380
rect 55850 81310 56150 81380
rect 56350 81310 56650 81380
rect 56850 81310 57150 81380
rect 57350 81310 57650 81380
rect 57850 81310 58150 81380
rect 58350 81310 58650 81380
rect 58850 81310 59150 81380
rect 59350 81310 59650 81380
rect 59850 81310 60150 81380
rect 60350 81310 60650 81380
rect 60850 81310 61150 81380
rect 61350 81310 61650 81380
rect 61850 81310 62150 81380
rect 62350 81310 62650 81380
rect 62850 81310 63150 81380
rect 63350 81310 63650 81380
rect 63850 81310 64150 81380
rect 64350 81310 64650 81380
rect 64850 81310 65150 81380
rect 65350 81310 65650 81380
rect 65850 81310 66150 81380
rect 66350 81310 66650 81380
rect 66850 81310 67150 81380
rect 67350 81310 67650 81380
rect 67850 81310 68150 81380
rect 68350 81310 68650 81380
rect 68850 81310 69150 81380
rect 69350 81310 69650 81380
rect 69850 81310 70150 81380
rect 70350 81310 70650 81380
rect 70850 81310 71150 81380
rect 71350 81310 71650 81380
rect 71850 81310 72150 81380
rect 72350 81310 72650 81380
rect 72850 81310 73150 81380
rect 73350 81310 73650 81380
rect 73850 81310 74150 81380
rect 74350 81310 74650 81380
rect 74850 81310 75150 81380
rect 75350 81310 75650 81380
rect 75850 81310 76150 81380
rect 76350 81310 76650 81380
rect 76850 81310 77150 81380
rect 77350 81310 77650 81380
rect 77850 81310 78150 81380
rect 78350 81310 78650 81380
rect 78850 81310 79150 81380
rect 79350 81310 79650 81380
rect 79850 81310 80150 81380
rect 80350 81310 80650 81380
rect 80850 81310 81150 81380
rect 81350 81310 81650 81380
rect 81850 81310 82150 81380
rect 82350 81310 82650 81380
rect 82850 81310 83150 81380
rect 83350 81310 83650 81380
rect 83850 81310 84150 81380
rect 84350 81310 84650 81380
rect 84850 81310 85150 81380
rect 85350 81310 85650 81380
rect 85850 81310 86150 81380
rect 86350 81310 86650 81380
rect 86850 81310 87150 81380
rect 87350 81310 87650 81380
rect 87850 81310 88150 81380
rect 88350 81310 88650 81380
rect 88850 81310 89150 81380
rect 89350 81310 89650 81380
rect 89850 81310 90150 81380
rect 90350 81310 90650 81380
rect 90850 81310 91150 81380
rect 91350 81310 91650 81380
rect 91850 81310 92150 81380
rect 92350 81310 92650 81380
rect 92850 81310 93150 81380
rect 93350 81310 93650 81380
rect 93850 81310 94150 81380
rect 94350 81310 94650 81380
rect 94850 81310 95150 81380
rect 95350 81310 95650 81380
rect 95850 81310 96150 81380
rect 96350 81310 96650 81380
rect 96850 81310 97150 81380
rect 97350 81310 97650 81380
rect 97850 81310 98150 81380
rect 98350 81310 98650 81380
rect 98850 81310 99150 81380
rect 99350 81310 99650 81380
rect 99850 81310 100150 81380
rect 100350 81310 100500 81380
rect -83500 81300 100500 81310
rect -83500 81280 -83380 81300
rect -83120 81280 -82880 81300
rect -82620 81280 -82380 81300
rect -82120 81280 -81880 81300
rect -81620 81280 -81380 81300
rect -81120 81280 -80880 81300
rect -80620 81280 -80380 81300
rect -80120 81280 -79880 81300
rect -79620 81280 -79380 81300
rect -79120 81280 -78880 81300
rect -78620 81280 -78380 81300
rect -78120 81280 -77880 81300
rect -77620 81280 -77380 81300
rect -77120 81280 -76880 81300
rect -76620 81280 -76380 81300
rect -76120 81280 -75880 81300
rect -75620 81280 -75380 81300
rect -75120 81280 -74880 81300
rect -74620 81280 -74380 81300
rect -74120 81280 -73880 81300
rect -73620 81280 -73380 81300
rect -73120 81280 -72880 81300
rect -72620 81280 -72380 81300
rect -72120 81280 -71880 81300
rect -71620 81280 -71380 81300
rect -71120 81280 -70880 81300
rect -70620 81280 -70380 81300
rect -70120 81280 -69880 81300
rect -69620 81280 -69380 81300
rect -69120 81280 -68880 81300
rect -68620 81280 -68380 81300
rect -68120 81280 -67880 81300
rect -67620 81280 -67380 81300
rect -67120 81280 -66880 81300
rect -66620 81280 -66380 81300
rect -66120 81280 -65880 81300
rect -65620 81280 -65380 81300
rect -65120 81280 -64880 81300
rect -64620 81280 -64380 81300
rect -64120 81280 -63880 81300
rect -63620 81280 -63380 81300
rect -63120 81280 -62880 81300
rect -62620 81280 -62380 81300
rect -62120 81280 -61880 81300
rect -61620 81280 -61380 81300
rect -61120 81280 -60880 81300
rect -60620 81280 -60380 81300
rect -60120 81280 -59880 81300
rect -59620 81280 -59380 81300
rect -59120 81280 -58880 81300
rect -58620 81280 -58380 81300
rect -58120 81280 -57880 81300
rect -57620 81280 -57380 81300
rect -57120 81280 -56880 81300
rect -56620 81280 -56380 81300
rect -56120 81280 -55880 81300
rect -55620 81280 -55380 81300
rect -55120 81280 -54880 81300
rect -54620 81280 -54380 81300
rect -54120 81280 -53880 81300
rect -53620 81280 -53380 81300
rect -53120 81280 -52880 81300
rect -52620 81280 -52380 81300
rect -52120 81280 -51880 81300
rect -51620 81280 -51380 81300
rect -51120 81280 -50880 81300
rect -50620 81280 -50380 81300
rect -50120 81280 -49880 81300
rect -49620 81280 -49380 81300
rect -49120 81280 -48880 81300
rect -48620 81280 -48380 81300
rect -48120 81280 -47880 81300
rect -47620 81280 -47380 81300
rect -47120 81280 -46880 81300
rect -46620 81280 -46380 81300
rect -46120 81280 -45880 81300
rect -45620 81280 -45380 81300
rect -45120 81280 -44880 81300
rect -44620 81280 -44380 81300
rect -44120 81280 -43880 81300
rect -43620 81280 -43380 81300
rect -43120 81280 -42880 81300
rect -42620 81280 -42380 81300
rect -42120 81280 -41880 81300
rect -41620 81280 -41380 81300
rect -41120 81280 -40880 81300
rect -40620 81280 -40380 81300
rect -40120 81280 -39880 81300
rect -39620 81280 -39380 81300
rect -39120 81280 -38880 81300
rect -38620 81280 -38380 81300
rect -38120 81280 -37880 81300
rect -37620 81280 -37380 81300
rect -37120 81280 -36880 81300
rect -36620 81280 -36380 81300
rect -36120 81280 -35880 81300
rect -35620 81280 -35380 81300
rect -35120 81280 -34880 81300
rect -34620 81280 -34380 81300
rect -34120 81280 -33880 81300
rect -33620 81280 -33380 81300
rect -33120 81280 -32880 81300
rect -32620 81280 -32380 81300
rect -32120 81280 -31880 81300
rect -31620 81280 -31380 81300
rect -31120 81280 -30880 81300
rect -30620 81280 -30380 81300
rect -30120 81280 -29880 81300
rect -29620 81280 -29380 81300
rect -29120 81280 -28880 81300
rect -28620 81280 -28380 81300
rect -28120 81280 -27880 81300
rect -27620 81280 -27380 81300
rect -27120 81280 -26880 81300
rect -26620 81280 -26380 81300
rect -26120 81280 -25880 81300
rect -25620 81280 -25380 81300
rect -25120 81280 -24880 81300
rect -24620 81280 -24380 81300
rect -24120 81280 -23880 81300
rect -23620 81280 -23380 81300
rect -23120 81280 -22880 81300
rect -22620 81280 -22380 81300
rect -22120 81280 -21880 81300
rect -21620 81280 -21380 81300
rect -21120 81280 -20880 81300
rect -20620 81280 -20380 81300
rect -20120 81280 -19880 81300
rect -19620 81280 -19380 81300
rect -19120 81280 -18880 81300
rect -18620 81280 -18380 81300
rect -18120 81280 -17880 81300
rect -17620 81280 -17380 81300
rect -17120 81280 -16880 81300
rect -16620 81280 -16380 81300
rect -16120 81280 -15880 81300
rect -15620 81280 -15380 81300
rect -15120 81280 -14880 81300
rect -14620 81280 -14380 81300
rect -14120 81280 -13880 81300
rect -13620 81280 -13380 81300
rect -13120 81280 -12880 81300
rect -12620 81280 -12380 81300
rect -12120 81280 -11880 81300
rect -11620 81280 -11380 81300
rect -11120 81280 -10880 81300
rect -10620 81280 -10380 81300
rect -10120 81280 -9880 81300
rect -9620 81280 -9380 81300
rect -9120 81280 -8880 81300
rect -8620 81280 -8380 81300
rect -8120 81280 -7880 81300
rect -7620 81280 -7380 81300
rect -7120 81280 -6880 81300
rect -6620 81280 -6380 81300
rect -6120 81280 -5880 81300
rect -5620 81280 -5380 81300
rect -5120 81280 -4880 81300
rect -4620 81280 -4380 81300
rect -4120 81280 -3880 81300
rect -3620 81280 -3380 81300
rect -3120 81280 -2880 81300
rect -2620 81280 -2380 81300
rect -2120 81280 -1880 81300
rect -1620 81280 -1380 81300
rect -1120 81280 -880 81300
rect -620 81280 -380 81300
rect -120 81280 120 81300
rect 380 81280 620 81300
rect 880 81280 1120 81300
rect 1380 81280 1620 81300
rect 1880 81280 2120 81300
rect 2380 81280 2620 81300
rect 2880 81280 3120 81300
rect 3380 81280 3620 81300
rect 3880 81280 4120 81300
rect 4380 81280 4620 81300
rect 4880 81280 5120 81300
rect 5380 81280 5620 81300
rect 5880 81280 6120 81300
rect 6380 81280 6620 81300
rect 6880 81280 7120 81300
rect 7380 81280 7620 81300
rect 7880 81280 8120 81300
rect 8380 81280 8620 81300
rect 8880 81280 9120 81300
rect 9380 81280 9620 81300
rect 9880 81280 10120 81300
rect 10380 81280 10620 81300
rect 10880 81280 11120 81300
rect 11380 81280 11620 81300
rect 11880 81280 12120 81300
rect 12380 81280 12620 81300
rect 12880 81280 13120 81300
rect 13380 81280 13620 81300
rect 13880 81280 14120 81300
rect 14380 81280 14620 81300
rect 14880 81280 15120 81300
rect 15380 81280 15620 81300
rect 15880 81280 16120 81300
rect 16380 81280 16620 81300
rect 16880 81280 17120 81300
rect 17380 81280 17620 81300
rect 17880 81280 18120 81300
rect 18380 81280 18620 81300
rect 18880 81280 19120 81300
rect 19380 81280 19620 81300
rect 19880 81280 20120 81300
rect 20380 81280 20620 81300
rect 20880 81280 21120 81300
rect 21380 81280 21620 81300
rect 21880 81280 22120 81300
rect 22380 81280 22620 81300
rect 22880 81280 23120 81300
rect 23380 81280 23620 81300
rect 23880 81280 24120 81300
rect 24380 81280 24620 81300
rect 24880 81280 25120 81300
rect 25380 81280 25620 81300
rect 25880 81280 26120 81300
rect 26380 81280 26620 81300
rect 26880 81280 27120 81300
rect 27380 81280 27620 81300
rect 27880 81280 28120 81300
rect 28380 81280 28620 81300
rect 28880 81280 29120 81300
rect 29380 81280 29620 81300
rect 29880 81280 30120 81300
rect 30380 81280 30620 81300
rect 30880 81280 31120 81300
rect 31380 81280 31620 81300
rect 31880 81280 32120 81300
rect 32380 81280 32620 81300
rect 32880 81280 33120 81300
rect 33380 81280 33620 81300
rect 33880 81280 34120 81300
rect 34380 81280 34620 81300
rect 34880 81280 35120 81300
rect 35380 81280 35620 81300
rect 35880 81280 36120 81300
rect 36380 81280 36620 81300
rect 36880 81280 37120 81300
rect 37380 81280 37620 81300
rect 37880 81280 38120 81300
rect 38380 81280 38620 81300
rect 38880 81280 39120 81300
rect 39380 81280 39620 81300
rect 39880 81280 40120 81300
rect 40380 81280 40620 81300
rect 40880 81280 41120 81300
rect 41380 81280 41620 81300
rect 41880 81280 42120 81300
rect 42380 81280 42620 81300
rect 42880 81280 43120 81300
rect 43380 81280 43620 81300
rect 43880 81280 44120 81300
rect 44380 81280 44620 81300
rect 44880 81280 45120 81300
rect 45380 81280 45620 81300
rect 45880 81280 46120 81300
rect 46380 81280 46620 81300
rect 46880 81280 47120 81300
rect 47380 81280 47620 81300
rect 47880 81280 48120 81300
rect 48380 81280 48620 81300
rect 48880 81280 49120 81300
rect 49380 81280 49620 81300
rect 49880 81280 50120 81300
rect 50380 81280 50620 81300
rect 50880 81280 51120 81300
rect 51380 81280 51620 81300
rect 51880 81280 52120 81300
rect 52380 81280 52620 81300
rect 52880 81280 53120 81300
rect 53380 81280 53620 81300
rect 53880 81280 54120 81300
rect 54380 81280 54620 81300
rect 54880 81280 55120 81300
rect 55380 81280 55620 81300
rect 55880 81280 56120 81300
rect 56380 81280 56620 81300
rect 56880 81280 57120 81300
rect 57380 81280 57620 81300
rect 57880 81280 58120 81300
rect 58380 81280 58620 81300
rect 58880 81280 59120 81300
rect 59380 81280 59620 81300
rect 59880 81280 60120 81300
rect 60380 81280 60620 81300
rect 60880 81280 61120 81300
rect 61380 81280 61620 81300
rect 61880 81280 62120 81300
rect 62380 81280 62620 81300
rect 62880 81280 63120 81300
rect 63380 81280 63620 81300
rect 63880 81280 64120 81300
rect 64380 81280 64620 81300
rect 64880 81280 65120 81300
rect 65380 81280 65620 81300
rect 65880 81280 66120 81300
rect 66380 81280 66620 81300
rect 66880 81280 67120 81300
rect 67380 81280 67620 81300
rect 67880 81280 68120 81300
rect 68380 81280 68620 81300
rect 68880 81280 69120 81300
rect 69380 81280 69620 81300
rect 69880 81280 70120 81300
rect 70380 81280 70620 81300
rect 70880 81280 71120 81300
rect 71380 81280 71620 81300
rect 71880 81280 72120 81300
rect 72380 81280 72620 81300
rect 72880 81280 73120 81300
rect 73380 81280 73620 81300
rect 73880 81280 74120 81300
rect 74380 81280 74620 81300
rect 74880 81280 75120 81300
rect 75380 81280 75620 81300
rect 75880 81280 76120 81300
rect 76380 81280 76620 81300
rect 76880 81280 77120 81300
rect 77380 81280 77620 81300
rect 77880 81280 78120 81300
rect 78380 81280 78620 81300
rect 78880 81280 79120 81300
rect 79380 81280 79620 81300
rect 79880 81280 80120 81300
rect 80380 81280 80620 81300
rect 80880 81280 81120 81300
rect 81380 81280 81620 81300
rect 81880 81280 82120 81300
rect 82380 81280 82620 81300
rect 82880 81280 83120 81300
rect 83380 81280 83620 81300
rect 83880 81280 84120 81300
rect 84380 81280 84620 81300
rect 84880 81280 85120 81300
rect 85380 81280 85620 81300
rect 85880 81280 86120 81300
rect 86380 81280 86620 81300
rect 86880 81280 87120 81300
rect 87380 81280 87620 81300
rect 87880 81280 88120 81300
rect 88380 81280 88620 81300
rect 88880 81280 89120 81300
rect 89380 81280 89620 81300
rect 89880 81280 90120 81300
rect 90380 81280 90620 81300
rect 90880 81280 91120 81300
rect 91380 81280 91620 81300
rect 91880 81280 92120 81300
rect 92380 81280 92620 81300
rect 92880 81280 93120 81300
rect 93380 81280 93620 81300
rect 93880 81280 94120 81300
rect 94380 81280 94620 81300
rect 94880 81280 95120 81300
rect 95380 81280 95620 81300
rect 95880 81280 96120 81300
rect 96380 81280 96620 81300
rect 96880 81280 97120 81300
rect 97380 81280 97620 81300
rect 97880 81280 98120 81300
rect 98380 81280 98620 81300
rect 98880 81280 99120 81300
rect 99380 81280 99620 81300
rect 99880 81280 100120 81300
rect 100380 81280 100500 81300
rect -83500 81250 -83400 81280
rect -83500 81050 -83480 81250
rect -83410 81050 -83400 81250
rect -83500 81020 -83400 81050
rect -83100 81250 -82900 81280
rect -83100 81050 -83090 81250
rect -83020 81050 -82980 81250
rect -82910 81050 -82900 81250
rect -83100 81020 -82900 81050
rect -82600 81250 -82400 81280
rect -82600 81050 -82590 81250
rect -82520 81050 -82480 81250
rect -82410 81050 -82400 81250
rect -82600 81020 -82400 81050
rect -82100 81250 -81900 81280
rect -82100 81050 -82090 81250
rect -82020 81050 -81980 81250
rect -81910 81050 -81900 81250
rect -82100 81020 -81900 81050
rect -81600 81250 -81400 81280
rect -81600 81050 -81590 81250
rect -81520 81050 -81480 81250
rect -81410 81050 -81400 81250
rect -81600 81020 -81400 81050
rect -81100 81250 -80900 81280
rect -81100 81050 -81090 81250
rect -81020 81050 -80980 81250
rect -80910 81050 -80900 81250
rect -81100 81020 -80900 81050
rect -80600 81250 -80400 81280
rect -80600 81050 -80590 81250
rect -80520 81050 -80480 81250
rect -80410 81050 -80400 81250
rect -80600 81020 -80400 81050
rect -80100 81250 -79900 81280
rect -80100 81050 -80090 81250
rect -80020 81050 -79980 81250
rect -79910 81050 -79900 81250
rect -80100 81020 -79900 81050
rect -79600 81250 -79400 81280
rect -79600 81050 -79590 81250
rect -79520 81050 -79480 81250
rect -79410 81050 -79400 81250
rect -79600 81020 -79400 81050
rect -79100 81250 -78900 81280
rect -79100 81050 -79090 81250
rect -79020 81050 -78980 81250
rect -78910 81050 -78900 81250
rect -79100 81020 -78900 81050
rect -78600 81250 -78400 81280
rect -78600 81050 -78590 81250
rect -78520 81050 -78480 81250
rect -78410 81050 -78400 81250
rect -78600 81020 -78400 81050
rect -78100 81250 -77900 81280
rect -78100 81050 -78090 81250
rect -78020 81050 -77980 81250
rect -77910 81050 -77900 81250
rect -78100 81020 -77900 81050
rect -77600 81250 -77400 81280
rect -77600 81050 -77590 81250
rect -77520 81050 -77480 81250
rect -77410 81050 -77400 81250
rect -77600 81020 -77400 81050
rect -77100 81250 -76900 81280
rect -77100 81050 -77090 81250
rect -77020 81050 -76980 81250
rect -76910 81050 -76900 81250
rect -77100 81020 -76900 81050
rect -76600 81250 -76400 81280
rect -76600 81050 -76590 81250
rect -76520 81050 -76480 81250
rect -76410 81050 -76400 81250
rect -76600 81020 -76400 81050
rect -76100 81250 -75900 81280
rect -76100 81050 -76090 81250
rect -76020 81050 -75980 81250
rect -75910 81050 -75900 81250
rect -76100 81020 -75900 81050
rect -75600 81250 -75400 81280
rect -75600 81050 -75590 81250
rect -75520 81050 -75480 81250
rect -75410 81050 -75400 81250
rect -75600 81020 -75400 81050
rect -75100 81250 -74900 81280
rect -75100 81050 -75090 81250
rect -75020 81050 -74980 81250
rect -74910 81050 -74900 81250
rect -75100 81020 -74900 81050
rect -74600 81250 -74400 81280
rect -74600 81050 -74590 81250
rect -74520 81050 -74480 81250
rect -74410 81050 -74400 81250
rect -74600 81020 -74400 81050
rect -74100 81250 -73900 81280
rect -74100 81050 -74090 81250
rect -74020 81050 -73980 81250
rect -73910 81050 -73900 81250
rect -74100 81020 -73900 81050
rect -73600 81250 -73400 81280
rect -73600 81050 -73590 81250
rect -73520 81050 -73480 81250
rect -73410 81050 -73400 81250
rect -73600 81020 -73400 81050
rect -73100 81250 -72900 81280
rect -73100 81050 -73090 81250
rect -73020 81050 -72980 81250
rect -72910 81050 -72900 81250
rect -73100 81020 -72900 81050
rect -72600 81250 -72400 81280
rect -72600 81050 -72590 81250
rect -72520 81050 -72480 81250
rect -72410 81050 -72400 81250
rect -72600 81020 -72400 81050
rect -72100 81250 -71900 81280
rect -72100 81050 -72090 81250
rect -72020 81050 -71980 81250
rect -71910 81050 -71900 81250
rect -72100 81020 -71900 81050
rect -71600 81250 -71400 81280
rect -71600 81050 -71590 81250
rect -71520 81050 -71480 81250
rect -71410 81050 -71400 81250
rect -71600 81020 -71400 81050
rect -71100 81250 -70900 81280
rect -71100 81050 -71090 81250
rect -71020 81050 -70980 81250
rect -70910 81050 -70900 81250
rect -71100 81020 -70900 81050
rect -70600 81250 -70400 81280
rect -70600 81050 -70590 81250
rect -70520 81050 -70480 81250
rect -70410 81050 -70400 81250
rect -70600 81020 -70400 81050
rect -70100 81250 -69900 81280
rect -70100 81050 -70090 81250
rect -70020 81050 -69980 81250
rect -69910 81050 -69900 81250
rect -70100 81020 -69900 81050
rect -69600 81250 -69400 81280
rect -69600 81050 -69590 81250
rect -69520 81050 -69480 81250
rect -69410 81050 -69400 81250
rect -69600 81020 -69400 81050
rect -69100 81250 -68900 81280
rect -69100 81050 -69090 81250
rect -69020 81050 -68980 81250
rect -68910 81050 -68900 81250
rect -69100 81020 -68900 81050
rect -68600 81250 -68400 81280
rect -68600 81050 -68590 81250
rect -68520 81050 -68480 81250
rect -68410 81050 -68400 81250
rect -68600 81020 -68400 81050
rect -68100 81250 -67900 81280
rect -68100 81050 -68090 81250
rect -68020 81050 -67980 81250
rect -67910 81050 -67900 81250
rect -68100 81020 -67900 81050
rect -67600 81250 -67400 81280
rect -67600 81050 -67590 81250
rect -67520 81050 -67480 81250
rect -67410 81050 -67400 81250
rect -67600 81020 -67400 81050
rect -67100 81250 -66900 81280
rect -67100 81050 -67090 81250
rect -67020 81050 -66980 81250
rect -66910 81050 -66900 81250
rect -67100 81020 -66900 81050
rect -66600 81250 -66400 81280
rect -66600 81050 -66590 81250
rect -66520 81050 -66480 81250
rect -66410 81050 -66400 81250
rect -66600 81020 -66400 81050
rect -66100 81250 -65900 81280
rect -66100 81050 -66090 81250
rect -66020 81050 -65980 81250
rect -65910 81050 -65900 81250
rect -66100 81020 -65900 81050
rect -65600 81250 -65400 81280
rect -65600 81050 -65590 81250
rect -65520 81050 -65480 81250
rect -65410 81050 -65400 81250
rect -65600 81020 -65400 81050
rect -65100 81250 -64900 81280
rect -65100 81050 -65090 81250
rect -65020 81050 -64980 81250
rect -64910 81050 -64900 81250
rect -65100 81020 -64900 81050
rect -64600 81250 -64400 81280
rect -64600 81050 -64590 81250
rect -64520 81050 -64480 81250
rect -64410 81050 -64400 81250
rect -64600 81020 -64400 81050
rect -64100 81250 -63900 81280
rect -64100 81050 -64090 81250
rect -64020 81050 -63980 81250
rect -63910 81050 -63900 81250
rect -64100 81020 -63900 81050
rect -63600 81250 -63400 81280
rect -63600 81050 -63590 81250
rect -63520 81050 -63480 81250
rect -63410 81050 -63400 81250
rect -63600 81020 -63400 81050
rect -63100 81250 -62900 81280
rect -63100 81050 -63090 81250
rect -63020 81050 -62980 81250
rect -62910 81050 -62900 81250
rect -63100 81020 -62900 81050
rect -62600 81250 -62400 81280
rect -62600 81050 -62590 81250
rect -62520 81050 -62480 81250
rect -62410 81050 -62400 81250
rect -62600 81020 -62400 81050
rect -62100 81250 -61900 81280
rect -62100 81050 -62090 81250
rect -62020 81050 -61980 81250
rect -61910 81050 -61900 81250
rect -62100 81020 -61900 81050
rect -61600 81250 -61400 81280
rect -61600 81050 -61590 81250
rect -61520 81050 -61480 81250
rect -61410 81050 -61400 81250
rect -61600 81020 -61400 81050
rect -61100 81250 -60900 81280
rect -61100 81050 -61090 81250
rect -61020 81050 -60980 81250
rect -60910 81050 -60900 81250
rect -61100 81020 -60900 81050
rect -60600 81250 -60400 81280
rect -60600 81050 -60590 81250
rect -60520 81050 -60480 81250
rect -60410 81050 -60400 81250
rect -60600 81020 -60400 81050
rect -60100 81250 -59900 81280
rect -60100 81050 -60090 81250
rect -60020 81050 -59980 81250
rect -59910 81050 -59900 81250
rect -60100 81020 -59900 81050
rect -59600 81250 -59400 81280
rect -59600 81050 -59590 81250
rect -59520 81050 -59480 81250
rect -59410 81050 -59400 81250
rect -59600 81020 -59400 81050
rect -59100 81250 -58900 81280
rect -59100 81050 -59090 81250
rect -59020 81050 -58980 81250
rect -58910 81050 -58900 81250
rect -59100 81020 -58900 81050
rect -58600 81250 -58400 81280
rect -58600 81050 -58590 81250
rect -58520 81050 -58480 81250
rect -58410 81050 -58400 81250
rect -58600 81020 -58400 81050
rect -58100 81250 -57900 81280
rect -58100 81050 -58090 81250
rect -58020 81050 -57980 81250
rect -57910 81050 -57900 81250
rect -58100 81020 -57900 81050
rect -57600 81250 -57400 81280
rect -57600 81050 -57590 81250
rect -57520 81050 -57480 81250
rect -57410 81050 -57400 81250
rect -57600 81020 -57400 81050
rect -57100 81250 -56900 81280
rect -57100 81050 -57090 81250
rect -57020 81050 -56980 81250
rect -56910 81050 -56900 81250
rect -57100 81020 -56900 81050
rect -56600 81250 -56400 81280
rect -56600 81050 -56590 81250
rect -56520 81050 -56480 81250
rect -56410 81050 -56400 81250
rect -56600 81020 -56400 81050
rect -56100 81250 -55900 81280
rect -56100 81050 -56090 81250
rect -56020 81050 -55980 81250
rect -55910 81050 -55900 81250
rect -56100 81020 -55900 81050
rect -55600 81250 -55400 81280
rect -55600 81050 -55590 81250
rect -55520 81050 -55480 81250
rect -55410 81050 -55400 81250
rect -55600 81020 -55400 81050
rect -55100 81250 -54900 81280
rect -55100 81050 -55090 81250
rect -55020 81050 -54980 81250
rect -54910 81050 -54900 81250
rect -55100 81020 -54900 81050
rect -54600 81250 -54400 81280
rect -54600 81050 -54590 81250
rect -54520 81050 -54480 81250
rect -54410 81050 -54400 81250
rect -54600 81020 -54400 81050
rect -54100 81250 -53900 81280
rect -54100 81050 -54090 81250
rect -54020 81050 -53980 81250
rect -53910 81050 -53900 81250
rect -54100 81020 -53900 81050
rect -53600 81250 -53400 81280
rect -53600 81050 -53590 81250
rect -53520 81050 -53480 81250
rect -53410 81050 -53400 81250
rect -53600 81020 -53400 81050
rect -53100 81250 -52900 81280
rect -53100 81050 -53090 81250
rect -53020 81050 -52980 81250
rect -52910 81050 -52900 81250
rect -53100 81020 -52900 81050
rect -52600 81250 -52400 81280
rect -52600 81050 -52590 81250
rect -52520 81050 -52480 81250
rect -52410 81050 -52400 81250
rect -52600 81020 -52400 81050
rect -52100 81250 -51900 81280
rect -52100 81050 -52090 81250
rect -52020 81050 -51980 81250
rect -51910 81050 -51900 81250
rect -52100 81020 -51900 81050
rect -51600 81250 -51400 81280
rect -51600 81050 -51590 81250
rect -51520 81050 -51480 81250
rect -51410 81050 -51400 81250
rect -51600 81020 -51400 81050
rect -51100 81250 -50900 81280
rect -51100 81050 -51090 81250
rect -51020 81050 -50980 81250
rect -50910 81050 -50900 81250
rect -51100 81020 -50900 81050
rect -50600 81250 -50400 81280
rect -50600 81050 -50590 81250
rect -50520 81050 -50480 81250
rect -50410 81050 -50400 81250
rect -50600 81020 -50400 81050
rect -50100 81250 -49900 81280
rect -50100 81050 -50090 81250
rect -50020 81050 -49980 81250
rect -49910 81050 -49900 81250
rect -50100 81020 -49900 81050
rect -49600 81250 -49400 81280
rect -49600 81050 -49590 81250
rect -49520 81050 -49480 81250
rect -49410 81050 -49400 81250
rect -49600 81020 -49400 81050
rect -49100 81250 -48900 81280
rect -49100 81050 -49090 81250
rect -49020 81050 -48980 81250
rect -48910 81050 -48900 81250
rect -49100 81020 -48900 81050
rect -48600 81250 -48400 81280
rect -48600 81050 -48590 81250
rect -48520 81050 -48480 81250
rect -48410 81050 -48400 81250
rect -48600 81020 -48400 81050
rect -48100 81250 -47900 81280
rect -48100 81050 -48090 81250
rect -48020 81050 -47980 81250
rect -47910 81050 -47900 81250
rect -48100 81020 -47900 81050
rect -47600 81250 -47400 81280
rect -47600 81050 -47590 81250
rect -47520 81050 -47480 81250
rect -47410 81050 -47400 81250
rect -47600 81020 -47400 81050
rect -47100 81250 -46900 81280
rect -47100 81050 -47090 81250
rect -47020 81050 -46980 81250
rect -46910 81050 -46900 81250
rect -47100 81020 -46900 81050
rect -46600 81250 -46400 81280
rect -46600 81050 -46590 81250
rect -46520 81050 -46480 81250
rect -46410 81050 -46400 81250
rect -46600 81020 -46400 81050
rect -46100 81250 -45900 81280
rect -46100 81050 -46090 81250
rect -46020 81050 -45980 81250
rect -45910 81050 -45900 81250
rect -46100 81020 -45900 81050
rect -45600 81250 -45400 81280
rect -45600 81050 -45590 81250
rect -45520 81050 -45480 81250
rect -45410 81050 -45400 81250
rect -45600 81020 -45400 81050
rect -45100 81250 -44900 81280
rect -45100 81050 -45090 81250
rect -45020 81050 -44980 81250
rect -44910 81050 -44900 81250
rect -45100 81020 -44900 81050
rect -44600 81250 -44400 81280
rect -44600 81050 -44590 81250
rect -44520 81050 -44480 81250
rect -44410 81050 -44400 81250
rect -44600 81020 -44400 81050
rect -44100 81250 -43900 81280
rect -44100 81050 -44090 81250
rect -44020 81050 -43980 81250
rect -43910 81050 -43900 81250
rect -44100 81020 -43900 81050
rect -43600 81250 -43400 81280
rect -43600 81050 -43590 81250
rect -43520 81050 -43480 81250
rect -43410 81050 -43400 81250
rect -43600 81020 -43400 81050
rect -43100 81250 -42900 81280
rect -43100 81050 -43090 81250
rect -43020 81050 -42980 81250
rect -42910 81050 -42900 81250
rect -43100 81020 -42900 81050
rect -42600 81250 -42400 81280
rect -42600 81050 -42590 81250
rect -42520 81050 -42480 81250
rect -42410 81050 -42400 81250
rect -42600 81020 -42400 81050
rect -42100 81250 -41900 81280
rect -42100 81050 -42090 81250
rect -42020 81050 -41980 81250
rect -41910 81050 -41900 81250
rect -42100 81020 -41900 81050
rect -41600 81250 -41400 81280
rect -41600 81050 -41590 81250
rect -41520 81050 -41480 81250
rect -41410 81050 -41400 81250
rect -41600 81020 -41400 81050
rect -41100 81250 -40900 81280
rect -41100 81050 -41090 81250
rect -41020 81050 -40980 81250
rect -40910 81050 -40900 81250
rect -41100 81020 -40900 81050
rect -40600 81250 -40400 81280
rect -40600 81050 -40590 81250
rect -40520 81050 -40480 81250
rect -40410 81050 -40400 81250
rect -40600 81020 -40400 81050
rect -40100 81250 -39900 81280
rect -40100 81050 -40090 81250
rect -40020 81050 -39980 81250
rect -39910 81050 -39900 81250
rect -40100 81020 -39900 81050
rect -39600 81250 -39400 81280
rect -39600 81050 -39590 81250
rect -39520 81050 -39480 81250
rect -39410 81050 -39400 81250
rect -39600 81020 -39400 81050
rect -39100 81250 -38900 81280
rect -39100 81050 -39090 81250
rect -39020 81050 -38980 81250
rect -38910 81050 -38900 81250
rect -39100 81020 -38900 81050
rect -38600 81250 -38400 81280
rect -38600 81050 -38590 81250
rect -38520 81050 -38480 81250
rect -38410 81050 -38400 81250
rect -38600 81020 -38400 81050
rect -38100 81250 -37900 81280
rect -38100 81050 -38090 81250
rect -38020 81050 -37980 81250
rect -37910 81050 -37900 81250
rect -38100 81020 -37900 81050
rect -37600 81250 -37400 81280
rect -37600 81050 -37590 81250
rect -37520 81050 -37480 81250
rect -37410 81050 -37400 81250
rect -37600 81020 -37400 81050
rect -37100 81250 -36900 81280
rect -37100 81050 -37090 81250
rect -37020 81050 -36980 81250
rect -36910 81050 -36900 81250
rect -37100 81020 -36900 81050
rect -36600 81250 -36400 81280
rect -36600 81050 -36590 81250
rect -36520 81050 -36480 81250
rect -36410 81050 -36400 81250
rect -36600 81020 -36400 81050
rect -36100 81250 -35900 81280
rect -36100 81050 -36090 81250
rect -36020 81050 -35980 81250
rect -35910 81050 -35900 81250
rect -36100 81020 -35900 81050
rect -35600 81250 -35400 81280
rect -35600 81050 -35590 81250
rect -35520 81050 -35480 81250
rect -35410 81050 -35400 81250
rect -35600 81020 -35400 81050
rect -35100 81250 -34900 81280
rect -35100 81050 -35090 81250
rect -35020 81050 -34980 81250
rect -34910 81050 -34900 81250
rect -35100 81020 -34900 81050
rect -34600 81250 -34400 81280
rect -34600 81050 -34590 81250
rect -34520 81050 -34480 81250
rect -34410 81050 -34400 81250
rect -34600 81020 -34400 81050
rect -34100 81250 -33900 81280
rect -34100 81050 -34090 81250
rect -34020 81050 -33980 81250
rect -33910 81050 -33900 81250
rect -34100 81020 -33900 81050
rect -33600 81250 -33400 81280
rect -33600 81050 -33590 81250
rect -33520 81050 -33480 81250
rect -33410 81050 -33400 81250
rect -33600 81020 -33400 81050
rect -33100 81250 -32900 81280
rect -33100 81050 -33090 81250
rect -33020 81050 -32980 81250
rect -32910 81050 -32900 81250
rect -33100 81020 -32900 81050
rect -32600 81250 -32400 81280
rect -32600 81050 -32590 81250
rect -32520 81050 -32480 81250
rect -32410 81050 -32400 81250
rect -32600 81020 -32400 81050
rect -32100 81250 -31900 81280
rect -32100 81050 -32090 81250
rect -32020 81050 -31980 81250
rect -31910 81050 -31900 81250
rect -32100 81020 -31900 81050
rect -31600 81250 -31400 81280
rect -31600 81050 -31590 81250
rect -31520 81050 -31480 81250
rect -31410 81050 -31400 81250
rect -31600 81020 -31400 81050
rect -31100 81250 -30900 81280
rect -31100 81050 -31090 81250
rect -31020 81050 -30980 81250
rect -30910 81050 -30900 81250
rect -31100 81020 -30900 81050
rect -30600 81250 -30400 81280
rect -30600 81050 -30590 81250
rect -30520 81050 -30480 81250
rect -30410 81050 -30400 81250
rect -30600 81020 -30400 81050
rect -30100 81250 -29900 81280
rect -30100 81050 -30090 81250
rect -30020 81050 -29980 81250
rect -29910 81050 -29900 81250
rect -30100 81020 -29900 81050
rect -29600 81250 -29400 81280
rect -29600 81050 -29590 81250
rect -29520 81050 -29480 81250
rect -29410 81050 -29400 81250
rect -29600 81020 -29400 81050
rect -29100 81250 -28900 81280
rect -29100 81050 -29090 81250
rect -29020 81050 -28980 81250
rect -28910 81050 -28900 81250
rect -29100 81020 -28900 81050
rect -28600 81250 -28400 81280
rect -28600 81050 -28590 81250
rect -28520 81050 -28480 81250
rect -28410 81050 -28400 81250
rect -28600 81020 -28400 81050
rect -28100 81250 -27900 81280
rect -28100 81050 -28090 81250
rect -28020 81050 -27980 81250
rect -27910 81050 -27900 81250
rect -28100 81020 -27900 81050
rect -27600 81250 -27400 81280
rect -27600 81050 -27590 81250
rect -27520 81050 -27480 81250
rect -27410 81050 -27400 81250
rect -27600 81020 -27400 81050
rect -27100 81250 -26900 81280
rect -27100 81050 -27090 81250
rect -27020 81050 -26980 81250
rect -26910 81050 -26900 81250
rect -27100 81020 -26900 81050
rect -26600 81250 -26400 81280
rect -26600 81050 -26590 81250
rect -26520 81050 -26480 81250
rect -26410 81050 -26400 81250
rect -26600 81020 -26400 81050
rect -26100 81250 -25900 81280
rect -26100 81050 -26090 81250
rect -26020 81050 -25980 81250
rect -25910 81050 -25900 81250
rect -26100 81020 -25900 81050
rect -25600 81250 -25400 81280
rect -25600 81050 -25590 81250
rect -25520 81050 -25480 81250
rect -25410 81050 -25400 81250
rect -25600 81020 -25400 81050
rect -25100 81250 -24900 81280
rect -25100 81050 -25090 81250
rect -25020 81050 -24980 81250
rect -24910 81050 -24900 81250
rect -25100 81020 -24900 81050
rect -24600 81250 -24400 81280
rect -24600 81050 -24590 81250
rect -24520 81050 -24480 81250
rect -24410 81050 -24400 81250
rect -24600 81020 -24400 81050
rect -24100 81250 -23900 81280
rect -24100 81050 -24090 81250
rect -24020 81050 -23980 81250
rect -23910 81050 -23900 81250
rect -24100 81020 -23900 81050
rect -23600 81250 -23400 81280
rect -23600 81050 -23590 81250
rect -23520 81050 -23480 81250
rect -23410 81050 -23400 81250
rect -23600 81020 -23400 81050
rect -23100 81250 -22900 81280
rect -23100 81050 -23090 81250
rect -23020 81050 -22980 81250
rect -22910 81050 -22900 81250
rect -23100 81020 -22900 81050
rect -22600 81250 -22400 81280
rect -22600 81050 -22590 81250
rect -22520 81050 -22480 81250
rect -22410 81050 -22400 81250
rect -22600 81020 -22400 81050
rect -22100 81250 -21900 81280
rect -22100 81050 -22090 81250
rect -22020 81050 -21980 81250
rect -21910 81050 -21900 81250
rect -22100 81020 -21900 81050
rect -21600 81250 -21400 81280
rect -21600 81050 -21590 81250
rect -21520 81050 -21480 81250
rect -21410 81050 -21400 81250
rect -21600 81020 -21400 81050
rect -21100 81250 -20900 81280
rect -21100 81050 -21090 81250
rect -21020 81050 -20980 81250
rect -20910 81050 -20900 81250
rect -21100 81020 -20900 81050
rect -20600 81250 -20400 81280
rect -20600 81050 -20590 81250
rect -20520 81050 -20480 81250
rect -20410 81050 -20400 81250
rect -20600 81020 -20400 81050
rect -20100 81250 -19900 81280
rect -20100 81050 -20090 81250
rect -20020 81050 -19980 81250
rect -19910 81050 -19900 81250
rect -20100 81020 -19900 81050
rect -19600 81250 -19400 81280
rect -19600 81050 -19590 81250
rect -19520 81050 -19480 81250
rect -19410 81050 -19400 81250
rect -19600 81020 -19400 81050
rect -19100 81250 -18900 81280
rect -19100 81050 -19090 81250
rect -19020 81050 -18980 81250
rect -18910 81050 -18900 81250
rect -19100 81020 -18900 81050
rect -18600 81250 -18400 81280
rect -18600 81050 -18590 81250
rect -18520 81050 -18480 81250
rect -18410 81050 -18400 81250
rect -18600 81020 -18400 81050
rect -18100 81250 -17900 81280
rect -18100 81050 -18090 81250
rect -18020 81050 -17980 81250
rect -17910 81050 -17900 81250
rect -18100 81020 -17900 81050
rect -17600 81250 -17400 81280
rect -17600 81050 -17590 81250
rect -17520 81050 -17480 81250
rect -17410 81050 -17400 81250
rect -17600 81020 -17400 81050
rect -17100 81250 -16900 81280
rect -17100 81050 -17090 81250
rect -17020 81050 -16980 81250
rect -16910 81050 -16900 81250
rect -17100 81020 -16900 81050
rect -16600 81250 -16400 81280
rect -16600 81050 -16590 81250
rect -16520 81050 -16480 81250
rect -16410 81050 -16400 81250
rect -16600 81020 -16400 81050
rect -16100 81250 -15900 81280
rect -16100 81050 -16090 81250
rect -16020 81050 -15980 81250
rect -15910 81050 -15900 81250
rect -16100 81020 -15900 81050
rect -15600 81250 -15400 81280
rect -15600 81050 -15590 81250
rect -15520 81050 -15480 81250
rect -15410 81050 -15400 81250
rect -15600 81020 -15400 81050
rect -15100 81250 -14900 81280
rect -15100 81050 -15090 81250
rect -15020 81050 -14980 81250
rect -14910 81050 -14900 81250
rect -15100 81020 -14900 81050
rect -14600 81250 -14400 81280
rect -14600 81050 -14590 81250
rect -14520 81050 -14480 81250
rect -14410 81050 -14400 81250
rect -14600 81020 -14400 81050
rect -14100 81250 -13900 81280
rect -14100 81050 -14090 81250
rect -14020 81050 -13980 81250
rect -13910 81050 -13900 81250
rect -14100 81020 -13900 81050
rect -13600 81250 -13400 81280
rect -13600 81050 -13590 81250
rect -13520 81050 -13480 81250
rect -13410 81050 -13400 81250
rect -13600 81020 -13400 81050
rect -13100 81250 -12900 81280
rect -13100 81050 -13090 81250
rect -13020 81050 -12980 81250
rect -12910 81050 -12900 81250
rect -13100 81020 -12900 81050
rect -12600 81250 -12400 81280
rect -12600 81050 -12590 81250
rect -12520 81050 -12480 81250
rect -12410 81050 -12400 81250
rect -12600 81020 -12400 81050
rect -12100 81250 -11900 81280
rect -12100 81050 -12090 81250
rect -12020 81050 -11980 81250
rect -11910 81050 -11900 81250
rect -12100 81020 -11900 81050
rect -11600 81250 -11400 81280
rect -11600 81050 -11590 81250
rect -11520 81050 -11480 81250
rect -11410 81050 -11400 81250
rect -11600 81020 -11400 81050
rect -11100 81250 -10900 81280
rect -11100 81050 -11090 81250
rect -11020 81050 -10980 81250
rect -10910 81050 -10900 81250
rect -11100 81020 -10900 81050
rect -10600 81250 -10400 81280
rect -10600 81050 -10590 81250
rect -10520 81050 -10480 81250
rect -10410 81050 -10400 81250
rect -10600 81020 -10400 81050
rect -10100 81250 -9900 81280
rect -10100 81050 -10090 81250
rect -10020 81050 -9980 81250
rect -9910 81050 -9900 81250
rect -10100 81020 -9900 81050
rect -9600 81250 -9400 81280
rect -9600 81050 -9590 81250
rect -9520 81050 -9480 81250
rect -9410 81050 -9400 81250
rect -9600 81020 -9400 81050
rect -9100 81250 -8900 81280
rect -9100 81050 -9090 81250
rect -9020 81050 -8980 81250
rect -8910 81050 -8900 81250
rect -9100 81020 -8900 81050
rect -8600 81250 -8400 81280
rect -8600 81050 -8590 81250
rect -8520 81050 -8480 81250
rect -8410 81050 -8400 81250
rect -8600 81020 -8400 81050
rect -8100 81250 -7900 81280
rect -8100 81050 -8090 81250
rect -8020 81050 -7980 81250
rect -7910 81050 -7900 81250
rect -8100 81020 -7900 81050
rect -7600 81250 -7400 81280
rect -7600 81050 -7590 81250
rect -7520 81050 -7480 81250
rect -7410 81050 -7400 81250
rect -7600 81020 -7400 81050
rect -7100 81250 -6900 81280
rect -7100 81050 -7090 81250
rect -7020 81050 -6980 81250
rect -6910 81050 -6900 81250
rect -7100 81020 -6900 81050
rect -6600 81250 -6400 81280
rect -6600 81050 -6590 81250
rect -6520 81050 -6480 81250
rect -6410 81050 -6400 81250
rect -6600 81020 -6400 81050
rect -6100 81250 -5900 81280
rect -6100 81050 -6090 81250
rect -6020 81050 -5980 81250
rect -5910 81050 -5900 81250
rect -6100 81020 -5900 81050
rect -5600 81250 -5400 81280
rect -5600 81050 -5590 81250
rect -5520 81050 -5480 81250
rect -5410 81050 -5400 81250
rect -5600 81020 -5400 81050
rect -5100 81250 -4900 81280
rect -5100 81050 -5090 81250
rect -5020 81050 -4980 81250
rect -4910 81050 -4900 81250
rect -5100 81020 -4900 81050
rect -4600 81250 -4400 81280
rect -4600 81050 -4590 81250
rect -4520 81050 -4480 81250
rect -4410 81050 -4400 81250
rect -4600 81020 -4400 81050
rect -4100 81250 -3900 81280
rect -4100 81050 -4090 81250
rect -4020 81050 -3980 81250
rect -3910 81050 -3900 81250
rect -4100 81020 -3900 81050
rect -3600 81250 -3400 81280
rect -3600 81050 -3590 81250
rect -3520 81050 -3480 81250
rect -3410 81050 -3400 81250
rect -3600 81020 -3400 81050
rect -3100 81250 -2900 81280
rect -3100 81050 -3090 81250
rect -3020 81050 -2980 81250
rect -2910 81050 -2900 81250
rect -3100 81020 -2900 81050
rect -2600 81250 -2400 81280
rect -2600 81050 -2590 81250
rect -2520 81050 -2480 81250
rect -2410 81050 -2400 81250
rect -2600 81020 -2400 81050
rect -2100 81250 -1900 81280
rect -2100 81050 -2090 81250
rect -2020 81050 -1980 81250
rect -1910 81050 -1900 81250
rect -2100 81020 -1900 81050
rect -1600 81250 -1400 81280
rect -1600 81050 -1590 81250
rect -1520 81050 -1480 81250
rect -1410 81050 -1400 81250
rect -1600 81020 -1400 81050
rect -1100 81250 -900 81280
rect -1100 81050 -1090 81250
rect -1020 81050 -980 81250
rect -910 81050 -900 81250
rect -1100 81020 -900 81050
rect -600 81250 -400 81280
rect -600 81050 -590 81250
rect -520 81050 -480 81250
rect -410 81050 -400 81250
rect -600 81020 -400 81050
rect -100 81250 100 81280
rect -100 81050 -90 81250
rect -20 81050 20 81250
rect 90 81050 100 81250
rect -100 81020 100 81050
rect 400 81250 600 81280
rect 400 81050 410 81250
rect 480 81050 520 81250
rect 590 81050 600 81250
rect 400 81020 600 81050
rect 900 81250 1100 81280
rect 900 81050 910 81250
rect 980 81050 1020 81250
rect 1090 81050 1100 81250
rect 900 81020 1100 81050
rect 1400 81250 1600 81280
rect 1400 81050 1410 81250
rect 1480 81050 1520 81250
rect 1590 81050 1600 81250
rect 1400 81020 1600 81050
rect 1900 81250 2100 81280
rect 1900 81050 1910 81250
rect 1980 81050 2020 81250
rect 2090 81050 2100 81250
rect 1900 81020 2100 81050
rect 2400 81250 2600 81280
rect 2400 81050 2410 81250
rect 2480 81050 2520 81250
rect 2590 81050 2600 81250
rect 2400 81020 2600 81050
rect 2900 81250 3100 81280
rect 2900 81050 2910 81250
rect 2980 81050 3020 81250
rect 3090 81050 3100 81250
rect 2900 81020 3100 81050
rect 3400 81250 3600 81280
rect 3400 81050 3410 81250
rect 3480 81050 3520 81250
rect 3590 81050 3600 81250
rect 3400 81020 3600 81050
rect 3900 81250 4100 81280
rect 3900 81050 3910 81250
rect 3980 81050 4020 81250
rect 4090 81050 4100 81250
rect 3900 81020 4100 81050
rect 4400 81250 4600 81280
rect 4400 81050 4410 81250
rect 4480 81050 4520 81250
rect 4590 81050 4600 81250
rect 4400 81020 4600 81050
rect 4900 81250 5100 81280
rect 4900 81050 4910 81250
rect 4980 81050 5020 81250
rect 5090 81050 5100 81250
rect 4900 81020 5100 81050
rect 5400 81250 5600 81280
rect 5400 81050 5410 81250
rect 5480 81050 5520 81250
rect 5590 81050 5600 81250
rect 5400 81020 5600 81050
rect 5900 81250 6100 81280
rect 5900 81050 5910 81250
rect 5980 81050 6020 81250
rect 6090 81050 6100 81250
rect 5900 81020 6100 81050
rect 6400 81250 6600 81280
rect 6400 81050 6410 81250
rect 6480 81050 6520 81250
rect 6590 81050 6600 81250
rect 6400 81020 6600 81050
rect 6900 81250 7100 81280
rect 6900 81050 6910 81250
rect 6980 81050 7020 81250
rect 7090 81050 7100 81250
rect 6900 81020 7100 81050
rect 7400 81250 7600 81280
rect 7400 81050 7410 81250
rect 7480 81050 7520 81250
rect 7590 81050 7600 81250
rect 7400 81020 7600 81050
rect 7900 81250 8100 81280
rect 7900 81050 7910 81250
rect 7980 81050 8020 81250
rect 8090 81050 8100 81250
rect 7900 81020 8100 81050
rect 8400 81250 8600 81280
rect 8400 81050 8410 81250
rect 8480 81050 8520 81250
rect 8590 81050 8600 81250
rect 8400 81020 8600 81050
rect 8900 81250 9100 81280
rect 8900 81050 8910 81250
rect 8980 81050 9020 81250
rect 9090 81050 9100 81250
rect 8900 81020 9100 81050
rect 9400 81250 9600 81280
rect 9400 81050 9410 81250
rect 9480 81050 9520 81250
rect 9590 81050 9600 81250
rect 9400 81020 9600 81050
rect 9900 81250 10100 81280
rect 9900 81050 9910 81250
rect 9980 81050 10020 81250
rect 10090 81050 10100 81250
rect 9900 81020 10100 81050
rect 10400 81250 10600 81280
rect 10400 81050 10410 81250
rect 10480 81050 10520 81250
rect 10590 81050 10600 81250
rect 10400 81020 10600 81050
rect 10900 81250 11100 81280
rect 10900 81050 10910 81250
rect 10980 81050 11020 81250
rect 11090 81050 11100 81250
rect 10900 81020 11100 81050
rect 11400 81250 11600 81280
rect 11400 81050 11410 81250
rect 11480 81050 11520 81250
rect 11590 81050 11600 81250
rect 11400 81020 11600 81050
rect 11900 81250 12100 81280
rect 11900 81050 11910 81250
rect 11980 81050 12020 81250
rect 12090 81050 12100 81250
rect 11900 81020 12100 81050
rect 12400 81250 12600 81280
rect 12400 81050 12410 81250
rect 12480 81050 12520 81250
rect 12590 81050 12600 81250
rect 12400 81020 12600 81050
rect 12900 81250 13100 81280
rect 12900 81050 12910 81250
rect 12980 81050 13020 81250
rect 13090 81050 13100 81250
rect 12900 81020 13100 81050
rect 13400 81250 13600 81280
rect 13400 81050 13410 81250
rect 13480 81050 13520 81250
rect 13590 81050 13600 81250
rect 13400 81020 13600 81050
rect 13900 81250 14100 81280
rect 13900 81050 13910 81250
rect 13980 81050 14020 81250
rect 14090 81050 14100 81250
rect 13900 81020 14100 81050
rect 14400 81250 14600 81280
rect 14400 81050 14410 81250
rect 14480 81050 14520 81250
rect 14590 81050 14600 81250
rect 14400 81020 14600 81050
rect 14900 81250 15100 81280
rect 14900 81050 14910 81250
rect 14980 81050 15020 81250
rect 15090 81050 15100 81250
rect 14900 81020 15100 81050
rect 15400 81250 15600 81280
rect 15400 81050 15410 81250
rect 15480 81050 15520 81250
rect 15590 81050 15600 81250
rect 15400 81020 15600 81050
rect 15900 81250 16100 81280
rect 15900 81050 15910 81250
rect 15980 81050 16020 81250
rect 16090 81050 16100 81250
rect 15900 81020 16100 81050
rect 16400 81250 16600 81280
rect 16400 81050 16410 81250
rect 16480 81050 16520 81250
rect 16590 81050 16600 81250
rect 16400 81020 16600 81050
rect 16900 81250 17100 81280
rect 16900 81050 16910 81250
rect 16980 81050 17020 81250
rect 17090 81050 17100 81250
rect 16900 81020 17100 81050
rect 17400 81250 17600 81280
rect 17400 81050 17410 81250
rect 17480 81050 17520 81250
rect 17590 81050 17600 81250
rect 17400 81020 17600 81050
rect 17900 81250 18100 81280
rect 17900 81050 17910 81250
rect 17980 81050 18020 81250
rect 18090 81050 18100 81250
rect 17900 81020 18100 81050
rect 18400 81250 18600 81280
rect 18400 81050 18410 81250
rect 18480 81050 18520 81250
rect 18590 81050 18600 81250
rect 18400 81020 18600 81050
rect 18900 81250 19100 81280
rect 18900 81050 18910 81250
rect 18980 81050 19020 81250
rect 19090 81050 19100 81250
rect 18900 81020 19100 81050
rect 19400 81250 19600 81280
rect 19400 81050 19410 81250
rect 19480 81050 19520 81250
rect 19590 81050 19600 81250
rect 19400 81020 19600 81050
rect 19900 81250 20100 81280
rect 19900 81050 19910 81250
rect 19980 81050 20020 81250
rect 20090 81050 20100 81250
rect 19900 81020 20100 81050
rect 20400 81250 20600 81280
rect 20400 81050 20410 81250
rect 20480 81050 20520 81250
rect 20590 81050 20600 81250
rect 20400 81020 20600 81050
rect 20900 81250 21100 81280
rect 20900 81050 20910 81250
rect 20980 81050 21020 81250
rect 21090 81050 21100 81250
rect 20900 81020 21100 81050
rect 21400 81250 21600 81280
rect 21400 81050 21410 81250
rect 21480 81050 21520 81250
rect 21590 81050 21600 81250
rect 21400 81020 21600 81050
rect 21900 81250 22100 81280
rect 21900 81050 21910 81250
rect 21980 81050 22020 81250
rect 22090 81050 22100 81250
rect 21900 81020 22100 81050
rect 22400 81250 22600 81280
rect 22400 81050 22410 81250
rect 22480 81050 22520 81250
rect 22590 81050 22600 81250
rect 22400 81020 22600 81050
rect 22900 81250 23100 81280
rect 22900 81050 22910 81250
rect 22980 81050 23020 81250
rect 23090 81050 23100 81250
rect 22900 81020 23100 81050
rect 23400 81250 23600 81280
rect 23400 81050 23410 81250
rect 23480 81050 23520 81250
rect 23590 81050 23600 81250
rect 23400 81020 23600 81050
rect 23900 81250 24100 81280
rect 23900 81050 23910 81250
rect 23980 81050 24020 81250
rect 24090 81050 24100 81250
rect 23900 81020 24100 81050
rect 24400 81250 24600 81280
rect 24400 81050 24410 81250
rect 24480 81050 24520 81250
rect 24590 81050 24600 81250
rect 24400 81020 24600 81050
rect 24900 81250 25100 81280
rect 24900 81050 24910 81250
rect 24980 81050 25020 81250
rect 25090 81050 25100 81250
rect 24900 81020 25100 81050
rect 25400 81250 25600 81280
rect 25400 81050 25410 81250
rect 25480 81050 25520 81250
rect 25590 81050 25600 81250
rect 25400 81020 25600 81050
rect 25900 81250 26100 81280
rect 25900 81050 25910 81250
rect 25980 81050 26020 81250
rect 26090 81050 26100 81250
rect 25900 81020 26100 81050
rect 26400 81250 26600 81280
rect 26400 81050 26410 81250
rect 26480 81050 26520 81250
rect 26590 81050 26600 81250
rect 26400 81020 26600 81050
rect 26900 81250 27100 81280
rect 26900 81050 26910 81250
rect 26980 81050 27020 81250
rect 27090 81050 27100 81250
rect 26900 81020 27100 81050
rect 27400 81250 27600 81280
rect 27400 81050 27410 81250
rect 27480 81050 27520 81250
rect 27590 81050 27600 81250
rect 27400 81020 27600 81050
rect 27900 81250 28100 81280
rect 27900 81050 27910 81250
rect 27980 81050 28020 81250
rect 28090 81050 28100 81250
rect 27900 81020 28100 81050
rect 28400 81250 28600 81280
rect 28400 81050 28410 81250
rect 28480 81050 28520 81250
rect 28590 81050 28600 81250
rect 28400 81020 28600 81050
rect 28900 81250 29100 81280
rect 28900 81050 28910 81250
rect 28980 81050 29020 81250
rect 29090 81050 29100 81250
rect 28900 81020 29100 81050
rect 29400 81250 29600 81280
rect 29400 81050 29410 81250
rect 29480 81050 29520 81250
rect 29590 81050 29600 81250
rect 29400 81020 29600 81050
rect 29900 81250 30100 81280
rect 29900 81050 29910 81250
rect 29980 81050 30020 81250
rect 30090 81050 30100 81250
rect 29900 81020 30100 81050
rect 30400 81250 30600 81280
rect 30400 81050 30410 81250
rect 30480 81050 30520 81250
rect 30590 81050 30600 81250
rect 30400 81020 30600 81050
rect 30900 81250 31100 81280
rect 30900 81050 30910 81250
rect 30980 81050 31020 81250
rect 31090 81050 31100 81250
rect 30900 81020 31100 81050
rect 31400 81250 31600 81280
rect 31400 81050 31410 81250
rect 31480 81050 31520 81250
rect 31590 81050 31600 81250
rect 31400 81020 31600 81050
rect 31900 81250 32100 81280
rect 31900 81050 31910 81250
rect 31980 81050 32020 81250
rect 32090 81050 32100 81250
rect 31900 81020 32100 81050
rect 32400 81250 32600 81280
rect 32400 81050 32410 81250
rect 32480 81050 32520 81250
rect 32590 81050 32600 81250
rect 32400 81020 32600 81050
rect 32900 81250 33100 81280
rect 32900 81050 32910 81250
rect 32980 81050 33020 81250
rect 33090 81050 33100 81250
rect 32900 81020 33100 81050
rect 33400 81250 33600 81280
rect 33400 81050 33410 81250
rect 33480 81050 33520 81250
rect 33590 81050 33600 81250
rect 33400 81020 33600 81050
rect 33900 81250 34100 81280
rect 33900 81050 33910 81250
rect 33980 81050 34020 81250
rect 34090 81050 34100 81250
rect 33900 81020 34100 81050
rect 34400 81250 34600 81280
rect 34400 81050 34410 81250
rect 34480 81050 34520 81250
rect 34590 81050 34600 81250
rect 34400 81020 34600 81050
rect 34900 81250 35100 81280
rect 34900 81050 34910 81250
rect 34980 81050 35020 81250
rect 35090 81050 35100 81250
rect 34900 81020 35100 81050
rect 35400 81250 35600 81280
rect 35400 81050 35410 81250
rect 35480 81050 35520 81250
rect 35590 81050 35600 81250
rect 35400 81020 35600 81050
rect 35900 81250 36100 81280
rect 35900 81050 35910 81250
rect 35980 81050 36020 81250
rect 36090 81050 36100 81250
rect 35900 81020 36100 81050
rect 36400 81250 36600 81280
rect 36400 81050 36410 81250
rect 36480 81050 36520 81250
rect 36590 81050 36600 81250
rect 36400 81020 36600 81050
rect 36900 81250 37100 81280
rect 36900 81050 36910 81250
rect 36980 81050 37020 81250
rect 37090 81050 37100 81250
rect 36900 81020 37100 81050
rect 37400 81250 37600 81280
rect 37400 81050 37410 81250
rect 37480 81050 37520 81250
rect 37590 81050 37600 81250
rect 37400 81020 37600 81050
rect 37900 81250 38100 81280
rect 37900 81050 37910 81250
rect 37980 81050 38020 81250
rect 38090 81050 38100 81250
rect 37900 81020 38100 81050
rect 38400 81250 38600 81280
rect 38400 81050 38410 81250
rect 38480 81050 38520 81250
rect 38590 81050 38600 81250
rect 38400 81020 38600 81050
rect 38900 81250 39100 81280
rect 38900 81050 38910 81250
rect 38980 81050 39020 81250
rect 39090 81050 39100 81250
rect 38900 81020 39100 81050
rect 39400 81250 39600 81280
rect 39400 81050 39410 81250
rect 39480 81050 39520 81250
rect 39590 81050 39600 81250
rect 39400 81020 39600 81050
rect 39900 81250 40100 81280
rect 39900 81050 39910 81250
rect 39980 81050 40020 81250
rect 40090 81050 40100 81250
rect 39900 81020 40100 81050
rect 40400 81250 40600 81280
rect 40400 81050 40410 81250
rect 40480 81050 40520 81250
rect 40590 81050 40600 81250
rect 40400 81020 40600 81050
rect 40900 81250 41100 81280
rect 40900 81050 40910 81250
rect 40980 81050 41020 81250
rect 41090 81050 41100 81250
rect 40900 81020 41100 81050
rect 41400 81250 41600 81280
rect 41400 81050 41410 81250
rect 41480 81050 41520 81250
rect 41590 81050 41600 81250
rect 41400 81020 41600 81050
rect 41900 81250 42100 81280
rect 41900 81050 41910 81250
rect 41980 81050 42020 81250
rect 42090 81050 42100 81250
rect 41900 81020 42100 81050
rect 42400 81250 42600 81280
rect 42400 81050 42410 81250
rect 42480 81050 42520 81250
rect 42590 81050 42600 81250
rect 42400 81020 42600 81050
rect 42900 81250 43100 81280
rect 42900 81050 42910 81250
rect 42980 81050 43020 81250
rect 43090 81050 43100 81250
rect 42900 81020 43100 81050
rect 43400 81250 43600 81280
rect 43400 81050 43410 81250
rect 43480 81050 43520 81250
rect 43590 81050 43600 81250
rect 43400 81020 43600 81050
rect 43900 81250 44100 81280
rect 43900 81050 43910 81250
rect 43980 81050 44020 81250
rect 44090 81050 44100 81250
rect 43900 81020 44100 81050
rect 44400 81250 44600 81280
rect 44400 81050 44410 81250
rect 44480 81050 44520 81250
rect 44590 81050 44600 81250
rect 44400 81020 44600 81050
rect 44900 81250 45100 81280
rect 44900 81050 44910 81250
rect 44980 81050 45020 81250
rect 45090 81050 45100 81250
rect 44900 81020 45100 81050
rect 45400 81250 45600 81280
rect 45400 81050 45410 81250
rect 45480 81050 45520 81250
rect 45590 81050 45600 81250
rect 45400 81020 45600 81050
rect 45900 81250 46100 81280
rect 45900 81050 45910 81250
rect 45980 81050 46020 81250
rect 46090 81050 46100 81250
rect 45900 81020 46100 81050
rect 46400 81250 46600 81280
rect 46400 81050 46410 81250
rect 46480 81050 46520 81250
rect 46590 81050 46600 81250
rect 46400 81020 46600 81050
rect 46900 81250 47100 81280
rect 46900 81050 46910 81250
rect 46980 81050 47020 81250
rect 47090 81050 47100 81250
rect 46900 81020 47100 81050
rect 47400 81250 47600 81280
rect 47400 81050 47410 81250
rect 47480 81050 47520 81250
rect 47590 81050 47600 81250
rect 47400 81020 47600 81050
rect 47900 81250 48100 81280
rect 47900 81050 47910 81250
rect 47980 81050 48020 81250
rect 48090 81050 48100 81250
rect 47900 81020 48100 81050
rect 48400 81250 48600 81280
rect 48400 81050 48410 81250
rect 48480 81050 48520 81250
rect 48590 81050 48600 81250
rect 48400 81020 48600 81050
rect 48900 81250 49100 81280
rect 48900 81050 48910 81250
rect 48980 81050 49020 81250
rect 49090 81050 49100 81250
rect 48900 81020 49100 81050
rect 49400 81250 49600 81280
rect 49400 81050 49410 81250
rect 49480 81050 49520 81250
rect 49590 81050 49600 81250
rect 49400 81020 49600 81050
rect 49900 81250 50100 81280
rect 49900 81050 49910 81250
rect 49980 81050 50020 81250
rect 50090 81050 50100 81250
rect 49900 81020 50100 81050
rect 50400 81250 50600 81280
rect 50400 81050 50410 81250
rect 50480 81050 50520 81250
rect 50590 81050 50600 81250
rect 50400 81020 50600 81050
rect 50900 81250 51100 81280
rect 50900 81050 50910 81250
rect 50980 81050 51020 81250
rect 51090 81050 51100 81250
rect 50900 81020 51100 81050
rect 51400 81250 51600 81280
rect 51400 81050 51410 81250
rect 51480 81050 51520 81250
rect 51590 81050 51600 81250
rect 51400 81020 51600 81050
rect 51900 81250 52100 81280
rect 51900 81050 51910 81250
rect 51980 81050 52020 81250
rect 52090 81050 52100 81250
rect 51900 81020 52100 81050
rect 52400 81250 52600 81280
rect 52400 81050 52410 81250
rect 52480 81050 52520 81250
rect 52590 81050 52600 81250
rect 52400 81020 52600 81050
rect 52900 81250 53100 81280
rect 52900 81050 52910 81250
rect 52980 81050 53020 81250
rect 53090 81050 53100 81250
rect 52900 81020 53100 81050
rect 53400 81250 53600 81280
rect 53400 81050 53410 81250
rect 53480 81050 53520 81250
rect 53590 81050 53600 81250
rect 53400 81020 53600 81050
rect 53900 81250 54100 81280
rect 53900 81050 53910 81250
rect 53980 81050 54020 81250
rect 54090 81050 54100 81250
rect 53900 81020 54100 81050
rect 54400 81250 54600 81280
rect 54400 81050 54410 81250
rect 54480 81050 54520 81250
rect 54590 81050 54600 81250
rect 54400 81020 54600 81050
rect 54900 81250 55100 81280
rect 54900 81050 54910 81250
rect 54980 81050 55020 81250
rect 55090 81050 55100 81250
rect 54900 81020 55100 81050
rect 55400 81250 55600 81280
rect 55400 81050 55410 81250
rect 55480 81050 55520 81250
rect 55590 81050 55600 81250
rect 55400 81020 55600 81050
rect 55900 81250 56100 81280
rect 55900 81050 55910 81250
rect 55980 81050 56020 81250
rect 56090 81050 56100 81250
rect 55900 81020 56100 81050
rect 56400 81250 56600 81280
rect 56400 81050 56410 81250
rect 56480 81050 56520 81250
rect 56590 81050 56600 81250
rect 56400 81020 56600 81050
rect 56900 81250 57100 81280
rect 56900 81050 56910 81250
rect 56980 81050 57020 81250
rect 57090 81050 57100 81250
rect 56900 81020 57100 81050
rect 57400 81250 57600 81280
rect 57400 81050 57410 81250
rect 57480 81050 57520 81250
rect 57590 81050 57600 81250
rect 57400 81020 57600 81050
rect 57900 81250 58100 81280
rect 57900 81050 57910 81250
rect 57980 81050 58020 81250
rect 58090 81050 58100 81250
rect 57900 81020 58100 81050
rect 58400 81250 58600 81280
rect 58400 81050 58410 81250
rect 58480 81050 58520 81250
rect 58590 81050 58600 81250
rect 58400 81020 58600 81050
rect 58900 81250 59100 81280
rect 58900 81050 58910 81250
rect 58980 81050 59020 81250
rect 59090 81050 59100 81250
rect 58900 81020 59100 81050
rect 59400 81250 59600 81280
rect 59400 81050 59410 81250
rect 59480 81050 59520 81250
rect 59590 81050 59600 81250
rect 59400 81020 59600 81050
rect 59900 81250 60100 81280
rect 59900 81050 59910 81250
rect 59980 81050 60020 81250
rect 60090 81050 60100 81250
rect 59900 81020 60100 81050
rect 60400 81250 60600 81280
rect 60400 81050 60410 81250
rect 60480 81050 60520 81250
rect 60590 81050 60600 81250
rect 60400 81020 60600 81050
rect 60900 81250 61100 81280
rect 60900 81050 60910 81250
rect 60980 81050 61020 81250
rect 61090 81050 61100 81250
rect 60900 81020 61100 81050
rect 61400 81250 61600 81280
rect 61400 81050 61410 81250
rect 61480 81050 61520 81250
rect 61590 81050 61600 81250
rect 61400 81020 61600 81050
rect 61900 81250 62100 81280
rect 61900 81050 61910 81250
rect 61980 81050 62020 81250
rect 62090 81050 62100 81250
rect 61900 81020 62100 81050
rect 62400 81250 62600 81280
rect 62400 81050 62410 81250
rect 62480 81050 62520 81250
rect 62590 81050 62600 81250
rect 62400 81020 62600 81050
rect 62900 81250 63100 81280
rect 62900 81050 62910 81250
rect 62980 81050 63020 81250
rect 63090 81050 63100 81250
rect 62900 81020 63100 81050
rect 63400 81250 63600 81280
rect 63400 81050 63410 81250
rect 63480 81050 63520 81250
rect 63590 81050 63600 81250
rect 63400 81020 63600 81050
rect 63900 81250 64100 81280
rect 63900 81050 63910 81250
rect 63980 81050 64020 81250
rect 64090 81050 64100 81250
rect 63900 81020 64100 81050
rect 64400 81250 64600 81280
rect 64400 81050 64410 81250
rect 64480 81050 64520 81250
rect 64590 81050 64600 81250
rect 64400 81020 64600 81050
rect 64900 81250 65100 81280
rect 64900 81050 64910 81250
rect 64980 81050 65020 81250
rect 65090 81050 65100 81250
rect 64900 81020 65100 81050
rect 65400 81250 65600 81280
rect 65400 81050 65410 81250
rect 65480 81050 65520 81250
rect 65590 81050 65600 81250
rect 65400 81020 65600 81050
rect 65900 81250 66100 81280
rect 65900 81050 65910 81250
rect 65980 81050 66020 81250
rect 66090 81050 66100 81250
rect 65900 81020 66100 81050
rect 66400 81250 66600 81280
rect 66400 81050 66410 81250
rect 66480 81050 66520 81250
rect 66590 81050 66600 81250
rect 66400 81020 66600 81050
rect 66900 81250 67100 81280
rect 66900 81050 66910 81250
rect 66980 81050 67020 81250
rect 67090 81050 67100 81250
rect 66900 81020 67100 81050
rect 67400 81250 67600 81280
rect 67400 81050 67410 81250
rect 67480 81050 67520 81250
rect 67590 81050 67600 81250
rect 67400 81020 67600 81050
rect 67900 81250 68100 81280
rect 67900 81050 67910 81250
rect 67980 81050 68020 81250
rect 68090 81050 68100 81250
rect 67900 81020 68100 81050
rect 68400 81250 68600 81280
rect 68400 81050 68410 81250
rect 68480 81050 68520 81250
rect 68590 81050 68600 81250
rect 68400 81020 68600 81050
rect 68900 81250 69100 81280
rect 68900 81050 68910 81250
rect 68980 81050 69020 81250
rect 69090 81050 69100 81250
rect 68900 81020 69100 81050
rect 69400 81250 69600 81280
rect 69400 81050 69410 81250
rect 69480 81050 69520 81250
rect 69590 81050 69600 81250
rect 69400 81020 69600 81050
rect 69900 81250 70100 81280
rect 69900 81050 69910 81250
rect 69980 81050 70020 81250
rect 70090 81050 70100 81250
rect 69900 81020 70100 81050
rect 70400 81250 70600 81280
rect 70400 81050 70410 81250
rect 70480 81050 70520 81250
rect 70590 81050 70600 81250
rect 70400 81020 70600 81050
rect 70900 81250 71100 81280
rect 70900 81050 70910 81250
rect 70980 81050 71020 81250
rect 71090 81050 71100 81250
rect 70900 81020 71100 81050
rect 71400 81250 71600 81280
rect 71400 81050 71410 81250
rect 71480 81050 71520 81250
rect 71590 81050 71600 81250
rect 71400 81020 71600 81050
rect 71900 81250 72100 81280
rect 71900 81050 71910 81250
rect 71980 81050 72020 81250
rect 72090 81050 72100 81250
rect 71900 81020 72100 81050
rect 72400 81250 72600 81280
rect 72400 81050 72410 81250
rect 72480 81050 72520 81250
rect 72590 81050 72600 81250
rect 72400 81020 72600 81050
rect 72900 81250 73100 81280
rect 72900 81050 72910 81250
rect 72980 81050 73020 81250
rect 73090 81050 73100 81250
rect 72900 81020 73100 81050
rect 73400 81250 73600 81280
rect 73400 81050 73410 81250
rect 73480 81050 73520 81250
rect 73590 81050 73600 81250
rect 73400 81020 73600 81050
rect 73900 81250 74100 81280
rect 73900 81050 73910 81250
rect 73980 81050 74020 81250
rect 74090 81050 74100 81250
rect 73900 81020 74100 81050
rect 74400 81250 74600 81280
rect 74400 81050 74410 81250
rect 74480 81050 74520 81250
rect 74590 81050 74600 81250
rect 74400 81020 74600 81050
rect 74900 81250 75100 81280
rect 74900 81050 74910 81250
rect 74980 81050 75020 81250
rect 75090 81050 75100 81250
rect 74900 81020 75100 81050
rect 75400 81250 75600 81280
rect 75400 81050 75410 81250
rect 75480 81050 75520 81250
rect 75590 81050 75600 81250
rect 75400 81020 75600 81050
rect 75900 81250 76100 81280
rect 75900 81050 75910 81250
rect 75980 81050 76020 81250
rect 76090 81050 76100 81250
rect 75900 81020 76100 81050
rect 76400 81250 76600 81280
rect 76400 81050 76410 81250
rect 76480 81050 76520 81250
rect 76590 81050 76600 81250
rect 76400 81020 76600 81050
rect 76900 81250 77100 81280
rect 76900 81050 76910 81250
rect 76980 81050 77020 81250
rect 77090 81050 77100 81250
rect 76900 81020 77100 81050
rect 77400 81250 77600 81280
rect 77400 81050 77410 81250
rect 77480 81050 77520 81250
rect 77590 81050 77600 81250
rect 77400 81020 77600 81050
rect 77900 81250 78100 81280
rect 77900 81050 77910 81250
rect 77980 81050 78020 81250
rect 78090 81050 78100 81250
rect 77900 81020 78100 81050
rect 78400 81250 78600 81280
rect 78400 81050 78410 81250
rect 78480 81050 78520 81250
rect 78590 81050 78600 81250
rect 78400 81020 78600 81050
rect 78900 81250 79100 81280
rect 78900 81050 78910 81250
rect 78980 81050 79020 81250
rect 79090 81050 79100 81250
rect 78900 81020 79100 81050
rect 79400 81250 79600 81280
rect 79400 81050 79410 81250
rect 79480 81050 79520 81250
rect 79590 81050 79600 81250
rect 79400 81020 79600 81050
rect 79900 81250 80100 81280
rect 79900 81050 79910 81250
rect 79980 81050 80020 81250
rect 80090 81050 80100 81250
rect 79900 81020 80100 81050
rect 80400 81250 80600 81280
rect 80400 81050 80410 81250
rect 80480 81050 80520 81250
rect 80590 81050 80600 81250
rect 80400 81020 80600 81050
rect 80900 81250 81100 81280
rect 80900 81050 80910 81250
rect 80980 81050 81020 81250
rect 81090 81050 81100 81250
rect 80900 81020 81100 81050
rect 81400 81250 81600 81280
rect 81400 81050 81410 81250
rect 81480 81050 81520 81250
rect 81590 81050 81600 81250
rect 81400 81020 81600 81050
rect 81900 81250 82100 81280
rect 81900 81050 81910 81250
rect 81980 81050 82020 81250
rect 82090 81050 82100 81250
rect 81900 81020 82100 81050
rect 82400 81250 82600 81280
rect 82400 81050 82410 81250
rect 82480 81050 82520 81250
rect 82590 81050 82600 81250
rect 82400 81020 82600 81050
rect 82900 81250 83100 81280
rect 82900 81050 82910 81250
rect 82980 81050 83020 81250
rect 83090 81050 83100 81250
rect 82900 81020 83100 81050
rect 83400 81250 83600 81280
rect 83400 81050 83410 81250
rect 83480 81050 83520 81250
rect 83590 81050 83600 81250
rect 83400 81020 83600 81050
rect 83900 81250 84100 81280
rect 83900 81050 83910 81250
rect 83980 81050 84020 81250
rect 84090 81050 84100 81250
rect 83900 81020 84100 81050
rect 84400 81250 84600 81280
rect 84400 81050 84410 81250
rect 84480 81050 84520 81250
rect 84590 81050 84600 81250
rect 84400 81020 84600 81050
rect 84900 81250 85100 81280
rect 84900 81050 84910 81250
rect 84980 81050 85020 81250
rect 85090 81050 85100 81250
rect 84900 81020 85100 81050
rect 85400 81250 85600 81280
rect 85400 81050 85410 81250
rect 85480 81050 85520 81250
rect 85590 81050 85600 81250
rect 85400 81020 85600 81050
rect 85900 81250 86100 81280
rect 85900 81050 85910 81250
rect 85980 81050 86020 81250
rect 86090 81050 86100 81250
rect 85900 81020 86100 81050
rect 86400 81250 86600 81280
rect 86400 81050 86410 81250
rect 86480 81050 86520 81250
rect 86590 81050 86600 81250
rect 86400 81020 86600 81050
rect 86900 81250 87100 81280
rect 86900 81050 86910 81250
rect 86980 81050 87020 81250
rect 87090 81050 87100 81250
rect 86900 81020 87100 81050
rect 87400 81250 87600 81280
rect 87400 81050 87410 81250
rect 87480 81050 87520 81250
rect 87590 81050 87600 81250
rect 87400 81020 87600 81050
rect 87900 81250 88100 81280
rect 87900 81050 87910 81250
rect 87980 81050 88020 81250
rect 88090 81050 88100 81250
rect 87900 81020 88100 81050
rect 88400 81250 88600 81280
rect 88400 81050 88410 81250
rect 88480 81050 88520 81250
rect 88590 81050 88600 81250
rect 88400 81020 88600 81050
rect 88900 81250 89100 81280
rect 88900 81050 88910 81250
rect 88980 81050 89020 81250
rect 89090 81050 89100 81250
rect 88900 81020 89100 81050
rect 89400 81250 89600 81280
rect 89400 81050 89410 81250
rect 89480 81050 89520 81250
rect 89590 81050 89600 81250
rect 89400 81020 89600 81050
rect 89900 81250 90100 81280
rect 89900 81050 89910 81250
rect 89980 81050 90020 81250
rect 90090 81050 90100 81250
rect 89900 81020 90100 81050
rect 90400 81250 90600 81280
rect 90400 81050 90410 81250
rect 90480 81050 90520 81250
rect 90590 81050 90600 81250
rect 90400 81020 90600 81050
rect 90900 81250 91100 81280
rect 90900 81050 90910 81250
rect 90980 81050 91020 81250
rect 91090 81050 91100 81250
rect 90900 81020 91100 81050
rect 91400 81250 91600 81280
rect 91400 81050 91410 81250
rect 91480 81050 91520 81250
rect 91590 81050 91600 81250
rect 91400 81020 91600 81050
rect 91900 81250 92100 81280
rect 91900 81050 91910 81250
rect 91980 81050 92020 81250
rect 92090 81050 92100 81250
rect 91900 81020 92100 81050
rect 92400 81250 92600 81280
rect 92400 81050 92410 81250
rect 92480 81050 92520 81250
rect 92590 81050 92600 81250
rect 92400 81020 92600 81050
rect 92900 81250 93100 81280
rect 92900 81050 92910 81250
rect 92980 81050 93020 81250
rect 93090 81050 93100 81250
rect 92900 81020 93100 81050
rect 93400 81250 93600 81280
rect 93400 81050 93410 81250
rect 93480 81050 93520 81250
rect 93590 81050 93600 81250
rect 93400 81020 93600 81050
rect 93900 81250 94100 81280
rect 93900 81050 93910 81250
rect 93980 81050 94020 81250
rect 94090 81050 94100 81250
rect 93900 81020 94100 81050
rect 94400 81250 94600 81280
rect 94400 81050 94410 81250
rect 94480 81050 94520 81250
rect 94590 81050 94600 81250
rect 94400 81020 94600 81050
rect 94900 81250 95100 81280
rect 94900 81050 94910 81250
rect 94980 81050 95020 81250
rect 95090 81050 95100 81250
rect 94900 81020 95100 81050
rect 95400 81250 95600 81280
rect 95400 81050 95410 81250
rect 95480 81050 95520 81250
rect 95590 81050 95600 81250
rect 95400 81020 95600 81050
rect 95900 81250 96100 81280
rect 95900 81050 95910 81250
rect 95980 81050 96020 81250
rect 96090 81050 96100 81250
rect 95900 81020 96100 81050
rect 96400 81250 96600 81280
rect 96400 81050 96410 81250
rect 96480 81050 96520 81250
rect 96590 81050 96600 81250
rect 96400 81020 96600 81050
rect 96900 81250 97100 81280
rect 96900 81050 96910 81250
rect 96980 81050 97020 81250
rect 97090 81050 97100 81250
rect 96900 81020 97100 81050
rect 97400 81250 97600 81280
rect 97400 81050 97410 81250
rect 97480 81050 97520 81250
rect 97590 81050 97600 81250
rect 97400 81020 97600 81050
rect 97900 81250 98100 81280
rect 97900 81050 97910 81250
rect 97980 81050 98020 81250
rect 98090 81050 98100 81250
rect 97900 81020 98100 81050
rect 98400 81250 98600 81280
rect 98400 81050 98410 81250
rect 98480 81050 98520 81250
rect 98590 81050 98600 81250
rect 98400 81020 98600 81050
rect 98900 81250 99100 81280
rect 98900 81050 98910 81250
rect 98980 81050 99020 81250
rect 99090 81050 99100 81250
rect 98900 81020 99100 81050
rect 99400 81250 99600 81280
rect 99400 81050 99410 81250
rect 99480 81050 99520 81250
rect 99590 81050 99600 81250
rect 99400 81020 99600 81050
rect 99900 81250 100100 81280
rect 99900 81050 99910 81250
rect 99980 81050 100020 81250
rect 100090 81050 100100 81250
rect 99900 81020 100100 81050
rect 100400 81250 100500 81280
rect 100400 81050 100410 81250
rect 100480 81050 100500 81250
rect 100400 81020 100500 81050
rect -83500 81000 -83380 81020
rect -83120 81000 -82880 81020
rect -82620 81000 -82380 81020
rect -82120 81000 -81880 81020
rect -81620 81000 -81380 81020
rect -81120 81000 -80880 81020
rect -80620 81000 -80380 81020
rect -80120 81000 -79880 81020
rect -79620 81000 -79380 81020
rect -79120 81000 -78880 81020
rect -78620 81000 -78380 81020
rect -78120 81000 -77880 81020
rect -77620 81000 -77380 81020
rect -77120 81000 -76880 81020
rect -76620 81000 -76380 81020
rect -76120 81000 -75880 81020
rect -75620 81000 -75380 81020
rect -75120 81000 -74880 81020
rect -74620 81000 -74380 81020
rect -74120 81000 -73880 81020
rect -73620 81000 -73380 81020
rect -73120 81000 -72880 81020
rect -72620 81000 -72380 81020
rect -72120 81000 -71880 81020
rect -71620 81000 -71380 81020
rect -71120 81000 -70880 81020
rect -70620 81000 -70380 81020
rect -70120 81000 -69880 81020
rect -69620 81000 -69380 81020
rect -69120 81000 -68880 81020
rect -68620 81000 -68380 81020
rect -68120 81000 -67880 81020
rect -67620 81000 -67380 81020
rect -67120 81000 -66880 81020
rect -66620 81000 -66380 81020
rect -66120 81000 -65880 81020
rect -65620 81000 -65380 81020
rect -65120 81000 -64880 81020
rect -64620 81000 -64380 81020
rect -64120 81000 -63880 81020
rect -63620 81000 -63380 81020
rect -63120 81000 -62880 81020
rect -62620 81000 -62380 81020
rect -62120 81000 -61880 81020
rect -61620 81000 -61380 81020
rect -61120 81000 -60880 81020
rect -60620 81000 -60380 81020
rect -60120 81000 -59880 81020
rect -59620 81000 -59380 81020
rect -59120 81000 -58880 81020
rect -58620 81000 -58380 81020
rect -58120 81000 -57880 81020
rect -57620 81000 -57380 81020
rect -57120 81000 -56880 81020
rect -56620 81000 -56380 81020
rect -56120 81000 -55880 81020
rect -55620 81000 -55380 81020
rect -55120 81000 -54880 81020
rect -54620 81000 -54380 81020
rect -54120 81000 -53880 81020
rect -53620 81000 -53380 81020
rect -53120 81000 -52880 81020
rect -52620 81000 -52380 81020
rect -52120 81000 -51880 81020
rect -51620 81000 -51380 81020
rect -51120 81000 -50880 81020
rect -50620 81000 -50380 81020
rect -50120 81000 -49880 81020
rect -49620 81000 -49380 81020
rect -49120 81000 -48880 81020
rect -48620 81000 -48380 81020
rect -48120 81000 -47880 81020
rect -47620 81000 -47380 81020
rect -47120 81000 -46880 81020
rect -46620 81000 -46380 81020
rect -46120 81000 -45880 81020
rect -45620 81000 -45380 81020
rect -45120 81000 -44880 81020
rect -44620 81000 -44380 81020
rect -44120 81000 -43880 81020
rect -43620 81000 -43380 81020
rect -43120 81000 -42880 81020
rect -42620 81000 -42380 81020
rect -42120 81000 -41880 81020
rect -41620 81000 -41380 81020
rect -41120 81000 -40880 81020
rect -40620 81000 -40380 81020
rect -40120 81000 -39880 81020
rect -39620 81000 -39380 81020
rect -39120 81000 -38880 81020
rect -38620 81000 -38380 81020
rect -38120 81000 -37880 81020
rect -37620 81000 -37380 81020
rect -37120 81000 -36880 81020
rect -36620 81000 -36380 81020
rect -36120 81000 -35880 81020
rect -35620 81000 -35380 81020
rect -35120 81000 -34880 81020
rect -34620 81000 -34380 81020
rect -34120 81000 -33880 81020
rect -33620 81000 -33380 81020
rect -33120 81000 -32880 81020
rect -32620 81000 -32380 81020
rect -32120 81000 -31880 81020
rect -31620 81000 -31380 81020
rect -31120 81000 -30880 81020
rect -30620 81000 -30380 81020
rect -30120 81000 -29880 81020
rect -29620 81000 -29380 81020
rect -29120 81000 -28880 81020
rect -28620 81000 -28380 81020
rect -28120 81000 -27880 81020
rect -27620 81000 -27380 81020
rect -27120 81000 -26880 81020
rect -26620 81000 -26380 81020
rect -26120 81000 -25880 81020
rect -25620 81000 -25380 81020
rect -25120 81000 -24880 81020
rect -24620 81000 -24380 81020
rect -24120 81000 -23880 81020
rect -23620 81000 -23380 81020
rect -23120 81000 -22880 81020
rect -22620 81000 -22380 81020
rect -22120 81000 -21880 81020
rect -21620 81000 -21380 81020
rect -21120 81000 -20880 81020
rect -20620 81000 -20380 81020
rect -20120 81000 -19880 81020
rect -19620 81000 -19380 81020
rect -19120 81000 -18880 81020
rect -18620 81000 -18380 81020
rect -18120 81000 -17880 81020
rect -17620 81000 -17380 81020
rect -17120 81000 -16880 81020
rect -16620 81000 -16380 81020
rect -16120 81000 -15880 81020
rect -15620 81000 -15380 81020
rect -15120 81000 -14880 81020
rect -14620 81000 -14380 81020
rect -14120 81000 -13880 81020
rect -13620 81000 -13380 81020
rect -13120 81000 -12880 81020
rect -12620 81000 -12380 81020
rect -12120 81000 -11880 81020
rect -11620 81000 -11380 81020
rect -11120 81000 -10880 81020
rect -10620 81000 -10380 81020
rect -10120 81000 -9880 81020
rect -9620 81000 -9380 81020
rect -9120 81000 -8880 81020
rect -8620 81000 -8380 81020
rect -8120 81000 -7880 81020
rect -7620 81000 -7380 81020
rect -7120 81000 -6880 81020
rect -6620 81000 -6380 81020
rect -6120 81000 -5880 81020
rect -5620 81000 -5380 81020
rect -5120 81000 -4880 81020
rect -4620 81000 -4380 81020
rect -4120 81000 -3880 81020
rect -3620 81000 -3380 81020
rect -3120 81000 -2880 81020
rect -2620 81000 -2380 81020
rect -2120 81000 -1880 81020
rect -1620 81000 -1380 81020
rect -1120 81000 -880 81020
rect -620 81000 -380 81020
rect -120 81000 120 81020
rect 380 81000 620 81020
rect 880 81000 1120 81020
rect 1380 81000 1620 81020
rect 1880 81000 2120 81020
rect 2380 81000 2620 81020
rect 2880 81000 3120 81020
rect 3380 81000 3620 81020
rect 3880 81000 4120 81020
rect 4380 81000 4620 81020
rect 4880 81000 5120 81020
rect 5380 81000 5620 81020
rect 5880 81000 6120 81020
rect 6380 81000 6620 81020
rect 6880 81000 7120 81020
rect 7380 81000 7620 81020
rect 7880 81000 8120 81020
rect 8380 81000 8620 81020
rect 8880 81000 9120 81020
rect 9380 81000 9620 81020
rect 9880 81000 10120 81020
rect 10380 81000 10620 81020
rect 10880 81000 11120 81020
rect 11380 81000 11620 81020
rect 11880 81000 12120 81020
rect 12380 81000 12620 81020
rect 12880 81000 13120 81020
rect 13380 81000 13620 81020
rect 13880 81000 14120 81020
rect 14380 81000 14620 81020
rect 14880 81000 15120 81020
rect 15380 81000 15620 81020
rect 15880 81000 16120 81020
rect 16380 81000 16620 81020
rect 16880 81000 17120 81020
rect 17380 81000 17620 81020
rect 17880 81000 18120 81020
rect 18380 81000 18620 81020
rect 18880 81000 19120 81020
rect 19380 81000 19620 81020
rect 19880 81000 20120 81020
rect 20380 81000 20620 81020
rect 20880 81000 21120 81020
rect 21380 81000 21620 81020
rect 21880 81000 22120 81020
rect 22380 81000 22620 81020
rect 22880 81000 23120 81020
rect 23380 81000 23620 81020
rect 23880 81000 24120 81020
rect 24380 81000 24620 81020
rect 24880 81000 25120 81020
rect 25380 81000 25620 81020
rect 25880 81000 26120 81020
rect 26380 81000 26620 81020
rect 26880 81000 27120 81020
rect 27380 81000 27620 81020
rect 27880 81000 28120 81020
rect 28380 81000 28620 81020
rect 28880 81000 29120 81020
rect 29380 81000 29620 81020
rect 29880 81000 30120 81020
rect 30380 81000 30620 81020
rect 30880 81000 31120 81020
rect 31380 81000 31620 81020
rect 31880 81000 32120 81020
rect 32380 81000 32620 81020
rect 32880 81000 33120 81020
rect 33380 81000 33620 81020
rect 33880 81000 34120 81020
rect 34380 81000 34620 81020
rect 34880 81000 35120 81020
rect 35380 81000 35620 81020
rect 35880 81000 36120 81020
rect 36380 81000 36620 81020
rect 36880 81000 37120 81020
rect 37380 81000 37620 81020
rect 37880 81000 38120 81020
rect 38380 81000 38620 81020
rect 38880 81000 39120 81020
rect 39380 81000 39620 81020
rect 39880 81000 40120 81020
rect 40380 81000 40620 81020
rect 40880 81000 41120 81020
rect 41380 81000 41620 81020
rect 41880 81000 42120 81020
rect 42380 81000 42620 81020
rect 42880 81000 43120 81020
rect 43380 81000 43620 81020
rect 43880 81000 44120 81020
rect 44380 81000 44620 81020
rect 44880 81000 45120 81020
rect 45380 81000 45620 81020
rect 45880 81000 46120 81020
rect 46380 81000 46620 81020
rect 46880 81000 47120 81020
rect 47380 81000 47620 81020
rect 47880 81000 48120 81020
rect 48380 81000 48620 81020
rect 48880 81000 49120 81020
rect 49380 81000 49620 81020
rect 49880 81000 50120 81020
rect 50380 81000 50620 81020
rect 50880 81000 51120 81020
rect 51380 81000 51620 81020
rect 51880 81000 52120 81020
rect 52380 81000 52620 81020
rect 52880 81000 53120 81020
rect 53380 81000 53620 81020
rect 53880 81000 54120 81020
rect 54380 81000 54620 81020
rect 54880 81000 55120 81020
rect 55380 81000 55620 81020
rect 55880 81000 56120 81020
rect 56380 81000 56620 81020
rect 56880 81000 57120 81020
rect 57380 81000 57620 81020
rect 57880 81000 58120 81020
rect 58380 81000 58620 81020
rect 58880 81000 59120 81020
rect 59380 81000 59620 81020
rect 59880 81000 60120 81020
rect 60380 81000 60620 81020
rect 60880 81000 61120 81020
rect 61380 81000 61620 81020
rect 61880 81000 62120 81020
rect 62380 81000 62620 81020
rect 62880 81000 63120 81020
rect 63380 81000 63620 81020
rect 63880 81000 64120 81020
rect 64380 81000 64620 81020
rect 64880 81000 65120 81020
rect 65380 81000 65620 81020
rect 65880 81000 66120 81020
rect 66380 81000 66620 81020
rect 66880 81000 67120 81020
rect 67380 81000 67620 81020
rect 67880 81000 68120 81020
rect 68380 81000 68620 81020
rect 68880 81000 69120 81020
rect 69380 81000 69620 81020
rect 69880 81000 70120 81020
rect 70380 81000 70620 81020
rect 70880 81000 71120 81020
rect 71380 81000 71620 81020
rect 71880 81000 72120 81020
rect 72380 81000 72620 81020
rect 72880 81000 73120 81020
rect 73380 81000 73620 81020
rect 73880 81000 74120 81020
rect 74380 81000 74620 81020
rect 74880 81000 75120 81020
rect 75380 81000 75620 81020
rect 75880 81000 76120 81020
rect 76380 81000 76620 81020
rect 76880 81000 77120 81020
rect 77380 81000 77620 81020
rect 77880 81000 78120 81020
rect 78380 81000 78620 81020
rect 78880 81000 79120 81020
rect 79380 81000 79620 81020
rect 79880 81000 80120 81020
rect 80380 81000 80620 81020
rect 80880 81000 81120 81020
rect 81380 81000 81620 81020
rect 81880 81000 82120 81020
rect 82380 81000 82620 81020
rect 82880 81000 83120 81020
rect 83380 81000 83620 81020
rect 83880 81000 84120 81020
rect 84380 81000 84620 81020
rect 84880 81000 85120 81020
rect 85380 81000 85620 81020
rect 85880 81000 86120 81020
rect 86380 81000 86620 81020
rect 86880 81000 87120 81020
rect 87380 81000 87620 81020
rect 87880 81000 88120 81020
rect 88380 81000 88620 81020
rect 88880 81000 89120 81020
rect 89380 81000 89620 81020
rect 89880 81000 90120 81020
rect 90380 81000 90620 81020
rect 90880 81000 91120 81020
rect 91380 81000 91620 81020
rect 91880 81000 92120 81020
rect 92380 81000 92620 81020
rect 92880 81000 93120 81020
rect 93380 81000 93620 81020
rect 93880 81000 94120 81020
rect 94380 81000 94620 81020
rect 94880 81000 95120 81020
rect 95380 81000 95620 81020
rect 95880 81000 96120 81020
rect 96380 81000 96620 81020
rect 96880 81000 97120 81020
rect 97380 81000 97620 81020
rect 97880 81000 98120 81020
rect 98380 81000 98620 81020
rect 98880 81000 99120 81020
rect 99380 81000 99620 81020
rect 99880 81000 100120 81020
rect 100380 81000 100500 81020
rect -83500 80990 100500 81000
rect -83500 80920 -83350 80990
rect -83150 80920 -82850 80990
rect -82650 80920 -82350 80990
rect -82150 80920 -81850 80990
rect -81650 80920 -81350 80990
rect -81150 80920 -80850 80990
rect -80650 80920 -80350 80990
rect -80150 80920 -79850 80990
rect -79650 80920 -79350 80990
rect -79150 80920 -78850 80990
rect -78650 80920 -78350 80990
rect -78150 80920 -77850 80990
rect -77650 80920 -77350 80990
rect -77150 80920 -76850 80990
rect -76650 80920 -76350 80990
rect -76150 80920 -75850 80990
rect -75650 80920 -75350 80990
rect -75150 80920 -74850 80990
rect -74650 80920 -74350 80990
rect -74150 80920 -73850 80990
rect -73650 80920 -73350 80990
rect -73150 80920 -72850 80990
rect -72650 80920 -72350 80990
rect -72150 80920 -71850 80990
rect -71650 80920 -71350 80990
rect -71150 80920 -70850 80990
rect -70650 80920 -70350 80990
rect -70150 80920 -69850 80990
rect -69650 80920 -69350 80990
rect -69150 80920 -68850 80990
rect -68650 80920 -68350 80990
rect -68150 80920 -67850 80990
rect -67650 80920 -67350 80990
rect -67150 80920 -66850 80990
rect -66650 80920 -66350 80990
rect -66150 80920 -65850 80990
rect -65650 80920 -65350 80990
rect -65150 80920 -64850 80990
rect -64650 80920 -64350 80990
rect -64150 80920 -63850 80990
rect -63650 80920 -63350 80990
rect -63150 80920 -62850 80990
rect -62650 80920 -62350 80990
rect -62150 80920 -61850 80990
rect -61650 80920 -61350 80990
rect -61150 80920 -60850 80990
rect -60650 80920 -60350 80990
rect -60150 80920 -59850 80990
rect -59650 80920 -59350 80990
rect -59150 80920 -58850 80990
rect -58650 80920 -58350 80990
rect -58150 80920 -57850 80990
rect -57650 80920 -57350 80990
rect -57150 80920 -56850 80990
rect -56650 80920 -56350 80990
rect -56150 80920 -55850 80990
rect -55650 80920 -55350 80990
rect -55150 80920 -54850 80990
rect -54650 80920 -54350 80990
rect -54150 80920 -53850 80990
rect -53650 80920 -53350 80990
rect -53150 80920 -52850 80990
rect -52650 80920 -52350 80990
rect -52150 80920 -51850 80990
rect -51650 80920 -51350 80990
rect -51150 80920 -50850 80990
rect -50650 80920 -50350 80990
rect -50150 80920 -49850 80990
rect -49650 80920 -49350 80990
rect -49150 80920 -48850 80990
rect -48650 80920 -48350 80990
rect -48150 80920 -47850 80990
rect -47650 80920 -47350 80990
rect -47150 80920 -46850 80990
rect -46650 80920 -46350 80990
rect -46150 80920 -45850 80990
rect -45650 80920 -45350 80990
rect -45150 80920 -44850 80990
rect -44650 80920 -44350 80990
rect -44150 80920 -43850 80990
rect -43650 80920 -43350 80990
rect -43150 80920 -42850 80990
rect -42650 80920 -42350 80990
rect -42150 80920 -41850 80990
rect -41650 80920 -41350 80990
rect -41150 80920 -40850 80990
rect -40650 80920 -40350 80990
rect -40150 80920 -39850 80990
rect -39650 80920 -39350 80990
rect -39150 80920 -38850 80990
rect -38650 80920 -38350 80990
rect -38150 80920 -37850 80990
rect -37650 80920 -37350 80990
rect -37150 80920 -36850 80990
rect -36650 80920 -36350 80990
rect -36150 80920 -35850 80990
rect -35650 80920 -35350 80990
rect -35150 80920 -34850 80990
rect -34650 80920 -34350 80990
rect -34150 80920 -33850 80990
rect -33650 80920 -33350 80990
rect -33150 80920 -32850 80990
rect -32650 80920 -32350 80990
rect -32150 80920 -31850 80990
rect -31650 80920 -31350 80990
rect -31150 80920 -30850 80990
rect -30650 80920 -30350 80990
rect -30150 80920 -29850 80990
rect -29650 80920 -29350 80990
rect -29150 80920 -28850 80990
rect -28650 80920 -28350 80990
rect -28150 80920 -27850 80990
rect -27650 80920 -27350 80990
rect -27150 80920 -26850 80990
rect -26650 80920 -26350 80990
rect -26150 80920 -25850 80990
rect -25650 80920 -25350 80990
rect -25150 80920 -24850 80990
rect -24650 80920 -24350 80990
rect -24150 80920 -23850 80990
rect -23650 80920 -23350 80990
rect -23150 80920 -22850 80990
rect -22650 80920 -22350 80990
rect -22150 80920 -21850 80990
rect -21650 80920 -21350 80990
rect -21150 80920 -20850 80990
rect -20650 80920 -20350 80990
rect -20150 80920 -19850 80990
rect -19650 80920 -19350 80990
rect -19150 80920 -18850 80990
rect -18650 80920 -18350 80990
rect -18150 80920 -17850 80990
rect -17650 80920 -17350 80990
rect -17150 80920 -16850 80990
rect -16650 80920 -16350 80990
rect -16150 80920 -15850 80990
rect -15650 80920 -15350 80990
rect -15150 80920 -14850 80990
rect -14650 80920 -14350 80990
rect -14150 80920 -13850 80990
rect -13650 80920 -13350 80990
rect -13150 80920 -12850 80990
rect -12650 80920 -12350 80990
rect -12150 80920 -11850 80990
rect -11650 80920 -11350 80990
rect -11150 80920 -10850 80990
rect -10650 80920 -10350 80990
rect -10150 80920 -9850 80990
rect -9650 80920 -9350 80990
rect -9150 80920 -8850 80990
rect -8650 80920 -8350 80990
rect -8150 80920 -7850 80990
rect -7650 80920 -7350 80990
rect -7150 80920 -6850 80990
rect -6650 80920 -6350 80990
rect -6150 80920 -5850 80990
rect -5650 80920 -5350 80990
rect -5150 80920 -4850 80990
rect -4650 80920 -4350 80990
rect -4150 80920 -3850 80990
rect -3650 80920 -3350 80990
rect -3150 80920 -2850 80990
rect -2650 80920 -2350 80990
rect -2150 80920 -1850 80990
rect -1650 80920 -1350 80990
rect -1150 80920 -850 80990
rect -650 80920 -350 80990
rect -150 80920 150 80990
rect 350 80920 650 80990
rect 850 80920 1150 80990
rect 1350 80920 1650 80990
rect 1850 80920 2150 80990
rect 2350 80920 2650 80990
rect 2850 80920 3150 80990
rect 3350 80920 3650 80990
rect 3850 80920 4150 80990
rect 4350 80920 4650 80990
rect 4850 80920 5150 80990
rect 5350 80920 5650 80990
rect 5850 80920 6150 80990
rect 6350 80920 6650 80990
rect 6850 80920 7150 80990
rect 7350 80920 7650 80990
rect 7850 80920 8150 80990
rect 8350 80920 8650 80990
rect 8850 80920 9150 80990
rect 9350 80920 9650 80990
rect 9850 80920 10150 80990
rect 10350 80920 10650 80990
rect 10850 80920 11150 80990
rect 11350 80920 11650 80990
rect 11850 80920 12150 80990
rect 12350 80920 12650 80990
rect 12850 80920 13150 80990
rect 13350 80920 13650 80990
rect 13850 80920 14150 80990
rect 14350 80920 14650 80990
rect 14850 80920 15150 80990
rect 15350 80920 15650 80990
rect 15850 80920 16150 80990
rect 16350 80920 16650 80990
rect 16850 80920 17150 80990
rect 17350 80920 17650 80990
rect 17850 80920 18150 80990
rect 18350 80920 18650 80990
rect 18850 80920 19150 80990
rect 19350 80920 19650 80990
rect 19850 80920 20150 80990
rect 20350 80920 20650 80990
rect 20850 80920 21150 80990
rect 21350 80920 21650 80990
rect 21850 80920 22150 80990
rect 22350 80920 22650 80990
rect 22850 80920 23150 80990
rect 23350 80920 23650 80990
rect 23850 80920 24150 80990
rect 24350 80920 24650 80990
rect 24850 80920 25150 80990
rect 25350 80920 25650 80990
rect 25850 80920 26150 80990
rect 26350 80920 26650 80990
rect 26850 80920 27150 80990
rect 27350 80920 27650 80990
rect 27850 80920 28150 80990
rect 28350 80920 28650 80990
rect 28850 80920 29150 80990
rect 29350 80920 29650 80990
rect 29850 80920 30150 80990
rect 30350 80920 30650 80990
rect 30850 80920 31150 80990
rect 31350 80920 31650 80990
rect 31850 80920 32150 80990
rect 32350 80920 32650 80990
rect 32850 80920 33150 80990
rect 33350 80920 33650 80990
rect 33850 80920 34150 80990
rect 34350 80920 34650 80990
rect 34850 80920 35150 80990
rect 35350 80920 35650 80990
rect 35850 80920 36150 80990
rect 36350 80920 36650 80990
rect 36850 80920 37150 80990
rect 37350 80920 37650 80990
rect 37850 80920 38150 80990
rect 38350 80920 38650 80990
rect 38850 80920 39150 80990
rect 39350 80920 39650 80990
rect 39850 80920 40150 80990
rect 40350 80920 40650 80990
rect 40850 80920 41150 80990
rect 41350 80920 41650 80990
rect 41850 80920 42150 80990
rect 42350 80920 42650 80990
rect 42850 80920 43150 80990
rect 43350 80920 43650 80990
rect 43850 80920 44150 80990
rect 44350 80920 44650 80990
rect 44850 80920 45150 80990
rect 45350 80920 45650 80990
rect 45850 80920 46150 80990
rect 46350 80920 46650 80990
rect 46850 80920 47150 80990
rect 47350 80920 47650 80990
rect 47850 80920 48150 80990
rect 48350 80920 48650 80990
rect 48850 80920 49150 80990
rect 49350 80920 49650 80990
rect 49850 80920 50150 80990
rect 50350 80920 50650 80990
rect 50850 80920 51150 80990
rect 51350 80920 51650 80990
rect 51850 80920 52150 80990
rect 52350 80920 52650 80990
rect 52850 80920 53150 80990
rect 53350 80920 53650 80990
rect 53850 80920 54150 80990
rect 54350 80920 54650 80990
rect 54850 80920 55150 80990
rect 55350 80920 55650 80990
rect 55850 80920 56150 80990
rect 56350 80920 56650 80990
rect 56850 80920 57150 80990
rect 57350 80920 57650 80990
rect 57850 80920 58150 80990
rect 58350 80920 58650 80990
rect 58850 80920 59150 80990
rect 59350 80920 59650 80990
rect 59850 80920 60150 80990
rect 60350 80920 60650 80990
rect 60850 80920 61150 80990
rect 61350 80920 61650 80990
rect 61850 80920 62150 80990
rect 62350 80920 62650 80990
rect 62850 80920 63150 80990
rect 63350 80920 63650 80990
rect 63850 80920 64150 80990
rect 64350 80920 64650 80990
rect 64850 80920 65150 80990
rect 65350 80920 65650 80990
rect 65850 80920 66150 80990
rect 66350 80920 66650 80990
rect 66850 80920 67150 80990
rect 67350 80920 67650 80990
rect 67850 80920 68150 80990
rect 68350 80920 68650 80990
rect 68850 80920 69150 80990
rect 69350 80920 69650 80990
rect 69850 80920 70150 80990
rect 70350 80920 70650 80990
rect 70850 80920 71150 80990
rect 71350 80920 71650 80990
rect 71850 80920 72150 80990
rect 72350 80920 72650 80990
rect 72850 80920 73150 80990
rect 73350 80920 73650 80990
rect 73850 80920 74150 80990
rect 74350 80920 74650 80990
rect 74850 80920 75150 80990
rect 75350 80920 75650 80990
rect 75850 80920 76150 80990
rect 76350 80920 76650 80990
rect 76850 80920 77150 80990
rect 77350 80920 77650 80990
rect 77850 80920 78150 80990
rect 78350 80920 78650 80990
rect 78850 80920 79150 80990
rect 79350 80920 79650 80990
rect 79850 80920 80150 80990
rect 80350 80920 80650 80990
rect 80850 80920 81150 80990
rect 81350 80920 81650 80990
rect 81850 80920 82150 80990
rect 82350 80920 82650 80990
rect 82850 80920 83150 80990
rect 83350 80920 83650 80990
rect 83850 80920 84150 80990
rect 84350 80920 84650 80990
rect 84850 80920 85150 80990
rect 85350 80920 85650 80990
rect 85850 80920 86150 80990
rect 86350 80920 86650 80990
rect 86850 80920 87150 80990
rect 87350 80920 87650 80990
rect 87850 80920 88150 80990
rect 88350 80920 88650 80990
rect 88850 80920 89150 80990
rect 89350 80920 89650 80990
rect 89850 80920 90150 80990
rect 90350 80920 90650 80990
rect 90850 80920 91150 80990
rect 91350 80920 91650 80990
rect 91850 80920 92150 80990
rect 92350 80920 92650 80990
rect 92850 80920 93150 80990
rect 93350 80920 93650 80990
rect 93850 80920 94150 80990
rect 94350 80920 94650 80990
rect 94850 80920 95150 80990
rect 95350 80920 95650 80990
rect 95850 80920 96150 80990
rect 96350 80920 96650 80990
rect 96850 80920 97150 80990
rect 97350 80920 97650 80990
rect 97850 80920 98150 80990
rect 98350 80920 98650 80990
rect 98850 80920 99150 80990
rect 99350 80920 99650 80990
rect 99850 80920 100150 80990
rect 100350 80920 100500 80990
rect -83500 80880 100500 80920
rect -83500 80810 -83350 80880
rect -83150 80810 -82850 80880
rect -82650 80810 -82350 80880
rect -82150 80810 -81850 80880
rect -81650 80810 -81350 80880
rect -81150 80810 -80850 80880
rect -80650 80810 -80350 80880
rect -80150 80810 -79850 80880
rect -79650 80810 -79350 80880
rect -79150 80810 -78850 80880
rect -78650 80810 -78350 80880
rect -78150 80810 -77850 80880
rect -77650 80810 -77350 80880
rect -77150 80810 -76850 80880
rect -76650 80810 -76350 80880
rect -76150 80810 -75850 80880
rect -75650 80810 -75350 80880
rect -75150 80810 -74850 80880
rect -74650 80810 -74350 80880
rect -74150 80810 -73850 80880
rect -73650 80810 -73350 80880
rect -73150 80810 -72850 80880
rect -72650 80810 -72350 80880
rect -72150 80810 -71850 80880
rect -71650 80810 -71350 80880
rect -71150 80810 -70850 80880
rect -70650 80810 -70350 80880
rect -70150 80810 -69850 80880
rect -69650 80810 -69350 80880
rect -69150 80810 -68850 80880
rect -68650 80810 -68350 80880
rect -68150 80810 -67850 80880
rect -67650 80810 -67350 80880
rect -67150 80810 -66850 80880
rect -66650 80810 -66350 80880
rect -66150 80810 -65850 80880
rect -65650 80810 -65350 80880
rect -65150 80810 -64850 80880
rect -64650 80810 -64350 80880
rect -64150 80810 -63850 80880
rect -63650 80810 -63350 80880
rect -63150 80810 -62850 80880
rect -62650 80810 -62350 80880
rect -62150 80810 -61850 80880
rect -61650 80810 -61350 80880
rect -61150 80810 -60850 80880
rect -60650 80810 -60350 80880
rect -60150 80810 -59850 80880
rect -59650 80810 -59350 80880
rect -59150 80810 -58850 80880
rect -58650 80810 -58350 80880
rect -58150 80810 -57850 80880
rect -57650 80810 -57350 80880
rect -57150 80810 -56850 80880
rect -56650 80810 -56350 80880
rect -56150 80810 -55850 80880
rect -55650 80810 -55350 80880
rect -55150 80810 -54850 80880
rect -54650 80810 -54350 80880
rect -54150 80810 -53850 80880
rect -53650 80810 -53350 80880
rect -53150 80810 -52850 80880
rect -52650 80810 -52350 80880
rect -52150 80810 -51850 80880
rect -51650 80810 -51350 80880
rect -51150 80810 -50850 80880
rect -50650 80810 -50350 80880
rect -50150 80810 -49850 80880
rect -49650 80810 -49350 80880
rect -49150 80810 -48850 80880
rect -48650 80810 -48350 80880
rect -48150 80810 -47850 80880
rect -47650 80810 -47350 80880
rect -47150 80810 -46850 80880
rect -46650 80810 -46350 80880
rect -46150 80810 -45850 80880
rect -45650 80810 -45350 80880
rect -45150 80810 -44850 80880
rect -44650 80810 -44350 80880
rect -44150 80810 -43850 80880
rect -43650 80810 -43350 80880
rect -43150 80810 -42850 80880
rect -42650 80810 -42350 80880
rect -42150 80810 -41850 80880
rect -41650 80810 -41350 80880
rect -41150 80810 -40850 80880
rect -40650 80810 -40350 80880
rect -40150 80810 -39850 80880
rect -39650 80810 -39350 80880
rect -39150 80810 -38850 80880
rect -38650 80810 -38350 80880
rect -38150 80810 -37850 80880
rect -37650 80810 -37350 80880
rect -37150 80810 -36850 80880
rect -36650 80810 -36350 80880
rect -36150 80810 -35850 80880
rect -35650 80810 -35350 80880
rect -35150 80810 -34850 80880
rect -34650 80810 -34350 80880
rect -34150 80810 -33850 80880
rect -33650 80810 -33350 80880
rect -33150 80810 -32850 80880
rect -32650 80810 -32350 80880
rect -32150 80810 -31850 80880
rect -31650 80810 -31350 80880
rect -31150 80810 -30850 80880
rect -30650 80810 -30350 80880
rect -30150 80810 -29850 80880
rect -29650 80810 -29350 80880
rect -29150 80810 -28850 80880
rect -28650 80810 -28350 80880
rect -28150 80810 -27850 80880
rect -27650 80810 -27350 80880
rect -27150 80810 -26850 80880
rect -26650 80810 -26350 80880
rect -26150 80810 -25850 80880
rect -25650 80810 -25350 80880
rect -25150 80810 -24850 80880
rect -24650 80810 -24350 80880
rect -24150 80810 -23850 80880
rect -23650 80810 -23350 80880
rect -23150 80810 -22850 80880
rect -22650 80810 -22350 80880
rect -22150 80810 -21850 80880
rect -21650 80810 -21350 80880
rect -21150 80810 -20850 80880
rect -20650 80810 -20350 80880
rect -20150 80810 -19850 80880
rect -19650 80810 -19350 80880
rect -19150 80810 -18850 80880
rect -18650 80810 -18350 80880
rect -18150 80810 -17850 80880
rect -17650 80810 -17350 80880
rect -17150 80810 -16850 80880
rect -16650 80810 -16350 80880
rect -16150 80810 -15850 80880
rect -15650 80810 -15350 80880
rect -15150 80810 -14850 80880
rect -14650 80810 -14350 80880
rect -14150 80810 -13850 80880
rect -13650 80810 -13350 80880
rect -13150 80810 -12850 80880
rect -12650 80810 -12350 80880
rect -12150 80810 -11850 80880
rect -11650 80810 -11350 80880
rect -11150 80810 -10850 80880
rect -10650 80810 -10350 80880
rect -10150 80810 -9850 80880
rect -9650 80810 -9350 80880
rect -9150 80810 -8850 80880
rect -8650 80810 -8350 80880
rect -8150 80810 -7850 80880
rect -7650 80810 -7350 80880
rect -7150 80810 -6850 80880
rect -6650 80810 -6350 80880
rect -6150 80810 -5850 80880
rect -5650 80810 -5350 80880
rect -5150 80810 -4850 80880
rect -4650 80810 -4350 80880
rect -4150 80810 -3850 80880
rect -3650 80810 -3350 80880
rect -3150 80810 -2850 80880
rect -2650 80810 -2350 80880
rect -2150 80810 -1850 80880
rect -1650 80810 -1350 80880
rect -1150 80810 -850 80880
rect -650 80810 -350 80880
rect -150 80810 150 80880
rect 350 80810 650 80880
rect 850 80810 1150 80880
rect 1350 80810 1650 80880
rect 1850 80810 2150 80880
rect 2350 80810 2650 80880
rect 2850 80810 3150 80880
rect 3350 80810 3650 80880
rect 3850 80810 4150 80880
rect 4350 80810 4650 80880
rect 4850 80810 5150 80880
rect 5350 80810 5650 80880
rect 5850 80810 6150 80880
rect 6350 80810 6650 80880
rect 6850 80810 7150 80880
rect 7350 80810 7650 80880
rect 7850 80810 8150 80880
rect 8350 80810 8650 80880
rect 8850 80810 9150 80880
rect 9350 80810 9650 80880
rect 9850 80810 10150 80880
rect 10350 80810 10650 80880
rect 10850 80810 11150 80880
rect 11350 80810 11650 80880
rect 11850 80810 12150 80880
rect 12350 80810 12650 80880
rect 12850 80810 13150 80880
rect 13350 80810 13650 80880
rect 13850 80810 14150 80880
rect 14350 80810 14650 80880
rect 14850 80810 15150 80880
rect 15350 80810 15650 80880
rect 15850 80810 16150 80880
rect 16350 80810 16650 80880
rect 16850 80810 17150 80880
rect 17350 80810 17650 80880
rect 17850 80810 18150 80880
rect 18350 80810 18650 80880
rect 18850 80810 19150 80880
rect 19350 80810 19650 80880
rect 19850 80810 20150 80880
rect 20350 80810 20650 80880
rect 20850 80810 21150 80880
rect 21350 80810 21650 80880
rect 21850 80810 22150 80880
rect 22350 80810 22650 80880
rect 22850 80810 23150 80880
rect 23350 80810 23650 80880
rect 23850 80810 24150 80880
rect 24350 80810 24650 80880
rect 24850 80810 25150 80880
rect 25350 80810 25650 80880
rect 25850 80810 26150 80880
rect 26350 80810 26650 80880
rect 26850 80810 27150 80880
rect 27350 80810 27650 80880
rect 27850 80810 28150 80880
rect 28350 80810 28650 80880
rect 28850 80810 29150 80880
rect 29350 80810 29650 80880
rect 29850 80810 30150 80880
rect 30350 80810 30650 80880
rect 30850 80810 31150 80880
rect 31350 80810 31650 80880
rect 31850 80810 32150 80880
rect 32350 80810 32650 80880
rect 32850 80810 33150 80880
rect 33350 80810 33650 80880
rect 33850 80810 34150 80880
rect 34350 80810 34650 80880
rect 34850 80810 35150 80880
rect 35350 80810 35650 80880
rect 35850 80810 36150 80880
rect 36350 80810 36650 80880
rect 36850 80810 37150 80880
rect 37350 80810 37650 80880
rect 37850 80810 38150 80880
rect 38350 80810 38650 80880
rect 38850 80810 39150 80880
rect 39350 80810 39650 80880
rect 39850 80810 40150 80880
rect 40350 80810 40650 80880
rect 40850 80810 41150 80880
rect 41350 80810 41650 80880
rect 41850 80810 42150 80880
rect 42350 80810 42650 80880
rect 42850 80810 43150 80880
rect 43350 80810 43650 80880
rect 43850 80810 44150 80880
rect 44350 80810 44650 80880
rect 44850 80810 45150 80880
rect 45350 80810 45650 80880
rect 45850 80810 46150 80880
rect 46350 80810 46650 80880
rect 46850 80810 47150 80880
rect 47350 80810 47650 80880
rect 47850 80810 48150 80880
rect 48350 80810 48650 80880
rect 48850 80810 49150 80880
rect 49350 80810 49650 80880
rect 49850 80810 50150 80880
rect 50350 80810 50650 80880
rect 50850 80810 51150 80880
rect 51350 80810 51650 80880
rect 51850 80810 52150 80880
rect 52350 80810 52650 80880
rect 52850 80810 53150 80880
rect 53350 80810 53650 80880
rect 53850 80810 54150 80880
rect 54350 80810 54650 80880
rect 54850 80810 55150 80880
rect 55350 80810 55650 80880
rect 55850 80810 56150 80880
rect 56350 80810 56650 80880
rect 56850 80810 57150 80880
rect 57350 80810 57650 80880
rect 57850 80810 58150 80880
rect 58350 80810 58650 80880
rect 58850 80810 59150 80880
rect 59350 80810 59650 80880
rect 59850 80810 60150 80880
rect 60350 80810 60650 80880
rect 60850 80810 61150 80880
rect 61350 80810 61650 80880
rect 61850 80810 62150 80880
rect 62350 80810 62650 80880
rect 62850 80810 63150 80880
rect 63350 80810 63650 80880
rect 63850 80810 64150 80880
rect 64350 80810 64650 80880
rect 64850 80810 65150 80880
rect 65350 80810 65650 80880
rect 65850 80810 66150 80880
rect 66350 80810 66650 80880
rect 66850 80810 67150 80880
rect 67350 80810 67650 80880
rect 67850 80810 68150 80880
rect 68350 80810 68650 80880
rect 68850 80810 69150 80880
rect 69350 80810 69650 80880
rect 69850 80810 70150 80880
rect 70350 80810 70650 80880
rect 70850 80810 71150 80880
rect 71350 80810 71650 80880
rect 71850 80810 72150 80880
rect 72350 80810 72650 80880
rect 72850 80810 73150 80880
rect 73350 80810 73650 80880
rect 73850 80810 74150 80880
rect 74350 80810 74650 80880
rect 74850 80810 75150 80880
rect 75350 80810 75650 80880
rect 75850 80810 76150 80880
rect 76350 80810 76650 80880
rect 76850 80810 77150 80880
rect 77350 80810 77650 80880
rect 77850 80810 78150 80880
rect 78350 80810 78650 80880
rect 78850 80810 79150 80880
rect 79350 80810 79650 80880
rect 79850 80810 80150 80880
rect 80350 80810 80650 80880
rect 80850 80810 81150 80880
rect 81350 80810 81650 80880
rect 81850 80810 82150 80880
rect 82350 80810 82650 80880
rect 82850 80810 83150 80880
rect 83350 80810 83650 80880
rect 83850 80810 84150 80880
rect 84350 80810 84650 80880
rect 84850 80810 85150 80880
rect 85350 80810 85650 80880
rect 85850 80810 86150 80880
rect 86350 80810 86650 80880
rect 86850 80810 87150 80880
rect 87350 80810 87650 80880
rect 87850 80810 88150 80880
rect 88350 80810 88650 80880
rect 88850 80810 89150 80880
rect 89350 80810 89650 80880
rect 89850 80810 90150 80880
rect 90350 80810 90650 80880
rect 90850 80810 91150 80880
rect 91350 80810 91650 80880
rect 91850 80810 92150 80880
rect 92350 80810 92650 80880
rect 92850 80810 93150 80880
rect 93350 80810 93650 80880
rect 93850 80810 94150 80880
rect 94350 80810 94650 80880
rect 94850 80810 95150 80880
rect 95350 80810 95650 80880
rect 95850 80810 96150 80880
rect 96350 80810 96650 80880
rect 96850 80810 97150 80880
rect 97350 80810 97650 80880
rect 97850 80810 98150 80880
rect 98350 80810 98650 80880
rect 98850 80810 99150 80880
rect 99350 80810 99650 80880
rect 99850 80810 100150 80880
rect 100350 80810 100500 80880
rect -83500 80800 100500 80810
rect -83500 80780 -83380 80800
rect -83120 80780 -82880 80800
rect -82620 80780 -82380 80800
rect -82120 80780 -81880 80800
rect -81620 80780 -81380 80800
rect -81120 80780 -80880 80800
rect -80620 80780 -80380 80800
rect -80120 80780 -79880 80800
rect -79620 80780 -79380 80800
rect -79120 80780 -78880 80800
rect -78620 80780 -78380 80800
rect -78120 80780 -77880 80800
rect -77620 80780 -77380 80800
rect -77120 80780 -76880 80800
rect -76620 80780 -76380 80800
rect -76120 80780 -75880 80800
rect -75620 80780 -75380 80800
rect -75120 80780 -74880 80800
rect -74620 80780 -74380 80800
rect -74120 80780 -73880 80800
rect -73620 80780 -73380 80800
rect -73120 80780 -72880 80800
rect -72620 80780 -72380 80800
rect -72120 80780 -71880 80800
rect -71620 80780 -71380 80800
rect -71120 80780 -70880 80800
rect -70620 80780 -70380 80800
rect -70120 80780 -69880 80800
rect -69620 80780 -69380 80800
rect -69120 80780 -68880 80800
rect -68620 80780 -68380 80800
rect -68120 80780 -67880 80800
rect -67620 80780 -67380 80800
rect -67120 80780 -66880 80800
rect -66620 80780 -66380 80800
rect -66120 80780 -65880 80800
rect -65620 80780 -65380 80800
rect -65120 80780 -64880 80800
rect -64620 80780 -64380 80800
rect -64120 80780 -63880 80800
rect -63620 80780 -63380 80800
rect -63120 80780 -62880 80800
rect -62620 80780 -62380 80800
rect -62120 80780 -61880 80800
rect -61620 80780 -61380 80800
rect -61120 80780 -60880 80800
rect -60620 80780 -60380 80800
rect -60120 80780 -59880 80800
rect -59620 80780 -59380 80800
rect -59120 80780 -58880 80800
rect -58620 80780 -58380 80800
rect -58120 80780 -57880 80800
rect -57620 80780 -57380 80800
rect -57120 80780 -56880 80800
rect -56620 80780 -56380 80800
rect -56120 80780 -55880 80800
rect -55620 80780 -55380 80800
rect -55120 80780 -54880 80800
rect -54620 80780 -54380 80800
rect -54120 80780 -53880 80800
rect -53620 80780 -53380 80800
rect -53120 80780 -52880 80800
rect -52620 80780 -52380 80800
rect -52120 80780 -51880 80800
rect -51620 80780 -51380 80800
rect -51120 80780 -50880 80800
rect -50620 80780 -50380 80800
rect -50120 80780 -49880 80800
rect -49620 80780 -49380 80800
rect -49120 80780 -48880 80800
rect -48620 80780 -48380 80800
rect -48120 80780 -47880 80800
rect -47620 80780 -47380 80800
rect -47120 80780 -46880 80800
rect -46620 80780 -46380 80800
rect -46120 80780 -45880 80800
rect -45620 80780 -45380 80800
rect -45120 80780 -44880 80800
rect -44620 80780 -44380 80800
rect -44120 80780 -43880 80800
rect -43620 80780 -43380 80800
rect -43120 80780 -42880 80800
rect -42620 80780 -42380 80800
rect -42120 80780 -41880 80800
rect -41620 80780 -41380 80800
rect -41120 80780 -40880 80800
rect -40620 80780 -40380 80800
rect -40120 80780 -39880 80800
rect -39620 80780 -39380 80800
rect -39120 80780 -38880 80800
rect -38620 80780 -38380 80800
rect -38120 80780 -37880 80800
rect -37620 80780 -37380 80800
rect -37120 80780 -36880 80800
rect -36620 80780 -36380 80800
rect -36120 80780 -35880 80800
rect -35620 80780 -35380 80800
rect -35120 80780 -34880 80800
rect -34620 80780 -34380 80800
rect -34120 80780 -33880 80800
rect -33620 80780 -33380 80800
rect -33120 80780 -32880 80800
rect -32620 80780 -32380 80800
rect -32120 80780 -31880 80800
rect -31620 80780 -31380 80800
rect -31120 80780 -30880 80800
rect -30620 80780 -30380 80800
rect -30120 80780 -29880 80800
rect -29620 80780 -29380 80800
rect -29120 80780 -28880 80800
rect -28620 80780 -28380 80800
rect -28120 80780 -27880 80800
rect -27620 80780 -27380 80800
rect -27120 80780 -26880 80800
rect -26620 80780 -26380 80800
rect -26120 80780 -25880 80800
rect -25620 80780 -25380 80800
rect -25120 80780 -24880 80800
rect -24620 80780 -24380 80800
rect -24120 80780 -23880 80800
rect -23620 80780 -23380 80800
rect -23120 80780 -22880 80800
rect -22620 80780 -22380 80800
rect -22120 80780 -21880 80800
rect -21620 80780 -21380 80800
rect -21120 80780 -20880 80800
rect -20620 80780 -20380 80800
rect -20120 80780 -19880 80800
rect -19620 80780 -19380 80800
rect -19120 80780 -18880 80800
rect -18620 80780 -18380 80800
rect -18120 80780 -17880 80800
rect -17620 80780 -17380 80800
rect -17120 80780 -16880 80800
rect -16620 80780 -16380 80800
rect -16120 80780 -15880 80800
rect -15620 80780 -15380 80800
rect -15120 80780 -14880 80800
rect -14620 80780 -14380 80800
rect -14120 80780 -13880 80800
rect -13620 80780 -13380 80800
rect -13120 80780 -12880 80800
rect -12620 80780 -12380 80800
rect -12120 80780 -11880 80800
rect -11620 80780 -11380 80800
rect -11120 80780 -10880 80800
rect -10620 80780 -10380 80800
rect -10120 80780 -9880 80800
rect -9620 80780 -9380 80800
rect -9120 80780 -8880 80800
rect -8620 80780 -8380 80800
rect -8120 80780 -7880 80800
rect -7620 80780 -7380 80800
rect -7120 80780 -6880 80800
rect -6620 80780 -6380 80800
rect -6120 80780 -5880 80800
rect -5620 80780 -5380 80800
rect -5120 80780 -4880 80800
rect -4620 80780 -4380 80800
rect -4120 80780 -3880 80800
rect -3620 80780 -3380 80800
rect -3120 80780 -2880 80800
rect -2620 80780 -2380 80800
rect -2120 80780 -1880 80800
rect -1620 80780 -1380 80800
rect -1120 80780 -880 80800
rect -620 80780 -380 80800
rect -120 80780 120 80800
rect 380 80780 620 80800
rect 880 80780 1120 80800
rect 1380 80780 1620 80800
rect 1880 80780 2120 80800
rect 2380 80780 2620 80800
rect 2880 80780 3120 80800
rect 3380 80780 3620 80800
rect 3880 80780 4120 80800
rect 4380 80780 4620 80800
rect 4880 80780 5120 80800
rect 5380 80780 5620 80800
rect 5880 80780 6120 80800
rect 6380 80780 6620 80800
rect 6880 80780 7120 80800
rect 7380 80780 7620 80800
rect 7880 80780 8120 80800
rect 8380 80780 8620 80800
rect 8880 80780 9120 80800
rect 9380 80780 9620 80800
rect 9880 80780 10120 80800
rect 10380 80780 10620 80800
rect 10880 80780 11120 80800
rect 11380 80780 11620 80800
rect 11880 80780 12120 80800
rect 12380 80780 12620 80800
rect 12880 80780 13120 80800
rect 13380 80780 13620 80800
rect 13880 80780 14120 80800
rect 14380 80780 14620 80800
rect 14880 80780 15120 80800
rect 15380 80780 15620 80800
rect 15880 80780 16120 80800
rect 16380 80780 16620 80800
rect 16880 80780 17120 80800
rect 17380 80780 17620 80800
rect 17880 80780 18120 80800
rect 18380 80780 18620 80800
rect 18880 80780 19120 80800
rect 19380 80780 19620 80800
rect 19880 80780 20120 80800
rect 20380 80780 20620 80800
rect 20880 80780 21120 80800
rect 21380 80780 21620 80800
rect 21880 80780 22120 80800
rect 22380 80780 22620 80800
rect 22880 80780 23120 80800
rect 23380 80780 23620 80800
rect 23880 80780 24120 80800
rect 24380 80780 24620 80800
rect 24880 80780 25120 80800
rect 25380 80780 25620 80800
rect 25880 80780 26120 80800
rect 26380 80780 26620 80800
rect 26880 80780 27120 80800
rect 27380 80780 27620 80800
rect 27880 80780 28120 80800
rect 28380 80780 28620 80800
rect 28880 80780 29120 80800
rect 29380 80780 29620 80800
rect 29880 80780 30120 80800
rect 30380 80780 30620 80800
rect 30880 80780 31120 80800
rect 31380 80780 31620 80800
rect 31880 80780 32120 80800
rect 32380 80780 32620 80800
rect 32880 80780 33120 80800
rect 33380 80780 33620 80800
rect 33880 80780 34120 80800
rect 34380 80780 34620 80800
rect 34880 80780 35120 80800
rect 35380 80780 35620 80800
rect 35880 80780 36120 80800
rect 36380 80780 36620 80800
rect 36880 80780 37120 80800
rect 37380 80780 37620 80800
rect 37880 80780 38120 80800
rect 38380 80780 38620 80800
rect 38880 80780 39120 80800
rect 39380 80780 39620 80800
rect 39880 80780 40120 80800
rect 40380 80780 40620 80800
rect 40880 80780 41120 80800
rect 41380 80780 41620 80800
rect 41880 80780 42120 80800
rect 42380 80780 42620 80800
rect 42880 80780 43120 80800
rect 43380 80780 43620 80800
rect 43880 80780 44120 80800
rect 44380 80780 44620 80800
rect 44880 80780 45120 80800
rect 45380 80780 45620 80800
rect 45880 80780 46120 80800
rect 46380 80780 46620 80800
rect 46880 80780 47120 80800
rect 47380 80780 47620 80800
rect 47880 80780 48120 80800
rect 48380 80780 48620 80800
rect 48880 80780 49120 80800
rect 49380 80780 49620 80800
rect 49880 80780 50120 80800
rect 50380 80780 50620 80800
rect 50880 80780 51120 80800
rect 51380 80780 51620 80800
rect 51880 80780 52120 80800
rect 52380 80780 52620 80800
rect 52880 80780 53120 80800
rect 53380 80780 53620 80800
rect 53880 80780 54120 80800
rect 54380 80780 54620 80800
rect 54880 80780 55120 80800
rect 55380 80780 55620 80800
rect 55880 80780 56120 80800
rect 56380 80780 56620 80800
rect 56880 80780 57120 80800
rect 57380 80780 57620 80800
rect 57880 80780 58120 80800
rect 58380 80780 58620 80800
rect 58880 80780 59120 80800
rect 59380 80780 59620 80800
rect 59880 80780 60120 80800
rect 60380 80780 60620 80800
rect 60880 80780 61120 80800
rect 61380 80780 61620 80800
rect 61880 80780 62120 80800
rect 62380 80780 62620 80800
rect 62880 80780 63120 80800
rect 63380 80780 63620 80800
rect 63880 80780 64120 80800
rect 64380 80780 64620 80800
rect 64880 80780 65120 80800
rect 65380 80780 65620 80800
rect 65880 80780 66120 80800
rect 66380 80780 66620 80800
rect 66880 80780 67120 80800
rect 67380 80780 67620 80800
rect 67880 80780 68120 80800
rect 68380 80780 68620 80800
rect 68880 80780 69120 80800
rect 69380 80780 69620 80800
rect 69880 80780 70120 80800
rect 70380 80780 70620 80800
rect 70880 80780 71120 80800
rect 71380 80780 71620 80800
rect 71880 80780 72120 80800
rect 72380 80780 72620 80800
rect 72880 80780 73120 80800
rect 73380 80780 73620 80800
rect 73880 80780 74120 80800
rect 74380 80780 74620 80800
rect 74880 80780 75120 80800
rect 75380 80780 75620 80800
rect 75880 80780 76120 80800
rect 76380 80780 76620 80800
rect 76880 80780 77120 80800
rect 77380 80780 77620 80800
rect 77880 80780 78120 80800
rect 78380 80780 78620 80800
rect 78880 80780 79120 80800
rect 79380 80780 79620 80800
rect 79880 80780 80120 80800
rect 80380 80780 80620 80800
rect 80880 80780 81120 80800
rect 81380 80780 81620 80800
rect 81880 80780 82120 80800
rect 82380 80780 82620 80800
rect 82880 80780 83120 80800
rect 83380 80780 83620 80800
rect 83880 80780 84120 80800
rect 84380 80780 84620 80800
rect 84880 80780 85120 80800
rect 85380 80780 85620 80800
rect 85880 80780 86120 80800
rect 86380 80780 86620 80800
rect 86880 80780 87120 80800
rect 87380 80780 87620 80800
rect 87880 80780 88120 80800
rect 88380 80780 88620 80800
rect 88880 80780 89120 80800
rect 89380 80780 89620 80800
rect 89880 80780 90120 80800
rect 90380 80780 90620 80800
rect 90880 80780 91120 80800
rect 91380 80780 91620 80800
rect 91880 80780 92120 80800
rect 92380 80780 92620 80800
rect 92880 80780 93120 80800
rect 93380 80780 93620 80800
rect 93880 80780 94120 80800
rect 94380 80780 94620 80800
rect 94880 80780 95120 80800
rect 95380 80780 95620 80800
rect 95880 80780 96120 80800
rect 96380 80780 96620 80800
rect 96880 80780 97120 80800
rect 97380 80780 97620 80800
rect 97880 80780 98120 80800
rect 98380 80780 98620 80800
rect 98880 80780 99120 80800
rect 99380 80780 99620 80800
rect 99880 80780 100120 80800
rect 100380 80780 100500 80800
rect -83500 80750 -83400 80780
rect -83500 80550 -83480 80750
rect -83410 80550 -83400 80750
rect -83500 80520 -83400 80550
rect -83100 80750 -82900 80780
rect -83100 80550 -83090 80750
rect -83020 80550 -82980 80750
rect -82910 80550 -82900 80750
rect -83100 80520 -82900 80550
rect -82600 80750 -82400 80780
rect -82600 80550 -82590 80750
rect -82520 80550 -82480 80750
rect -82410 80550 -82400 80750
rect -82600 80520 -82400 80550
rect -82100 80750 -81900 80780
rect -82100 80550 -82090 80750
rect -82020 80550 -81980 80750
rect -81910 80550 -81900 80750
rect -82100 80520 -81900 80550
rect -81600 80750 -81400 80780
rect -81600 80550 -81590 80750
rect -81520 80550 -81480 80750
rect -81410 80550 -81400 80750
rect -81600 80520 -81400 80550
rect -81100 80750 -80900 80780
rect -81100 80550 -81090 80750
rect -81020 80550 -80980 80750
rect -80910 80550 -80900 80750
rect -81100 80520 -80900 80550
rect -80600 80750 -80400 80780
rect -80600 80550 -80590 80750
rect -80520 80550 -80480 80750
rect -80410 80550 -80400 80750
rect -80600 80520 -80400 80550
rect -80100 80750 -79900 80780
rect -80100 80550 -80090 80750
rect -80020 80550 -79980 80750
rect -79910 80550 -79900 80750
rect -80100 80520 -79900 80550
rect -79600 80750 -79400 80780
rect -79600 80550 -79590 80750
rect -79520 80550 -79480 80750
rect -79410 80550 -79400 80750
rect -79600 80520 -79400 80550
rect -79100 80750 -78900 80780
rect -79100 80550 -79090 80750
rect -79020 80550 -78980 80750
rect -78910 80550 -78900 80750
rect -79100 80520 -78900 80550
rect -78600 80750 -78400 80780
rect -78600 80550 -78590 80750
rect -78520 80550 -78480 80750
rect -78410 80550 -78400 80750
rect -78600 80520 -78400 80550
rect -78100 80750 -77900 80780
rect -78100 80550 -78090 80750
rect -78020 80550 -77980 80750
rect -77910 80550 -77900 80750
rect -78100 80520 -77900 80550
rect -77600 80750 -77400 80780
rect -77600 80550 -77590 80750
rect -77520 80550 -77480 80750
rect -77410 80550 -77400 80750
rect -77600 80520 -77400 80550
rect -77100 80750 -76900 80780
rect -77100 80550 -77090 80750
rect -77020 80550 -76980 80750
rect -76910 80550 -76900 80750
rect -77100 80520 -76900 80550
rect -76600 80750 -76400 80780
rect -76600 80550 -76590 80750
rect -76520 80550 -76480 80750
rect -76410 80550 -76400 80750
rect -76600 80520 -76400 80550
rect -76100 80750 -75900 80780
rect -76100 80550 -76090 80750
rect -76020 80550 -75980 80750
rect -75910 80550 -75900 80750
rect -76100 80520 -75900 80550
rect -75600 80750 -75400 80780
rect -75600 80550 -75590 80750
rect -75520 80550 -75480 80750
rect -75410 80550 -75400 80750
rect -75600 80520 -75400 80550
rect -75100 80750 -74900 80780
rect -75100 80550 -75090 80750
rect -75020 80550 -74980 80750
rect -74910 80550 -74900 80750
rect -75100 80520 -74900 80550
rect -74600 80750 -74400 80780
rect -74600 80550 -74590 80750
rect -74520 80550 -74480 80750
rect -74410 80550 -74400 80750
rect -74600 80520 -74400 80550
rect -74100 80750 -73900 80780
rect -74100 80550 -74090 80750
rect -74020 80550 -73980 80750
rect -73910 80550 -73900 80750
rect -74100 80520 -73900 80550
rect -73600 80750 -73400 80780
rect -73600 80550 -73590 80750
rect -73520 80550 -73480 80750
rect -73410 80550 -73400 80750
rect -73600 80520 -73400 80550
rect -73100 80750 -72900 80780
rect -73100 80550 -73090 80750
rect -73020 80550 -72980 80750
rect -72910 80550 -72900 80750
rect -73100 80520 -72900 80550
rect -72600 80750 -72400 80780
rect -72600 80550 -72590 80750
rect -72520 80550 -72480 80750
rect -72410 80550 -72400 80750
rect -72600 80520 -72400 80550
rect -72100 80750 -71900 80780
rect -72100 80550 -72090 80750
rect -72020 80550 -71980 80750
rect -71910 80550 -71900 80750
rect -72100 80520 -71900 80550
rect -71600 80750 -71400 80780
rect -71600 80550 -71590 80750
rect -71520 80550 -71480 80750
rect -71410 80550 -71400 80750
rect -71600 80520 -71400 80550
rect -71100 80750 -70900 80780
rect -71100 80550 -71090 80750
rect -71020 80550 -70980 80750
rect -70910 80550 -70900 80750
rect -71100 80520 -70900 80550
rect -70600 80750 -70400 80780
rect -70600 80550 -70590 80750
rect -70520 80550 -70480 80750
rect -70410 80550 -70400 80750
rect -70600 80520 -70400 80550
rect -70100 80750 -69900 80780
rect -70100 80550 -70090 80750
rect -70020 80550 -69980 80750
rect -69910 80550 -69900 80750
rect -70100 80520 -69900 80550
rect -69600 80750 -69400 80780
rect -69600 80550 -69590 80750
rect -69520 80550 -69480 80750
rect -69410 80550 -69400 80750
rect -69600 80520 -69400 80550
rect -69100 80750 -68900 80780
rect -69100 80550 -69090 80750
rect -69020 80550 -68980 80750
rect -68910 80550 -68900 80750
rect -69100 80520 -68900 80550
rect -68600 80750 -68400 80780
rect -68600 80550 -68590 80750
rect -68520 80550 -68480 80750
rect -68410 80550 -68400 80750
rect -68600 80520 -68400 80550
rect -68100 80750 -67900 80780
rect -68100 80550 -68090 80750
rect -68020 80550 -67980 80750
rect -67910 80550 -67900 80750
rect -68100 80520 -67900 80550
rect -67600 80750 -67400 80780
rect -67600 80550 -67590 80750
rect -67520 80550 -67480 80750
rect -67410 80550 -67400 80750
rect -67600 80520 -67400 80550
rect -67100 80750 -66900 80780
rect -67100 80550 -67090 80750
rect -67020 80550 -66980 80750
rect -66910 80550 -66900 80750
rect -67100 80520 -66900 80550
rect -66600 80750 -66400 80780
rect -66600 80550 -66590 80750
rect -66520 80550 -66480 80750
rect -66410 80550 -66400 80750
rect -66600 80520 -66400 80550
rect -66100 80750 -65900 80780
rect -66100 80550 -66090 80750
rect -66020 80550 -65980 80750
rect -65910 80550 -65900 80750
rect -66100 80520 -65900 80550
rect -65600 80750 -65400 80780
rect -65600 80550 -65590 80750
rect -65520 80550 -65480 80750
rect -65410 80550 -65400 80750
rect -65600 80520 -65400 80550
rect -65100 80750 -64900 80780
rect -65100 80550 -65090 80750
rect -65020 80550 -64980 80750
rect -64910 80550 -64900 80750
rect -65100 80520 -64900 80550
rect -64600 80750 -64400 80780
rect -64600 80550 -64590 80750
rect -64520 80550 -64480 80750
rect -64410 80550 -64400 80750
rect -64600 80520 -64400 80550
rect -64100 80750 -63900 80780
rect -64100 80550 -64090 80750
rect -64020 80550 -63980 80750
rect -63910 80550 -63900 80750
rect -64100 80520 -63900 80550
rect -63600 80750 -63400 80780
rect -63600 80550 -63590 80750
rect -63520 80550 -63480 80750
rect -63410 80550 -63400 80750
rect -63600 80520 -63400 80550
rect -63100 80750 -62900 80780
rect -63100 80550 -63090 80750
rect -63020 80550 -62980 80750
rect -62910 80550 -62900 80750
rect -63100 80520 -62900 80550
rect -62600 80750 -62400 80780
rect -62600 80550 -62590 80750
rect -62520 80550 -62480 80750
rect -62410 80550 -62400 80750
rect -62600 80520 -62400 80550
rect -62100 80750 -61900 80780
rect -62100 80550 -62090 80750
rect -62020 80550 -61980 80750
rect -61910 80550 -61900 80750
rect -62100 80520 -61900 80550
rect -61600 80750 -61400 80780
rect -61600 80550 -61590 80750
rect -61520 80550 -61480 80750
rect -61410 80550 -61400 80750
rect -61600 80520 -61400 80550
rect -61100 80750 -60900 80780
rect -61100 80550 -61090 80750
rect -61020 80550 -60980 80750
rect -60910 80550 -60900 80750
rect -61100 80520 -60900 80550
rect -60600 80750 -60400 80780
rect -60600 80550 -60590 80750
rect -60520 80550 -60480 80750
rect -60410 80550 -60400 80750
rect -60600 80520 -60400 80550
rect -60100 80750 -59900 80780
rect -60100 80550 -60090 80750
rect -60020 80550 -59980 80750
rect -59910 80550 -59900 80750
rect -60100 80520 -59900 80550
rect -59600 80750 -59400 80780
rect -59600 80550 -59590 80750
rect -59520 80550 -59480 80750
rect -59410 80550 -59400 80750
rect -59600 80520 -59400 80550
rect -59100 80750 -58900 80780
rect -59100 80550 -59090 80750
rect -59020 80550 -58980 80750
rect -58910 80550 -58900 80750
rect -59100 80520 -58900 80550
rect -58600 80750 -58400 80780
rect -58600 80550 -58590 80750
rect -58520 80550 -58480 80750
rect -58410 80550 -58400 80750
rect -58600 80520 -58400 80550
rect -58100 80750 -57900 80780
rect -58100 80550 -58090 80750
rect -58020 80550 -57980 80750
rect -57910 80550 -57900 80750
rect -58100 80520 -57900 80550
rect -57600 80750 -57400 80780
rect -57600 80550 -57590 80750
rect -57520 80550 -57480 80750
rect -57410 80550 -57400 80750
rect -57600 80520 -57400 80550
rect -57100 80750 -56900 80780
rect -57100 80550 -57090 80750
rect -57020 80550 -56980 80750
rect -56910 80550 -56900 80750
rect -57100 80520 -56900 80550
rect -56600 80750 -56400 80780
rect -56600 80550 -56590 80750
rect -56520 80550 -56480 80750
rect -56410 80550 -56400 80750
rect -56600 80520 -56400 80550
rect -56100 80750 -55900 80780
rect -56100 80550 -56090 80750
rect -56020 80550 -55980 80750
rect -55910 80550 -55900 80750
rect -56100 80520 -55900 80550
rect -55600 80750 -55400 80780
rect -55600 80550 -55590 80750
rect -55520 80550 -55480 80750
rect -55410 80550 -55400 80750
rect -55600 80520 -55400 80550
rect -55100 80750 -54900 80780
rect -55100 80550 -55090 80750
rect -55020 80550 -54980 80750
rect -54910 80550 -54900 80750
rect -55100 80520 -54900 80550
rect -54600 80750 -54400 80780
rect -54600 80550 -54590 80750
rect -54520 80550 -54480 80750
rect -54410 80550 -54400 80750
rect -54600 80520 -54400 80550
rect -54100 80750 -53900 80780
rect -54100 80550 -54090 80750
rect -54020 80550 -53980 80750
rect -53910 80550 -53900 80750
rect -54100 80520 -53900 80550
rect -53600 80750 -53400 80780
rect -53600 80550 -53590 80750
rect -53520 80550 -53480 80750
rect -53410 80550 -53400 80750
rect -53600 80520 -53400 80550
rect -53100 80750 -52900 80780
rect -53100 80550 -53090 80750
rect -53020 80550 -52980 80750
rect -52910 80550 -52900 80750
rect -53100 80520 -52900 80550
rect -52600 80750 -52400 80780
rect -52600 80550 -52590 80750
rect -52520 80550 -52480 80750
rect -52410 80550 -52400 80750
rect -52600 80520 -52400 80550
rect -52100 80750 -51900 80780
rect -52100 80550 -52090 80750
rect -52020 80550 -51980 80750
rect -51910 80550 -51900 80750
rect -52100 80520 -51900 80550
rect -51600 80750 -51400 80780
rect -51600 80550 -51590 80750
rect -51520 80550 -51480 80750
rect -51410 80550 -51400 80750
rect -51600 80520 -51400 80550
rect -51100 80750 -50900 80780
rect -51100 80550 -51090 80750
rect -51020 80550 -50980 80750
rect -50910 80550 -50900 80750
rect -51100 80520 -50900 80550
rect -50600 80750 -50400 80780
rect -50600 80550 -50590 80750
rect -50520 80550 -50480 80750
rect -50410 80550 -50400 80750
rect -50600 80520 -50400 80550
rect -50100 80750 -49900 80780
rect -50100 80550 -50090 80750
rect -50020 80550 -49980 80750
rect -49910 80550 -49900 80750
rect -50100 80520 -49900 80550
rect -49600 80750 -49400 80780
rect -49600 80550 -49590 80750
rect -49520 80550 -49480 80750
rect -49410 80550 -49400 80750
rect -49600 80520 -49400 80550
rect -49100 80750 -48900 80780
rect -49100 80550 -49090 80750
rect -49020 80550 -48980 80750
rect -48910 80550 -48900 80750
rect -49100 80520 -48900 80550
rect -48600 80750 -48400 80780
rect -48600 80550 -48590 80750
rect -48520 80550 -48480 80750
rect -48410 80550 -48400 80750
rect -48600 80520 -48400 80550
rect -48100 80750 -47900 80780
rect -48100 80550 -48090 80750
rect -48020 80550 -47980 80750
rect -47910 80550 -47900 80750
rect -48100 80520 -47900 80550
rect -47600 80750 -47400 80780
rect -47600 80550 -47590 80750
rect -47520 80550 -47480 80750
rect -47410 80550 -47400 80750
rect -47600 80520 -47400 80550
rect -47100 80750 -46900 80780
rect -47100 80550 -47090 80750
rect -47020 80550 -46980 80750
rect -46910 80550 -46900 80750
rect -47100 80520 -46900 80550
rect -46600 80750 -46400 80780
rect -46600 80550 -46590 80750
rect -46520 80550 -46480 80750
rect -46410 80550 -46400 80750
rect -46600 80520 -46400 80550
rect -46100 80750 -45900 80780
rect -46100 80550 -46090 80750
rect -46020 80550 -45980 80750
rect -45910 80550 -45900 80750
rect -46100 80520 -45900 80550
rect -45600 80750 -45400 80780
rect -45600 80550 -45590 80750
rect -45520 80550 -45480 80750
rect -45410 80550 -45400 80750
rect -45600 80520 -45400 80550
rect -45100 80750 -44900 80780
rect -45100 80550 -45090 80750
rect -45020 80550 -44980 80750
rect -44910 80550 -44900 80750
rect -45100 80520 -44900 80550
rect -44600 80750 -44400 80780
rect -44600 80550 -44590 80750
rect -44520 80550 -44480 80750
rect -44410 80550 -44400 80750
rect -44600 80520 -44400 80550
rect -44100 80750 -43900 80780
rect -44100 80550 -44090 80750
rect -44020 80550 -43980 80750
rect -43910 80550 -43900 80750
rect -44100 80520 -43900 80550
rect -43600 80750 -43400 80780
rect -43600 80550 -43590 80750
rect -43520 80550 -43480 80750
rect -43410 80550 -43400 80750
rect -43600 80520 -43400 80550
rect -43100 80750 -42900 80780
rect -43100 80550 -43090 80750
rect -43020 80550 -42980 80750
rect -42910 80550 -42900 80750
rect -43100 80520 -42900 80550
rect -42600 80750 -42400 80780
rect -42600 80550 -42590 80750
rect -42520 80550 -42480 80750
rect -42410 80550 -42400 80750
rect -42600 80520 -42400 80550
rect -42100 80750 -41900 80780
rect -42100 80550 -42090 80750
rect -42020 80550 -41980 80750
rect -41910 80550 -41900 80750
rect -42100 80520 -41900 80550
rect -41600 80750 -41400 80780
rect -41600 80550 -41590 80750
rect -41520 80550 -41480 80750
rect -41410 80550 -41400 80750
rect -41600 80520 -41400 80550
rect -41100 80750 -40900 80780
rect -41100 80550 -41090 80750
rect -41020 80550 -40980 80750
rect -40910 80550 -40900 80750
rect -41100 80520 -40900 80550
rect -40600 80750 -40400 80780
rect -40600 80550 -40590 80750
rect -40520 80550 -40480 80750
rect -40410 80550 -40400 80750
rect -40600 80520 -40400 80550
rect -40100 80750 -39900 80780
rect -40100 80550 -40090 80750
rect -40020 80550 -39980 80750
rect -39910 80550 -39900 80750
rect -40100 80520 -39900 80550
rect -39600 80750 -39400 80780
rect -39600 80550 -39590 80750
rect -39520 80550 -39480 80750
rect -39410 80550 -39400 80750
rect -39600 80520 -39400 80550
rect -39100 80750 -38900 80780
rect -39100 80550 -39090 80750
rect -39020 80550 -38980 80750
rect -38910 80550 -38900 80750
rect -39100 80520 -38900 80550
rect -38600 80750 -38400 80780
rect -38600 80550 -38590 80750
rect -38520 80550 -38480 80750
rect -38410 80550 -38400 80750
rect -38600 80520 -38400 80550
rect -38100 80750 -37900 80780
rect -38100 80550 -38090 80750
rect -38020 80550 -37980 80750
rect -37910 80550 -37900 80750
rect -38100 80520 -37900 80550
rect -37600 80750 -37400 80780
rect -37600 80550 -37590 80750
rect -37520 80550 -37480 80750
rect -37410 80550 -37400 80750
rect -37600 80520 -37400 80550
rect -37100 80750 -36900 80780
rect -37100 80550 -37090 80750
rect -37020 80550 -36980 80750
rect -36910 80550 -36900 80750
rect -37100 80520 -36900 80550
rect -36600 80750 -36400 80780
rect -36600 80550 -36590 80750
rect -36520 80550 -36480 80750
rect -36410 80550 -36400 80750
rect -36600 80520 -36400 80550
rect -36100 80750 -35900 80780
rect -36100 80550 -36090 80750
rect -36020 80550 -35980 80750
rect -35910 80550 -35900 80750
rect -36100 80520 -35900 80550
rect -35600 80750 -35400 80780
rect -35600 80550 -35590 80750
rect -35520 80550 -35480 80750
rect -35410 80550 -35400 80750
rect -35600 80520 -35400 80550
rect -35100 80750 -34900 80780
rect -35100 80550 -35090 80750
rect -35020 80550 -34980 80750
rect -34910 80550 -34900 80750
rect -35100 80520 -34900 80550
rect -34600 80750 -34400 80780
rect -34600 80550 -34590 80750
rect -34520 80550 -34480 80750
rect -34410 80550 -34400 80750
rect -34600 80520 -34400 80550
rect -34100 80750 -33900 80780
rect -34100 80550 -34090 80750
rect -34020 80550 -33980 80750
rect -33910 80550 -33900 80750
rect -34100 80520 -33900 80550
rect -33600 80750 -33400 80780
rect -33600 80550 -33590 80750
rect -33520 80550 -33480 80750
rect -33410 80550 -33400 80750
rect -33600 80520 -33400 80550
rect -33100 80750 -32900 80780
rect -33100 80550 -33090 80750
rect -33020 80550 -32980 80750
rect -32910 80550 -32900 80750
rect -33100 80520 -32900 80550
rect -32600 80750 -32400 80780
rect -32600 80550 -32590 80750
rect -32520 80550 -32480 80750
rect -32410 80550 -32400 80750
rect -32600 80520 -32400 80550
rect -32100 80750 -31900 80780
rect -32100 80550 -32090 80750
rect -32020 80550 -31980 80750
rect -31910 80550 -31900 80750
rect -32100 80520 -31900 80550
rect -31600 80750 -31400 80780
rect -31600 80550 -31590 80750
rect -31520 80550 -31480 80750
rect -31410 80550 -31400 80750
rect -31600 80520 -31400 80550
rect -31100 80750 -30900 80780
rect -31100 80550 -31090 80750
rect -31020 80550 -30980 80750
rect -30910 80550 -30900 80750
rect -31100 80520 -30900 80550
rect -30600 80750 -30400 80780
rect -30600 80550 -30590 80750
rect -30520 80550 -30480 80750
rect -30410 80550 -30400 80750
rect -30600 80520 -30400 80550
rect -30100 80750 -29900 80780
rect -30100 80550 -30090 80750
rect -30020 80550 -29980 80750
rect -29910 80550 -29900 80750
rect -30100 80520 -29900 80550
rect -29600 80750 -29400 80780
rect -29600 80550 -29590 80750
rect -29520 80550 -29480 80750
rect -29410 80550 -29400 80750
rect -29600 80520 -29400 80550
rect -29100 80750 -28900 80780
rect -29100 80550 -29090 80750
rect -29020 80550 -28980 80750
rect -28910 80550 -28900 80750
rect -29100 80520 -28900 80550
rect -28600 80750 -28400 80780
rect -28600 80550 -28590 80750
rect -28520 80550 -28480 80750
rect -28410 80550 -28400 80750
rect -28600 80520 -28400 80550
rect -28100 80750 -27900 80780
rect -28100 80550 -28090 80750
rect -28020 80550 -27980 80750
rect -27910 80550 -27900 80750
rect -28100 80520 -27900 80550
rect -27600 80750 -27400 80780
rect -27600 80550 -27590 80750
rect -27520 80550 -27480 80750
rect -27410 80550 -27400 80750
rect -27600 80520 -27400 80550
rect -27100 80750 -26900 80780
rect -27100 80550 -27090 80750
rect -27020 80550 -26980 80750
rect -26910 80550 -26900 80750
rect -27100 80520 -26900 80550
rect -26600 80750 -26400 80780
rect -26600 80550 -26590 80750
rect -26520 80550 -26480 80750
rect -26410 80550 -26400 80750
rect -26600 80520 -26400 80550
rect -26100 80750 -25900 80780
rect -26100 80550 -26090 80750
rect -26020 80550 -25980 80750
rect -25910 80550 -25900 80750
rect -26100 80520 -25900 80550
rect -25600 80750 -25400 80780
rect -25600 80550 -25590 80750
rect -25520 80550 -25480 80750
rect -25410 80550 -25400 80750
rect -25600 80520 -25400 80550
rect -25100 80750 -24900 80780
rect -25100 80550 -25090 80750
rect -25020 80550 -24980 80750
rect -24910 80550 -24900 80750
rect -25100 80520 -24900 80550
rect -24600 80750 -24400 80780
rect -24600 80550 -24590 80750
rect -24520 80550 -24480 80750
rect -24410 80550 -24400 80750
rect -24600 80520 -24400 80550
rect -24100 80750 -23900 80780
rect -24100 80550 -24090 80750
rect -24020 80550 -23980 80750
rect -23910 80550 -23900 80750
rect -24100 80520 -23900 80550
rect -23600 80750 -23400 80780
rect -23600 80550 -23590 80750
rect -23520 80550 -23480 80750
rect -23410 80550 -23400 80750
rect -23600 80520 -23400 80550
rect -23100 80750 -22900 80780
rect -23100 80550 -23090 80750
rect -23020 80550 -22980 80750
rect -22910 80550 -22900 80750
rect -23100 80520 -22900 80550
rect -22600 80750 -22400 80780
rect -22600 80550 -22590 80750
rect -22520 80550 -22480 80750
rect -22410 80550 -22400 80750
rect -22600 80520 -22400 80550
rect -22100 80750 -21900 80780
rect -22100 80550 -22090 80750
rect -22020 80550 -21980 80750
rect -21910 80550 -21900 80750
rect -22100 80520 -21900 80550
rect -21600 80750 -21400 80780
rect -21600 80550 -21590 80750
rect -21520 80550 -21480 80750
rect -21410 80550 -21400 80750
rect -21600 80520 -21400 80550
rect -21100 80750 -20900 80780
rect -21100 80550 -21090 80750
rect -21020 80550 -20980 80750
rect -20910 80550 -20900 80750
rect -21100 80520 -20900 80550
rect -20600 80750 -20400 80780
rect -20600 80550 -20590 80750
rect -20520 80550 -20480 80750
rect -20410 80550 -20400 80750
rect -20600 80520 -20400 80550
rect -20100 80750 -19900 80780
rect -20100 80550 -20090 80750
rect -20020 80550 -19980 80750
rect -19910 80550 -19900 80750
rect -20100 80520 -19900 80550
rect -19600 80750 -19400 80780
rect -19600 80550 -19590 80750
rect -19520 80550 -19480 80750
rect -19410 80550 -19400 80750
rect -19600 80520 -19400 80550
rect -19100 80750 -18900 80780
rect -19100 80550 -19090 80750
rect -19020 80550 -18980 80750
rect -18910 80550 -18900 80750
rect -19100 80520 -18900 80550
rect -18600 80750 -18400 80780
rect -18600 80550 -18590 80750
rect -18520 80550 -18480 80750
rect -18410 80550 -18400 80750
rect -18600 80520 -18400 80550
rect -18100 80750 -17900 80780
rect -18100 80550 -18090 80750
rect -18020 80550 -17980 80750
rect -17910 80550 -17900 80750
rect -18100 80520 -17900 80550
rect -17600 80750 -17400 80780
rect -17600 80550 -17590 80750
rect -17520 80550 -17480 80750
rect -17410 80550 -17400 80750
rect -17600 80520 -17400 80550
rect -17100 80750 -16900 80780
rect -17100 80550 -17090 80750
rect -17020 80550 -16980 80750
rect -16910 80550 -16900 80750
rect -17100 80520 -16900 80550
rect -16600 80750 -16400 80780
rect -16600 80550 -16590 80750
rect -16520 80550 -16480 80750
rect -16410 80550 -16400 80750
rect -16600 80520 -16400 80550
rect -16100 80750 -15900 80780
rect -16100 80550 -16090 80750
rect -16020 80550 -15980 80750
rect -15910 80550 -15900 80750
rect -16100 80520 -15900 80550
rect -15600 80750 -15400 80780
rect -15600 80550 -15590 80750
rect -15520 80550 -15480 80750
rect -15410 80550 -15400 80750
rect -15600 80520 -15400 80550
rect -15100 80750 -14900 80780
rect -15100 80550 -15090 80750
rect -15020 80550 -14980 80750
rect -14910 80550 -14900 80750
rect -15100 80520 -14900 80550
rect -14600 80750 -14400 80780
rect -14600 80550 -14590 80750
rect -14520 80550 -14480 80750
rect -14410 80550 -14400 80750
rect -14600 80520 -14400 80550
rect -14100 80750 -13900 80780
rect -14100 80550 -14090 80750
rect -14020 80550 -13980 80750
rect -13910 80550 -13900 80750
rect -14100 80520 -13900 80550
rect -13600 80750 -13400 80780
rect -13600 80550 -13590 80750
rect -13520 80550 -13480 80750
rect -13410 80550 -13400 80750
rect -13600 80520 -13400 80550
rect -13100 80750 -12900 80780
rect -13100 80550 -13090 80750
rect -13020 80550 -12980 80750
rect -12910 80550 -12900 80750
rect -13100 80520 -12900 80550
rect -12600 80750 -12400 80780
rect -12600 80550 -12590 80750
rect -12520 80550 -12480 80750
rect -12410 80550 -12400 80750
rect -12600 80520 -12400 80550
rect -12100 80750 -11900 80780
rect -12100 80550 -12090 80750
rect -12020 80550 -11980 80750
rect -11910 80550 -11900 80750
rect -12100 80520 -11900 80550
rect -11600 80750 -11400 80780
rect -11600 80550 -11590 80750
rect -11520 80550 -11480 80750
rect -11410 80550 -11400 80750
rect -11600 80520 -11400 80550
rect -11100 80750 -10900 80780
rect -11100 80550 -11090 80750
rect -11020 80550 -10980 80750
rect -10910 80550 -10900 80750
rect -11100 80520 -10900 80550
rect -10600 80750 -10400 80780
rect -10600 80550 -10590 80750
rect -10520 80550 -10480 80750
rect -10410 80550 -10400 80750
rect -10600 80520 -10400 80550
rect -10100 80750 -9900 80780
rect -10100 80550 -10090 80750
rect -10020 80550 -9980 80750
rect -9910 80550 -9900 80750
rect -10100 80520 -9900 80550
rect -9600 80750 -9400 80780
rect -9600 80550 -9590 80750
rect -9520 80550 -9480 80750
rect -9410 80550 -9400 80750
rect -9600 80520 -9400 80550
rect -9100 80750 -8900 80780
rect -9100 80550 -9090 80750
rect -9020 80550 -8980 80750
rect -8910 80550 -8900 80750
rect -9100 80520 -8900 80550
rect -8600 80750 -8400 80780
rect -8600 80550 -8590 80750
rect -8520 80550 -8480 80750
rect -8410 80550 -8400 80750
rect -8600 80520 -8400 80550
rect -8100 80750 -7900 80780
rect -8100 80550 -8090 80750
rect -8020 80550 -7980 80750
rect -7910 80550 -7900 80750
rect -8100 80520 -7900 80550
rect -7600 80750 -7400 80780
rect -7600 80550 -7590 80750
rect -7520 80550 -7480 80750
rect -7410 80550 -7400 80750
rect -7600 80520 -7400 80550
rect -7100 80750 -6900 80780
rect -7100 80550 -7090 80750
rect -7020 80550 -6980 80750
rect -6910 80550 -6900 80750
rect -7100 80520 -6900 80550
rect -6600 80750 -6400 80780
rect -6600 80550 -6590 80750
rect -6520 80550 -6480 80750
rect -6410 80550 -6400 80750
rect -6600 80520 -6400 80550
rect -6100 80750 -5900 80780
rect -6100 80550 -6090 80750
rect -6020 80550 -5980 80750
rect -5910 80550 -5900 80750
rect -6100 80520 -5900 80550
rect -5600 80750 -5400 80780
rect -5600 80550 -5590 80750
rect -5520 80550 -5480 80750
rect -5410 80550 -5400 80750
rect -5600 80520 -5400 80550
rect -5100 80750 -4900 80780
rect -5100 80550 -5090 80750
rect -5020 80550 -4980 80750
rect -4910 80550 -4900 80750
rect -5100 80520 -4900 80550
rect -4600 80750 -4400 80780
rect -4600 80550 -4590 80750
rect -4520 80550 -4480 80750
rect -4410 80550 -4400 80750
rect -4600 80520 -4400 80550
rect -4100 80750 -3900 80780
rect -4100 80550 -4090 80750
rect -4020 80550 -3980 80750
rect -3910 80550 -3900 80750
rect -4100 80520 -3900 80550
rect -3600 80750 -3400 80780
rect -3600 80550 -3590 80750
rect -3520 80550 -3480 80750
rect -3410 80550 -3400 80750
rect -3600 80520 -3400 80550
rect -3100 80750 -2900 80780
rect -3100 80550 -3090 80750
rect -3020 80550 -2980 80750
rect -2910 80550 -2900 80750
rect -3100 80520 -2900 80550
rect -2600 80750 -2400 80780
rect -2600 80550 -2590 80750
rect -2520 80550 -2480 80750
rect -2410 80550 -2400 80750
rect -2600 80520 -2400 80550
rect -2100 80750 -1900 80780
rect -2100 80550 -2090 80750
rect -2020 80550 -1980 80750
rect -1910 80550 -1900 80750
rect -2100 80520 -1900 80550
rect -1600 80750 -1400 80780
rect -1600 80550 -1590 80750
rect -1520 80550 -1480 80750
rect -1410 80550 -1400 80750
rect -1600 80520 -1400 80550
rect -1100 80750 -900 80780
rect -1100 80550 -1090 80750
rect -1020 80550 -980 80750
rect -910 80550 -900 80750
rect -1100 80520 -900 80550
rect -600 80750 -400 80780
rect -600 80550 -590 80750
rect -520 80550 -480 80750
rect -410 80550 -400 80750
rect -600 80520 -400 80550
rect -100 80750 100 80780
rect -100 80550 -90 80750
rect -20 80550 20 80750
rect 90 80550 100 80750
rect -100 80520 100 80550
rect 400 80750 600 80780
rect 400 80550 410 80750
rect 480 80550 520 80750
rect 590 80550 600 80750
rect 400 80520 600 80550
rect 900 80750 1100 80780
rect 900 80550 910 80750
rect 980 80550 1020 80750
rect 1090 80550 1100 80750
rect 900 80520 1100 80550
rect 1400 80750 1600 80780
rect 1400 80550 1410 80750
rect 1480 80550 1520 80750
rect 1590 80550 1600 80750
rect 1400 80520 1600 80550
rect 1900 80750 2100 80780
rect 1900 80550 1910 80750
rect 1980 80550 2020 80750
rect 2090 80550 2100 80750
rect 1900 80520 2100 80550
rect 2400 80750 2600 80780
rect 2400 80550 2410 80750
rect 2480 80550 2520 80750
rect 2590 80550 2600 80750
rect 2400 80520 2600 80550
rect 2900 80750 3100 80780
rect 2900 80550 2910 80750
rect 2980 80550 3020 80750
rect 3090 80550 3100 80750
rect 2900 80520 3100 80550
rect 3400 80750 3600 80780
rect 3400 80550 3410 80750
rect 3480 80550 3520 80750
rect 3590 80550 3600 80750
rect 3400 80520 3600 80550
rect 3900 80750 4100 80780
rect 3900 80550 3910 80750
rect 3980 80550 4020 80750
rect 4090 80550 4100 80750
rect 3900 80520 4100 80550
rect 4400 80750 4600 80780
rect 4400 80550 4410 80750
rect 4480 80550 4520 80750
rect 4590 80550 4600 80750
rect 4400 80520 4600 80550
rect 4900 80750 5100 80780
rect 4900 80550 4910 80750
rect 4980 80550 5020 80750
rect 5090 80550 5100 80750
rect 4900 80520 5100 80550
rect 5400 80750 5600 80780
rect 5400 80550 5410 80750
rect 5480 80550 5520 80750
rect 5590 80550 5600 80750
rect 5400 80520 5600 80550
rect 5900 80750 6100 80780
rect 5900 80550 5910 80750
rect 5980 80550 6020 80750
rect 6090 80550 6100 80750
rect 5900 80520 6100 80550
rect 6400 80750 6600 80780
rect 6400 80550 6410 80750
rect 6480 80550 6520 80750
rect 6590 80550 6600 80750
rect 6400 80520 6600 80550
rect 6900 80750 7100 80780
rect 6900 80550 6910 80750
rect 6980 80550 7020 80750
rect 7090 80550 7100 80750
rect 6900 80520 7100 80550
rect 7400 80750 7600 80780
rect 7400 80550 7410 80750
rect 7480 80550 7520 80750
rect 7590 80550 7600 80750
rect 7400 80520 7600 80550
rect 7900 80750 8100 80780
rect 7900 80550 7910 80750
rect 7980 80550 8020 80750
rect 8090 80550 8100 80750
rect 7900 80520 8100 80550
rect 8400 80750 8600 80780
rect 8400 80550 8410 80750
rect 8480 80550 8520 80750
rect 8590 80550 8600 80750
rect 8400 80520 8600 80550
rect 8900 80750 9100 80780
rect 8900 80550 8910 80750
rect 8980 80550 9020 80750
rect 9090 80550 9100 80750
rect 8900 80520 9100 80550
rect 9400 80750 9600 80780
rect 9400 80550 9410 80750
rect 9480 80550 9520 80750
rect 9590 80550 9600 80750
rect 9400 80520 9600 80550
rect 9900 80750 10100 80780
rect 9900 80550 9910 80750
rect 9980 80550 10020 80750
rect 10090 80550 10100 80750
rect 9900 80520 10100 80550
rect 10400 80750 10600 80780
rect 10400 80550 10410 80750
rect 10480 80550 10520 80750
rect 10590 80550 10600 80750
rect 10400 80520 10600 80550
rect 10900 80750 11100 80780
rect 10900 80550 10910 80750
rect 10980 80550 11020 80750
rect 11090 80550 11100 80750
rect 10900 80520 11100 80550
rect 11400 80750 11600 80780
rect 11400 80550 11410 80750
rect 11480 80550 11520 80750
rect 11590 80550 11600 80750
rect 11400 80520 11600 80550
rect 11900 80750 12100 80780
rect 11900 80550 11910 80750
rect 11980 80550 12020 80750
rect 12090 80550 12100 80750
rect 11900 80520 12100 80550
rect 12400 80750 12600 80780
rect 12400 80550 12410 80750
rect 12480 80550 12520 80750
rect 12590 80550 12600 80750
rect 12400 80520 12600 80550
rect 12900 80750 13100 80780
rect 12900 80550 12910 80750
rect 12980 80550 13020 80750
rect 13090 80550 13100 80750
rect 12900 80520 13100 80550
rect 13400 80750 13600 80780
rect 13400 80550 13410 80750
rect 13480 80550 13520 80750
rect 13590 80550 13600 80750
rect 13400 80520 13600 80550
rect 13900 80750 14100 80780
rect 13900 80550 13910 80750
rect 13980 80550 14020 80750
rect 14090 80550 14100 80750
rect 13900 80520 14100 80550
rect 14400 80750 14600 80780
rect 14400 80550 14410 80750
rect 14480 80550 14520 80750
rect 14590 80550 14600 80750
rect 14400 80520 14600 80550
rect 14900 80750 15100 80780
rect 14900 80550 14910 80750
rect 14980 80550 15020 80750
rect 15090 80550 15100 80750
rect 14900 80520 15100 80550
rect 15400 80750 15600 80780
rect 15400 80550 15410 80750
rect 15480 80550 15520 80750
rect 15590 80550 15600 80750
rect 15400 80520 15600 80550
rect 15900 80750 16100 80780
rect 15900 80550 15910 80750
rect 15980 80550 16020 80750
rect 16090 80550 16100 80750
rect 15900 80520 16100 80550
rect 16400 80750 16600 80780
rect 16400 80550 16410 80750
rect 16480 80550 16520 80750
rect 16590 80550 16600 80750
rect 16400 80520 16600 80550
rect 16900 80750 17100 80780
rect 16900 80550 16910 80750
rect 16980 80550 17020 80750
rect 17090 80550 17100 80750
rect 16900 80520 17100 80550
rect 17400 80750 17600 80780
rect 17400 80550 17410 80750
rect 17480 80550 17520 80750
rect 17590 80550 17600 80750
rect 17400 80520 17600 80550
rect 17900 80750 18100 80780
rect 17900 80550 17910 80750
rect 17980 80550 18020 80750
rect 18090 80550 18100 80750
rect 17900 80520 18100 80550
rect 18400 80750 18600 80780
rect 18400 80550 18410 80750
rect 18480 80550 18520 80750
rect 18590 80550 18600 80750
rect 18400 80520 18600 80550
rect 18900 80750 19100 80780
rect 18900 80550 18910 80750
rect 18980 80550 19020 80750
rect 19090 80550 19100 80750
rect 18900 80520 19100 80550
rect 19400 80750 19600 80780
rect 19400 80550 19410 80750
rect 19480 80550 19520 80750
rect 19590 80550 19600 80750
rect 19400 80520 19600 80550
rect 19900 80750 20100 80780
rect 19900 80550 19910 80750
rect 19980 80550 20020 80750
rect 20090 80550 20100 80750
rect 19900 80520 20100 80550
rect 20400 80750 20600 80780
rect 20400 80550 20410 80750
rect 20480 80550 20520 80750
rect 20590 80550 20600 80750
rect 20400 80520 20600 80550
rect 20900 80750 21100 80780
rect 20900 80550 20910 80750
rect 20980 80550 21020 80750
rect 21090 80550 21100 80750
rect 20900 80520 21100 80550
rect 21400 80750 21600 80780
rect 21400 80550 21410 80750
rect 21480 80550 21520 80750
rect 21590 80550 21600 80750
rect 21400 80520 21600 80550
rect 21900 80750 22100 80780
rect 21900 80550 21910 80750
rect 21980 80550 22020 80750
rect 22090 80550 22100 80750
rect 21900 80520 22100 80550
rect 22400 80750 22600 80780
rect 22400 80550 22410 80750
rect 22480 80550 22520 80750
rect 22590 80550 22600 80750
rect 22400 80520 22600 80550
rect 22900 80750 23100 80780
rect 22900 80550 22910 80750
rect 22980 80550 23020 80750
rect 23090 80550 23100 80750
rect 22900 80520 23100 80550
rect 23400 80750 23600 80780
rect 23400 80550 23410 80750
rect 23480 80550 23520 80750
rect 23590 80550 23600 80750
rect 23400 80520 23600 80550
rect 23900 80750 24100 80780
rect 23900 80550 23910 80750
rect 23980 80550 24020 80750
rect 24090 80550 24100 80750
rect 23900 80520 24100 80550
rect 24400 80750 24600 80780
rect 24400 80550 24410 80750
rect 24480 80550 24520 80750
rect 24590 80550 24600 80750
rect 24400 80520 24600 80550
rect 24900 80750 25100 80780
rect 24900 80550 24910 80750
rect 24980 80550 25020 80750
rect 25090 80550 25100 80750
rect 24900 80520 25100 80550
rect 25400 80750 25600 80780
rect 25400 80550 25410 80750
rect 25480 80550 25520 80750
rect 25590 80550 25600 80750
rect 25400 80520 25600 80550
rect 25900 80750 26100 80780
rect 25900 80550 25910 80750
rect 25980 80550 26020 80750
rect 26090 80550 26100 80750
rect 25900 80520 26100 80550
rect 26400 80750 26600 80780
rect 26400 80550 26410 80750
rect 26480 80550 26520 80750
rect 26590 80550 26600 80750
rect 26400 80520 26600 80550
rect 26900 80750 27100 80780
rect 26900 80550 26910 80750
rect 26980 80550 27020 80750
rect 27090 80550 27100 80750
rect 26900 80520 27100 80550
rect 27400 80750 27600 80780
rect 27400 80550 27410 80750
rect 27480 80550 27520 80750
rect 27590 80550 27600 80750
rect 27400 80520 27600 80550
rect 27900 80750 28100 80780
rect 27900 80550 27910 80750
rect 27980 80550 28020 80750
rect 28090 80550 28100 80750
rect 27900 80520 28100 80550
rect 28400 80750 28600 80780
rect 28400 80550 28410 80750
rect 28480 80550 28520 80750
rect 28590 80550 28600 80750
rect 28400 80520 28600 80550
rect 28900 80750 29100 80780
rect 28900 80550 28910 80750
rect 28980 80550 29020 80750
rect 29090 80550 29100 80750
rect 28900 80520 29100 80550
rect 29400 80750 29600 80780
rect 29400 80550 29410 80750
rect 29480 80550 29520 80750
rect 29590 80550 29600 80750
rect 29400 80520 29600 80550
rect 29900 80750 30100 80780
rect 29900 80550 29910 80750
rect 29980 80550 30020 80750
rect 30090 80550 30100 80750
rect 29900 80520 30100 80550
rect 30400 80750 30600 80780
rect 30400 80550 30410 80750
rect 30480 80550 30520 80750
rect 30590 80550 30600 80750
rect 30400 80520 30600 80550
rect 30900 80750 31100 80780
rect 30900 80550 30910 80750
rect 30980 80550 31020 80750
rect 31090 80550 31100 80750
rect 30900 80520 31100 80550
rect 31400 80750 31600 80780
rect 31400 80550 31410 80750
rect 31480 80550 31520 80750
rect 31590 80550 31600 80750
rect 31400 80520 31600 80550
rect 31900 80750 32100 80780
rect 31900 80550 31910 80750
rect 31980 80550 32020 80750
rect 32090 80550 32100 80750
rect 31900 80520 32100 80550
rect 32400 80750 32600 80780
rect 32400 80550 32410 80750
rect 32480 80550 32520 80750
rect 32590 80550 32600 80750
rect 32400 80520 32600 80550
rect 32900 80750 33100 80780
rect 32900 80550 32910 80750
rect 32980 80550 33020 80750
rect 33090 80550 33100 80750
rect 32900 80520 33100 80550
rect 33400 80750 33600 80780
rect 33400 80550 33410 80750
rect 33480 80550 33520 80750
rect 33590 80550 33600 80750
rect 33400 80520 33600 80550
rect 33900 80750 34100 80780
rect 33900 80550 33910 80750
rect 33980 80550 34020 80750
rect 34090 80550 34100 80750
rect 33900 80520 34100 80550
rect 34400 80750 34600 80780
rect 34400 80550 34410 80750
rect 34480 80550 34520 80750
rect 34590 80550 34600 80750
rect 34400 80520 34600 80550
rect 34900 80750 35100 80780
rect 34900 80550 34910 80750
rect 34980 80550 35020 80750
rect 35090 80550 35100 80750
rect 34900 80520 35100 80550
rect 35400 80750 35600 80780
rect 35400 80550 35410 80750
rect 35480 80550 35520 80750
rect 35590 80550 35600 80750
rect 35400 80520 35600 80550
rect 35900 80750 36100 80780
rect 35900 80550 35910 80750
rect 35980 80550 36020 80750
rect 36090 80550 36100 80750
rect 35900 80520 36100 80550
rect 36400 80750 36600 80780
rect 36400 80550 36410 80750
rect 36480 80550 36520 80750
rect 36590 80550 36600 80750
rect 36400 80520 36600 80550
rect 36900 80750 37100 80780
rect 36900 80550 36910 80750
rect 36980 80550 37020 80750
rect 37090 80550 37100 80750
rect 36900 80520 37100 80550
rect 37400 80750 37600 80780
rect 37400 80550 37410 80750
rect 37480 80550 37520 80750
rect 37590 80550 37600 80750
rect 37400 80520 37600 80550
rect 37900 80750 38100 80780
rect 37900 80550 37910 80750
rect 37980 80550 38020 80750
rect 38090 80550 38100 80750
rect 37900 80520 38100 80550
rect 38400 80750 38600 80780
rect 38400 80550 38410 80750
rect 38480 80550 38520 80750
rect 38590 80550 38600 80750
rect 38400 80520 38600 80550
rect 38900 80750 39100 80780
rect 38900 80550 38910 80750
rect 38980 80550 39020 80750
rect 39090 80550 39100 80750
rect 38900 80520 39100 80550
rect 39400 80750 39600 80780
rect 39400 80550 39410 80750
rect 39480 80550 39520 80750
rect 39590 80550 39600 80750
rect 39400 80520 39600 80550
rect 39900 80750 40100 80780
rect 39900 80550 39910 80750
rect 39980 80550 40020 80750
rect 40090 80550 40100 80750
rect 39900 80520 40100 80550
rect 40400 80750 40600 80780
rect 40400 80550 40410 80750
rect 40480 80550 40520 80750
rect 40590 80550 40600 80750
rect 40400 80520 40600 80550
rect 40900 80750 41100 80780
rect 40900 80550 40910 80750
rect 40980 80550 41020 80750
rect 41090 80550 41100 80750
rect 40900 80520 41100 80550
rect 41400 80750 41600 80780
rect 41400 80550 41410 80750
rect 41480 80550 41520 80750
rect 41590 80550 41600 80750
rect 41400 80520 41600 80550
rect 41900 80750 42100 80780
rect 41900 80550 41910 80750
rect 41980 80550 42020 80750
rect 42090 80550 42100 80750
rect 41900 80520 42100 80550
rect 42400 80750 42600 80780
rect 42400 80550 42410 80750
rect 42480 80550 42520 80750
rect 42590 80550 42600 80750
rect 42400 80520 42600 80550
rect 42900 80750 43100 80780
rect 42900 80550 42910 80750
rect 42980 80550 43020 80750
rect 43090 80550 43100 80750
rect 42900 80520 43100 80550
rect 43400 80750 43600 80780
rect 43400 80550 43410 80750
rect 43480 80550 43520 80750
rect 43590 80550 43600 80750
rect 43400 80520 43600 80550
rect 43900 80750 44100 80780
rect 43900 80550 43910 80750
rect 43980 80550 44020 80750
rect 44090 80550 44100 80750
rect 43900 80520 44100 80550
rect 44400 80750 44600 80780
rect 44400 80550 44410 80750
rect 44480 80550 44520 80750
rect 44590 80550 44600 80750
rect 44400 80520 44600 80550
rect 44900 80750 45100 80780
rect 44900 80550 44910 80750
rect 44980 80550 45020 80750
rect 45090 80550 45100 80750
rect 44900 80520 45100 80550
rect 45400 80750 45600 80780
rect 45400 80550 45410 80750
rect 45480 80550 45520 80750
rect 45590 80550 45600 80750
rect 45400 80520 45600 80550
rect 45900 80750 46100 80780
rect 45900 80550 45910 80750
rect 45980 80550 46020 80750
rect 46090 80550 46100 80750
rect 45900 80520 46100 80550
rect 46400 80750 46600 80780
rect 46400 80550 46410 80750
rect 46480 80550 46520 80750
rect 46590 80550 46600 80750
rect 46400 80520 46600 80550
rect 46900 80750 47100 80780
rect 46900 80550 46910 80750
rect 46980 80550 47020 80750
rect 47090 80550 47100 80750
rect 46900 80520 47100 80550
rect 47400 80750 47600 80780
rect 47400 80550 47410 80750
rect 47480 80550 47520 80750
rect 47590 80550 47600 80750
rect 47400 80520 47600 80550
rect 47900 80750 48100 80780
rect 47900 80550 47910 80750
rect 47980 80550 48020 80750
rect 48090 80550 48100 80750
rect 47900 80520 48100 80550
rect 48400 80750 48600 80780
rect 48400 80550 48410 80750
rect 48480 80550 48520 80750
rect 48590 80550 48600 80750
rect 48400 80520 48600 80550
rect 48900 80750 49100 80780
rect 48900 80550 48910 80750
rect 48980 80550 49020 80750
rect 49090 80550 49100 80750
rect 48900 80520 49100 80550
rect 49400 80750 49600 80780
rect 49400 80550 49410 80750
rect 49480 80550 49520 80750
rect 49590 80550 49600 80750
rect 49400 80520 49600 80550
rect 49900 80750 50100 80780
rect 49900 80550 49910 80750
rect 49980 80550 50020 80750
rect 50090 80550 50100 80750
rect 49900 80520 50100 80550
rect 50400 80750 50600 80780
rect 50400 80550 50410 80750
rect 50480 80550 50520 80750
rect 50590 80550 50600 80750
rect 50400 80520 50600 80550
rect 50900 80750 51100 80780
rect 50900 80550 50910 80750
rect 50980 80550 51020 80750
rect 51090 80550 51100 80750
rect 50900 80520 51100 80550
rect 51400 80750 51600 80780
rect 51400 80550 51410 80750
rect 51480 80550 51520 80750
rect 51590 80550 51600 80750
rect 51400 80520 51600 80550
rect 51900 80750 52100 80780
rect 51900 80550 51910 80750
rect 51980 80550 52020 80750
rect 52090 80550 52100 80750
rect 51900 80520 52100 80550
rect 52400 80750 52600 80780
rect 52400 80550 52410 80750
rect 52480 80550 52520 80750
rect 52590 80550 52600 80750
rect 52400 80520 52600 80550
rect 52900 80750 53100 80780
rect 52900 80550 52910 80750
rect 52980 80550 53020 80750
rect 53090 80550 53100 80750
rect 52900 80520 53100 80550
rect 53400 80750 53600 80780
rect 53400 80550 53410 80750
rect 53480 80550 53520 80750
rect 53590 80550 53600 80750
rect 53400 80520 53600 80550
rect 53900 80750 54100 80780
rect 53900 80550 53910 80750
rect 53980 80550 54020 80750
rect 54090 80550 54100 80750
rect 53900 80520 54100 80550
rect 54400 80750 54600 80780
rect 54400 80550 54410 80750
rect 54480 80550 54520 80750
rect 54590 80550 54600 80750
rect 54400 80520 54600 80550
rect 54900 80750 55100 80780
rect 54900 80550 54910 80750
rect 54980 80550 55020 80750
rect 55090 80550 55100 80750
rect 54900 80520 55100 80550
rect 55400 80750 55600 80780
rect 55400 80550 55410 80750
rect 55480 80550 55520 80750
rect 55590 80550 55600 80750
rect 55400 80520 55600 80550
rect 55900 80750 56100 80780
rect 55900 80550 55910 80750
rect 55980 80550 56020 80750
rect 56090 80550 56100 80750
rect 55900 80520 56100 80550
rect 56400 80750 56600 80780
rect 56400 80550 56410 80750
rect 56480 80550 56520 80750
rect 56590 80550 56600 80750
rect 56400 80520 56600 80550
rect 56900 80750 57100 80780
rect 56900 80550 56910 80750
rect 56980 80550 57020 80750
rect 57090 80550 57100 80750
rect 56900 80520 57100 80550
rect 57400 80750 57600 80780
rect 57400 80550 57410 80750
rect 57480 80550 57520 80750
rect 57590 80550 57600 80750
rect 57400 80520 57600 80550
rect 57900 80750 58100 80780
rect 57900 80550 57910 80750
rect 57980 80550 58020 80750
rect 58090 80550 58100 80750
rect 57900 80520 58100 80550
rect 58400 80750 58600 80780
rect 58400 80550 58410 80750
rect 58480 80550 58520 80750
rect 58590 80550 58600 80750
rect 58400 80520 58600 80550
rect 58900 80750 59100 80780
rect 58900 80550 58910 80750
rect 58980 80550 59020 80750
rect 59090 80550 59100 80750
rect 58900 80520 59100 80550
rect 59400 80750 59600 80780
rect 59400 80550 59410 80750
rect 59480 80550 59520 80750
rect 59590 80550 59600 80750
rect 59400 80520 59600 80550
rect 59900 80750 60100 80780
rect 59900 80550 59910 80750
rect 59980 80550 60020 80750
rect 60090 80550 60100 80750
rect 59900 80520 60100 80550
rect 60400 80750 60600 80780
rect 60400 80550 60410 80750
rect 60480 80550 60520 80750
rect 60590 80550 60600 80750
rect 60400 80520 60600 80550
rect 60900 80750 61100 80780
rect 60900 80550 60910 80750
rect 60980 80550 61020 80750
rect 61090 80550 61100 80750
rect 60900 80520 61100 80550
rect 61400 80750 61600 80780
rect 61400 80550 61410 80750
rect 61480 80550 61520 80750
rect 61590 80550 61600 80750
rect 61400 80520 61600 80550
rect 61900 80750 62100 80780
rect 61900 80550 61910 80750
rect 61980 80550 62020 80750
rect 62090 80550 62100 80750
rect 61900 80520 62100 80550
rect 62400 80750 62600 80780
rect 62400 80550 62410 80750
rect 62480 80550 62520 80750
rect 62590 80550 62600 80750
rect 62400 80520 62600 80550
rect 62900 80750 63100 80780
rect 62900 80550 62910 80750
rect 62980 80550 63020 80750
rect 63090 80550 63100 80750
rect 62900 80520 63100 80550
rect 63400 80750 63600 80780
rect 63400 80550 63410 80750
rect 63480 80550 63520 80750
rect 63590 80550 63600 80750
rect 63400 80520 63600 80550
rect 63900 80750 64100 80780
rect 63900 80550 63910 80750
rect 63980 80550 64020 80750
rect 64090 80550 64100 80750
rect 63900 80520 64100 80550
rect 64400 80750 64600 80780
rect 64400 80550 64410 80750
rect 64480 80550 64520 80750
rect 64590 80550 64600 80750
rect 64400 80520 64600 80550
rect 64900 80750 65100 80780
rect 64900 80550 64910 80750
rect 64980 80550 65020 80750
rect 65090 80550 65100 80750
rect 64900 80520 65100 80550
rect 65400 80750 65600 80780
rect 65400 80550 65410 80750
rect 65480 80550 65520 80750
rect 65590 80550 65600 80750
rect 65400 80520 65600 80550
rect 65900 80750 66100 80780
rect 65900 80550 65910 80750
rect 65980 80550 66020 80750
rect 66090 80550 66100 80750
rect 65900 80520 66100 80550
rect 66400 80750 66600 80780
rect 66400 80550 66410 80750
rect 66480 80550 66520 80750
rect 66590 80550 66600 80750
rect 66400 80520 66600 80550
rect 66900 80750 67100 80780
rect 66900 80550 66910 80750
rect 66980 80550 67020 80750
rect 67090 80550 67100 80750
rect 66900 80520 67100 80550
rect 67400 80750 67600 80780
rect 67400 80550 67410 80750
rect 67480 80550 67520 80750
rect 67590 80550 67600 80750
rect 67400 80520 67600 80550
rect 67900 80750 68100 80780
rect 67900 80550 67910 80750
rect 67980 80550 68020 80750
rect 68090 80550 68100 80750
rect 67900 80520 68100 80550
rect 68400 80750 68600 80780
rect 68400 80550 68410 80750
rect 68480 80550 68520 80750
rect 68590 80550 68600 80750
rect 68400 80520 68600 80550
rect 68900 80750 69100 80780
rect 68900 80550 68910 80750
rect 68980 80550 69020 80750
rect 69090 80550 69100 80750
rect 68900 80520 69100 80550
rect 69400 80750 69600 80780
rect 69400 80550 69410 80750
rect 69480 80550 69520 80750
rect 69590 80550 69600 80750
rect 69400 80520 69600 80550
rect 69900 80750 70100 80780
rect 69900 80550 69910 80750
rect 69980 80550 70020 80750
rect 70090 80550 70100 80750
rect 69900 80520 70100 80550
rect 70400 80750 70600 80780
rect 70400 80550 70410 80750
rect 70480 80550 70520 80750
rect 70590 80550 70600 80750
rect 70400 80520 70600 80550
rect 70900 80750 71100 80780
rect 70900 80550 70910 80750
rect 70980 80550 71020 80750
rect 71090 80550 71100 80750
rect 70900 80520 71100 80550
rect 71400 80750 71600 80780
rect 71400 80550 71410 80750
rect 71480 80550 71520 80750
rect 71590 80550 71600 80750
rect 71400 80520 71600 80550
rect 71900 80750 72100 80780
rect 71900 80550 71910 80750
rect 71980 80550 72020 80750
rect 72090 80550 72100 80750
rect 71900 80520 72100 80550
rect 72400 80750 72600 80780
rect 72400 80550 72410 80750
rect 72480 80550 72520 80750
rect 72590 80550 72600 80750
rect 72400 80520 72600 80550
rect 72900 80750 73100 80780
rect 72900 80550 72910 80750
rect 72980 80550 73020 80750
rect 73090 80550 73100 80750
rect 72900 80520 73100 80550
rect 73400 80750 73600 80780
rect 73400 80550 73410 80750
rect 73480 80550 73520 80750
rect 73590 80550 73600 80750
rect 73400 80520 73600 80550
rect 73900 80750 74100 80780
rect 73900 80550 73910 80750
rect 73980 80550 74020 80750
rect 74090 80550 74100 80750
rect 73900 80520 74100 80550
rect 74400 80750 74600 80780
rect 74400 80550 74410 80750
rect 74480 80550 74520 80750
rect 74590 80550 74600 80750
rect 74400 80520 74600 80550
rect 74900 80750 75100 80780
rect 74900 80550 74910 80750
rect 74980 80550 75020 80750
rect 75090 80550 75100 80750
rect 74900 80520 75100 80550
rect 75400 80750 75600 80780
rect 75400 80550 75410 80750
rect 75480 80550 75520 80750
rect 75590 80550 75600 80750
rect 75400 80520 75600 80550
rect 75900 80750 76100 80780
rect 75900 80550 75910 80750
rect 75980 80550 76020 80750
rect 76090 80550 76100 80750
rect 75900 80520 76100 80550
rect 76400 80750 76600 80780
rect 76400 80550 76410 80750
rect 76480 80550 76520 80750
rect 76590 80550 76600 80750
rect 76400 80520 76600 80550
rect 76900 80750 77100 80780
rect 76900 80550 76910 80750
rect 76980 80550 77020 80750
rect 77090 80550 77100 80750
rect 76900 80520 77100 80550
rect 77400 80750 77600 80780
rect 77400 80550 77410 80750
rect 77480 80550 77520 80750
rect 77590 80550 77600 80750
rect 77400 80520 77600 80550
rect 77900 80750 78100 80780
rect 77900 80550 77910 80750
rect 77980 80550 78020 80750
rect 78090 80550 78100 80750
rect 77900 80520 78100 80550
rect 78400 80750 78600 80780
rect 78400 80550 78410 80750
rect 78480 80550 78520 80750
rect 78590 80550 78600 80750
rect 78400 80520 78600 80550
rect 78900 80750 79100 80780
rect 78900 80550 78910 80750
rect 78980 80550 79020 80750
rect 79090 80550 79100 80750
rect 78900 80520 79100 80550
rect 79400 80750 79600 80780
rect 79400 80550 79410 80750
rect 79480 80550 79520 80750
rect 79590 80550 79600 80750
rect 79400 80520 79600 80550
rect 79900 80750 80100 80780
rect 79900 80550 79910 80750
rect 79980 80550 80020 80750
rect 80090 80550 80100 80750
rect 79900 80520 80100 80550
rect 80400 80750 80600 80780
rect 80400 80550 80410 80750
rect 80480 80550 80520 80750
rect 80590 80550 80600 80750
rect 80400 80520 80600 80550
rect 80900 80750 81100 80780
rect 80900 80550 80910 80750
rect 80980 80550 81020 80750
rect 81090 80550 81100 80750
rect 80900 80520 81100 80550
rect 81400 80750 81600 80780
rect 81400 80550 81410 80750
rect 81480 80550 81520 80750
rect 81590 80550 81600 80750
rect 81400 80520 81600 80550
rect 81900 80750 82100 80780
rect 81900 80550 81910 80750
rect 81980 80550 82020 80750
rect 82090 80550 82100 80750
rect 81900 80520 82100 80550
rect 82400 80750 82600 80780
rect 82400 80550 82410 80750
rect 82480 80550 82520 80750
rect 82590 80550 82600 80750
rect 82400 80520 82600 80550
rect 82900 80750 83100 80780
rect 82900 80550 82910 80750
rect 82980 80550 83020 80750
rect 83090 80550 83100 80750
rect 82900 80520 83100 80550
rect 83400 80750 83600 80780
rect 83400 80550 83410 80750
rect 83480 80550 83520 80750
rect 83590 80550 83600 80750
rect 83400 80520 83600 80550
rect 83900 80750 84100 80780
rect 83900 80550 83910 80750
rect 83980 80550 84020 80750
rect 84090 80550 84100 80750
rect 83900 80520 84100 80550
rect 84400 80750 84600 80780
rect 84400 80550 84410 80750
rect 84480 80550 84520 80750
rect 84590 80550 84600 80750
rect 84400 80520 84600 80550
rect 84900 80750 85100 80780
rect 84900 80550 84910 80750
rect 84980 80550 85020 80750
rect 85090 80550 85100 80750
rect 84900 80520 85100 80550
rect 85400 80750 85600 80780
rect 85400 80550 85410 80750
rect 85480 80550 85520 80750
rect 85590 80550 85600 80750
rect 85400 80520 85600 80550
rect 85900 80750 86100 80780
rect 85900 80550 85910 80750
rect 85980 80550 86020 80750
rect 86090 80550 86100 80750
rect 85900 80520 86100 80550
rect 86400 80750 86600 80780
rect 86400 80550 86410 80750
rect 86480 80550 86520 80750
rect 86590 80550 86600 80750
rect 86400 80520 86600 80550
rect 86900 80750 87100 80780
rect 86900 80550 86910 80750
rect 86980 80550 87020 80750
rect 87090 80550 87100 80750
rect 86900 80520 87100 80550
rect 87400 80750 87600 80780
rect 87400 80550 87410 80750
rect 87480 80550 87520 80750
rect 87590 80550 87600 80750
rect 87400 80520 87600 80550
rect 87900 80750 88100 80780
rect 87900 80550 87910 80750
rect 87980 80550 88020 80750
rect 88090 80550 88100 80750
rect 87900 80520 88100 80550
rect 88400 80750 88600 80780
rect 88400 80550 88410 80750
rect 88480 80550 88520 80750
rect 88590 80550 88600 80750
rect 88400 80520 88600 80550
rect 88900 80750 89100 80780
rect 88900 80550 88910 80750
rect 88980 80550 89020 80750
rect 89090 80550 89100 80750
rect 88900 80520 89100 80550
rect 89400 80750 89600 80780
rect 89400 80550 89410 80750
rect 89480 80550 89520 80750
rect 89590 80550 89600 80750
rect 89400 80520 89600 80550
rect 89900 80750 90100 80780
rect 89900 80550 89910 80750
rect 89980 80550 90020 80750
rect 90090 80550 90100 80750
rect 89900 80520 90100 80550
rect 90400 80750 90600 80780
rect 90400 80550 90410 80750
rect 90480 80550 90520 80750
rect 90590 80550 90600 80750
rect 90400 80520 90600 80550
rect 90900 80750 91100 80780
rect 90900 80550 90910 80750
rect 90980 80550 91020 80750
rect 91090 80550 91100 80750
rect 90900 80520 91100 80550
rect 91400 80750 91600 80780
rect 91400 80550 91410 80750
rect 91480 80550 91520 80750
rect 91590 80550 91600 80750
rect 91400 80520 91600 80550
rect 91900 80750 92100 80780
rect 91900 80550 91910 80750
rect 91980 80550 92020 80750
rect 92090 80550 92100 80750
rect 91900 80520 92100 80550
rect 92400 80750 92600 80780
rect 92400 80550 92410 80750
rect 92480 80550 92520 80750
rect 92590 80550 92600 80750
rect 92400 80520 92600 80550
rect 92900 80750 93100 80780
rect 92900 80550 92910 80750
rect 92980 80550 93020 80750
rect 93090 80550 93100 80750
rect 92900 80520 93100 80550
rect 93400 80750 93600 80780
rect 93400 80550 93410 80750
rect 93480 80550 93520 80750
rect 93590 80550 93600 80750
rect 93400 80520 93600 80550
rect 93900 80750 94100 80780
rect 93900 80550 93910 80750
rect 93980 80550 94020 80750
rect 94090 80550 94100 80750
rect 93900 80520 94100 80550
rect 94400 80750 94600 80780
rect 94400 80550 94410 80750
rect 94480 80550 94520 80750
rect 94590 80550 94600 80750
rect 94400 80520 94600 80550
rect 94900 80750 95100 80780
rect 94900 80550 94910 80750
rect 94980 80550 95020 80750
rect 95090 80550 95100 80750
rect 94900 80520 95100 80550
rect 95400 80750 95600 80780
rect 95400 80550 95410 80750
rect 95480 80550 95520 80750
rect 95590 80550 95600 80750
rect 95400 80520 95600 80550
rect 95900 80750 96100 80780
rect 95900 80550 95910 80750
rect 95980 80550 96020 80750
rect 96090 80550 96100 80750
rect 95900 80520 96100 80550
rect 96400 80750 96600 80780
rect 96400 80550 96410 80750
rect 96480 80550 96520 80750
rect 96590 80550 96600 80750
rect 96400 80520 96600 80550
rect 96900 80750 97100 80780
rect 96900 80550 96910 80750
rect 96980 80550 97020 80750
rect 97090 80550 97100 80750
rect 96900 80520 97100 80550
rect 97400 80750 97600 80780
rect 97400 80550 97410 80750
rect 97480 80550 97520 80750
rect 97590 80550 97600 80750
rect 97400 80520 97600 80550
rect 97900 80750 98100 80780
rect 97900 80550 97910 80750
rect 97980 80550 98020 80750
rect 98090 80550 98100 80750
rect 97900 80520 98100 80550
rect 98400 80750 98600 80780
rect 98400 80550 98410 80750
rect 98480 80550 98520 80750
rect 98590 80550 98600 80750
rect 98400 80520 98600 80550
rect 98900 80750 99100 80780
rect 98900 80550 98910 80750
rect 98980 80550 99020 80750
rect 99090 80550 99100 80750
rect 98900 80520 99100 80550
rect 99400 80750 99600 80780
rect 99400 80550 99410 80750
rect 99480 80550 99520 80750
rect 99590 80550 99600 80750
rect 99400 80520 99600 80550
rect 99900 80750 100100 80780
rect 99900 80550 99910 80750
rect 99980 80550 100020 80750
rect 100090 80550 100100 80750
rect 99900 80520 100100 80550
rect 100400 80750 100500 80780
rect 100400 80550 100410 80750
rect 100480 80550 100500 80750
rect 100400 80520 100500 80550
rect -83500 80500 -83380 80520
rect -83120 80500 -82880 80520
rect -82620 80500 -82380 80520
rect -82120 80500 -81880 80520
rect -81620 80500 -81380 80520
rect -81120 80500 -80880 80520
rect -80620 80500 -80380 80520
rect -80120 80500 -79880 80520
rect -79620 80500 -79380 80520
rect -79120 80500 -78880 80520
rect -78620 80500 -78380 80520
rect -78120 80500 -77880 80520
rect -77620 80500 -77380 80520
rect -77120 80500 -76880 80520
rect -76620 80500 -76380 80520
rect -76120 80500 -75880 80520
rect -75620 80500 -75380 80520
rect -75120 80500 -74880 80520
rect -74620 80500 -74380 80520
rect -74120 80500 -73880 80520
rect -73620 80500 -73380 80520
rect -73120 80500 -72880 80520
rect -72620 80500 -72380 80520
rect -72120 80500 -71880 80520
rect -71620 80500 -71380 80520
rect -71120 80500 -70880 80520
rect -70620 80500 -70380 80520
rect -70120 80500 -69880 80520
rect -69620 80500 -69380 80520
rect -69120 80500 -68880 80520
rect -68620 80500 -68380 80520
rect -68120 80500 -67880 80520
rect -67620 80500 -67380 80520
rect -67120 80500 -66880 80520
rect -66620 80500 -66380 80520
rect -66120 80500 -65880 80520
rect -65620 80500 -65380 80520
rect -65120 80500 -64880 80520
rect -64620 80500 -64380 80520
rect -64120 80500 -63880 80520
rect -63620 80500 -63380 80520
rect -63120 80500 -62880 80520
rect -62620 80500 -62380 80520
rect -62120 80500 -61880 80520
rect -61620 80500 -61380 80520
rect -61120 80500 -60880 80520
rect -60620 80500 -60380 80520
rect -60120 80500 -59880 80520
rect -59620 80500 -59380 80520
rect -59120 80500 -58880 80520
rect -58620 80500 -58380 80520
rect -58120 80500 -57880 80520
rect -57620 80500 -57380 80520
rect -57120 80500 -56880 80520
rect -56620 80500 -56380 80520
rect -56120 80500 -55880 80520
rect -55620 80500 -55380 80520
rect -55120 80500 -54880 80520
rect -54620 80500 -54380 80520
rect -54120 80500 -53880 80520
rect -53620 80500 -53380 80520
rect -53120 80500 -52880 80520
rect -52620 80500 -52380 80520
rect -52120 80500 -51880 80520
rect -51620 80500 -51380 80520
rect -51120 80500 -50880 80520
rect -50620 80500 -50380 80520
rect -50120 80500 -49880 80520
rect -49620 80500 -49380 80520
rect -49120 80500 -48880 80520
rect -48620 80500 -48380 80520
rect -48120 80500 -47880 80520
rect -47620 80500 -47380 80520
rect -47120 80500 -46880 80520
rect -46620 80500 -46380 80520
rect -46120 80500 -45880 80520
rect -45620 80500 -45380 80520
rect -45120 80500 -44880 80520
rect -44620 80500 -44380 80520
rect -44120 80500 -43880 80520
rect -43620 80500 -43380 80520
rect -43120 80500 -42880 80520
rect -42620 80500 -42380 80520
rect -42120 80500 -41880 80520
rect -41620 80500 -41380 80520
rect -41120 80500 -40880 80520
rect -40620 80500 -40380 80520
rect -40120 80500 -39880 80520
rect -39620 80500 -39380 80520
rect -39120 80500 -38880 80520
rect -38620 80500 -38380 80520
rect -38120 80500 -37880 80520
rect -37620 80500 -37380 80520
rect -37120 80500 -36880 80520
rect -36620 80500 -36380 80520
rect -36120 80500 -35880 80520
rect -35620 80500 -35380 80520
rect -35120 80500 -34880 80520
rect -34620 80500 -34380 80520
rect -34120 80500 -33880 80520
rect -33620 80500 -33380 80520
rect -33120 80500 -32880 80520
rect -32620 80500 -32380 80520
rect -32120 80500 -31880 80520
rect -31620 80500 -31380 80520
rect -31120 80500 -30880 80520
rect -30620 80500 -30380 80520
rect -30120 80500 -29880 80520
rect -29620 80500 -29380 80520
rect -29120 80500 -28880 80520
rect -28620 80500 -28380 80520
rect -28120 80500 -27880 80520
rect -27620 80500 -27380 80520
rect -27120 80500 -26880 80520
rect -26620 80500 -26380 80520
rect -26120 80500 -25880 80520
rect -25620 80500 -25380 80520
rect -25120 80500 -24880 80520
rect -24620 80500 -24380 80520
rect -24120 80500 -23880 80520
rect -23620 80500 -23380 80520
rect -23120 80500 -22880 80520
rect -22620 80500 -22380 80520
rect -22120 80500 -21880 80520
rect -21620 80500 -21380 80520
rect -21120 80500 -20880 80520
rect -20620 80500 -20380 80520
rect -20120 80500 -19880 80520
rect -19620 80500 -19380 80520
rect -19120 80500 -18880 80520
rect -18620 80500 -18380 80520
rect -18120 80500 -17880 80520
rect -17620 80500 -17380 80520
rect -17120 80500 -16880 80520
rect -16620 80500 -16380 80520
rect -16120 80500 -15880 80520
rect -15620 80500 -15380 80520
rect -15120 80500 -14880 80520
rect -14620 80500 -14380 80520
rect -14120 80500 -13880 80520
rect -13620 80500 -13380 80520
rect -13120 80500 -12880 80520
rect -12620 80500 -12380 80520
rect -12120 80500 -11880 80520
rect -11620 80500 -11380 80520
rect -11120 80500 -10880 80520
rect -10620 80500 -10380 80520
rect -10120 80500 -9880 80520
rect -9620 80500 -9380 80520
rect -9120 80500 -8880 80520
rect -8620 80500 -8380 80520
rect -8120 80500 -7880 80520
rect -7620 80500 -7380 80520
rect -7120 80500 -6880 80520
rect -6620 80500 -6380 80520
rect -6120 80500 -5880 80520
rect -5620 80500 -5380 80520
rect -5120 80500 -4880 80520
rect -4620 80500 -4380 80520
rect -4120 80500 -3880 80520
rect -3620 80500 -3380 80520
rect -3120 80500 -2880 80520
rect -2620 80500 -2380 80520
rect -2120 80500 -1880 80520
rect -1620 80500 -1380 80520
rect -1120 80500 -880 80520
rect -620 80500 -380 80520
rect -120 80500 120 80520
rect 380 80500 620 80520
rect 880 80500 1120 80520
rect 1380 80500 1620 80520
rect 1880 80500 2120 80520
rect 2380 80500 2620 80520
rect 2880 80500 3120 80520
rect 3380 80500 3620 80520
rect 3880 80500 4120 80520
rect 4380 80500 4620 80520
rect 4880 80500 5120 80520
rect 5380 80500 5620 80520
rect 5880 80500 6120 80520
rect 6380 80500 6620 80520
rect 6880 80500 7120 80520
rect 7380 80500 7620 80520
rect 7880 80500 8120 80520
rect 8380 80500 8620 80520
rect 8880 80500 9120 80520
rect 9380 80500 9620 80520
rect 9880 80500 10120 80520
rect 10380 80500 10620 80520
rect 10880 80500 11120 80520
rect 11380 80500 11620 80520
rect 11880 80500 12120 80520
rect 12380 80500 12620 80520
rect 12880 80500 13120 80520
rect 13380 80500 13620 80520
rect 13880 80500 14120 80520
rect 14380 80500 14620 80520
rect 14880 80500 15120 80520
rect 15380 80500 15620 80520
rect 15880 80500 16120 80520
rect 16380 80500 16620 80520
rect 16880 80500 17120 80520
rect 17380 80500 17620 80520
rect 17880 80500 18120 80520
rect 18380 80500 18620 80520
rect 18880 80500 19120 80520
rect 19380 80500 19620 80520
rect 19880 80500 20120 80520
rect 20380 80500 20620 80520
rect 20880 80500 21120 80520
rect 21380 80500 21620 80520
rect 21880 80500 22120 80520
rect 22380 80500 22620 80520
rect 22880 80500 23120 80520
rect 23380 80500 23620 80520
rect 23880 80500 24120 80520
rect 24380 80500 24620 80520
rect 24880 80500 25120 80520
rect 25380 80500 25620 80520
rect 25880 80500 26120 80520
rect 26380 80500 26620 80520
rect 26880 80500 27120 80520
rect 27380 80500 27620 80520
rect 27880 80500 28120 80520
rect 28380 80500 28620 80520
rect 28880 80500 29120 80520
rect 29380 80500 29620 80520
rect 29880 80500 30120 80520
rect 30380 80500 30620 80520
rect 30880 80500 31120 80520
rect 31380 80500 31620 80520
rect 31880 80500 32120 80520
rect 32380 80500 32620 80520
rect 32880 80500 33120 80520
rect 33380 80500 33620 80520
rect 33880 80500 34120 80520
rect 34380 80500 34620 80520
rect 34880 80500 35120 80520
rect 35380 80500 35620 80520
rect 35880 80500 36120 80520
rect 36380 80500 36620 80520
rect 36880 80500 37120 80520
rect 37380 80500 37620 80520
rect 37880 80500 38120 80520
rect 38380 80500 38620 80520
rect 38880 80500 39120 80520
rect 39380 80500 39620 80520
rect 39880 80500 40120 80520
rect 40380 80500 40620 80520
rect 40880 80500 41120 80520
rect 41380 80500 41620 80520
rect 41880 80500 42120 80520
rect 42380 80500 42620 80520
rect 42880 80500 43120 80520
rect 43380 80500 43620 80520
rect 43880 80500 44120 80520
rect 44380 80500 44620 80520
rect 44880 80500 45120 80520
rect 45380 80500 45620 80520
rect 45880 80500 46120 80520
rect 46380 80500 46620 80520
rect 46880 80500 47120 80520
rect 47380 80500 47620 80520
rect 47880 80500 48120 80520
rect 48380 80500 48620 80520
rect 48880 80500 49120 80520
rect 49380 80500 49620 80520
rect 49880 80500 50120 80520
rect 50380 80500 50620 80520
rect 50880 80500 51120 80520
rect 51380 80500 51620 80520
rect 51880 80500 52120 80520
rect 52380 80500 52620 80520
rect 52880 80500 53120 80520
rect 53380 80500 53620 80520
rect 53880 80500 54120 80520
rect 54380 80500 54620 80520
rect 54880 80500 55120 80520
rect 55380 80500 55620 80520
rect 55880 80500 56120 80520
rect 56380 80500 56620 80520
rect 56880 80500 57120 80520
rect 57380 80500 57620 80520
rect 57880 80500 58120 80520
rect 58380 80500 58620 80520
rect 58880 80500 59120 80520
rect 59380 80500 59620 80520
rect 59880 80500 60120 80520
rect 60380 80500 60620 80520
rect 60880 80500 61120 80520
rect 61380 80500 61620 80520
rect 61880 80500 62120 80520
rect 62380 80500 62620 80520
rect 62880 80500 63120 80520
rect 63380 80500 63620 80520
rect 63880 80500 64120 80520
rect 64380 80500 64620 80520
rect 64880 80500 65120 80520
rect 65380 80500 65620 80520
rect 65880 80500 66120 80520
rect 66380 80500 66620 80520
rect 66880 80500 67120 80520
rect 67380 80500 67620 80520
rect 67880 80500 68120 80520
rect 68380 80500 68620 80520
rect 68880 80500 69120 80520
rect 69380 80500 69620 80520
rect 69880 80500 70120 80520
rect 70380 80500 70620 80520
rect 70880 80500 71120 80520
rect 71380 80500 71620 80520
rect 71880 80500 72120 80520
rect 72380 80500 72620 80520
rect 72880 80500 73120 80520
rect 73380 80500 73620 80520
rect 73880 80500 74120 80520
rect 74380 80500 74620 80520
rect 74880 80500 75120 80520
rect 75380 80500 75620 80520
rect 75880 80500 76120 80520
rect 76380 80500 76620 80520
rect 76880 80500 77120 80520
rect 77380 80500 77620 80520
rect 77880 80500 78120 80520
rect 78380 80500 78620 80520
rect 78880 80500 79120 80520
rect 79380 80500 79620 80520
rect 79880 80500 80120 80520
rect 80380 80500 80620 80520
rect 80880 80500 81120 80520
rect 81380 80500 81620 80520
rect 81880 80500 82120 80520
rect 82380 80500 82620 80520
rect 82880 80500 83120 80520
rect 83380 80500 83620 80520
rect 83880 80500 84120 80520
rect 84380 80500 84620 80520
rect 84880 80500 85120 80520
rect 85380 80500 85620 80520
rect 85880 80500 86120 80520
rect 86380 80500 86620 80520
rect 86880 80500 87120 80520
rect 87380 80500 87620 80520
rect 87880 80500 88120 80520
rect 88380 80500 88620 80520
rect 88880 80500 89120 80520
rect 89380 80500 89620 80520
rect 89880 80500 90120 80520
rect 90380 80500 90620 80520
rect 90880 80500 91120 80520
rect 91380 80500 91620 80520
rect 91880 80500 92120 80520
rect 92380 80500 92620 80520
rect 92880 80500 93120 80520
rect 93380 80500 93620 80520
rect 93880 80500 94120 80520
rect 94380 80500 94620 80520
rect 94880 80500 95120 80520
rect 95380 80500 95620 80520
rect 95880 80500 96120 80520
rect 96380 80500 96620 80520
rect 96880 80500 97120 80520
rect 97380 80500 97620 80520
rect 97880 80500 98120 80520
rect 98380 80500 98620 80520
rect 98880 80500 99120 80520
rect 99380 80500 99620 80520
rect 99880 80500 100120 80520
rect 100380 80500 100500 80520
rect -83500 80490 100500 80500
rect -83500 80420 -83350 80490
rect -83150 80420 -82850 80490
rect -82650 80420 -82350 80490
rect -82150 80420 -81850 80490
rect -81650 80420 -81350 80490
rect -81150 80420 -80850 80490
rect -80650 80420 -80350 80490
rect -80150 80420 -79850 80490
rect -79650 80420 -79350 80490
rect -79150 80420 -78850 80490
rect -78650 80420 -78350 80490
rect -78150 80420 -77850 80490
rect -77650 80420 -77350 80490
rect -77150 80420 -76850 80490
rect -76650 80420 -76350 80490
rect -76150 80420 -75850 80490
rect -75650 80420 -75350 80490
rect -75150 80420 -74850 80490
rect -74650 80420 -74350 80490
rect -74150 80420 -73850 80490
rect -73650 80420 -73350 80490
rect -73150 80420 -72850 80490
rect -72650 80420 -72350 80490
rect -72150 80420 -71850 80490
rect -71650 80420 -71350 80490
rect -71150 80420 -70850 80490
rect -70650 80420 -70350 80490
rect -70150 80420 -69850 80490
rect -69650 80420 -69350 80490
rect -69150 80420 -68850 80490
rect -68650 80420 -68350 80490
rect -68150 80420 -67850 80490
rect -67650 80420 -67350 80490
rect -67150 80420 -66850 80490
rect -66650 80420 -66350 80490
rect -66150 80420 -65850 80490
rect -65650 80420 -65350 80490
rect -65150 80420 -64850 80490
rect -64650 80420 -64350 80490
rect -64150 80420 -63850 80490
rect -63650 80420 -63350 80490
rect -63150 80420 -62850 80490
rect -62650 80420 -62350 80490
rect -62150 80420 -61850 80490
rect -61650 80420 -61350 80490
rect -61150 80420 -60850 80490
rect -60650 80420 -60350 80490
rect -60150 80420 -59850 80490
rect -59650 80420 -59350 80490
rect -59150 80420 -58850 80490
rect -58650 80420 -58350 80490
rect -58150 80420 -57850 80490
rect -57650 80420 -57350 80490
rect -57150 80420 -56850 80490
rect -56650 80420 -56350 80490
rect -56150 80420 -55850 80490
rect -55650 80420 -55350 80490
rect -55150 80420 -54850 80490
rect -54650 80420 -54350 80490
rect -54150 80420 -53850 80490
rect -53650 80420 -53350 80490
rect -53150 80420 -52850 80490
rect -52650 80420 -52350 80490
rect -52150 80420 -51850 80490
rect -51650 80420 -51350 80490
rect -51150 80420 -50850 80490
rect -50650 80420 -50350 80490
rect -50150 80420 -49850 80490
rect -49650 80420 -49350 80490
rect -49150 80420 -48850 80490
rect -48650 80420 -48350 80490
rect -48150 80420 -47850 80490
rect -47650 80420 -47350 80490
rect -47150 80420 -46850 80490
rect -46650 80420 -46350 80490
rect -46150 80420 -45850 80490
rect -45650 80420 -45350 80490
rect -45150 80420 -44850 80490
rect -44650 80420 -44350 80490
rect -44150 80420 -43850 80490
rect -43650 80420 -43350 80490
rect -43150 80420 -42850 80490
rect -42650 80420 -42350 80490
rect -42150 80420 -41850 80490
rect -41650 80420 -41350 80490
rect -41150 80420 -40850 80490
rect -40650 80420 -40350 80490
rect -40150 80420 -39850 80490
rect -39650 80420 -39350 80490
rect -39150 80420 -38850 80490
rect -38650 80420 -38350 80490
rect -38150 80420 -37850 80490
rect -37650 80420 -37350 80490
rect -37150 80420 -36850 80490
rect -36650 80420 -36350 80490
rect -36150 80420 -35850 80490
rect -35650 80420 -35350 80490
rect -35150 80420 -34850 80490
rect -34650 80420 -34350 80490
rect -34150 80420 -33850 80490
rect -33650 80420 -33350 80490
rect -33150 80420 -32850 80490
rect -32650 80420 -32350 80490
rect -32150 80420 -31850 80490
rect -31650 80420 -31350 80490
rect -31150 80420 -30850 80490
rect -30650 80420 -30350 80490
rect -30150 80420 -29850 80490
rect -29650 80420 -29350 80490
rect -29150 80420 -28850 80490
rect -28650 80420 -28350 80490
rect -28150 80420 -27850 80490
rect -27650 80420 -27350 80490
rect -27150 80420 -26850 80490
rect -26650 80420 -26350 80490
rect -26150 80420 -25850 80490
rect -25650 80420 -25350 80490
rect -25150 80420 -24850 80490
rect -24650 80420 -24350 80490
rect -24150 80420 -23850 80490
rect -23650 80420 -23350 80490
rect -23150 80420 -22850 80490
rect -22650 80420 -22350 80490
rect -22150 80420 -21850 80490
rect -21650 80420 -21350 80490
rect -21150 80420 -20850 80490
rect -20650 80420 -20350 80490
rect -20150 80420 -19850 80490
rect -19650 80420 -19350 80490
rect -19150 80420 -18850 80490
rect -18650 80420 -18350 80490
rect -18150 80420 -17850 80490
rect -17650 80420 -17350 80490
rect -17150 80420 -16850 80490
rect -16650 80420 -16350 80490
rect -16150 80420 -15850 80490
rect -15650 80420 -15350 80490
rect -15150 80420 -14850 80490
rect -14650 80420 -14350 80490
rect -14150 80420 -13850 80490
rect -13650 80420 -13350 80490
rect -13150 80420 -12850 80490
rect -12650 80420 -12350 80490
rect -12150 80420 -11850 80490
rect -11650 80420 -11350 80490
rect -11150 80420 -10850 80490
rect -10650 80420 -10350 80490
rect -10150 80420 -9850 80490
rect -9650 80420 -9350 80490
rect -9150 80420 -8850 80490
rect -8650 80420 -8350 80490
rect -8150 80420 -7850 80490
rect -7650 80420 -7350 80490
rect -7150 80420 -6850 80490
rect -6650 80420 -6350 80490
rect -6150 80420 -5850 80490
rect -5650 80420 -5350 80490
rect -5150 80420 -4850 80490
rect -4650 80420 -4350 80490
rect -4150 80420 -3850 80490
rect -3650 80420 -3350 80490
rect -3150 80420 -2850 80490
rect -2650 80420 -2350 80490
rect -2150 80420 -1850 80490
rect -1650 80420 -1350 80490
rect -1150 80420 -850 80490
rect -650 80420 -350 80490
rect -150 80420 150 80490
rect 350 80420 650 80490
rect 850 80420 1150 80490
rect 1350 80420 1650 80490
rect 1850 80420 2150 80490
rect 2350 80420 2650 80490
rect 2850 80420 3150 80490
rect 3350 80420 3650 80490
rect 3850 80420 4150 80490
rect 4350 80420 4650 80490
rect 4850 80420 5150 80490
rect 5350 80420 5650 80490
rect 5850 80420 6150 80490
rect 6350 80420 6650 80490
rect 6850 80420 7150 80490
rect 7350 80420 7650 80490
rect 7850 80420 8150 80490
rect 8350 80420 8650 80490
rect 8850 80420 9150 80490
rect 9350 80420 9650 80490
rect 9850 80420 10150 80490
rect 10350 80420 10650 80490
rect 10850 80420 11150 80490
rect 11350 80420 11650 80490
rect 11850 80420 12150 80490
rect 12350 80420 12650 80490
rect 12850 80420 13150 80490
rect 13350 80420 13650 80490
rect 13850 80420 14150 80490
rect 14350 80420 14650 80490
rect 14850 80420 15150 80490
rect 15350 80420 15650 80490
rect 15850 80420 16150 80490
rect 16350 80420 16650 80490
rect 16850 80420 17150 80490
rect 17350 80420 17650 80490
rect 17850 80420 18150 80490
rect 18350 80420 18650 80490
rect 18850 80420 19150 80490
rect 19350 80420 19650 80490
rect 19850 80420 20150 80490
rect 20350 80420 20650 80490
rect 20850 80420 21150 80490
rect 21350 80420 21650 80490
rect 21850 80420 22150 80490
rect 22350 80420 22650 80490
rect 22850 80420 23150 80490
rect 23350 80420 23650 80490
rect 23850 80420 24150 80490
rect 24350 80420 24650 80490
rect 24850 80420 25150 80490
rect 25350 80420 25650 80490
rect 25850 80420 26150 80490
rect 26350 80420 26650 80490
rect 26850 80420 27150 80490
rect 27350 80420 27650 80490
rect 27850 80420 28150 80490
rect 28350 80420 28650 80490
rect 28850 80420 29150 80490
rect 29350 80420 29650 80490
rect 29850 80420 30150 80490
rect 30350 80420 30650 80490
rect 30850 80420 31150 80490
rect 31350 80420 31650 80490
rect 31850 80420 32150 80490
rect 32350 80420 32650 80490
rect 32850 80420 33150 80490
rect 33350 80420 33650 80490
rect 33850 80420 34150 80490
rect 34350 80420 34650 80490
rect 34850 80420 35150 80490
rect 35350 80420 35650 80490
rect 35850 80420 36150 80490
rect 36350 80420 36650 80490
rect 36850 80420 37150 80490
rect 37350 80420 37650 80490
rect 37850 80420 38150 80490
rect 38350 80420 38650 80490
rect 38850 80420 39150 80490
rect 39350 80420 39650 80490
rect 39850 80420 40150 80490
rect 40350 80420 40650 80490
rect 40850 80420 41150 80490
rect 41350 80420 41650 80490
rect 41850 80420 42150 80490
rect 42350 80420 42650 80490
rect 42850 80420 43150 80490
rect 43350 80420 43650 80490
rect 43850 80420 44150 80490
rect 44350 80420 44650 80490
rect 44850 80420 45150 80490
rect 45350 80420 45650 80490
rect 45850 80420 46150 80490
rect 46350 80420 46650 80490
rect 46850 80420 47150 80490
rect 47350 80420 47650 80490
rect 47850 80420 48150 80490
rect 48350 80420 48650 80490
rect 48850 80420 49150 80490
rect 49350 80420 49650 80490
rect 49850 80420 50150 80490
rect 50350 80420 50650 80490
rect 50850 80420 51150 80490
rect 51350 80420 51650 80490
rect 51850 80420 52150 80490
rect 52350 80420 52650 80490
rect 52850 80420 53150 80490
rect 53350 80420 53650 80490
rect 53850 80420 54150 80490
rect 54350 80420 54650 80490
rect 54850 80420 55150 80490
rect 55350 80420 55650 80490
rect 55850 80420 56150 80490
rect 56350 80420 56650 80490
rect 56850 80420 57150 80490
rect 57350 80420 57650 80490
rect 57850 80420 58150 80490
rect 58350 80420 58650 80490
rect 58850 80420 59150 80490
rect 59350 80420 59650 80490
rect 59850 80420 60150 80490
rect 60350 80420 60650 80490
rect 60850 80420 61150 80490
rect 61350 80420 61650 80490
rect 61850 80420 62150 80490
rect 62350 80420 62650 80490
rect 62850 80420 63150 80490
rect 63350 80420 63650 80490
rect 63850 80420 64150 80490
rect 64350 80420 64650 80490
rect 64850 80420 65150 80490
rect 65350 80420 65650 80490
rect 65850 80420 66150 80490
rect 66350 80420 66650 80490
rect 66850 80420 67150 80490
rect 67350 80420 67650 80490
rect 67850 80420 68150 80490
rect 68350 80420 68650 80490
rect 68850 80420 69150 80490
rect 69350 80420 69650 80490
rect 69850 80420 70150 80490
rect 70350 80420 70650 80490
rect 70850 80420 71150 80490
rect 71350 80420 71650 80490
rect 71850 80420 72150 80490
rect 72350 80420 72650 80490
rect 72850 80420 73150 80490
rect 73350 80420 73650 80490
rect 73850 80420 74150 80490
rect 74350 80420 74650 80490
rect 74850 80420 75150 80490
rect 75350 80420 75650 80490
rect 75850 80420 76150 80490
rect 76350 80420 76650 80490
rect 76850 80420 77150 80490
rect 77350 80420 77650 80490
rect 77850 80420 78150 80490
rect 78350 80420 78650 80490
rect 78850 80420 79150 80490
rect 79350 80420 79650 80490
rect 79850 80420 80150 80490
rect 80350 80420 80650 80490
rect 80850 80420 81150 80490
rect 81350 80420 81650 80490
rect 81850 80420 82150 80490
rect 82350 80420 82650 80490
rect 82850 80420 83150 80490
rect 83350 80420 83650 80490
rect 83850 80420 84150 80490
rect 84350 80420 84650 80490
rect 84850 80420 85150 80490
rect 85350 80420 85650 80490
rect 85850 80420 86150 80490
rect 86350 80420 86650 80490
rect 86850 80420 87150 80490
rect 87350 80420 87650 80490
rect 87850 80420 88150 80490
rect 88350 80420 88650 80490
rect 88850 80420 89150 80490
rect 89350 80420 89650 80490
rect 89850 80420 90150 80490
rect 90350 80420 90650 80490
rect 90850 80420 91150 80490
rect 91350 80420 91650 80490
rect 91850 80420 92150 80490
rect 92350 80420 92650 80490
rect 92850 80420 93150 80490
rect 93350 80420 93650 80490
rect 93850 80420 94150 80490
rect 94350 80420 94650 80490
rect 94850 80420 95150 80490
rect 95350 80420 95650 80490
rect 95850 80420 96150 80490
rect 96350 80420 96650 80490
rect 96850 80420 97150 80490
rect 97350 80420 97650 80490
rect 97850 80420 98150 80490
rect 98350 80420 98650 80490
rect 98850 80420 99150 80490
rect 99350 80420 99650 80490
rect 99850 80420 100150 80490
rect 100350 80420 100500 80490
rect -83500 80380 100500 80420
rect -83500 80310 -83350 80380
rect -83150 80310 -82850 80380
rect -82650 80310 -82350 80380
rect -82150 80310 -81850 80380
rect -81650 80310 -81350 80380
rect -81150 80310 -80850 80380
rect -80650 80310 -80350 80380
rect -80150 80310 -79850 80380
rect -79650 80310 -79350 80380
rect -79150 80310 -78850 80380
rect -78650 80310 -78350 80380
rect -78150 80310 -77850 80380
rect -77650 80310 -77350 80380
rect -77150 80310 -76850 80380
rect -76650 80310 -76350 80380
rect -76150 80310 -75850 80380
rect -75650 80310 -75350 80380
rect -75150 80310 -74850 80380
rect -74650 80310 -74350 80380
rect -74150 80310 -73850 80380
rect -73650 80310 -73350 80380
rect -73150 80310 -72850 80380
rect -72650 80310 -72350 80380
rect -72150 80310 -71850 80380
rect -71650 80310 -71350 80380
rect -71150 80310 -70850 80380
rect -70650 80310 -70350 80380
rect -70150 80310 -69850 80380
rect -69650 80310 -69350 80380
rect -69150 80310 -68850 80380
rect -68650 80310 -68350 80380
rect -68150 80310 -67850 80380
rect -67650 80310 -67350 80380
rect -67150 80310 -66850 80380
rect -66650 80310 -66350 80380
rect -66150 80310 -65850 80380
rect -65650 80310 -65350 80380
rect -65150 80310 -64850 80380
rect -64650 80310 -64350 80380
rect -64150 80310 -63850 80380
rect -63650 80310 -63350 80380
rect -63150 80310 -62850 80380
rect -62650 80310 -62350 80380
rect -62150 80310 -61850 80380
rect -61650 80310 -61350 80380
rect -61150 80310 -60850 80380
rect -60650 80310 -60350 80380
rect -60150 80310 -59850 80380
rect -59650 80310 -59350 80380
rect -59150 80310 -58850 80380
rect -58650 80310 -58350 80380
rect -58150 80310 -57850 80380
rect -57650 80310 -57350 80380
rect -57150 80310 -56850 80380
rect -56650 80310 -56350 80380
rect -56150 80310 -55850 80380
rect -55650 80310 -55350 80380
rect -55150 80310 -54850 80380
rect -54650 80310 -54350 80380
rect -54150 80310 -53850 80380
rect -53650 80310 -53350 80380
rect -53150 80310 -52850 80380
rect -52650 80310 -52350 80380
rect -52150 80310 -51850 80380
rect -51650 80310 -51350 80380
rect -51150 80310 -50850 80380
rect -50650 80310 -50350 80380
rect -50150 80310 -49850 80380
rect -49650 80310 -49350 80380
rect -49150 80310 -48850 80380
rect -48650 80310 -48350 80380
rect -48150 80310 -47850 80380
rect -47650 80310 -47350 80380
rect -47150 80310 -46850 80380
rect -46650 80310 -46350 80380
rect -46150 80310 -45850 80380
rect -45650 80310 -45350 80380
rect -45150 80310 -44850 80380
rect -44650 80310 -44350 80380
rect -44150 80310 -43850 80380
rect -43650 80310 -43350 80380
rect -43150 80310 -42850 80380
rect -42650 80310 -42350 80380
rect -42150 80310 -41850 80380
rect -41650 80310 -41350 80380
rect -41150 80310 -40850 80380
rect -40650 80310 -40350 80380
rect -40150 80310 -39850 80380
rect -39650 80310 -39350 80380
rect -39150 80310 -38850 80380
rect -38650 80310 -38350 80380
rect -38150 80310 -37850 80380
rect -37650 80310 -37350 80380
rect -37150 80310 -36850 80380
rect -36650 80310 -36350 80380
rect -36150 80310 -35850 80380
rect -35650 80310 -35350 80380
rect -35150 80310 -34850 80380
rect -34650 80310 -34350 80380
rect -34150 80310 -33850 80380
rect -33650 80310 -33350 80380
rect -33150 80310 -32850 80380
rect -32650 80310 -32350 80380
rect -32150 80310 -31850 80380
rect -31650 80310 -31350 80380
rect -31150 80310 -30850 80380
rect -30650 80310 -30350 80380
rect -30150 80310 -29850 80380
rect -29650 80310 -29350 80380
rect -29150 80310 -28850 80380
rect -28650 80310 -28350 80380
rect -28150 80310 -27850 80380
rect -27650 80310 -27350 80380
rect -27150 80310 -26850 80380
rect -26650 80310 -26350 80380
rect -26150 80310 -25850 80380
rect -25650 80310 -25350 80380
rect -25150 80310 -24850 80380
rect -24650 80310 -24350 80380
rect -24150 80310 -23850 80380
rect -23650 80310 -23350 80380
rect -23150 80310 -22850 80380
rect -22650 80310 -22350 80380
rect -22150 80310 -21850 80380
rect -21650 80310 -21350 80380
rect -21150 80310 -20850 80380
rect -20650 80310 -20350 80380
rect -20150 80310 -19850 80380
rect -19650 80310 -19350 80380
rect -19150 80310 -18850 80380
rect -18650 80310 -18350 80380
rect -18150 80310 -17850 80380
rect -17650 80310 -17350 80380
rect -17150 80310 -16850 80380
rect -16650 80310 -16350 80380
rect -16150 80310 -15850 80380
rect -15650 80310 -15350 80380
rect -15150 80310 -14850 80380
rect -14650 80310 -14350 80380
rect -14150 80310 -13850 80380
rect -13650 80310 -13350 80380
rect -13150 80310 -12850 80380
rect -12650 80310 -12350 80380
rect -12150 80310 -11850 80380
rect -11650 80310 -11350 80380
rect -11150 80310 -10850 80380
rect -10650 80310 -10350 80380
rect -10150 80310 -9850 80380
rect -9650 80310 -9350 80380
rect -9150 80310 -8850 80380
rect -8650 80310 -8350 80380
rect -8150 80310 -7850 80380
rect -7650 80310 -7350 80380
rect -7150 80310 -6850 80380
rect -6650 80310 -6350 80380
rect -6150 80310 -5850 80380
rect -5650 80310 -5350 80380
rect -5150 80310 -4850 80380
rect -4650 80310 -4350 80380
rect -4150 80310 -3850 80380
rect -3650 80310 -3350 80380
rect -3150 80310 -2850 80380
rect -2650 80310 -2350 80380
rect -2150 80310 -1850 80380
rect -1650 80310 -1350 80380
rect -1150 80310 -850 80380
rect -650 80310 -350 80380
rect -150 80310 150 80380
rect 350 80310 650 80380
rect 850 80310 1150 80380
rect 1350 80310 1650 80380
rect 1850 80310 2150 80380
rect 2350 80310 2650 80380
rect 2850 80310 3150 80380
rect 3350 80310 3650 80380
rect 3850 80310 4150 80380
rect 4350 80310 4650 80380
rect 4850 80310 5150 80380
rect 5350 80310 5650 80380
rect 5850 80310 6150 80380
rect 6350 80310 6650 80380
rect 6850 80310 7150 80380
rect 7350 80310 7650 80380
rect 7850 80310 8150 80380
rect 8350 80310 8650 80380
rect 8850 80310 9150 80380
rect 9350 80310 9650 80380
rect 9850 80310 10150 80380
rect 10350 80310 10650 80380
rect 10850 80310 11150 80380
rect 11350 80310 11650 80380
rect 11850 80310 12150 80380
rect 12350 80310 12650 80380
rect 12850 80310 13150 80380
rect 13350 80310 13650 80380
rect 13850 80310 14150 80380
rect 14350 80310 14650 80380
rect 14850 80310 15150 80380
rect 15350 80310 15650 80380
rect 15850 80310 16150 80380
rect 16350 80310 16650 80380
rect 16850 80310 17150 80380
rect 17350 80310 17650 80380
rect 17850 80310 18150 80380
rect 18350 80310 18650 80380
rect 18850 80310 19150 80380
rect 19350 80310 19650 80380
rect 19850 80310 20150 80380
rect 20350 80310 20650 80380
rect 20850 80310 21150 80380
rect 21350 80310 21650 80380
rect 21850 80310 22150 80380
rect 22350 80310 22650 80380
rect 22850 80310 23150 80380
rect 23350 80310 23650 80380
rect 23850 80310 24150 80380
rect 24350 80310 24650 80380
rect 24850 80310 25150 80380
rect 25350 80310 25650 80380
rect 25850 80310 26150 80380
rect 26350 80310 26650 80380
rect 26850 80310 27150 80380
rect 27350 80310 27650 80380
rect 27850 80310 28150 80380
rect 28350 80310 28650 80380
rect 28850 80310 29150 80380
rect 29350 80310 29650 80380
rect 29850 80310 30150 80380
rect 30350 80310 30650 80380
rect 30850 80310 31150 80380
rect 31350 80310 31650 80380
rect 31850 80310 32150 80380
rect 32350 80310 32650 80380
rect 32850 80310 33150 80380
rect 33350 80310 33650 80380
rect 33850 80310 34150 80380
rect 34350 80310 34650 80380
rect 34850 80310 35150 80380
rect 35350 80310 35650 80380
rect 35850 80310 36150 80380
rect 36350 80310 36650 80380
rect 36850 80310 37150 80380
rect 37350 80310 37650 80380
rect 37850 80310 38150 80380
rect 38350 80310 38650 80380
rect 38850 80310 39150 80380
rect 39350 80310 39650 80380
rect 39850 80310 40150 80380
rect 40350 80310 40650 80380
rect 40850 80310 41150 80380
rect 41350 80310 41650 80380
rect 41850 80310 42150 80380
rect 42350 80310 42650 80380
rect 42850 80310 43150 80380
rect 43350 80310 43650 80380
rect 43850 80310 44150 80380
rect 44350 80310 44650 80380
rect 44850 80310 45150 80380
rect 45350 80310 45650 80380
rect 45850 80310 46150 80380
rect 46350 80310 46650 80380
rect 46850 80310 47150 80380
rect 47350 80310 47650 80380
rect 47850 80310 48150 80380
rect 48350 80310 48650 80380
rect 48850 80310 49150 80380
rect 49350 80310 49650 80380
rect 49850 80310 50150 80380
rect 50350 80310 50650 80380
rect 50850 80310 51150 80380
rect 51350 80310 51650 80380
rect 51850 80310 52150 80380
rect 52350 80310 52650 80380
rect 52850 80310 53150 80380
rect 53350 80310 53650 80380
rect 53850 80310 54150 80380
rect 54350 80310 54650 80380
rect 54850 80310 55150 80380
rect 55350 80310 55650 80380
rect 55850 80310 56150 80380
rect 56350 80310 56650 80380
rect 56850 80310 57150 80380
rect 57350 80310 57650 80380
rect 57850 80310 58150 80380
rect 58350 80310 58650 80380
rect 58850 80310 59150 80380
rect 59350 80310 59650 80380
rect 59850 80310 60150 80380
rect 60350 80310 60650 80380
rect 60850 80310 61150 80380
rect 61350 80310 61650 80380
rect 61850 80310 62150 80380
rect 62350 80310 62650 80380
rect 62850 80310 63150 80380
rect 63350 80310 63650 80380
rect 63850 80310 64150 80380
rect 64350 80310 64650 80380
rect 64850 80310 65150 80380
rect 65350 80310 65650 80380
rect 65850 80310 66150 80380
rect 66350 80310 66650 80380
rect 66850 80310 67150 80380
rect 67350 80310 67650 80380
rect 67850 80310 68150 80380
rect 68350 80310 68650 80380
rect 68850 80310 69150 80380
rect 69350 80310 69650 80380
rect 69850 80310 70150 80380
rect 70350 80310 70650 80380
rect 70850 80310 71150 80380
rect 71350 80310 71650 80380
rect 71850 80310 72150 80380
rect 72350 80310 72650 80380
rect 72850 80310 73150 80380
rect 73350 80310 73650 80380
rect 73850 80310 74150 80380
rect 74350 80310 74650 80380
rect 74850 80310 75150 80380
rect 75350 80310 75650 80380
rect 75850 80310 76150 80380
rect 76350 80310 76650 80380
rect 76850 80310 77150 80380
rect 77350 80310 77650 80380
rect 77850 80310 78150 80380
rect 78350 80310 78650 80380
rect 78850 80310 79150 80380
rect 79350 80310 79650 80380
rect 79850 80310 80150 80380
rect 80350 80310 80650 80380
rect 80850 80310 81150 80380
rect 81350 80310 81650 80380
rect 81850 80310 82150 80380
rect 82350 80310 82650 80380
rect 82850 80310 83150 80380
rect 83350 80310 83650 80380
rect 83850 80310 84150 80380
rect 84350 80310 84650 80380
rect 84850 80310 85150 80380
rect 85350 80310 85650 80380
rect 85850 80310 86150 80380
rect 86350 80310 86650 80380
rect 86850 80310 87150 80380
rect 87350 80310 87650 80380
rect 87850 80310 88150 80380
rect 88350 80310 88650 80380
rect 88850 80310 89150 80380
rect 89350 80310 89650 80380
rect 89850 80310 90150 80380
rect 90350 80310 90650 80380
rect 90850 80310 91150 80380
rect 91350 80310 91650 80380
rect 91850 80310 92150 80380
rect 92350 80310 92650 80380
rect 92850 80310 93150 80380
rect 93350 80310 93650 80380
rect 93850 80310 94150 80380
rect 94350 80310 94650 80380
rect 94850 80310 95150 80380
rect 95350 80310 95650 80380
rect 95850 80310 96150 80380
rect 96350 80310 96650 80380
rect 96850 80310 97150 80380
rect 97350 80310 97650 80380
rect 97850 80310 98150 80380
rect 98350 80310 98650 80380
rect 98850 80310 99150 80380
rect 99350 80310 99650 80380
rect 99850 80310 100150 80380
rect 100350 80310 100500 80380
rect -83500 80300 100500 80310
rect -83500 80280 -83380 80300
rect -83120 80280 -82880 80300
rect -82620 80280 -82380 80300
rect -82120 80280 -81880 80300
rect -81620 80280 -81380 80300
rect -81120 80280 -80880 80300
rect -80620 80280 -80380 80300
rect -80120 80280 -79880 80300
rect -79620 80280 -79380 80300
rect -79120 80280 -78880 80300
rect -78620 80280 -78380 80300
rect -78120 80280 -77880 80300
rect -77620 80280 -77380 80300
rect -77120 80280 -76880 80300
rect -76620 80280 -76380 80300
rect -76120 80280 -75880 80300
rect -75620 80280 -75380 80300
rect -75120 80280 -74880 80300
rect -74620 80280 -74380 80300
rect -74120 80280 -73880 80300
rect -73620 80280 -73380 80300
rect -73120 80280 -72880 80300
rect -72620 80280 -72380 80300
rect -72120 80280 -71880 80300
rect -71620 80280 -71380 80300
rect -71120 80280 -70880 80300
rect -70620 80280 -70380 80300
rect -70120 80280 -69880 80300
rect -69620 80280 -69380 80300
rect -69120 80280 -68880 80300
rect -68620 80280 -68380 80300
rect -68120 80280 -67880 80300
rect -67620 80280 -67380 80300
rect -67120 80280 -66880 80300
rect -66620 80280 -66380 80300
rect -66120 80280 -65880 80300
rect -65620 80280 -65380 80300
rect -65120 80280 -64880 80300
rect -64620 80280 -64380 80300
rect -64120 80280 -63880 80300
rect -63620 80280 -63380 80300
rect -63120 80280 -62880 80300
rect -62620 80280 -62380 80300
rect -62120 80280 -61880 80300
rect -61620 80280 -61380 80300
rect -61120 80280 -60880 80300
rect -60620 80280 -60380 80300
rect -60120 80280 -59880 80300
rect -59620 80280 -59380 80300
rect -59120 80280 -58880 80300
rect -58620 80280 -58380 80300
rect -58120 80280 -57880 80300
rect -57620 80280 -57380 80300
rect -57120 80280 -56880 80300
rect -56620 80280 -56380 80300
rect -56120 80280 -55880 80300
rect -55620 80280 -55380 80300
rect -55120 80280 -54880 80300
rect -54620 80280 -54380 80300
rect -54120 80280 -53880 80300
rect -53620 80280 -53380 80300
rect -53120 80280 -52880 80300
rect -52620 80280 -52380 80300
rect -52120 80280 -51880 80300
rect -51620 80280 -51380 80300
rect -51120 80280 -50880 80300
rect -50620 80280 -50380 80300
rect -50120 80280 -49880 80300
rect -49620 80280 -49380 80300
rect -49120 80280 -48880 80300
rect -48620 80280 -48380 80300
rect -48120 80280 -47880 80300
rect -47620 80280 -47380 80300
rect -47120 80280 -46880 80300
rect -46620 80280 -46380 80300
rect -46120 80280 -45880 80300
rect -45620 80280 -45380 80300
rect -45120 80280 -44880 80300
rect -44620 80280 -44380 80300
rect -44120 80280 -43880 80300
rect -43620 80280 -43380 80300
rect -43120 80280 -42880 80300
rect -42620 80280 -42380 80300
rect -42120 80280 -41880 80300
rect -41620 80280 -41380 80300
rect -41120 80280 -40880 80300
rect -40620 80280 -40380 80300
rect -40120 80280 -39880 80300
rect -39620 80280 -39380 80300
rect -39120 80280 -38880 80300
rect -38620 80280 -38380 80300
rect -38120 80280 -37880 80300
rect -37620 80280 -37380 80300
rect -37120 80280 -36880 80300
rect -36620 80280 -36380 80300
rect -36120 80280 -35880 80300
rect -35620 80280 -35380 80300
rect -35120 80280 -34880 80300
rect -34620 80280 -34380 80300
rect -34120 80280 -33880 80300
rect -33620 80280 -33380 80300
rect -33120 80280 -32880 80300
rect -32620 80280 -32380 80300
rect -32120 80280 -31880 80300
rect -31620 80280 -31380 80300
rect -31120 80280 -30880 80300
rect -30620 80280 -30380 80300
rect -30120 80280 -29880 80300
rect -29620 80280 -29380 80300
rect -29120 80280 -28880 80300
rect -28620 80280 -28380 80300
rect -28120 80280 -27880 80300
rect -27620 80280 -27380 80300
rect -27120 80280 -26880 80300
rect -26620 80280 -26380 80300
rect -26120 80280 -25880 80300
rect -25620 80280 -25380 80300
rect -25120 80280 -24880 80300
rect -24620 80280 -24380 80300
rect -24120 80280 -23880 80300
rect -23620 80280 -23380 80300
rect -23120 80280 -22880 80300
rect -22620 80280 -22380 80300
rect -22120 80280 -21880 80300
rect -21620 80280 -21380 80300
rect -21120 80280 -20880 80300
rect -20620 80280 -20380 80300
rect -20120 80280 -19880 80300
rect -19620 80280 -19380 80300
rect -19120 80280 -18880 80300
rect -18620 80280 -18380 80300
rect -18120 80280 -17880 80300
rect -17620 80280 -17380 80300
rect -17120 80280 -16880 80300
rect -16620 80280 -16380 80300
rect -16120 80280 -15880 80300
rect -15620 80280 -15380 80300
rect -15120 80280 -14880 80300
rect -14620 80280 -14380 80300
rect -14120 80280 -13880 80300
rect -13620 80280 -13380 80300
rect -13120 80280 -12880 80300
rect -12620 80280 -12380 80300
rect -12120 80280 -11880 80300
rect -11620 80280 -11380 80300
rect -11120 80280 -10880 80300
rect -10620 80280 -10380 80300
rect -10120 80280 -9880 80300
rect -9620 80280 -9380 80300
rect -9120 80280 -8880 80300
rect -8620 80280 -8380 80300
rect -8120 80280 -7880 80300
rect -7620 80280 -7380 80300
rect -7120 80280 -6880 80300
rect -6620 80280 -6380 80300
rect -6120 80280 -5880 80300
rect -5620 80280 -5380 80300
rect -5120 80280 -4880 80300
rect -4620 80280 -4380 80300
rect -4120 80280 -3880 80300
rect -3620 80280 -3380 80300
rect -3120 80280 -2880 80300
rect -2620 80280 -2380 80300
rect -2120 80280 -1880 80300
rect -1620 80280 -1380 80300
rect -1120 80280 -880 80300
rect -620 80280 -380 80300
rect -120 80280 120 80300
rect 380 80280 620 80300
rect 880 80280 1120 80300
rect 1380 80280 1620 80300
rect 1880 80280 2120 80300
rect 2380 80280 2620 80300
rect 2880 80280 3120 80300
rect 3380 80280 3620 80300
rect 3880 80280 4120 80300
rect 4380 80280 4620 80300
rect 4880 80280 5120 80300
rect 5380 80280 5620 80300
rect 5880 80280 6120 80300
rect 6380 80280 6620 80300
rect 6880 80280 7120 80300
rect 7380 80280 7620 80300
rect 7880 80280 8120 80300
rect 8380 80280 8620 80300
rect 8880 80280 9120 80300
rect 9380 80280 9620 80300
rect 9880 80280 10120 80300
rect 10380 80280 10620 80300
rect 10880 80280 11120 80300
rect 11380 80280 11620 80300
rect 11880 80280 12120 80300
rect 12380 80280 12620 80300
rect 12880 80280 13120 80300
rect 13380 80280 13620 80300
rect 13880 80280 14120 80300
rect 14380 80280 14620 80300
rect 14880 80280 15120 80300
rect 15380 80280 15620 80300
rect 15880 80280 16120 80300
rect 16380 80280 16620 80300
rect 16880 80280 17120 80300
rect 17380 80280 17620 80300
rect 17880 80280 18120 80300
rect 18380 80280 18620 80300
rect 18880 80280 19120 80300
rect 19380 80280 19620 80300
rect 19880 80280 20120 80300
rect 20380 80280 20620 80300
rect 20880 80280 21120 80300
rect 21380 80280 21620 80300
rect 21880 80280 22120 80300
rect 22380 80280 22620 80300
rect 22880 80280 23120 80300
rect 23380 80280 23620 80300
rect 23880 80280 24120 80300
rect 24380 80280 24620 80300
rect 24880 80280 25120 80300
rect 25380 80280 25620 80300
rect 25880 80280 26120 80300
rect 26380 80280 26620 80300
rect 26880 80280 27120 80300
rect 27380 80280 27620 80300
rect 27880 80280 28120 80300
rect 28380 80280 28620 80300
rect 28880 80280 29120 80300
rect 29380 80280 29620 80300
rect 29880 80280 30120 80300
rect 30380 80280 30620 80300
rect 30880 80280 31120 80300
rect 31380 80280 31620 80300
rect 31880 80280 32120 80300
rect 32380 80280 32620 80300
rect 32880 80280 33120 80300
rect 33380 80280 33620 80300
rect 33880 80280 34120 80300
rect 34380 80280 34620 80300
rect 34880 80280 35120 80300
rect 35380 80280 35620 80300
rect 35880 80280 36120 80300
rect 36380 80280 36620 80300
rect 36880 80280 37120 80300
rect 37380 80280 37620 80300
rect 37880 80280 38120 80300
rect 38380 80280 38620 80300
rect 38880 80280 39120 80300
rect 39380 80280 39620 80300
rect 39880 80280 40120 80300
rect 40380 80280 40620 80300
rect 40880 80280 41120 80300
rect 41380 80280 41620 80300
rect 41880 80280 42120 80300
rect 42380 80280 42620 80300
rect 42880 80280 43120 80300
rect 43380 80280 43620 80300
rect 43880 80280 44120 80300
rect 44380 80280 44620 80300
rect 44880 80280 45120 80300
rect 45380 80280 45620 80300
rect 45880 80280 46120 80300
rect 46380 80280 46620 80300
rect 46880 80280 47120 80300
rect 47380 80280 47620 80300
rect 47880 80280 48120 80300
rect 48380 80280 48620 80300
rect 48880 80280 49120 80300
rect 49380 80280 49620 80300
rect 49880 80280 50120 80300
rect 50380 80280 50620 80300
rect 50880 80280 51120 80300
rect 51380 80280 51620 80300
rect 51880 80280 52120 80300
rect 52380 80280 52620 80300
rect 52880 80280 53120 80300
rect 53380 80280 53620 80300
rect 53880 80280 54120 80300
rect 54380 80280 54620 80300
rect 54880 80280 55120 80300
rect 55380 80280 55620 80300
rect 55880 80280 56120 80300
rect 56380 80280 56620 80300
rect 56880 80280 57120 80300
rect 57380 80280 57620 80300
rect 57880 80280 58120 80300
rect 58380 80280 58620 80300
rect 58880 80280 59120 80300
rect 59380 80280 59620 80300
rect 59880 80280 60120 80300
rect 60380 80280 60620 80300
rect 60880 80280 61120 80300
rect 61380 80280 61620 80300
rect 61880 80280 62120 80300
rect 62380 80280 62620 80300
rect 62880 80280 63120 80300
rect 63380 80280 63620 80300
rect 63880 80280 64120 80300
rect 64380 80280 64620 80300
rect 64880 80280 65120 80300
rect 65380 80280 65620 80300
rect 65880 80280 66120 80300
rect 66380 80280 66620 80300
rect 66880 80280 67120 80300
rect 67380 80280 67620 80300
rect 67880 80280 68120 80300
rect 68380 80280 68620 80300
rect 68880 80280 69120 80300
rect 69380 80280 69620 80300
rect 69880 80280 70120 80300
rect 70380 80280 70620 80300
rect 70880 80280 71120 80300
rect 71380 80280 71620 80300
rect 71880 80280 72120 80300
rect 72380 80280 72620 80300
rect 72880 80280 73120 80300
rect 73380 80280 73620 80300
rect 73880 80280 74120 80300
rect 74380 80280 74620 80300
rect 74880 80280 75120 80300
rect 75380 80280 75620 80300
rect 75880 80280 76120 80300
rect 76380 80280 76620 80300
rect 76880 80280 77120 80300
rect 77380 80280 77620 80300
rect 77880 80280 78120 80300
rect 78380 80280 78620 80300
rect 78880 80280 79120 80300
rect 79380 80280 79620 80300
rect 79880 80280 80120 80300
rect 80380 80280 80620 80300
rect 80880 80280 81120 80300
rect 81380 80280 81620 80300
rect 81880 80280 82120 80300
rect 82380 80280 82620 80300
rect 82880 80280 83120 80300
rect 83380 80280 83620 80300
rect 83880 80280 84120 80300
rect 84380 80280 84620 80300
rect 84880 80280 85120 80300
rect 85380 80280 85620 80300
rect 85880 80280 86120 80300
rect 86380 80280 86620 80300
rect 86880 80280 87120 80300
rect 87380 80280 87620 80300
rect 87880 80280 88120 80300
rect 88380 80280 88620 80300
rect 88880 80280 89120 80300
rect 89380 80280 89620 80300
rect 89880 80280 90120 80300
rect 90380 80280 90620 80300
rect 90880 80280 91120 80300
rect 91380 80280 91620 80300
rect 91880 80280 92120 80300
rect 92380 80280 92620 80300
rect 92880 80280 93120 80300
rect 93380 80280 93620 80300
rect 93880 80280 94120 80300
rect 94380 80280 94620 80300
rect 94880 80280 95120 80300
rect 95380 80280 95620 80300
rect 95880 80280 96120 80300
rect 96380 80280 96620 80300
rect 96880 80280 97120 80300
rect 97380 80280 97620 80300
rect 97880 80280 98120 80300
rect 98380 80280 98620 80300
rect 98880 80280 99120 80300
rect 99380 80280 99620 80300
rect 99880 80280 100120 80300
rect 100380 80280 100500 80300
rect -83500 80250 -83400 80280
rect -83500 80050 -83480 80250
rect -83410 80050 -83400 80250
rect -83500 80020 -83400 80050
rect -83100 80250 -82900 80280
rect -83100 80050 -83090 80250
rect -83020 80050 -82980 80250
rect -82910 80050 -82900 80250
rect -83100 80020 -82900 80050
rect -82600 80250 -82400 80280
rect -82600 80050 -82590 80250
rect -82520 80050 -82480 80250
rect -82410 80050 -82400 80250
rect -82600 80020 -82400 80050
rect -82100 80250 -81900 80280
rect -82100 80050 -82090 80250
rect -82020 80050 -81980 80250
rect -81910 80050 -81900 80250
rect -82100 80020 -81900 80050
rect -81600 80250 -81400 80280
rect -81600 80050 -81590 80250
rect -81520 80050 -81480 80250
rect -81410 80050 -81400 80250
rect -81600 80020 -81400 80050
rect -81100 80250 -80900 80280
rect -81100 80050 -81090 80250
rect -81020 80050 -80980 80250
rect -80910 80050 -80900 80250
rect -81100 80020 -80900 80050
rect -80600 80250 -80400 80280
rect -80600 80050 -80590 80250
rect -80520 80050 -80480 80250
rect -80410 80050 -80400 80250
rect -80600 80020 -80400 80050
rect -80100 80250 -79900 80280
rect -80100 80050 -80090 80250
rect -80020 80050 -79980 80250
rect -79910 80050 -79900 80250
rect -80100 80020 -79900 80050
rect -79600 80250 -79400 80280
rect -79600 80050 -79590 80250
rect -79520 80050 -79480 80250
rect -79410 80050 -79400 80250
rect -79600 80020 -79400 80050
rect -79100 80250 -78900 80280
rect -79100 80050 -79090 80250
rect -79020 80050 -78980 80250
rect -78910 80050 -78900 80250
rect -79100 80020 -78900 80050
rect -78600 80250 -78400 80280
rect -78600 80050 -78590 80250
rect -78520 80050 -78480 80250
rect -78410 80050 -78400 80250
rect -78600 80020 -78400 80050
rect -78100 80250 -77900 80280
rect -78100 80050 -78090 80250
rect -78020 80050 -77980 80250
rect -77910 80050 -77900 80250
rect -78100 80020 -77900 80050
rect -77600 80250 -77400 80280
rect -77600 80050 -77590 80250
rect -77520 80050 -77480 80250
rect -77410 80050 -77400 80250
rect -77600 80020 -77400 80050
rect -77100 80250 -76900 80280
rect -77100 80050 -77090 80250
rect -77020 80050 -76980 80250
rect -76910 80050 -76900 80250
rect -77100 80020 -76900 80050
rect -76600 80250 -76400 80280
rect -76600 80050 -76590 80250
rect -76520 80050 -76480 80250
rect -76410 80050 -76400 80250
rect -76600 80020 -76400 80050
rect -76100 80250 -75900 80280
rect -76100 80050 -76090 80250
rect -76020 80050 -75980 80250
rect -75910 80050 -75900 80250
rect -76100 80020 -75900 80050
rect -75600 80250 -75400 80280
rect -75600 80050 -75590 80250
rect -75520 80050 -75480 80250
rect -75410 80050 -75400 80250
rect -75600 80020 -75400 80050
rect -75100 80250 -74900 80280
rect -75100 80050 -75090 80250
rect -75020 80050 -74980 80250
rect -74910 80050 -74900 80250
rect -75100 80020 -74900 80050
rect -74600 80250 -74400 80280
rect -74600 80050 -74590 80250
rect -74520 80050 -74480 80250
rect -74410 80050 -74400 80250
rect -74600 80020 -74400 80050
rect -74100 80250 -73900 80280
rect -74100 80050 -74090 80250
rect -74020 80050 -73980 80250
rect -73910 80050 -73900 80250
rect -74100 80020 -73900 80050
rect -73600 80250 -73400 80280
rect -73600 80050 -73590 80250
rect -73520 80050 -73480 80250
rect -73410 80050 -73400 80250
rect -73600 80020 -73400 80050
rect -73100 80250 -72900 80280
rect -73100 80050 -73090 80250
rect -73020 80050 -72980 80250
rect -72910 80050 -72900 80250
rect -73100 80020 -72900 80050
rect -72600 80250 -72400 80280
rect -72600 80050 -72590 80250
rect -72520 80050 -72480 80250
rect -72410 80050 -72400 80250
rect -72600 80020 -72400 80050
rect -72100 80250 -71900 80280
rect -72100 80050 -72090 80250
rect -72020 80050 -71980 80250
rect -71910 80050 -71900 80250
rect -72100 80020 -71900 80050
rect -71600 80250 -71400 80280
rect -71600 80050 -71590 80250
rect -71520 80050 -71480 80250
rect -71410 80050 -71400 80250
rect -71600 80020 -71400 80050
rect -71100 80250 -70900 80280
rect -71100 80050 -71090 80250
rect -71020 80050 -70980 80250
rect -70910 80050 -70900 80250
rect -71100 80020 -70900 80050
rect -70600 80250 -70400 80280
rect -70600 80050 -70590 80250
rect -70520 80050 -70480 80250
rect -70410 80050 -70400 80250
rect -70600 80020 -70400 80050
rect -70100 80250 -69900 80280
rect -70100 80050 -70090 80250
rect -70020 80050 -69980 80250
rect -69910 80050 -69900 80250
rect -70100 80020 -69900 80050
rect -69600 80250 -69400 80280
rect -69600 80050 -69590 80250
rect -69520 80050 -69480 80250
rect -69410 80050 -69400 80250
rect -69600 80020 -69400 80050
rect -69100 80250 -68900 80280
rect -69100 80050 -69090 80250
rect -69020 80050 -68980 80250
rect -68910 80050 -68900 80250
rect -69100 80020 -68900 80050
rect -68600 80250 -68400 80280
rect -68600 80050 -68590 80250
rect -68520 80050 -68480 80250
rect -68410 80050 -68400 80250
rect -68600 80020 -68400 80050
rect -68100 80250 -67900 80280
rect -68100 80050 -68090 80250
rect -68020 80050 -67980 80250
rect -67910 80050 -67900 80250
rect -68100 80020 -67900 80050
rect -67600 80250 -67400 80280
rect -67600 80050 -67590 80250
rect -67520 80050 -67480 80250
rect -67410 80050 -67400 80250
rect -67600 80020 -67400 80050
rect -67100 80250 -66900 80280
rect -67100 80050 -67090 80250
rect -67020 80050 -66980 80250
rect -66910 80050 -66900 80250
rect -67100 80020 -66900 80050
rect -66600 80250 -66400 80280
rect -66600 80050 -66590 80250
rect -66520 80050 -66480 80250
rect -66410 80050 -66400 80250
rect -66600 80020 -66400 80050
rect -66100 80250 -65900 80280
rect -66100 80050 -66090 80250
rect -66020 80050 -65980 80250
rect -65910 80050 -65900 80250
rect -66100 80020 -65900 80050
rect -65600 80250 -65400 80280
rect -65600 80050 -65590 80250
rect -65520 80050 -65480 80250
rect -65410 80050 -65400 80250
rect -65600 80020 -65400 80050
rect -65100 80250 -64900 80280
rect -65100 80050 -65090 80250
rect -65020 80050 -64980 80250
rect -64910 80050 -64900 80250
rect -65100 80020 -64900 80050
rect -64600 80250 -64400 80280
rect -64600 80050 -64590 80250
rect -64520 80050 -64480 80250
rect -64410 80050 -64400 80250
rect -64600 80020 -64400 80050
rect -64100 80250 -63900 80280
rect -64100 80050 -64090 80250
rect -64020 80050 -63980 80250
rect -63910 80050 -63900 80250
rect -64100 80020 -63900 80050
rect -63600 80250 -63400 80280
rect -63600 80050 -63590 80250
rect -63520 80050 -63480 80250
rect -63410 80050 -63400 80250
rect -63600 80020 -63400 80050
rect -63100 80250 -62900 80280
rect -63100 80050 -63090 80250
rect -63020 80050 -62980 80250
rect -62910 80050 -62900 80250
rect -63100 80020 -62900 80050
rect -62600 80250 -62400 80280
rect -62600 80050 -62590 80250
rect -62520 80050 -62480 80250
rect -62410 80050 -62400 80250
rect -62600 80020 -62400 80050
rect -62100 80250 -61900 80280
rect -62100 80050 -62090 80250
rect -62020 80050 -61980 80250
rect -61910 80050 -61900 80250
rect -62100 80020 -61900 80050
rect -61600 80250 -61400 80280
rect -61600 80050 -61590 80250
rect -61520 80050 -61480 80250
rect -61410 80050 -61400 80250
rect -61600 80020 -61400 80050
rect -61100 80250 -60900 80280
rect -61100 80050 -61090 80250
rect -61020 80050 -60980 80250
rect -60910 80050 -60900 80250
rect -61100 80020 -60900 80050
rect -60600 80250 -60400 80280
rect -60600 80050 -60590 80250
rect -60520 80050 -60480 80250
rect -60410 80050 -60400 80250
rect -60600 80020 -60400 80050
rect -60100 80250 -59900 80280
rect -60100 80050 -60090 80250
rect -60020 80050 -59980 80250
rect -59910 80050 -59900 80250
rect -60100 80020 -59900 80050
rect -59600 80250 -59400 80280
rect -59600 80050 -59590 80250
rect -59520 80050 -59480 80250
rect -59410 80050 -59400 80250
rect -59600 80020 -59400 80050
rect -59100 80250 -58900 80280
rect -59100 80050 -59090 80250
rect -59020 80050 -58980 80250
rect -58910 80050 -58900 80250
rect -59100 80020 -58900 80050
rect -58600 80250 -58400 80280
rect -58600 80050 -58590 80250
rect -58520 80050 -58480 80250
rect -58410 80050 -58400 80250
rect -58600 80020 -58400 80050
rect -58100 80250 -57900 80280
rect -58100 80050 -58090 80250
rect -58020 80050 -57980 80250
rect -57910 80050 -57900 80250
rect -58100 80020 -57900 80050
rect -57600 80250 -57400 80280
rect -57600 80050 -57590 80250
rect -57520 80050 -57480 80250
rect -57410 80050 -57400 80250
rect -57600 80020 -57400 80050
rect -57100 80250 -56900 80280
rect -57100 80050 -57090 80250
rect -57020 80050 -56980 80250
rect -56910 80050 -56900 80250
rect -57100 80020 -56900 80050
rect -56600 80250 -56400 80280
rect -56600 80050 -56590 80250
rect -56520 80050 -56480 80250
rect -56410 80050 -56400 80250
rect -56600 80020 -56400 80050
rect -56100 80250 -55900 80280
rect -56100 80050 -56090 80250
rect -56020 80050 -55980 80250
rect -55910 80050 -55900 80250
rect -56100 80020 -55900 80050
rect -55600 80250 -55400 80280
rect -55600 80050 -55590 80250
rect -55520 80050 -55480 80250
rect -55410 80050 -55400 80250
rect -55600 80020 -55400 80050
rect -55100 80250 -54900 80280
rect -55100 80050 -55090 80250
rect -55020 80050 -54980 80250
rect -54910 80050 -54900 80250
rect -55100 80020 -54900 80050
rect -54600 80250 -54400 80280
rect -54600 80050 -54590 80250
rect -54520 80050 -54480 80250
rect -54410 80050 -54400 80250
rect -54600 80020 -54400 80050
rect -54100 80250 -53900 80280
rect -54100 80050 -54090 80250
rect -54020 80050 -53980 80250
rect -53910 80050 -53900 80250
rect -54100 80020 -53900 80050
rect -53600 80250 -53400 80280
rect -53600 80050 -53590 80250
rect -53520 80050 -53480 80250
rect -53410 80050 -53400 80250
rect -53600 80020 -53400 80050
rect -53100 80250 -52900 80280
rect -53100 80050 -53090 80250
rect -53020 80050 -52980 80250
rect -52910 80050 -52900 80250
rect -53100 80020 -52900 80050
rect -52600 80250 -52400 80280
rect -52600 80050 -52590 80250
rect -52520 80050 -52480 80250
rect -52410 80050 -52400 80250
rect -52600 80020 -52400 80050
rect -52100 80250 -51900 80280
rect -52100 80050 -52090 80250
rect -52020 80050 -51980 80250
rect -51910 80050 -51900 80250
rect -52100 80020 -51900 80050
rect -51600 80250 -51400 80280
rect -51600 80050 -51590 80250
rect -51520 80050 -51480 80250
rect -51410 80050 -51400 80250
rect -51600 80020 -51400 80050
rect -51100 80250 -50900 80280
rect -51100 80050 -51090 80250
rect -51020 80050 -50980 80250
rect -50910 80050 -50900 80250
rect -51100 80020 -50900 80050
rect -50600 80250 -50400 80280
rect -50600 80050 -50590 80250
rect -50520 80050 -50480 80250
rect -50410 80050 -50400 80250
rect -50600 80020 -50400 80050
rect -50100 80250 -49900 80280
rect -50100 80050 -50090 80250
rect -50020 80050 -49980 80250
rect -49910 80050 -49900 80250
rect -50100 80020 -49900 80050
rect -49600 80250 -49400 80280
rect -49600 80050 -49590 80250
rect -49520 80050 -49480 80250
rect -49410 80050 -49400 80250
rect -49600 80020 -49400 80050
rect -49100 80250 -48900 80280
rect -49100 80050 -49090 80250
rect -49020 80050 -48980 80250
rect -48910 80050 -48900 80250
rect -49100 80020 -48900 80050
rect -48600 80250 -48400 80280
rect -48600 80050 -48590 80250
rect -48520 80050 -48480 80250
rect -48410 80050 -48400 80250
rect -48600 80020 -48400 80050
rect -48100 80250 -47900 80280
rect -48100 80050 -48090 80250
rect -48020 80050 -47980 80250
rect -47910 80050 -47900 80250
rect -48100 80020 -47900 80050
rect -47600 80250 -47400 80280
rect -47600 80050 -47590 80250
rect -47520 80050 -47480 80250
rect -47410 80050 -47400 80250
rect -47600 80020 -47400 80050
rect -47100 80250 -46900 80280
rect -47100 80050 -47090 80250
rect -47020 80050 -46980 80250
rect -46910 80050 -46900 80250
rect -47100 80020 -46900 80050
rect -46600 80250 -46400 80280
rect -46600 80050 -46590 80250
rect -46520 80050 -46480 80250
rect -46410 80050 -46400 80250
rect -46600 80020 -46400 80050
rect -46100 80250 -45900 80280
rect -46100 80050 -46090 80250
rect -46020 80050 -45980 80250
rect -45910 80050 -45900 80250
rect -46100 80020 -45900 80050
rect -45600 80250 -45400 80280
rect -45600 80050 -45590 80250
rect -45520 80050 -45480 80250
rect -45410 80050 -45400 80250
rect -45600 80020 -45400 80050
rect -45100 80250 -44900 80280
rect -45100 80050 -45090 80250
rect -45020 80050 -44980 80250
rect -44910 80050 -44900 80250
rect -45100 80020 -44900 80050
rect -44600 80250 -44400 80280
rect -44600 80050 -44590 80250
rect -44520 80050 -44480 80250
rect -44410 80050 -44400 80250
rect -44600 80020 -44400 80050
rect -44100 80250 -43900 80280
rect -44100 80050 -44090 80250
rect -44020 80050 -43980 80250
rect -43910 80050 -43900 80250
rect -44100 80020 -43900 80050
rect -43600 80250 -43400 80280
rect -43600 80050 -43590 80250
rect -43520 80050 -43480 80250
rect -43410 80050 -43400 80250
rect -43600 80020 -43400 80050
rect -43100 80250 -42900 80280
rect -43100 80050 -43090 80250
rect -43020 80050 -42980 80250
rect -42910 80050 -42900 80250
rect -43100 80020 -42900 80050
rect -42600 80250 -42400 80280
rect -42600 80050 -42590 80250
rect -42520 80050 -42480 80250
rect -42410 80050 -42400 80250
rect -42600 80020 -42400 80050
rect -42100 80250 -41900 80280
rect -42100 80050 -42090 80250
rect -42020 80050 -41980 80250
rect -41910 80050 -41900 80250
rect -42100 80020 -41900 80050
rect -41600 80250 -41400 80280
rect -41600 80050 -41590 80250
rect -41520 80050 -41480 80250
rect -41410 80050 -41400 80250
rect -41600 80020 -41400 80050
rect -41100 80250 -40900 80280
rect -41100 80050 -41090 80250
rect -41020 80050 -40980 80250
rect -40910 80050 -40900 80250
rect -41100 80020 -40900 80050
rect -40600 80250 -40400 80280
rect -40600 80050 -40590 80250
rect -40520 80050 -40480 80250
rect -40410 80050 -40400 80250
rect -40600 80020 -40400 80050
rect -40100 80250 -39900 80280
rect -40100 80050 -40090 80250
rect -40020 80050 -39980 80250
rect -39910 80050 -39900 80250
rect -40100 80020 -39900 80050
rect -39600 80250 -39400 80280
rect -39600 80050 -39590 80250
rect -39520 80050 -39480 80250
rect -39410 80050 -39400 80250
rect -39600 80020 -39400 80050
rect -39100 80250 -38900 80280
rect -39100 80050 -39090 80250
rect -39020 80050 -38980 80250
rect -38910 80050 -38900 80250
rect -39100 80020 -38900 80050
rect -38600 80250 -38400 80280
rect -38600 80050 -38590 80250
rect -38520 80050 -38480 80250
rect -38410 80050 -38400 80250
rect -38600 80020 -38400 80050
rect -38100 80250 -37900 80280
rect -38100 80050 -38090 80250
rect -38020 80050 -37980 80250
rect -37910 80050 -37900 80250
rect -38100 80020 -37900 80050
rect -37600 80250 -37400 80280
rect -37600 80050 -37590 80250
rect -37520 80050 -37480 80250
rect -37410 80050 -37400 80250
rect -37600 80020 -37400 80050
rect -37100 80250 -36900 80280
rect -37100 80050 -37090 80250
rect -37020 80050 -36980 80250
rect -36910 80050 -36900 80250
rect -37100 80020 -36900 80050
rect -36600 80250 -36400 80280
rect -36600 80050 -36590 80250
rect -36520 80050 -36480 80250
rect -36410 80050 -36400 80250
rect -36600 80020 -36400 80050
rect -36100 80250 -35900 80280
rect -36100 80050 -36090 80250
rect -36020 80050 -35980 80250
rect -35910 80050 -35900 80250
rect -36100 80020 -35900 80050
rect -35600 80250 -35400 80280
rect -35600 80050 -35590 80250
rect -35520 80050 -35480 80250
rect -35410 80050 -35400 80250
rect -35600 80020 -35400 80050
rect -35100 80250 -34900 80280
rect -35100 80050 -35090 80250
rect -35020 80050 -34980 80250
rect -34910 80050 -34900 80250
rect -35100 80020 -34900 80050
rect -34600 80250 -34400 80280
rect -34600 80050 -34590 80250
rect -34520 80050 -34480 80250
rect -34410 80050 -34400 80250
rect -34600 80020 -34400 80050
rect -34100 80250 -33900 80280
rect -34100 80050 -34090 80250
rect -34020 80050 -33980 80250
rect -33910 80050 -33900 80250
rect -34100 80020 -33900 80050
rect -33600 80250 -33400 80280
rect -33600 80050 -33590 80250
rect -33520 80050 -33480 80250
rect -33410 80050 -33400 80250
rect -33600 80020 -33400 80050
rect -33100 80250 -32900 80280
rect -33100 80050 -33090 80250
rect -33020 80050 -32980 80250
rect -32910 80050 -32900 80250
rect -33100 80020 -32900 80050
rect -32600 80250 -32400 80280
rect -32600 80050 -32590 80250
rect -32520 80050 -32480 80250
rect -32410 80050 -32400 80250
rect -32600 80020 -32400 80050
rect -32100 80250 -31900 80280
rect -32100 80050 -32090 80250
rect -32020 80050 -31980 80250
rect -31910 80050 -31900 80250
rect -32100 80020 -31900 80050
rect -31600 80250 -31400 80280
rect -31600 80050 -31590 80250
rect -31520 80050 -31480 80250
rect -31410 80050 -31400 80250
rect -31600 80020 -31400 80050
rect -31100 80250 -30900 80280
rect -31100 80050 -31090 80250
rect -31020 80050 -30980 80250
rect -30910 80050 -30900 80250
rect -31100 80020 -30900 80050
rect -30600 80250 -30400 80280
rect -30600 80050 -30590 80250
rect -30520 80050 -30480 80250
rect -30410 80050 -30400 80250
rect -30600 80020 -30400 80050
rect -30100 80250 -29900 80280
rect -30100 80050 -30090 80250
rect -30020 80050 -29980 80250
rect -29910 80050 -29900 80250
rect -30100 80020 -29900 80050
rect -29600 80250 -29400 80280
rect -29600 80050 -29590 80250
rect -29520 80050 -29480 80250
rect -29410 80050 -29400 80250
rect -29600 80020 -29400 80050
rect -29100 80250 -28900 80280
rect -29100 80050 -29090 80250
rect -29020 80050 -28980 80250
rect -28910 80050 -28900 80250
rect -29100 80020 -28900 80050
rect -28600 80250 -28400 80280
rect -28600 80050 -28590 80250
rect -28520 80050 -28480 80250
rect -28410 80050 -28400 80250
rect -28600 80020 -28400 80050
rect -28100 80250 -27900 80280
rect -28100 80050 -28090 80250
rect -28020 80050 -27980 80250
rect -27910 80050 -27900 80250
rect -28100 80020 -27900 80050
rect -27600 80250 -27400 80280
rect -27600 80050 -27590 80250
rect -27520 80050 -27480 80250
rect -27410 80050 -27400 80250
rect -27600 80020 -27400 80050
rect -27100 80250 -26900 80280
rect -27100 80050 -27090 80250
rect -27020 80050 -26980 80250
rect -26910 80050 -26900 80250
rect -27100 80020 -26900 80050
rect -26600 80250 -26400 80280
rect -26600 80050 -26590 80250
rect -26520 80050 -26480 80250
rect -26410 80050 -26400 80250
rect -26600 80020 -26400 80050
rect -26100 80250 -25900 80280
rect -26100 80050 -26090 80250
rect -26020 80050 -25980 80250
rect -25910 80050 -25900 80250
rect -26100 80020 -25900 80050
rect -25600 80250 -25400 80280
rect -25600 80050 -25590 80250
rect -25520 80050 -25480 80250
rect -25410 80050 -25400 80250
rect -25600 80020 -25400 80050
rect -25100 80250 -24900 80280
rect -25100 80050 -25090 80250
rect -25020 80050 -24980 80250
rect -24910 80050 -24900 80250
rect -25100 80020 -24900 80050
rect -24600 80250 -24400 80280
rect -24600 80050 -24590 80250
rect -24520 80050 -24480 80250
rect -24410 80050 -24400 80250
rect -24600 80020 -24400 80050
rect -24100 80250 -23900 80280
rect -24100 80050 -24090 80250
rect -24020 80050 -23980 80250
rect -23910 80050 -23900 80250
rect -24100 80020 -23900 80050
rect -23600 80250 -23400 80280
rect -23600 80050 -23590 80250
rect -23520 80050 -23480 80250
rect -23410 80050 -23400 80250
rect -23600 80020 -23400 80050
rect -23100 80250 -22900 80280
rect -23100 80050 -23090 80250
rect -23020 80050 -22980 80250
rect -22910 80050 -22900 80250
rect -23100 80020 -22900 80050
rect -22600 80250 -22400 80280
rect -22600 80050 -22590 80250
rect -22520 80050 -22480 80250
rect -22410 80050 -22400 80250
rect -22600 80020 -22400 80050
rect -22100 80250 -21900 80280
rect -22100 80050 -22090 80250
rect -22020 80050 -21980 80250
rect -21910 80050 -21900 80250
rect -22100 80020 -21900 80050
rect -21600 80250 -21400 80280
rect -21600 80050 -21590 80250
rect -21520 80050 -21480 80250
rect -21410 80050 -21400 80250
rect -21600 80020 -21400 80050
rect -21100 80250 -20900 80280
rect -21100 80050 -21090 80250
rect -21020 80050 -20980 80250
rect -20910 80050 -20900 80250
rect -21100 80020 -20900 80050
rect -20600 80250 -20400 80280
rect -20600 80050 -20590 80250
rect -20520 80050 -20480 80250
rect -20410 80050 -20400 80250
rect -20600 80020 -20400 80050
rect -20100 80250 -19900 80280
rect -20100 80050 -20090 80250
rect -20020 80050 -19980 80250
rect -19910 80050 -19900 80250
rect -20100 80020 -19900 80050
rect -19600 80250 -19400 80280
rect -19600 80050 -19590 80250
rect -19520 80050 -19480 80250
rect -19410 80050 -19400 80250
rect -19600 80020 -19400 80050
rect -19100 80250 -18900 80280
rect -19100 80050 -19090 80250
rect -19020 80050 -18980 80250
rect -18910 80050 -18900 80250
rect -19100 80020 -18900 80050
rect -18600 80250 -18400 80280
rect -18600 80050 -18590 80250
rect -18520 80050 -18480 80250
rect -18410 80050 -18400 80250
rect -18600 80020 -18400 80050
rect -18100 80250 -17900 80280
rect -18100 80050 -18090 80250
rect -18020 80050 -17980 80250
rect -17910 80050 -17900 80250
rect -18100 80020 -17900 80050
rect -17600 80250 -17400 80280
rect -17600 80050 -17590 80250
rect -17520 80050 -17480 80250
rect -17410 80050 -17400 80250
rect -17600 80020 -17400 80050
rect -17100 80250 -16900 80280
rect -17100 80050 -17090 80250
rect -17020 80050 -16980 80250
rect -16910 80050 -16900 80250
rect -17100 80020 -16900 80050
rect -16600 80250 -16400 80280
rect -16600 80050 -16590 80250
rect -16520 80050 -16480 80250
rect -16410 80050 -16400 80250
rect -16600 80020 -16400 80050
rect -16100 80250 -15900 80280
rect -16100 80050 -16090 80250
rect -16020 80050 -15980 80250
rect -15910 80050 -15900 80250
rect -16100 80020 -15900 80050
rect -15600 80250 -15400 80280
rect -15600 80050 -15590 80250
rect -15520 80050 -15480 80250
rect -15410 80050 -15400 80250
rect -15600 80020 -15400 80050
rect -15100 80250 -14900 80280
rect -15100 80050 -15090 80250
rect -15020 80050 -14980 80250
rect -14910 80050 -14900 80250
rect -15100 80020 -14900 80050
rect -14600 80250 -14400 80280
rect -14600 80050 -14590 80250
rect -14520 80050 -14480 80250
rect -14410 80050 -14400 80250
rect -14600 80020 -14400 80050
rect -14100 80250 -13900 80280
rect -14100 80050 -14090 80250
rect -14020 80050 -13980 80250
rect -13910 80050 -13900 80250
rect -14100 80020 -13900 80050
rect -13600 80250 -13400 80280
rect -13600 80050 -13590 80250
rect -13520 80050 -13480 80250
rect -13410 80050 -13400 80250
rect -13600 80020 -13400 80050
rect -13100 80250 -12900 80280
rect -13100 80050 -13090 80250
rect -13020 80050 -12980 80250
rect -12910 80050 -12900 80250
rect -13100 80020 -12900 80050
rect -12600 80250 -12400 80280
rect -12600 80050 -12590 80250
rect -12520 80050 -12480 80250
rect -12410 80050 -12400 80250
rect -12600 80020 -12400 80050
rect -12100 80250 -11900 80280
rect -12100 80050 -12090 80250
rect -12020 80050 -11980 80250
rect -11910 80050 -11900 80250
rect -12100 80020 -11900 80050
rect -11600 80250 -11400 80280
rect -11600 80050 -11590 80250
rect -11520 80050 -11480 80250
rect -11410 80050 -11400 80250
rect -11600 80020 -11400 80050
rect -11100 80250 -10900 80280
rect -11100 80050 -11090 80250
rect -11020 80050 -10980 80250
rect -10910 80050 -10900 80250
rect -11100 80020 -10900 80050
rect -10600 80250 -10400 80280
rect -10600 80050 -10590 80250
rect -10520 80050 -10480 80250
rect -10410 80050 -10400 80250
rect -10600 80020 -10400 80050
rect -10100 80250 -9900 80280
rect -10100 80050 -10090 80250
rect -10020 80050 -9980 80250
rect -9910 80050 -9900 80250
rect -10100 80020 -9900 80050
rect -9600 80250 -9400 80280
rect -9600 80050 -9590 80250
rect -9520 80050 -9480 80250
rect -9410 80050 -9400 80250
rect -9600 80020 -9400 80050
rect -9100 80250 -8900 80280
rect -9100 80050 -9090 80250
rect -9020 80050 -8980 80250
rect -8910 80050 -8900 80250
rect -9100 80020 -8900 80050
rect -8600 80250 -8400 80280
rect -8600 80050 -8590 80250
rect -8520 80050 -8480 80250
rect -8410 80050 -8400 80250
rect -8600 80020 -8400 80050
rect -8100 80250 -7900 80280
rect -8100 80050 -8090 80250
rect -8020 80050 -7980 80250
rect -7910 80050 -7900 80250
rect -8100 80020 -7900 80050
rect -7600 80250 -7400 80280
rect -7600 80050 -7590 80250
rect -7520 80050 -7480 80250
rect -7410 80050 -7400 80250
rect -7600 80020 -7400 80050
rect -7100 80250 -6900 80280
rect -7100 80050 -7090 80250
rect -7020 80050 -6980 80250
rect -6910 80050 -6900 80250
rect -7100 80020 -6900 80050
rect -6600 80250 -6400 80280
rect -6600 80050 -6590 80250
rect -6520 80050 -6480 80250
rect -6410 80050 -6400 80250
rect -6600 80020 -6400 80050
rect -6100 80250 -5900 80280
rect -6100 80050 -6090 80250
rect -6020 80050 -5980 80250
rect -5910 80050 -5900 80250
rect -6100 80020 -5900 80050
rect -5600 80250 -5400 80280
rect -5600 80050 -5590 80250
rect -5520 80050 -5480 80250
rect -5410 80050 -5400 80250
rect -5600 80020 -5400 80050
rect -5100 80250 -4900 80280
rect -5100 80050 -5090 80250
rect -5020 80050 -4980 80250
rect -4910 80050 -4900 80250
rect -5100 80020 -4900 80050
rect -4600 80250 -4400 80280
rect -4600 80050 -4590 80250
rect -4520 80050 -4480 80250
rect -4410 80050 -4400 80250
rect -4600 80020 -4400 80050
rect -4100 80250 -3900 80280
rect -4100 80050 -4090 80250
rect -4020 80050 -3980 80250
rect -3910 80050 -3900 80250
rect -4100 80020 -3900 80050
rect -3600 80250 -3400 80280
rect -3600 80050 -3590 80250
rect -3520 80050 -3480 80250
rect -3410 80050 -3400 80250
rect -3600 80020 -3400 80050
rect -3100 80250 -2900 80280
rect -3100 80050 -3090 80250
rect -3020 80050 -2980 80250
rect -2910 80050 -2900 80250
rect -3100 80020 -2900 80050
rect -2600 80250 -2400 80280
rect -2600 80050 -2590 80250
rect -2520 80050 -2480 80250
rect -2410 80050 -2400 80250
rect -2600 80020 -2400 80050
rect -2100 80250 -1900 80280
rect -2100 80050 -2090 80250
rect -2020 80050 -1980 80250
rect -1910 80050 -1900 80250
rect -2100 80020 -1900 80050
rect -1600 80250 -1400 80280
rect -1600 80050 -1590 80250
rect -1520 80050 -1480 80250
rect -1410 80050 -1400 80250
rect -1600 80020 -1400 80050
rect -1100 80250 -900 80280
rect -1100 80050 -1090 80250
rect -1020 80050 -980 80250
rect -910 80050 -900 80250
rect -1100 80020 -900 80050
rect -600 80250 -400 80280
rect -600 80050 -590 80250
rect -520 80050 -480 80250
rect -410 80050 -400 80250
rect -600 80020 -400 80050
rect -100 80250 100 80280
rect -100 80050 -90 80250
rect -20 80050 20 80250
rect 90 80050 100 80250
rect -100 80020 100 80050
rect 400 80250 600 80280
rect 400 80050 410 80250
rect 480 80050 520 80250
rect 590 80050 600 80250
rect 400 80020 600 80050
rect 900 80250 1100 80280
rect 900 80050 910 80250
rect 980 80050 1020 80250
rect 1090 80050 1100 80250
rect 900 80020 1100 80050
rect 1400 80250 1600 80280
rect 1400 80050 1410 80250
rect 1480 80050 1520 80250
rect 1590 80050 1600 80250
rect 1400 80020 1600 80050
rect 1900 80250 2100 80280
rect 1900 80050 1910 80250
rect 1980 80050 2020 80250
rect 2090 80050 2100 80250
rect 1900 80020 2100 80050
rect 2400 80250 2600 80280
rect 2400 80050 2410 80250
rect 2480 80050 2520 80250
rect 2590 80050 2600 80250
rect 2400 80020 2600 80050
rect 2900 80250 3100 80280
rect 2900 80050 2910 80250
rect 2980 80050 3020 80250
rect 3090 80050 3100 80250
rect 2900 80020 3100 80050
rect 3400 80250 3600 80280
rect 3400 80050 3410 80250
rect 3480 80050 3520 80250
rect 3590 80050 3600 80250
rect 3400 80020 3600 80050
rect 3900 80250 4100 80280
rect 3900 80050 3910 80250
rect 3980 80050 4020 80250
rect 4090 80050 4100 80250
rect 3900 80020 4100 80050
rect 4400 80250 4600 80280
rect 4400 80050 4410 80250
rect 4480 80050 4520 80250
rect 4590 80050 4600 80250
rect 4400 80020 4600 80050
rect 4900 80250 5100 80280
rect 4900 80050 4910 80250
rect 4980 80050 5020 80250
rect 5090 80050 5100 80250
rect 4900 80020 5100 80050
rect 5400 80250 5600 80280
rect 5400 80050 5410 80250
rect 5480 80050 5520 80250
rect 5590 80050 5600 80250
rect 5400 80020 5600 80050
rect 5900 80250 6100 80280
rect 5900 80050 5910 80250
rect 5980 80050 6020 80250
rect 6090 80050 6100 80250
rect 5900 80020 6100 80050
rect 6400 80250 6600 80280
rect 6400 80050 6410 80250
rect 6480 80050 6520 80250
rect 6590 80050 6600 80250
rect 6400 80020 6600 80050
rect 6900 80250 7100 80280
rect 6900 80050 6910 80250
rect 6980 80050 7020 80250
rect 7090 80050 7100 80250
rect 6900 80020 7100 80050
rect 7400 80250 7600 80280
rect 7400 80050 7410 80250
rect 7480 80050 7520 80250
rect 7590 80050 7600 80250
rect 7400 80020 7600 80050
rect 7900 80250 8100 80280
rect 7900 80050 7910 80250
rect 7980 80050 8020 80250
rect 8090 80050 8100 80250
rect 7900 80020 8100 80050
rect 8400 80250 8600 80280
rect 8400 80050 8410 80250
rect 8480 80050 8520 80250
rect 8590 80050 8600 80250
rect 8400 80020 8600 80050
rect 8900 80250 9100 80280
rect 8900 80050 8910 80250
rect 8980 80050 9020 80250
rect 9090 80050 9100 80250
rect 8900 80020 9100 80050
rect 9400 80250 9600 80280
rect 9400 80050 9410 80250
rect 9480 80050 9520 80250
rect 9590 80050 9600 80250
rect 9400 80020 9600 80050
rect 9900 80250 10100 80280
rect 9900 80050 9910 80250
rect 9980 80050 10020 80250
rect 10090 80050 10100 80250
rect 9900 80020 10100 80050
rect 10400 80250 10600 80280
rect 10400 80050 10410 80250
rect 10480 80050 10520 80250
rect 10590 80050 10600 80250
rect 10400 80020 10600 80050
rect 10900 80250 11100 80280
rect 10900 80050 10910 80250
rect 10980 80050 11020 80250
rect 11090 80050 11100 80250
rect 10900 80020 11100 80050
rect 11400 80250 11600 80280
rect 11400 80050 11410 80250
rect 11480 80050 11520 80250
rect 11590 80050 11600 80250
rect 11400 80020 11600 80050
rect 11900 80250 12100 80280
rect 11900 80050 11910 80250
rect 11980 80050 12020 80250
rect 12090 80050 12100 80250
rect 11900 80020 12100 80050
rect 12400 80250 12600 80280
rect 12400 80050 12410 80250
rect 12480 80050 12520 80250
rect 12590 80050 12600 80250
rect 12400 80020 12600 80050
rect 12900 80250 13100 80280
rect 12900 80050 12910 80250
rect 12980 80050 13020 80250
rect 13090 80050 13100 80250
rect 12900 80020 13100 80050
rect 13400 80250 13600 80280
rect 13400 80050 13410 80250
rect 13480 80050 13520 80250
rect 13590 80050 13600 80250
rect 13400 80020 13600 80050
rect 13900 80250 14100 80280
rect 13900 80050 13910 80250
rect 13980 80050 14020 80250
rect 14090 80050 14100 80250
rect 13900 80020 14100 80050
rect 14400 80250 14600 80280
rect 14400 80050 14410 80250
rect 14480 80050 14520 80250
rect 14590 80050 14600 80250
rect 14400 80020 14600 80050
rect 14900 80250 15100 80280
rect 14900 80050 14910 80250
rect 14980 80050 15020 80250
rect 15090 80050 15100 80250
rect 14900 80020 15100 80050
rect 15400 80250 15600 80280
rect 15400 80050 15410 80250
rect 15480 80050 15520 80250
rect 15590 80050 15600 80250
rect 15400 80020 15600 80050
rect 15900 80250 16100 80280
rect 15900 80050 15910 80250
rect 15980 80050 16020 80250
rect 16090 80050 16100 80250
rect 15900 80020 16100 80050
rect 16400 80250 16600 80280
rect 16400 80050 16410 80250
rect 16480 80050 16520 80250
rect 16590 80050 16600 80250
rect 16400 80020 16600 80050
rect 16900 80250 17100 80280
rect 16900 80050 16910 80250
rect 16980 80050 17020 80250
rect 17090 80050 17100 80250
rect 16900 80020 17100 80050
rect 17400 80250 17600 80280
rect 17400 80050 17410 80250
rect 17480 80050 17520 80250
rect 17590 80050 17600 80250
rect 17400 80020 17600 80050
rect 17900 80250 18100 80280
rect 17900 80050 17910 80250
rect 17980 80050 18020 80250
rect 18090 80050 18100 80250
rect 17900 80020 18100 80050
rect 18400 80250 18600 80280
rect 18400 80050 18410 80250
rect 18480 80050 18520 80250
rect 18590 80050 18600 80250
rect 18400 80020 18600 80050
rect 18900 80250 19100 80280
rect 18900 80050 18910 80250
rect 18980 80050 19020 80250
rect 19090 80050 19100 80250
rect 18900 80020 19100 80050
rect 19400 80250 19600 80280
rect 19400 80050 19410 80250
rect 19480 80050 19520 80250
rect 19590 80050 19600 80250
rect 19400 80020 19600 80050
rect 19900 80250 20100 80280
rect 19900 80050 19910 80250
rect 19980 80050 20020 80250
rect 20090 80050 20100 80250
rect 19900 80020 20100 80050
rect 20400 80250 20600 80280
rect 20400 80050 20410 80250
rect 20480 80050 20520 80250
rect 20590 80050 20600 80250
rect 20400 80020 20600 80050
rect 20900 80250 21100 80280
rect 20900 80050 20910 80250
rect 20980 80050 21020 80250
rect 21090 80050 21100 80250
rect 20900 80020 21100 80050
rect 21400 80250 21600 80280
rect 21400 80050 21410 80250
rect 21480 80050 21520 80250
rect 21590 80050 21600 80250
rect 21400 80020 21600 80050
rect 21900 80250 22100 80280
rect 21900 80050 21910 80250
rect 21980 80050 22020 80250
rect 22090 80050 22100 80250
rect 21900 80020 22100 80050
rect 22400 80250 22600 80280
rect 22400 80050 22410 80250
rect 22480 80050 22520 80250
rect 22590 80050 22600 80250
rect 22400 80020 22600 80050
rect 22900 80250 23100 80280
rect 22900 80050 22910 80250
rect 22980 80050 23020 80250
rect 23090 80050 23100 80250
rect 22900 80020 23100 80050
rect 23400 80250 23600 80280
rect 23400 80050 23410 80250
rect 23480 80050 23520 80250
rect 23590 80050 23600 80250
rect 23400 80020 23600 80050
rect 23900 80250 24100 80280
rect 23900 80050 23910 80250
rect 23980 80050 24020 80250
rect 24090 80050 24100 80250
rect 23900 80020 24100 80050
rect 24400 80250 24600 80280
rect 24400 80050 24410 80250
rect 24480 80050 24520 80250
rect 24590 80050 24600 80250
rect 24400 80020 24600 80050
rect 24900 80250 25100 80280
rect 24900 80050 24910 80250
rect 24980 80050 25020 80250
rect 25090 80050 25100 80250
rect 24900 80020 25100 80050
rect 25400 80250 25600 80280
rect 25400 80050 25410 80250
rect 25480 80050 25520 80250
rect 25590 80050 25600 80250
rect 25400 80020 25600 80050
rect 25900 80250 26100 80280
rect 25900 80050 25910 80250
rect 25980 80050 26020 80250
rect 26090 80050 26100 80250
rect 25900 80020 26100 80050
rect 26400 80250 26600 80280
rect 26400 80050 26410 80250
rect 26480 80050 26520 80250
rect 26590 80050 26600 80250
rect 26400 80020 26600 80050
rect 26900 80250 27100 80280
rect 26900 80050 26910 80250
rect 26980 80050 27020 80250
rect 27090 80050 27100 80250
rect 26900 80020 27100 80050
rect 27400 80250 27600 80280
rect 27400 80050 27410 80250
rect 27480 80050 27520 80250
rect 27590 80050 27600 80250
rect 27400 80020 27600 80050
rect 27900 80250 28100 80280
rect 27900 80050 27910 80250
rect 27980 80050 28020 80250
rect 28090 80050 28100 80250
rect 27900 80020 28100 80050
rect 28400 80250 28600 80280
rect 28400 80050 28410 80250
rect 28480 80050 28520 80250
rect 28590 80050 28600 80250
rect 28400 80020 28600 80050
rect 28900 80250 29100 80280
rect 28900 80050 28910 80250
rect 28980 80050 29020 80250
rect 29090 80050 29100 80250
rect 28900 80020 29100 80050
rect 29400 80250 29600 80280
rect 29400 80050 29410 80250
rect 29480 80050 29520 80250
rect 29590 80050 29600 80250
rect 29400 80020 29600 80050
rect 29900 80250 30100 80280
rect 29900 80050 29910 80250
rect 29980 80050 30020 80250
rect 30090 80050 30100 80250
rect 29900 80020 30100 80050
rect 30400 80250 30600 80280
rect 30400 80050 30410 80250
rect 30480 80050 30520 80250
rect 30590 80050 30600 80250
rect 30400 80020 30600 80050
rect 30900 80250 31100 80280
rect 30900 80050 30910 80250
rect 30980 80050 31020 80250
rect 31090 80050 31100 80250
rect 30900 80020 31100 80050
rect 31400 80250 31600 80280
rect 31400 80050 31410 80250
rect 31480 80050 31520 80250
rect 31590 80050 31600 80250
rect 31400 80020 31600 80050
rect 31900 80250 32100 80280
rect 31900 80050 31910 80250
rect 31980 80050 32020 80250
rect 32090 80050 32100 80250
rect 31900 80020 32100 80050
rect 32400 80250 32600 80280
rect 32400 80050 32410 80250
rect 32480 80050 32520 80250
rect 32590 80050 32600 80250
rect 32400 80020 32600 80050
rect 32900 80250 33100 80280
rect 32900 80050 32910 80250
rect 32980 80050 33020 80250
rect 33090 80050 33100 80250
rect 32900 80020 33100 80050
rect 33400 80250 33600 80280
rect 33400 80050 33410 80250
rect 33480 80050 33520 80250
rect 33590 80050 33600 80250
rect 33400 80020 33600 80050
rect 33900 80250 34100 80280
rect 33900 80050 33910 80250
rect 33980 80050 34020 80250
rect 34090 80050 34100 80250
rect 33900 80020 34100 80050
rect 34400 80250 34600 80280
rect 34400 80050 34410 80250
rect 34480 80050 34520 80250
rect 34590 80050 34600 80250
rect 34400 80020 34600 80050
rect 34900 80250 35100 80280
rect 34900 80050 34910 80250
rect 34980 80050 35020 80250
rect 35090 80050 35100 80250
rect 34900 80020 35100 80050
rect 35400 80250 35600 80280
rect 35400 80050 35410 80250
rect 35480 80050 35520 80250
rect 35590 80050 35600 80250
rect 35400 80020 35600 80050
rect 35900 80250 36100 80280
rect 35900 80050 35910 80250
rect 35980 80050 36020 80250
rect 36090 80050 36100 80250
rect 35900 80020 36100 80050
rect 36400 80250 36600 80280
rect 36400 80050 36410 80250
rect 36480 80050 36520 80250
rect 36590 80050 36600 80250
rect 36400 80020 36600 80050
rect 36900 80250 37100 80280
rect 36900 80050 36910 80250
rect 36980 80050 37020 80250
rect 37090 80050 37100 80250
rect 36900 80020 37100 80050
rect 37400 80250 37600 80280
rect 37400 80050 37410 80250
rect 37480 80050 37520 80250
rect 37590 80050 37600 80250
rect 37400 80020 37600 80050
rect 37900 80250 38100 80280
rect 37900 80050 37910 80250
rect 37980 80050 38020 80250
rect 38090 80050 38100 80250
rect 37900 80020 38100 80050
rect 38400 80250 38600 80280
rect 38400 80050 38410 80250
rect 38480 80050 38520 80250
rect 38590 80050 38600 80250
rect 38400 80020 38600 80050
rect 38900 80250 39100 80280
rect 38900 80050 38910 80250
rect 38980 80050 39020 80250
rect 39090 80050 39100 80250
rect 38900 80020 39100 80050
rect 39400 80250 39600 80280
rect 39400 80050 39410 80250
rect 39480 80050 39520 80250
rect 39590 80050 39600 80250
rect 39400 80020 39600 80050
rect 39900 80250 40100 80280
rect 39900 80050 39910 80250
rect 39980 80050 40020 80250
rect 40090 80050 40100 80250
rect 39900 80020 40100 80050
rect 40400 80250 40600 80280
rect 40400 80050 40410 80250
rect 40480 80050 40520 80250
rect 40590 80050 40600 80250
rect 40400 80020 40600 80050
rect 40900 80250 41100 80280
rect 40900 80050 40910 80250
rect 40980 80050 41020 80250
rect 41090 80050 41100 80250
rect 40900 80020 41100 80050
rect 41400 80250 41600 80280
rect 41400 80050 41410 80250
rect 41480 80050 41520 80250
rect 41590 80050 41600 80250
rect 41400 80020 41600 80050
rect 41900 80250 42100 80280
rect 41900 80050 41910 80250
rect 41980 80050 42020 80250
rect 42090 80050 42100 80250
rect 41900 80020 42100 80050
rect 42400 80250 42600 80280
rect 42400 80050 42410 80250
rect 42480 80050 42520 80250
rect 42590 80050 42600 80250
rect 42400 80020 42600 80050
rect 42900 80250 43100 80280
rect 42900 80050 42910 80250
rect 42980 80050 43020 80250
rect 43090 80050 43100 80250
rect 42900 80020 43100 80050
rect 43400 80250 43600 80280
rect 43400 80050 43410 80250
rect 43480 80050 43520 80250
rect 43590 80050 43600 80250
rect 43400 80020 43600 80050
rect 43900 80250 44100 80280
rect 43900 80050 43910 80250
rect 43980 80050 44020 80250
rect 44090 80050 44100 80250
rect 43900 80020 44100 80050
rect 44400 80250 44600 80280
rect 44400 80050 44410 80250
rect 44480 80050 44520 80250
rect 44590 80050 44600 80250
rect 44400 80020 44600 80050
rect 44900 80250 45100 80280
rect 44900 80050 44910 80250
rect 44980 80050 45020 80250
rect 45090 80050 45100 80250
rect 44900 80020 45100 80050
rect 45400 80250 45600 80280
rect 45400 80050 45410 80250
rect 45480 80050 45520 80250
rect 45590 80050 45600 80250
rect 45400 80020 45600 80050
rect 45900 80250 46100 80280
rect 45900 80050 45910 80250
rect 45980 80050 46020 80250
rect 46090 80050 46100 80250
rect 45900 80020 46100 80050
rect 46400 80250 46600 80280
rect 46400 80050 46410 80250
rect 46480 80050 46520 80250
rect 46590 80050 46600 80250
rect 46400 80020 46600 80050
rect 46900 80250 47100 80280
rect 46900 80050 46910 80250
rect 46980 80050 47020 80250
rect 47090 80050 47100 80250
rect 46900 80020 47100 80050
rect 47400 80250 47600 80280
rect 47400 80050 47410 80250
rect 47480 80050 47520 80250
rect 47590 80050 47600 80250
rect 47400 80020 47600 80050
rect 47900 80250 48100 80280
rect 47900 80050 47910 80250
rect 47980 80050 48020 80250
rect 48090 80050 48100 80250
rect 47900 80020 48100 80050
rect 48400 80250 48600 80280
rect 48400 80050 48410 80250
rect 48480 80050 48520 80250
rect 48590 80050 48600 80250
rect 48400 80020 48600 80050
rect 48900 80250 49100 80280
rect 48900 80050 48910 80250
rect 48980 80050 49020 80250
rect 49090 80050 49100 80250
rect 48900 80020 49100 80050
rect 49400 80250 49600 80280
rect 49400 80050 49410 80250
rect 49480 80050 49520 80250
rect 49590 80050 49600 80250
rect 49400 80020 49600 80050
rect 49900 80250 50100 80280
rect 49900 80050 49910 80250
rect 49980 80050 50020 80250
rect 50090 80050 50100 80250
rect 49900 80020 50100 80050
rect 50400 80250 50600 80280
rect 50400 80050 50410 80250
rect 50480 80050 50520 80250
rect 50590 80050 50600 80250
rect 50400 80020 50600 80050
rect 50900 80250 51100 80280
rect 50900 80050 50910 80250
rect 50980 80050 51020 80250
rect 51090 80050 51100 80250
rect 50900 80020 51100 80050
rect 51400 80250 51600 80280
rect 51400 80050 51410 80250
rect 51480 80050 51520 80250
rect 51590 80050 51600 80250
rect 51400 80020 51600 80050
rect 51900 80250 52100 80280
rect 51900 80050 51910 80250
rect 51980 80050 52020 80250
rect 52090 80050 52100 80250
rect 51900 80020 52100 80050
rect 52400 80250 52600 80280
rect 52400 80050 52410 80250
rect 52480 80050 52520 80250
rect 52590 80050 52600 80250
rect 52400 80020 52600 80050
rect 52900 80250 53100 80280
rect 52900 80050 52910 80250
rect 52980 80050 53020 80250
rect 53090 80050 53100 80250
rect 52900 80020 53100 80050
rect 53400 80250 53600 80280
rect 53400 80050 53410 80250
rect 53480 80050 53520 80250
rect 53590 80050 53600 80250
rect 53400 80020 53600 80050
rect 53900 80250 54100 80280
rect 53900 80050 53910 80250
rect 53980 80050 54020 80250
rect 54090 80050 54100 80250
rect 53900 80020 54100 80050
rect 54400 80250 54600 80280
rect 54400 80050 54410 80250
rect 54480 80050 54520 80250
rect 54590 80050 54600 80250
rect 54400 80020 54600 80050
rect 54900 80250 55100 80280
rect 54900 80050 54910 80250
rect 54980 80050 55020 80250
rect 55090 80050 55100 80250
rect 54900 80020 55100 80050
rect 55400 80250 55600 80280
rect 55400 80050 55410 80250
rect 55480 80050 55520 80250
rect 55590 80050 55600 80250
rect 55400 80020 55600 80050
rect 55900 80250 56100 80280
rect 55900 80050 55910 80250
rect 55980 80050 56020 80250
rect 56090 80050 56100 80250
rect 55900 80020 56100 80050
rect 56400 80250 56600 80280
rect 56400 80050 56410 80250
rect 56480 80050 56520 80250
rect 56590 80050 56600 80250
rect 56400 80020 56600 80050
rect 56900 80250 57100 80280
rect 56900 80050 56910 80250
rect 56980 80050 57020 80250
rect 57090 80050 57100 80250
rect 56900 80020 57100 80050
rect 57400 80250 57600 80280
rect 57400 80050 57410 80250
rect 57480 80050 57520 80250
rect 57590 80050 57600 80250
rect 57400 80020 57600 80050
rect 57900 80250 58100 80280
rect 57900 80050 57910 80250
rect 57980 80050 58020 80250
rect 58090 80050 58100 80250
rect 57900 80020 58100 80050
rect 58400 80250 58600 80280
rect 58400 80050 58410 80250
rect 58480 80050 58520 80250
rect 58590 80050 58600 80250
rect 58400 80020 58600 80050
rect 58900 80250 59100 80280
rect 58900 80050 58910 80250
rect 58980 80050 59020 80250
rect 59090 80050 59100 80250
rect 58900 80020 59100 80050
rect 59400 80250 59600 80280
rect 59400 80050 59410 80250
rect 59480 80050 59520 80250
rect 59590 80050 59600 80250
rect 59400 80020 59600 80050
rect 59900 80250 60100 80280
rect 59900 80050 59910 80250
rect 59980 80050 60020 80250
rect 60090 80050 60100 80250
rect 59900 80020 60100 80050
rect 60400 80250 60600 80280
rect 60400 80050 60410 80250
rect 60480 80050 60520 80250
rect 60590 80050 60600 80250
rect 60400 80020 60600 80050
rect 60900 80250 61100 80280
rect 60900 80050 60910 80250
rect 60980 80050 61020 80250
rect 61090 80050 61100 80250
rect 60900 80020 61100 80050
rect 61400 80250 61600 80280
rect 61400 80050 61410 80250
rect 61480 80050 61520 80250
rect 61590 80050 61600 80250
rect 61400 80020 61600 80050
rect 61900 80250 62100 80280
rect 61900 80050 61910 80250
rect 61980 80050 62020 80250
rect 62090 80050 62100 80250
rect 61900 80020 62100 80050
rect 62400 80250 62600 80280
rect 62400 80050 62410 80250
rect 62480 80050 62520 80250
rect 62590 80050 62600 80250
rect 62400 80020 62600 80050
rect 62900 80250 63100 80280
rect 62900 80050 62910 80250
rect 62980 80050 63020 80250
rect 63090 80050 63100 80250
rect 62900 80020 63100 80050
rect 63400 80250 63600 80280
rect 63400 80050 63410 80250
rect 63480 80050 63520 80250
rect 63590 80050 63600 80250
rect 63400 80020 63600 80050
rect 63900 80250 64100 80280
rect 63900 80050 63910 80250
rect 63980 80050 64020 80250
rect 64090 80050 64100 80250
rect 63900 80020 64100 80050
rect 64400 80250 64600 80280
rect 64400 80050 64410 80250
rect 64480 80050 64520 80250
rect 64590 80050 64600 80250
rect 64400 80020 64600 80050
rect 64900 80250 65100 80280
rect 64900 80050 64910 80250
rect 64980 80050 65020 80250
rect 65090 80050 65100 80250
rect 64900 80020 65100 80050
rect 65400 80250 65600 80280
rect 65400 80050 65410 80250
rect 65480 80050 65520 80250
rect 65590 80050 65600 80250
rect 65400 80020 65600 80050
rect 65900 80250 66100 80280
rect 65900 80050 65910 80250
rect 65980 80050 66020 80250
rect 66090 80050 66100 80250
rect 65900 80020 66100 80050
rect 66400 80250 66600 80280
rect 66400 80050 66410 80250
rect 66480 80050 66520 80250
rect 66590 80050 66600 80250
rect 66400 80020 66600 80050
rect 66900 80250 67100 80280
rect 66900 80050 66910 80250
rect 66980 80050 67020 80250
rect 67090 80050 67100 80250
rect 66900 80020 67100 80050
rect 67400 80250 67600 80280
rect 67400 80050 67410 80250
rect 67480 80050 67520 80250
rect 67590 80050 67600 80250
rect 67400 80020 67600 80050
rect 67900 80250 68100 80280
rect 67900 80050 67910 80250
rect 67980 80050 68020 80250
rect 68090 80050 68100 80250
rect 67900 80020 68100 80050
rect 68400 80250 68600 80280
rect 68400 80050 68410 80250
rect 68480 80050 68520 80250
rect 68590 80050 68600 80250
rect 68400 80020 68600 80050
rect 68900 80250 69100 80280
rect 68900 80050 68910 80250
rect 68980 80050 69020 80250
rect 69090 80050 69100 80250
rect 68900 80020 69100 80050
rect 69400 80250 69600 80280
rect 69400 80050 69410 80250
rect 69480 80050 69520 80250
rect 69590 80050 69600 80250
rect 69400 80020 69600 80050
rect 69900 80250 70100 80280
rect 69900 80050 69910 80250
rect 69980 80050 70020 80250
rect 70090 80050 70100 80250
rect 69900 80020 70100 80050
rect 70400 80250 70600 80280
rect 70400 80050 70410 80250
rect 70480 80050 70520 80250
rect 70590 80050 70600 80250
rect 70400 80020 70600 80050
rect 70900 80250 71100 80280
rect 70900 80050 70910 80250
rect 70980 80050 71020 80250
rect 71090 80050 71100 80250
rect 70900 80020 71100 80050
rect 71400 80250 71600 80280
rect 71400 80050 71410 80250
rect 71480 80050 71520 80250
rect 71590 80050 71600 80250
rect 71400 80020 71600 80050
rect 71900 80250 72100 80280
rect 71900 80050 71910 80250
rect 71980 80050 72020 80250
rect 72090 80050 72100 80250
rect 71900 80020 72100 80050
rect 72400 80250 72600 80280
rect 72400 80050 72410 80250
rect 72480 80050 72520 80250
rect 72590 80050 72600 80250
rect 72400 80020 72600 80050
rect 72900 80250 73100 80280
rect 72900 80050 72910 80250
rect 72980 80050 73020 80250
rect 73090 80050 73100 80250
rect 72900 80020 73100 80050
rect 73400 80250 73600 80280
rect 73400 80050 73410 80250
rect 73480 80050 73520 80250
rect 73590 80050 73600 80250
rect 73400 80020 73600 80050
rect 73900 80250 74100 80280
rect 73900 80050 73910 80250
rect 73980 80050 74020 80250
rect 74090 80050 74100 80250
rect 73900 80020 74100 80050
rect 74400 80250 74600 80280
rect 74400 80050 74410 80250
rect 74480 80050 74520 80250
rect 74590 80050 74600 80250
rect 74400 80020 74600 80050
rect 74900 80250 75100 80280
rect 74900 80050 74910 80250
rect 74980 80050 75020 80250
rect 75090 80050 75100 80250
rect 74900 80020 75100 80050
rect 75400 80250 75600 80280
rect 75400 80050 75410 80250
rect 75480 80050 75520 80250
rect 75590 80050 75600 80250
rect 75400 80020 75600 80050
rect 75900 80250 76100 80280
rect 75900 80050 75910 80250
rect 75980 80050 76020 80250
rect 76090 80050 76100 80250
rect 75900 80020 76100 80050
rect 76400 80250 76600 80280
rect 76400 80050 76410 80250
rect 76480 80050 76520 80250
rect 76590 80050 76600 80250
rect 76400 80020 76600 80050
rect 76900 80250 77100 80280
rect 76900 80050 76910 80250
rect 76980 80050 77020 80250
rect 77090 80050 77100 80250
rect 76900 80020 77100 80050
rect 77400 80250 77600 80280
rect 77400 80050 77410 80250
rect 77480 80050 77520 80250
rect 77590 80050 77600 80250
rect 77400 80020 77600 80050
rect 77900 80250 78100 80280
rect 77900 80050 77910 80250
rect 77980 80050 78020 80250
rect 78090 80050 78100 80250
rect 77900 80020 78100 80050
rect 78400 80250 78600 80280
rect 78400 80050 78410 80250
rect 78480 80050 78520 80250
rect 78590 80050 78600 80250
rect 78400 80020 78600 80050
rect 78900 80250 79100 80280
rect 78900 80050 78910 80250
rect 78980 80050 79020 80250
rect 79090 80050 79100 80250
rect 78900 80020 79100 80050
rect 79400 80250 79600 80280
rect 79400 80050 79410 80250
rect 79480 80050 79520 80250
rect 79590 80050 79600 80250
rect 79400 80020 79600 80050
rect 79900 80250 80100 80280
rect 79900 80050 79910 80250
rect 79980 80050 80020 80250
rect 80090 80050 80100 80250
rect 79900 80020 80100 80050
rect 80400 80250 80600 80280
rect 80400 80050 80410 80250
rect 80480 80050 80520 80250
rect 80590 80050 80600 80250
rect 80400 80020 80600 80050
rect 80900 80250 81100 80280
rect 80900 80050 80910 80250
rect 80980 80050 81020 80250
rect 81090 80050 81100 80250
rect 80900 80020 81100 80050
rect 81400 80250 81600 80280
rect 81400 80050 81410 80250
rect 81480 80050 81520 80250
rect 81590 80050 81600 80250
rect 81400 80020 81600 80050
rect 81900 80250 82100 80280
rect 81900 80050 81910 80250
rect 81980 80050 82020 80250
rect 82090 80050 82100 80250
rect 81900 80020 82100 80050
rect 82400 80250 82600 80280
rect 82400 80050 82410 80250
rect 82480 80050 82520 80250
rect 82590 80050 82600 80250
rect 82400 80020 82600 80050
rect 82900 80250 83100 80280
rect 82900 80050 82910 80250
rect 82980 80050 83020 80250
rect 83090 80050 83100 80250
rect 82900 80020 83100 80050
rect 83400 80250 83600 80280
rect 83400 80050 83410 80250
rect 83480 80050 83520 80250
rect 83590 80050 83600 80250
rect 83400 80020 83600 80050
rect 83900 80250 84100 80280
rect 83900 80050 83910 80250
rect 83980 80050 84020 80250
rect 84090 80050 84100 80250
rect 83900 80020 84100 80050
rect 84400 80250 84600 80280
rect 84400 80050 84410 80250
rect 84480 80050 84520 80250
rect 84590 80050 84600 80250
rect 84400 80020 84600 80050
rect 84900 80250 85100 80280
rect 84900 80050 84910 80250
rect 84980 80050 85020 80250
rect 85090 80050 85100 80250
rect 84900 80020 85100 80050
rect 85400 80250 85600 80280
rect 85400 80050 85410 80250
rect 85480 80050 85520 80250
rect 85590 80050 85600 80250
rect 85400 80020 85600 80050
rect 85900 80250 86100 80280
rect 85900 80050 85910 80250
rect 85980 80050 86020 80250
rect 86090 80050 86100 80250
rect 85900 80020 86100 80050
rect 86400 80250 86600 80280
rect 86400 80050 86410 80250
rect 86480 80050 86520 80250
rect 86590 80050 86600 80250
rect 86400 80020 86600 80050
rect 86900 80250 87100 80280
rect 86900 80050 86910 80250
rect 86980 80050 87020 80250
rect 87090 80050 87100 80250
rect 86900 80020 87100 80050
rect 87400 80250 87600 80280
rect 87400 80050 87410 80250
rect 87480 80050 87520 80250
rect 87590 80050 87600 80250
rect 87400 80020 87600 80050
rect 87900 80250 88100 80280
rect 87900 80050 87910 80250
rect 87980 80050 88020 80250
rect 88090 80050 88100 80250
rect 87900 80020 88100 80050
rect 88400 80250 88600 80280
rect 88400 80050 88410 80250
rect 88480 80050 88520 80250
rect 88590 80050 88600 80250
rect 88400 80020 88600 80050
rect 88900 80250 89100 80280
rect 88900 80050 88910 80250
rect 88980 80050 89020 80250
rect 89090 80050 89100 80250
rect 88900 80020 89100 80050
rect 89400 80250 89600 80280
rect 89400 80050 89410 80250
rect 89480 80050 89520 80250
rect 89590 80050 89600 80250
rect 89400 80020 89600 80050
rect 89900 80250 90100 80280
rect 89900 80050 89910 80250
rect 89980 80050 90020 80250
rect 90090 80050 90100 80250
rect 89900 80020 90100 80050
rect 90400 80250 90600 80280
rect 90400 80050 90410 80250
rect 90480 80050 90520 80250
rect 90590 80050 90600 80250
rect 90400 80020 90600 80050
rect 90900 80250 91100 80280
rect 90900 80050 90910 80250
rect 90980 80050 91020 80250
rect 91090 80050 91100 80250
rect 90900 80020 91100 80050
rect 91400 80250 91600 80280
rect 91400 80050 91410 80250
rect 91480 80050 91520 80250
rect 91590 80050 91600 80250
rect 91400 80020 91600 80050
rect 91900 80250 92100 80280
rect 91900 80050 91910 80250
rect 91980 80050 92020 80250
rect 92090 80050 92100 80250
rect 91900 80020 92100 80050
rect 92400 80250 92600 80280
rect 92400 80050 92410 80250
rect 92480 80050 92520 80250
rect 92590 80050 92600 80250
rect 92400 80020 92600 80050
rect 92900 80250 93100 80280
rect 92900 80050 92910 80250
rect 92980 80050 93020 80250
rect 93090 80050 93100 80250
rect 92900 80020 93100 80050
rect 93400 80250 93600 80280
rect 93400 80050 93410 80250
rect 93480 80050 93520 80250
rect 93590 80050 93600 80250
rect 93400 80020 93600 80050
rect 93900 80250 94100 80280
rect 93900 80050 93910 80250
rect 93980 80050 94020 80250
rect 94090 80050 94100 80250
rect 93900 80020 94100 80050
rect 94400 80250 94600 80280
rect 94400 80050 94410 80250
rect 94480 80050 94520 80250
rect 94590 80050 94600 80250
rect 94400 80020 94600 80050
rect 94900 80250 95100 80280
rect 94900 80050 94910 80250
rect 94980 80050 95020 80250
rect 95090 80050 95100 80250
rect 94900 80020 95100 80050
rect 95400 80250 95600 80280
rect 95400 80050 95410 80250
rect 95480 80050 95520 80250
rect 95590 80050 95600 80250
rect 95400 80020 95600 80050
rect 95900 80250 96100 80280
rect 95900 80050 95910 80250
rect 95980 80050 96020 80250
rect 96090 80050 96100 80250
rect 95900 80020 96100 80050
rect 96400 80250 96600 80280
rect 96400 80050 96410 80250
rect 96480 80050 96520 80250
rect 96590 80050 96600 80250
rect 96400 80020 96600 80050
rect 96900 80250 97100 80280
rect 96900 80050 96910 80250
rect 96980 80050 97020 80250
rect 97090 80050 97100 80250
rect 96900 80020 97100 80050
rect 97400 80250 97600 80280
rect 97400 80050 97410 80250
rect 97480 80050 97520 80250
rect 97590 80050 97600 80250
rect 97400 80020 97600 80050
rect 97900 80250 98100 80280
rect 97900 80050 97910 80250
rect 97980 80050 98020 80250
rect 98090 80050 98100 80250
rect 97900 80020 98100 80050
rect 98400 80250 98600 80280
rect 98400 80050 98410 80250
rect 98480 80050 98520 80250
rect 98590 80050 98600 80250
rect 98400 80020 98600 80050
rect 98900 80250 99100 80280
rect 98900 80050 98910 80250
rect 98980 80050 99020 80250
rect 99090 80050 99100 80250
rect 98900 80020 99100 80050
rect 99400 80250 99600 80280
rect 99400 80050 99410 80250
rect 99480 80050 99520 80250
rect 99590 80050 99600 80250
rect 99400 80020 99600 80050
rect 99900 80250 100100 80280
rect 99900 80050 99910 80250
rect 99980 80050 100020 80250
rect 100090 80050 100100 80250
rect 99900 80020 100100 80050
rect 100400 80250 100500 80280
rect 100400 80050 100410 80250
rect 100480 80050 100500 80250
rect 100400 80020 100500 80050
rect -83500 80000 -83380 80020
rect -83120 80000 -82880 80020
rect -82620 80000 -82380 80020
rect -82120 80000 -81880 80020
rect -81620 80000 -81380 80020
rect -81120 80000 -80880 80020
rect -80620 80000 -80380 80020
rect -80120 80000 -79880 80020
rect -79620 80000 -79380 80020
rect -79120 80000 -78880 80020
rect -78620 80000 -78380 80020
rect -78120 80000 -77880 80020
rect -77620 80000 -77380 80020
rect -77120 80000 -76880 80020
rect -76620 80000 -76380 80020
rect -76120 80000 -75880 80020
rect -75620 80000 -75380 80020
rect -75120 80000 -74880 80020
rect -74620 80000 -74380 80020
rect -74120 80000 -73880 80020
rect -73620 80000 -73380 80020
rect -73120 80000 -72880 80020
rect -72620 80000 -72380 80020
rect -72120 80000 -71880 80020
rect -71620 80000 -71380 80020
rect -71120 80000 -70880 80020
rect -70620 80000 -70380 80020
rect -70120 80000 -69880 80020
rect -69620 80000 -69380 80020
rect -69120 80000 -68880 80020
rect -68620 80000 -68380 80020
rect -68120 80000 -67880 80020
rect -67620 80000 -67380 80020
rect -67120 80000 -66880 80020
rect -66620 80000 -66380 80020
rect -66120 80000 -65880 80020
rect -65620 80000 -65380 80020
rect -65120 80000 -64880 80020
rect -64620 80000 -64380 80020
rect -64120 80000 -63880 80020
rect -63620 80000 -63380 80020
rect -63120 80000 -62880 80020
rect -62620 80000 -62380 80020
rect -62120 80000 -61880 80020
rect -61620 80000 -61380 80020
rect -61120 80000 -60880 80020
rect -60620 80000 -60380 80020
rect -60120 80000 -59880 80020
rect -59620 80000 -59380 80020
rect -59120 80000 -58880 80020
rect -58620 80000 -58380 80020
rect -58120 80000 -57880 80020
rect -57620 80000 -57380 80020
rect -57120 80000 -56880 80020
rect -56620 80000 -56380 80020
rect -56120 80000 -55880 80020
rect -55620 80000 -55380 80020
rect -55120 80000 -54880 80020
rect -54620 80000 -54380 80020
rect -54120 80000 -53880 80020
rect -53620 80000 -53380 80020
rect -53120 80000 -52880 80020
rect -52620 80000 -52380 80020
rect -52120 80000 -51880 80020
rect -51620 80000 -51380 80020
rect -51120 80000 -50880 80020
rect -50620 80000 -50380 80020
rect -50120 80000 -49880 80020
rect -49620 80000 -49380 80020
rect -49120 80000 -48880 80020
rect -48620 80000 -48380 80020
rect -48120 80000 -47880 80020
rect -47620 80000 -47380 80020
rect -47120 80000 -46880 80020
rect -46620 80000 -46380 80020
rect -46120 80000 -45880 80020
rect -45620 80000 -45380 80020
rect -45120 80000 -44880 80020
rect -44620 80000 -44380 80020
rect -44120 80000 -43880 80020
rect -43620 80000 -43380 80020
rect -43120 80000 -42880 80020
rect -42620 80000 -42380 80020
rect -42120 80000 -41880 80020
rect -41620 80000 -41380 80020
rect -41120 80000 -40880 80020
rect -40620 80000 -40380 80020
rect -40120 80000 -39880 80020
rect -39620 80000 -39380 80020
rect -39120 80000 -38880 80020
rect -38620 80000 -38380 80020
rect -38120 80000 -37880 80020
rect -37620 80000 -37380 80020
rect -37120 80000 -36880 80020
rect -36620 80000 -36380 80020
rect -36120 80000 -35880 80020
rect -35620 80000 -35380 80020
rect -35120 80000 -34880 80020
rect -34620 80000 -34380 80020
rect -34120 80000 -33880 80020
rect -33620 80000 -33380 80020
rect -33120 80000 -32880 80020
rect -32620 80000 -32380 80020
rect -32120 80000 -31880 80020
rect -31620 80000 -31380 80020
rect -31120 80000 -30880 80020
rect -30620 80000 -30380 80020
rect -30120 80000 -29880 80020
rect -29620 80000 -29380 80020
rect -29120 80000 -28880 80020
rect -28620 80000 -28380 80020
rect -28120 80000 -27880 80020
rect -27620 80000 -27380 80020
rect -27120 80000 -26880 80020
rect -26620 80000 -26380 80020
rect -26120 80000 -25880 80020
rect -25620 80000 -25380 80020
rect -25120 80000 -24880 80020
rect -24620 80000 -24380 80020
rect -24120 80000 -23880 80020
rect -23620 80000 -23380 80020
rect -23120 80000 -22880 80020
rect -22620 80000 -22380 80020
rect -22120 80000 -21880 80020
rect -21620 80000 -21380 80020
rect -21120 80000 -20880 80020
rect -20620 80000 -20380 80020
rect -20120 80000 -19880 80020
rect -19620 80000 -19380 80020
rect -19120 80000 -18880 80020
rect -18620 80000 -18380 80020
rect -18120 80000 -17880 80020
rect -17620 80000 -17380 80020
rect -17120 80000 -16880 80020
rect -16620 80000 -16380 80020
rect -16120 80000 -15880 80020
rect -15620 80000 -15380 80020
rect -15120 80000 -14880 80020
rect -14620 80000 -14380 80020
rect -14120 80000 -13880 80020
rect -13620 80000 -13380 80020
rect -13120 80000 -12880 80020
rect -12620 80000 -12380 80020
rect -12120 80000 -11880 80020
rect -11620 80000 -11380 80020
rect -11120 80000 -10880 80020
rect -10620 80000 -10380 80020
rect -10120 80000 -9880 80020
rect -9620 80000 -9380 80020
rect -9120 80000 -8880 80020
rect -8620 80000 -8380 80020
rect -8120 80000 -7880 80020
rect -7620 80000 -7380 80020
rect -7120 80000 -6880 80020
rect -6620 80000 -6380 80020
rect -6120 80000 -5880 80020
rect -5620 80000 -5380 80020
rect -5120 80000 -4880 80020
rect -4620 80000 -4380 80020
rect -4120 80000 -3880 80020
rect -3620 80000 -3380 80020
rect -3120 80000 -2880 80020
rect -2620 80000 -2380 80020
rect -2120 80000 -1880 80020
rect -1620 80000 -1380 80020
rect -1120 80000 -880 80020
rect -620 80000 -380 80020
rect -120 80000 120 80020
rect 380 80000 620 80020
rect 880 80000 1120 80020
rect 1380 80000 1620 80020
rect 1880 80000 2120 80020
rect 2380 80000 2620 80020
rect 2880 80000 3120 80020
rect 3380 80000 3620 80020
rect 3880 80000 4120 80020
rect 4380 80000 4620 80020
rect 4880 80000 5120 80020
rect 5380 80000 5620 80020
rect 5880 80000 6120 80020
rect 6380 80000 6620 80020
rect 6880 80000 7120 80020
rect 7380 80000 7620 80020
rect 7880 80000 8120 80020
rect 8380 80000 8620 80020
rect 8880 80000 9120 80020
rect 9380 80000 9620 80020
rect 9880 80000 10120 80020
rect 10380 80000 10620 80020
rect 10880 80000 11120 80020
rect 11380 80000 11620 80020
rect 11880 80000 12120 80020
rect 12380 80000 12620 80020
rect 12880 80000 13120 80020
rect 13380 80000 13620 80020
rect 13880 80000 14120 80020
rect 14380 80000 14620 80020
rect 14880 80000 15120 80020
rect 15380 80000 15620 80020
rect 15880 80000 16120 80020
rect 16380 80000 16620 80020
rect 16880 80000 17120 80020
rect 17380 80000 17620 80020
rect 17880 80000 18120 80020
rect 18380 80000 18620 80020
rect 18880 80000 19120 80020
rect 19380 80000 19620 80020
rect 19880 80000 20120 80020
rect 20380 80000 20620 80020
rect 20880 80000 21120 80020
rect 21380 80000 21620 80020
rect 21880 80000 22120 80020
rect 22380 80000 22620 80020
rect 22880 80000 23120 80020
rect 23380 80000 23620 80020
rect 23880 80000 24120 80020
rect 24380 80000 24620 80020
rect 24880 80000 25120 80020
rect 25380 80000 25620 80020
rect 25880 80000 26120 80020
rect 26380 80000 26620 80020
rect 26880 80000 27120 80020
rect 27380 80000 27620 80020
rect 27880 80000 28120 80020
rect 28380 80000 28620 80020
rect 28880 80000 29120 80020
rect 29380 80000 29620 80020
rect 29880 80000 30120 80020
rect 30380 80000 30620 80020
rect 30880 80000 31120 80020
rect 31380 80000 31620 80020
rect 31880 80000 32120 80020
rect 32380 80000 32620 80020
rect 32880 80000 33120 80020
rect 33380 80000 33620 80020
rect 33880 80000 34120 80020
rect 34380 80000 34620 80020
rect 34880 80000 35120 80020
rect 35380 80000 35620 80020
rect 35880 80000 36120 80020
rect 36380 80000 36620 80020
rect 36880 80000 37120 80020
rect 37380 80000 37620 80020
rect 37880 80000 38120 80020
rect 38380 80000 38620 80020
rect 38880 80000 39120 80020
rect 39380 80000 39620 80020
rect 39880 80000 40120 80020
rect 40380 80000 40620 80020
rect 40880 80000 41120 80020
rect 41380 80000 41620 80020
rect 41880 80000 42120 80020
rect 42380 80000 42620 80020
rect 42880 80000 43120 80020
rect 43380 80000 43620 80020
rect 43880 80000 44120 80020
rect 44380 80000 44620 80020
rect 44880 80000 45120 80020
rect 45380 80000 45620 80020
rect 45880 80000 46120 80020
rect 46380 80000 46620 80020
rect 46880 80000 47120 80020
rect 47380 80000 47620 80020
rect 47880 80000 48120 80020
rect 48380 80000 48620 80020
rect 48880 80000 49120 80020
rect 49380 80000 49620 80020
rect 49880 80000 50120 80020
rect 50380 80000 50620 80020
rect 50880 80000 51120 80020
rect 51380 80000 51620 80020
rect 51880 80000 52120 80020
rect 52380 80000 52620 80020
rect 52880 80000 53120 80020
rect 53380 80000 53620 80020
rect 53880 80000 54120 80020
rect 54380 80000 54620 80020
rect 54880 80000 55120 80020
rect 55380 80000 55620 80020
rect 55880 80000 56120 80020
rect 56380 80000 56620 80020
rect 56880 80000 57120 80020
rect 57380 80000 57620 80020
rect 57880 80000 58120 80020
rect 58380 80000 58620 80020
rect 58880 80000 59120 80020
rect 59380 80000 59620 80020
rect 59880 80000 60120 80020
rect 60380 80000 60620 80020
rect 60880 80000 61120 80020
rect 61380 80000 61620 80020
rect 61880 80000 62120 80020
rect 62380 80000 62620 80020
rect 62880 80000 63120 80020
rect 63380 80000 63620 80020
rect 63880 80000 64120 80020
rect 64380 80000 64620 80020
rect 64880 80000 65120 80020
rect 65380 80000 65620 80020
rect 65880 80000 66120 80020
rect 66380 80000 66620 80020
rect 66880 80000 67120 80020
rect 67380 80000 67620 80020
rect 67880 80000 68120 80020
rect 68380 80000 68620 80020
rect 68880 80000 69120 80020
rect 69380 80000 69620 80020
rect 69880 80000 70120 80020
rect 70380 80000 70620 80020
rect 70880 80000 71120 80020
rect 71380 80000 71620 80020
rect 71880 80000 72120 80020
rect 72380 80000 72620 80020
rect 72880 80000 73120 80020
rect 73380 80000 73620 80020
rect 73880 80000 74120 80020
rect 74380 80000 74620 80020
rect 74880 80000 75120 80020
rect 75380 80000 75620 80020
rect 75880 80000 76120 80020
rect 76380 80000 76620 80020
rect 76880 80000 77120 80020
rect 77380 80000 77620 80020
rect 77880 80000 78120 80020
rect 78380 80000 78620 80020
rect 78880 80000 79120 80020
rect 79380 80000 79620 80020
rect 79880 80000 80120 80020
rect 80380 80000 80620 80020
rect 80880 80000 81120 80020
rect 81380 80000 81620 80020
rect 81880 80000 82120 80020
rect 82380 80000 82620 80020
rect 82880 80000 83120 80020
rect 83380 80000 83620 80020
rect 83880 80000 84120 80020
rect 84380 80000 84620 80020
rect 84880 80000 85120 80020
rect 85380 80000 85620 80020
rect 85880 80000 86120 80020
rect 86380 80000 86620 80020
rect 86880 80000 87120 80020
rect 87380 80000 87620 80020
rect 87880 80000 88120 80020
rect 88380 80000 88620 80020
rect 88880 80000 89120 80020
rect 89380 80000 89620 80020
rect 89880 80000 90120 80020
rect 90380 80000 90620 80020
rect 90880 80000 91120 80020
rect 91380 80000 91620 80020
rect 91880 80000 92120 80020
rect 92380 80000 92620 80020
rect 92880 80000 93120 80020
rect 93380 80000 93620 80020
rect 93880 80000 94120 80020
rect 94380 80000 94620 80020
rect 94880 80000 95120 80020
rect 95380 80000 95620 80020
rect 95880 80000 96120 80020
rect 96380 80000 96620 80020
rect 96880 80000 97120 80020
rect 97380 80000 97620 80020
rect 97880 80000 98120 80020
rect 98380 80000 98620 80020
rect 98880 80000 99120 80020
rect 99380 80000 99620 80020
rect 99880 80000 100120 80020
rect 100380 80000 100500 80020
rect -83500 79990 100500 80000
rect -83500 79920 -83350 79990
rect -83150 79920 -82850 79990
rect -82650 79920 -82350 79990
rect -82150 79920 -81850 79990
rect -81650 79920 -81350 79990
rect -81150 79920 -80850 79990
rect -80650 79920 -80350 79990
rect -80150 79920 -79850 79990
rect -79650 79920 -79350 79990
rect -79150 79920 -78850 79990
rect -78650 79920 -78350 79990
rect -78150 79920 -77850 79990
rect -77650 79920 -77350 79990
rect -77150 79920 -76850 79990
rect -76650 79920 -76350 79990
rect -76150 79920 -75850 79990
rect -75650 79920 -75350 79990
rect -75150 79920 -74850 79990
rect -74650 79920 -74350 79990
rect -74150 79920 -73850 79990
rect -73650 79920 -73350 79990
rect -73150 79920 -72850 79990
rect -72650 79920 -72350 79990
rect -72150 79920 -71850 79990
rect -71650 79920 -71350 79990
rect -71150 79920 -70850 79990
rect -70650 79920 -70350 79990
rect -70150 79920 -69850 79990
rect -69650 79920 -69350 79990
rect -69150 79920 -68850 79990
rect -68650 79920 -68350 79990
rect -68150 79920 -67850 79990
rect -67650 79920 -67350 79990
rect -67150 79920 -66850 79990
rect -66650 79920 -66350 79990
rect -66150 79920 -65850 79990
rect -65650 79920 -65350 79990
rect -65150 79920 -64850 79990
rect -64650 79920 -64350 79990
rect -64150 79920 -63850 79990
rect -63650 79920 -63350 79990
rect -63150 79920 -62850 79990
rect -62650 79920 -62350 79990
rect -62150 79920 -61850 79990
rect -61650 79920 -61350 79990
rect -61150 79920 -60850 79990
rect -60650 79920 -60350 79990
rect -60150 79920 -59850 79990
rect -59650 79920 -59350 79990
rect -59150 79920 -58850 79990
rect -58650 79920 -58350 79990
rect -58150 79920 -57850 79990
rect -57650 79920 -57350 79990
rect -57150 79920 -56850 79990
rect -56650 79920 -56350 79990
rect -56150 79920 -55850 79990
rect -55650 79920 -55350 79990
rect -55150 79920 -54850 79990
rect -54650 79920 -54350 79990
rect -54150 79920 -53850 79990
rect -53650 79920 -53350 79990
rect -53150 79920 -52850 79990
rect -52650 79920 -52350 79990
rect -52150 79920 -51850 79990
rect -51650 79920 -51350 79990
rect -51150 79920 -50850 79990
rect -50650 79920 -50350 79990
rect -50150 79920 -49850 79990
rect -49650 79920 -49350 79990
rect -49150 79920 -48850 79990
rect -48650 79920 -48350 79990
rect -48150 79920 -47850 79990
rect -47650 79920 -47350 79990
rect -47150 79920 -46850 79990
rect -46650 79920 -46350 79990
rect -46150 79920 -45850 79990
rect -45650 79920 -45350 79990
rect -45150 79920 -44850 79990
rect -44650 79920 -44350 79990
rect -44150 79920 -43850 79990
rect -43650 79920 -43350 79990
rect -43150 79920 -42850 79990
rect -42650 79920 -42350 79990
rect -42150 79920 -41850 79990
rect -41650 79920 -41350 79990
rect -41150 79920 -40850 79990
rect -40650 79920 -40350 79990
rect -40150 79920 -39850 79990
rect -39650 79920 -39350 79990
rect -39150 79920 -38850 79990
rect -38650 79920 -38350 79990
rect -38150 79920 -37850 79990
rect -37650 79920 -37350 79990
rect -37150 79920 -36850 79990
rect -36650 79920 -36350 79990
rect -36150 79920 -35850 79990
rect -35650 79920 -35350 79990
rect -35150 79920 -34850 79990
rect -34650 79920 -34350 79990
rect -34150 79920 -33850 79990
rect -33650 79920 -33350 79990
rect -33150 79920 -32850 79990
rect -32650 79920 -32350 79990
rect -32150 79920 -31850 79990
rect -31650 79920 -31350 79990
rect -31150 79920 -30850 79990
rect -30650 79920 -30350 79990
rect -30150 79920 -29850 79990
rect -29650 79920 -29350 79990
rect -29150 79920 -28850 79990
rect -28650 79920 -28350 79990
rect -28150 79920 -27850 79990
rect -27650 79920 -27350 79990
rect -27150 79920 -26850 79990
rect -26650 79920 -26350 79990
rect -26150 79920 -25850 79990
rect -25650 79920 -25350 79990
rect -25150 79920 -24850 79990
rect -24650 79920 -24350 79990
rect -24150 79920 -23850 79990
rect -23650 79920 -23350 79990
rect -23150 79920 -22850 79990
rect -22650 79920 -22350 79990
rect -22150 79920 -21850 79990
rect -21650 79920 -21350 79990
rect -21150 79920 -20850 79990
rect -20650 79920 -20350 79990
rect -20150 79920 -19850 79990
rect -19650 79920 -19350 79990
rect -19150 79920 -18850 79990
rect -18650 79920 -18350 79990
rect -18150 79920 -17850 79990
rect -17650 79920 -17350 79990
rect -17150 79920 -16850 79990
rect -16650 79920 -16350 79990
rect -16150 79920 -15850 79990
rect -15650 79920 -15350 79990
rect -15150 79920 -14850 79990
rect -14650 79920 -14350 79990
rect -14150 79920 -13850 79990
rect -13650 79920 -13350 79990
rect -13150 79920 -12850 79990
rect -12650 79920 -12350 79990
rect -12150 79920 -11850 79990
rect -11650 79920 -11350 79990
rect -11150 79920 -10850 79990
rect -10650 79920 -10350 79990
rect -10150 79920 -9850 79990
rect -9650 79920 -9350 79990
rect -9150 79920 -8850 79990
rect -8650 79920 -8350 79990
rect -8150 79920 -7850 79990
rect -7650 79920 -7350 79990
rect -7150 79920 -6850 79990
rect -6650 79920 -6350 79990
rect -6150 79920 -5850 79990
rect -5650 79920 -5350 79990
rect -5150 79920 -4850 79990
rect -4650 79920 -4350 79990
rect -4150 79920 -3850 79990
rect -3650 79920 -3350 79990
rect -3150 79920 -2850 79990
rect -2650 79920 -2350 79990
rect -2150 79920 -1850 79990
rect -1650 79920 -1350 79990
rect -1150 79920 -850 79990
rect -650 79920 -350 79990
rect -150 79920 150 79990
rect 350 79920 650 79990
rect 850 79920 1150 79990
rect 1350 79920 1650 79990
rect 1850 79920 2150 79990
rect 2350 79920 2650 79990
rect 2850 79920 3150 79990
rect 3350 79920 3650 79990
rect 3850 79920 4150 79990
rect 4350 79920 4650 79990
rect 4850 79920 5150 79990
rect 5350 79920 5650 79990
rect 5850 79920 6150 79990
rect 6350 79920 6650 79990
rect 6850 79920 7150 79990
rect 7350 79920 7650 79990
rect 7850 79920 8150 79990
rect 8350 79920 8650 79990
rect 8850 79920 9150 79990
rect 9350 79920 9650 79990
rect 9850 79920 10150 79990
rect 10350 79920 10650 79990
rect 10850 79920 11150 79990
rect 11350 79920 11650 79990
rect 11850 79920 12150 79990
rect 12350 79920 12650 79990
rect 12850 79920 13150 79990
rect 13350 79920 13650 79990
rect 13850 79920 14150 79990
rect 14350 79920 14650 79990
rect 14850 79920 15150 79990
rect 15350 79920 15650 79990
rect 15850 79920 16150 79990
rect 16350 79920 16650 79990
rect 16850 79920 17150 79990
rect 17350 79920 17650 79990
rect 17850 79920 18150 79990
rect 18350 79920 18650 79990
rect 18850 79920 19150 79990
rect 19350 79920 19650 79990
rect 19850 79920 20150 79990
rect 20350 79920 20650 79990
rect 20850 79920 21150 79990
rect 21350 79920 21650 79990
rect 21850 79920 22150 79990
rect 22350 79920 22650 79990
rect 22850 79920 23150 79990
rect 23350 79920 23650 79990
rect 23850 79920 24150 79990
rect 24350 79920 24650 79990
rect 24850 79920 25150 79990
rect 25350 79920 25650 79990
rect 25850 79920 26150 79990
rect 26350 79920 26650 79990
rect 26850 79920 27150 79990
rect 27350 79920 27650 79990
rect 27850 79920 28150 79990
rect 28350 79920 28650 79990
rect 28850 79920 29150 79990
rect 29350 79920 29650 79990
rect 29850 79920 30150 79990
rect 30350 79920 30650 79990
rect 30850 79920 31150 79990
rect 31350 79920 31650 79990
rect 31850 79920 32150 79990
rect 32350 79920 32650 79990
rect 32850 79920 33150 79990
rect 33350 79920 33650 79990
rect 33850 79920 34150 79990
rect 34350 79920 34650 79990
rect 34850 79920 35150 79990
rect 35350 79920 35650 79990
rect 35850 79920 36150 79990
rect 36350 79920 36650 79990
rect 36850 79920 37150 79990
rect 37350 79920 37650 79990
rect 37850 79920 38150 79990
rect 38350 79920 38650 79990
rect 38850 79920 39150 79990
rect 39350 79920 39650 79990
rect 39850 79920 40150 79990
rect 40350 79920 40650 79990
rect 40850 79920 41150 79990
rect 41350 79920 41650 79990
rect 41850 79920 42150 79990
rect 42350 79920 42650 79990
rect 42850 79920 43150 79990
rect 43350 79920 43650 79990
rect 43850 79920 44150 79990
rect 44350 79920 44650 79990
rect 44850 79920 45150 79990
rect 45350 79920 45650 79990
rect 45850 79920 46150 79990
rect 46350 79920 46650 79990
rect 46850 79920 47150 79990
rect 47350 79920 47650 79990
rect 47850 79920 48150 79990
rect 48350 79920 48650 79990
rect 48850 79920 49150 79990
rect 49350 79920 49650 79990
rect 49850 79920 50150 79990
rect 50350 79920 50650 79990
rect 50850 79920 51150 79990
rect 51350 79920 51650 79990
rect 51850 79920 52150 79990
rect 52350 79920 52650 79990
rect 52850 79920 53150 79990
rect 53350 79920 53650 79990
rect 53850 79920 54150 79990
rect 54350 79920 54650 79990
rect 54850 79920 55150 79990
rect 55350 79920 55650 79990
rect 55850 79920 56150 79990
rect 56350 79920 56650 79990
rect 56850 79920 57150 79990
rect 57350 79920 57650 79990
rect 57850 79920 58150 79990
rect 58350 79920 58650 79990
rect 58850 79920 59150 79990
rect 59350 79920 59650 79990
rect 59850 79920 60150 79990
rect 60350 79920 60650 79990
rect 60850 79920 61150 79990
rect 61350 79920 61650 79990
rect 61850 79920 62150 79990
rect 62350 79920 62650 79990
rect 62850 79920 63150 79990
rect 63350 79920 63650 79990
rect 63850 79920 64150 79990
rect 64350 79920 64650 79990
rect 64850 79920 65150 79990
rect 65350 79920 65650 79990
rect 65850 79920 66150 79990
rect 66350 79920 66650 79990
rect 66850 79920 67150 79990
rect 67350 79920 67650 79990
rect 67850 79920 68150 79990
rect 68350 79920 68650 79990
rect 68850 79920 69150 79990
rect 69350 79920 69650 79990
rect 69850 79920 70150 79990
rect 70350 79920 70650 79990
rect 70850 79920 71150 79990
rect 71350 79920 71650 79990
rect 71850 79920 72150 79990
rect 72350 79920 72650 79990
rect 72850 79920 73150 79990
rect 73350 79920 73650 79990
rect 73850 79920 74150 79990
rect 74350 79920 74650 79990
rect 74850 79920 75150 79990
rect 75350 79920 75650 79990
rect 75850 79920 76150 79990
rect 76350 79920 76650 79990
rect 76850 79920 77150 79990
rect 77350 79920 77650 79990
rect 77850 79920 78150 79990
rect 78350 79920 78650 79990
rect 78850 79920 79150 79990
rect 79350 79920 79650 79990
rect 79850 79920 80150 79990
rect 80350 79920 80650 79990
rect 80850 79920 81150 79990
rect 81350 79920 81650 79990
rect 81850 79920 82150 79990
rect 82350 79920 82650 79990
rect 82850 79920 83150 79990
rect 83350 79920 83650 79990
rect 83850 79920 84150 79990
rect 84350 79920 84650 79990
rect 84850 79920 85150 79990
rect 85350 79920 85650 79990
rect 85850 79920 86150 79990
rect 86350 79920 86650 79990
rect 86850 79920 87150 79990
rect 87350 79920 87650 79990
rect 87850 79920 88150 79990
rect 88350 79920 88650 79990
rect 88850 79920 89150 79990
rect 89350 79920 89650 79990
rect 89850 79920 90150 79990
rect 90350 79920 90650 79990
rect 90850 79920 91150 79990
rect 91350 79920 91650 79990
rect 91850 79920 92150 79990
rect 92350 79920 92650 79990
rect 92850 79920 93150 79990
rect 93350 79920 93650 79990
rect 93850 79920 94150 79990
rect 94350 79920 94650 79990
rect 94850 79920 95150 79990
rect 95350 79920 95650 79990
rect 95850 79920 96150 79990
rect 96350 79920 96650 79990
rect 96850 79920 97150 79990
rect 97350 79920 97650 79990
rect 97850 79920 98150 79990
rect 98350 79920 98650 79990
rect 98850 79920 99150 79990
rect 99350 79920 99650 79990
rect 99850 79920 100150 79990
rect 100350 79920 100500 79990
rect -83500 79900 100500 79920
rect 128500 25800 143500 25900
rect 128500 25780 128620 25800
rect 128880 25780 129120 25800
rect 129380 25780 129620 25800
rect 129880 25780 130120 25800
rect 130380 25780 130620 25800
rect 130880 25780 131120 25800
rect 131380 25780 131620 25800
rect 131880 25780 132120 25800
rect 132380 25780 132620 25800
rect 132880 25780 133120 25800
rect 133380 25780 133620 25800
rect 133880 25780 134120 25800
rect 134380 25780 134620 25800
rect 134880 25780 135120 25800
rect 135380 25780 135620 25800
rect 135880 25780 136120 25800
rect 136380 25780 136620 25800
rect 136880 25780 137120 25800
rect 137380 25780 137620 25800
rect 137880 25780 138120 25800
rect 138380 25780 138620 25800
rect 138880 25780 139120 25800
rect 139380 25780 139620 25800
rect 139880 25780 140120 25800
rect 140380 25780 140620 25800
rect 140880 25780 141120 25800
rect 141380 25780 141620 25800
rect 141880 25780 142120 25800
rect 142380 25780 142620 25800
rect 142880 25780 143120 25800
rect 143380 25780 143500 25800
rect 128500 25520 128600 25780
rect 128900 25520 129100 25780
rect 129400 25520 129600 25780
rect 129900 25520 130100 25780
rect 130400 25520 130600 25780
rect 130900 25520 131100 25780
rect 131400 25520 131600 25780
rect 131900 25520 132100 25780
rect 132400 25520 132600 25780
rect 132900 25520 133100 25780
rect 133400 25520 133600 25780
rect 133900 25520 134100 25780
rect 134400 25520 134600 25780
rect 134900 25520 135100 25780
rect 135400 25520 135600 25780
rect 135900 25520 136100 25780
rect 136400 25520 136600 25780
rect 136900 25520 137100 25780
rect 137400 25520 137600 25780
rect 137900 25520 138100 25780
rect 138400 25520 138600 25780
rect 138900 25520 139100 25780
rect 139400 25520 139600 25780
rect 139900 25520 140100 25780
rect 140400 25520 140600 25780
rect 140900 25520 141100 25780
rect 141400 25520 141600 25780
rect 141900 25520 142100 25780
rect 142400 25520 142600 25780
rect 142900 25520 143100 25780
rect 143400 25520 143500 25780
rect 128500 25500 128620 25520
rect 128880 25500 129120 25520
rect 129380 25500 129620 25520
rect 129880 25500 130120 25520
rect 130380 25500 130620 25520
rect 130880 25500 131120 25520
rect 131380 25500 131620 25520
rect 131880 25500 132120 25520
rect 132380 25500 132620 25520
rect 132880 25500 133120 25520
rect 133380 25500 133620 25520
rect 133880 25500 134120 25520
rect 134380 25500 134620 25520
rect 134880 25500 135120 25520
rect 135380 25500 135620 25520
rect 135880 25500 136120 25520
rect 136380 25500 136620 25520
rect 136880 25500 137120 25520
rect 137380 25500 137620 25520
rect 137880 25500 138120 25520
rect 138380 25500 138620 25520
rect 138880 25500 139120 25520
rect 139380 25500 139620 25520
rect 139880 25500 140120 25520
rect 140380 25500 140620 25520
rect 140880 25500 141120 25520
rect 141380 25500 141620 25520
rect 141880 25500 142120 25520
rect 142380 25500 142620 25520
rect 142880 25500 143120 25520
rect 143380 25500 143500 25520
rect 128500 25300 143500 25500
rect 128500 25280 128620 25300
rect 128880 25280 129120 25300
rect 129380 25280 129620 25300
rect 129880 25280 130120 25300
rect 130380 25280 130620 25300
rect 130880 25280 131120 25300
rect 131380 25280 131620 25300
rect 131880 25280 132120 25300
rect 132380 25280 132620 25300
rect 132880 25280 133120 25300
rect 133380 25280 133620 25300
rect 133880 25280 134120 25300
rect 134380 25280 134620 25300
rect 134880 25280 135120 25300
rect 135380 25280 135620 25300
rect 135880 25280 136120 25300
rect 136380 25280 136620 25300
rect 136880 25280 137120 25300
rect 137380 25280 137620 25300
rect 137880 25280 138120 25300
rect 138380 25280 138620 25300
rect 138880 25280 139120 25300
rect 139380 25280 139620 25300
rect 139880 25280 140120 25300
rect 140380 25280 140620 25300
rect 140880 25280 141120 25300
rect 141380 25280 141620 25300
rect 141880 25280 142120 25300
rect 142380 25280 142620 25300
rect 142880 25280 143120 25300
rect 143380 25280 143500 25300
rect 128500 25020 128600 25280
rect 128900 25020 129100 25280
rect 129400 25020 129600 25280
rect 129900 25020 130100 25280
rect 130400 25020 130600 25280
rect 130900 25020 131100 25280
rect 131400 25020 131600 25280
rect 131900 25020 132100 25280
rect 132400 25020 132600 25280
rect 132900 25020 133100 25280
rect 133400 25020 133600 25280
rect 133900 25020 134100 25280
rect 134400 25020 134600 25280
rect 134900 25020 135100 25280
rect 135400 25020 135600 25280
rect 135900 25020 136100 25280
rect 136400 25020 136600 25280
rect 136900 25020 137100 25280
rect 137400 25020 137600 25280
rect 137900 25020 138100 25280
rect 138400 25020 138600 25280
rect 138900 25020 139100 25280
rect 139400 25020 139600 25280
rect 139900 25020 140100 25280
rect 140400 25020 140600 25280
rect 140900 25020 141100 25280
rect 141400 25020 141600 25280
rect 141900 25020 142100 25280
rect 142400 25020 142600 25280
rect 142900 25020 143100 25280
rect 143400 25020 143500 25280
rect 128500 25000 128620 25020
rect 128880 25000 129120 25020
rect 129380 25000 129620 25020
rect 129880 25000 130120 25020
rect 130380 25000 130620 25020
rect 130880 25000 131120 25020
rect 131380 25000 131620 25020
rect 131880 25000 132120 25020
rect 132380 25000 132620 25020
rect 132880 25000 133120 25020
rect 133380 25000 133620 25020
rect 133880 25000 134120 25020
rect 134380 25000 134620 25020
rect 134880 25000 135120 25020
rect 135380 25000 135620 25020
rect 135880 25000 136120 25020
rect 136380 25000 136620 25020
rect 136880 25000 137120 25020
rect 137380 25000 137620 25020
rect 137880 25000 138120 25020
rect 138380 25000 138620 25020
rect 138880 25000 139120 25020
rect 139380 25000 139620 25020
rect 139880 25000 140120 25020
rect 140380 25000 140620 25020
rect 140880 25000 141120 25020
rect 141380 25000 141620 25020
rect 141880 25000 142120 25020
rect 142380 25000 142620 25020
rect 142880 25000 143120 25020
rect 143380 25000 143500 25020
rect 128500 24800 143500 25000
rect 128500 24780 128620 24800
rect 128880 24780 129120 24800
rect 129380 24780 129620 24800
rect 129880 24780 130120 24800
rect 130380 24780 130620 24800
rect 130880 24780 131120 24800
rect 131380 24780 131620 24800
rect 131880 24780 132120 24800
rect 132380 24780 132620 24800
rect 132880 24780 133120 24800
rect 133380 24780 133620 24800
rect 133880 24780 134120 24800
rect 134380 24780 134620 24800
rect 134880 24780 135120 24800
rect 135380 24780 135620 24800
rect 135880 24780 136120 24800
rect 136380 24780 136620 24800
rect 136880 24780 137120 24800
rect 137380 24780 137620 24800
rect 137880 24780 138120 24800
rect 138380 24780 138620 24800
rect 138880 24780 139120 24800
rect 139380 24780 139620 24800
rect 139880 24780 140120 24800
rect 140380 24780 140620 24800
rect 140880 24780 141120 24800
rect 141380 24780 141620 24800
rect 141880 24780 142120 24800
rect 142380 24780 142620 24800
rect 142880 24780 143120 24800
rect 143380 24780 143500 24800
rect 128500 24520 128600 24780
rect 128900 24520 129100 24780
rect 129400 24520 129600 24780
rect 129900 24520 130100 24780
rect 130400 24520 130600 24780
rect 130900 24520 131100 24780
rect 131400 24520 131600 24780
rect 131900 24520 132100 24780
rect 132400 24520 132600 24780
rect 132900 24520 133100 24780
rect 133400 24520 133600 24780
rect 133900 24520 134100 24780
rect 134400 24520 134600 24780
rect 134900 24520 135100 24780
rect 135400 24520 135600 24780
rect 135900 24520 136100 24780
rect 136400 24520 136600 24780
rect 136900 24520 137100 24780
rect 137400 24520 137600 24780
rect 137900 24520 138100 24780
rect 138400 24520 138600 24780
rect 138900 24520 139100 24780
rect 139400 24520 139600 24780
rect 139900 24520 140100 24780
rect 140400 24520 140600 24780
rect 140900 24520 141100 24780
rect 141400 24520 141600 24780
rect 141900 24520 142100 24780
rect 142400 24520 142600 24780
rect 142900 24520 143100 24780
rect 143400 24520 143500 24780
rect 128500 24500 128620 24520
rect 128880 24500 129120 24520
rect 129380 24500 129620 24520
rect 129880 24500 130120 24520
rect 130380 24500 130620 24520
rect 130880 24500 131120 24520
rect 131380 24500 131620 24520
rect 131880 24500 132120 24520
rect 132380 24500 132620 24520
rect 132880 24500 133120 24520
rect 133380 24500 133620 24520
rect 133880 24500 134120 24520
rect 134380 24500 134620 24520
rect 134880 24500 135120 24520
rect 135380 24500 135620 24520
rect 135880 24500 136120 24520
rect 136380 24500 136620 24520
rect 136880 24500 137120 24520
rect 137380 24500 137620 24520
rect 137880 24500 138120 24520
rect 138380 24500 138620 24520
rect 138880 24500 139120 24520
rect 139380 24500 139620 24520
rect 139880 24500 140120 24520
rect 140380 24500 140620 24520
rect 140880 24500 141120 24520
rect 141380 24500 141620 24520
rect 141880 24500 142120 24520
rect 142380 24500 142620 24520
rect 142880 24500 143120 24520
rect 143380 24500 143500 24520
rect 128500 24300 143500 24500
rect 128500 24280 128620 24300
rect 128880 24280 129120 24300
rect 129380 24280 129620 24300
rect 129880 24280 130120 24300
rect 130380 24280 130620 24300
rect 130880 24280 131120 24300
rect 131380 24280 131620 24300
rect 131880 24280 132120 24300
rect 132380 24280 132620 24300
rect 132880 24280 133120 24300
rect 133380 24280 133620 24300
rect 133880 24280 134120 24300
rect 134380 24280 134620 24300
rect 134880 24280 135120 24300
rect 135380 24280 135620 24300
rect 135880 24280 136120 24300
rect 136380 24280 136620 24300
rect 136880 24280 137120 24300
rect 137380 24280 137620 24300
rect 137880 24280 138120 24300
rect 138380 24280 138620 24300
rect 138880 24280 139120 24300
rect 139380 24280 139620 24300
rect 139880 24280 140120 24300
rect 140380 24280 140620 24300
rect 140880 24280 141120 24300
rect 141380 24280 141620 24300
rect 141880 24280 142120 24300
rect 142380 24280 142620 24300
rect 142880 24280 143120 24300
rect 143380 24280 143500 24300
rect 128500 24020 128600 24280
rect 128900 24020 129100 24280
rect 129400 24020 129600 24280
rect 129900 24020 130100 24280
rect 130400 24020 130600 24280
rect 130900 24020 131100 24280
rect 131400 24020 131600 24280
rect 131900 24020 132100 24280
rect 132400 24020 132600 24280
rect 132900 24020 133100 24280
rect 133400 24020 133600 24280
rect 133900 24020 134100 24280
rect 134400 24020 134600 24280
rect 134900 24020 135100 24280
rect 135400 24020 135600 24280
rect 135900 24020 136100 24280
rect 136400 24020 136600 24280
rect 136900 24020 137100 24280
rect 137400 24020 137600 24280
rect 137900 24020 138100 24280
rect 138400 24020 138600 24280
rect 138900 24020 139100 24280
rect 139400 24020 139600 24280
rect 139900 24020 140100 24280
rect 140400 24020 140600 24280
rect 140900 24020 141100 24280
rect 141400 24020 141600 24280
rect 141900 24020 142100 24280
rect 142400 24020 142600 24280
rect 142900 24020 143100 24280
rect 143400 24020 143500 24280
rect 128500 24000 128620 24020
rect 128880 24000 129120 24020
rect 129380 24000 129620 24020
rect 129880 24000 130120 24020
rect 130380 24000 130620 24020
rect 130880 24000 131120 24020
rect 131380 24000 131620 24020
rect 131880 24000 132120 24020
rect 132380 24000 132620 24020
rect 132880 24000 133120 24020
rect 133380 24000 133620 24020
rect 133880 24000 134120 24020
rect 134380 24000 134620 24020
rect 134880 24000 135120 24020
rect 135380 24000 135620 24020
rect 135880 24000 136120 24020
rect 136380 24000 136620 24020
rect 136880 24000 137120 24020
rect 137380 24000 137620 24020
rect 137880 24000 138120 24020
rect 138380 24000 138620 24020
rect 138880 24000 139120 24020
rect 139380 24000 139620 24020
rect 139880 24000 140120 24020
rect 140380 24000 140620 24020
rect 140880 24000 141120 24020
rect 141380 24000 141620 24020
rect 141880 24000 142120 24020
rect 142380 24000 142620 24020
rect 142880 24000 143120 24020
rect 143380 24000 143500 24020
rect 128500 23900 143500 24000
rect 140500 23800 143500 23900
rect 140500 23780 140620 23800
rect 140880 23780 141120 23800
rect 141380 23780 141620 23800
rect 141880 23780 142120 23800
rect 142380 23780 142620 23800
rect 142880 23780 143120 23800
rect 143380 23780 143500 23800
rect 140500 23520 140600 23780
rect 140900 23520 141100 23780
rect 141400 23520 141600 23780
rect 141900 23520 142100 23780
rect 142400 23520 142600 23780
rect 142900 23520 143100 23780
rect 143400 23520 143500 23780
rect 140500 23500 140620 23520
rect 140880 23500 141120 23520
rect 141380 23500 141620 23520
rect 141880 23500 142120 23520
rect 142380 23500 142620 23520
rect 142880 23500 143120 23520
rect 143380 23500 143500 23520
rect 140500 23300 143500 23500
rect 140500 23280 140620 23300
rect 140880 23280 141120 23300
rect 141380 23280 141620 23300
rect 141880 23280 142120 23300
rect 142380 23280 142620 23300
rect 142880 23280 143120 23300
rect 143380 23280 143500 23300
rect 140500 23020 140600 23280
rect 140900 23020 141100 23280
rect 141400 23020 141600 23280
rect 141900 23020 142100 23280
rect 142400 23020 142600 23280
rect 142900 23020 143100 23280
rect 143400 23020 143500 23280
rect 140500 23000 140620 23020
rect 140880 23000 141120 23020
rect 141380 23000 141620 23020
rect 141880 23000 142120 23020
rect 142380 23000 142620 23020
rect 142880 23000 143120 23020
rect 143380 23000 143500 23020
rect 140500 22800 143500 23000
rect 140500 22780 140620 22800
rect 140880 22780 141120 22800
rect 141380 22780 141620 22800
rect 141880 22780 142120 22800
rect 142380 22780 142620 22800
rect 142880 22780 143120 22800
rect 143380 22780 143500 22800
rect 140500 22520 140600 22780
rect 140900 22520 141100 22780
rect 141400 22520 141600 22780
rect 141900 22520 142100 22780
rect 142400 22520 142600 22780
rect 142900 22520 143100 22780
rect 143400 22520 143500 22780
rect 140500 22500 140620 22520
rect 140880 22500 141120 22520
rect 141380 22500 141620 22520
rect 141880 22500 142120 22520
rect 142380 22500 142620 22520
rect 142880 22500 143120 22520
rect 143380 22500 143500 22520
rect 140500 22300 143500 22500
rect 140500 22280 140620 22300
rect 140880 22280 141120 22300
rect 141380 22280 141620 22300
rect 141880 22280 142120 22300
rect 142380 22280 142620 22300
rect 142880 22280 143120 22300
rect 143380 22280 143500 22300
rect 140500 22020 140600 22280
rect 140900 22020 141100 22280
rect 141400 22020 141600 22280
rect 141900 22020 142100 22280
rect 142400 22020 142600 22280
rect 142900 22020 143100 22280
rect 143400 22020 143500 22280
rect 140500 22000 140620 22020
rect 140880 22000 141120 22020
rect 141380 22000 141620 22020
rect 141880 22000 142120 22020
rect 142380 22000 142620 22020
rect 142880 22000 143120 22020
rect 143380 22000 143500 22020
rect 140500 21800 143500 22000
rect 140500 21780 140620 21800
rect 140880 21780 141120 21800
rect 141380 21780 141620 21800
rect 141880 21780 142120 21800
rect 142380 21780 142620 21800
rect 142880 21780 143120 21800
rect 143380 21780 143500 21800
rect 140500 21520 140600 21780
rect 140900 21520 141100 21780
rect 141400 21520 141600 21780
rect 141900 21520 142100 21780
rect 142400 21520 142600 21780
rect 142900 21520 143100 21780
rect 143400 21520 143500 21780
rect 140500 21500 140620 21520
rect 140880 21500 141120 21520
rect 141380 21500 141620 21520
rect 141880 21500 142120 21520
rect 142380 21500 142620 21520
rect 142880 21500 143120 21520
rect 143380 21500 143500 21520
rect 140500 21300 143500 21500
rect 140500 21280 140620 21300
rect 140880 21280 141120 21300
rect 141380 21280 141620 21300
rect 141880 21280 142120 21300
rect 142380 21280 142620 21300
rect 142880 21280 143120 21300
rect 143380 21280 143500 21300
rect 140500 21020 140600 21280
rect 140900 21020 141100 21280
rect 141400 21020 141600 21280
rect 141900 21020 142100 21280
rect 142400 21020 142600 21280
rect 142900 21020 143100 21280
rect 143400 21020 143500 21280
rect 140500 21000 140620 21020
rect 140880 21000 141120 21020
rect 141380 21000 141620 21020
rect 141880 21000 142120 21020
rect 142380 21000 142620 21020
rect 142880 21000 143120 21020
rect 143380 21000 143500 21020
rect 140500 20800 143500 21000
rect 140500 20780 140620 20800
rect 140880 20780 141120 20800
rect 141380 20780 141620 20800
rect 141880 20780 142120 20800
rect 142380 20780 142620 20800
rect 142880 20780 143120 20800
rect 143380 20780 143500 20800
rect 140500 20520 140600 20780
rect 140900 20520 141100 20780
rect 141400 20520 141600 20780
rect 141900 20520 142100 20780
rect 142400 20520 142600 20780
rect 142900 20520 143100 20780
rect 143400 20520 143500 20780
rect 140500 20500 140620 20520
rect 140880 20500 141120 20520
rect 141380 20500 141620 20520
rect 141880 20500 142120 20520
rect 142380 20500 142620 20520
rect 142880 20500 143120 20520
rect 143380 20500 143500 20520
rect 140500 20300 143500 20500
rect 140500 20280 140620 20300
rect 140880 20280 141120 20300
rect 141380 20280 141620 20300
rect 141880 20280 142120 20300
rect 142380 20280 142620 20300
rect 142880 20280 143120 20300
rect 143380 20280 143500 20300
rect 140500 20020 140600 20280
rect 140900 20020 141100 20280
rect 141400 20020 141600 20280
rect 141900 20020 142100 20280
rect 142400 20020 142600 20280
rect 142900 20020 143100 20280
rect 143400 20020 143500 20280
rect 140500 20000 140620 20020
rect 140880 20000 141120 20020
rect 141380 20000 141620 20020
rect 141880 20000 142120 20020
rect 142380 20000 142620 20020
rect 142880 20000 143120 20020
rect 143380 20000 143500 20020
rect 140500 19800 143500 20000
rect 140500 19780 140620 19800
rect 140880 19780 141120 19800
rect 141380 19780 141620 19800
rect 141880 19780 142120 19800
rect 142380 19780 142620 19800
rect 142880 19780 143120 19800
rect 143380 19780 143500 19800
rect 140500 19520 140600 19780
rect 140900 19520 141100 19780
rect 141400 19520 141600 19780
rect 141900 19520 142100 19780
rect 142400 19520 142600 19780
rect 142900 19520 143100 19780
rect 143400 19520 143500 19780
rect 140500 19500 140620 19520
rect 140880 19500 141120 19520
rect 141380 19500 141620 19520
rect 141880 19500 142120 19520
rect 142380 19500 142620 19520
rect 142880 19500 143120 19520
rect 143380 19500 143500 19520
rect 140500 19300 143500 19500
rect 140500 19280 140620 19300
rect 140880 19280 141120 19300
rect 141380 19280 141620 19300
rect 141880 19280 142120 19300
rect 142380 19280 142620 19300
rect 142880 19280 143120 19300
rect 143380 19280 143500 19300
rect 140500 19020 140600 19280
rect 140900 19020 141100 19280
rect 141400 19020 141600 19280
rect 141900 19020 142100 19280
rect 142400 19020 142600 19280
rect 142900 19020 143100 19280
rect 143400 19020 143500 19280
rect 140500 19000 140620 19020
rect 140880 19000 141120 19020
rect 141380 19000 141620 19020
rect 141880 19000 142120 19020
rect 142380 19000 142620 19020
rect 142880 19000 143120 19020
rect 143380 19000 143500 19020
rect 140500 18800 143500 19000
rect 140500 18780 140620 18800
rect 140880 18780 141120 18800
rect 141380 18780 141620 18800
rect 141880 18780 142120 18800
rect 142380 18780 142620 18800
rect 142880 18780 143120 18800
rect 143380 18780 143500 18800
rect 140500 18520 140600 18780
rect 140900 18520 141100 18780
rect 141400 18520 141600 18780
rect 141900 18520 142100 18780
rect 142400 18520 142600 18780
rect 142900 18520 143100 18780
rect 143400 18520 143500 18780
rect 140500 18500 140620 18520
rect 140880 18500 141120 18520
rect 141380 18500 141620 18520
rect 141880 18500 142120 18520
rect 142380 18500 142620 18520
rect 142880 18500 143120 18520
rect 143380 18500 143500 18520
rect 140500 18300 143500 18500
rect 140500 18280 140620 18300
rect 140880 18280 141120 18300
rect 141380 18280 141620 18300
rect 141880 18280 142120 18300
rect 142380 18280 142620 18300
rect 142880 18280 143120 18300
rect 143380 18280 143500 18300
rect 140500 18020 140600 18280
rect 140900 18020 141100 18280
rect 141400 18020 141600 18280
rect 141900 18020 142100 18280
rect 142400 18020 142600 18280
rect 142900 18020 143100 18280
rect 143400 18020 143500 18280
rect 140500 18000 140620 18020
rect 140880 18000 141120 18020
rect 141380 18000 141620 18020
rect 141880 18000 142120 18020
rect 142380 18000 142620 18020
rect 142880 18000 143120 18020
rect 143380 18000 143500 18020
rect 140500 17800 143500 18000
rect 140500 17780 140620 17800
rect 140880 17780 141120 17800
rect 141380 17780 141620 17800
rect 141880 17780 142120 17800
rect 142380 17780 142620 17800
rect 142880 17780 143120 17800
rect 143380 17780 143500 17800
rect 140500 17520 140600 17780
rect 140900 17520 141100 17780
rect 141400 17520 141600 17780
rect 141900 17520 142100 17780
rect 142400 17520 142600 17780
rect 142900 17520 143100 17780
rect 143400 17520 143500 17780
rect 140500 17500 140620 17520
rect 140880 17500 141120 17520
rect 141380 17500 141620 17520
rect 141880 17500 142120 17520
rect 142380 17500 142620 17520
rect 142880 17500 143120 17520
rect 143380 17500 143500 17520
rect 140500 17300 143500 17500
rect 140500 17280 140620 17300
rect 140880 17280 141120 17300
rect 141380 17280 141620 17300
rect 141880 17280 142120 17300
rect 142380 17280 142620 17300
rect 142880 17280 143120 17300
rect 143380 17280 143500 17300
rect 140500 17020 140600 17280
rect 140900 17020 141100 17280
rect 141400 17020 141600 17280
rect 141900 17020 142100 17280
rect 142400 17020 142600 17280
rect 142900 17020 143100 17280
rect 143400 17020 143500 17280
rect 140500 17000 140620 17020
rect 140880 17000 141120 17020
rect 141380 17000 141620 17020
rect 141880 17000 142120 17020
rect 142380 17000 142620 17020
rect 142880 17000 143120 17020
rect 143380 17000 143500 17020
rect 140500 16800 143500 17000
rect 140500 16780 140620 16800
rect 140880 16780 141120 16800
rect 141380 16780 141620 16800
rect 141880 16780 142120 16800
rect 142380 16780 142620 16800
rect 142880 16780 143120 16800
rect 143380 16780 143500 16800
rect 140500 16520 140600 16780
rect 140900 16520 141100 16780
rect 141400 16520 141600 16780
rect 141900 16520 142100 16780
rect 142400 16520 142600 16780
rect 142900 16520 143100 16780
rect 143400 16520 143500 16780
rect 140500 16500 140620 16520
rect 140880 16500 141120 16520
rect 141380 16500 141620 16520
rect 141880 16500 142120 16520
rect 142380 16500 142620 16520
rect 142880 16500 143120 16520
rect 143380 16500 143500 16520
rect 140500 16300 143500 16500
rect 140500 16280 140620 16300
rect 140880 16280 141120 16300
rect 141380 16280 141620 16300
rect 141880 16280 142120 16300
rect 142380 16280 142620 16300
rect 142880 16280 143120 16300
rect 143380 16280 143500 16300
rect 140500 16020 140600 16280
rect 140900 16020 141100 16280
rect 141400 16020 141600 16280
rect 141900 16020 142100 16280
rect 142400 16020 142600 16280
rect 142900 16020 143100 16280
rect 143400 16020 143500 16280
rect 140500 16000 140620 16020
rect 140880 16000 141120 16020
rect 141380 16000 141620 16020
rect 141880 16000 142120 16020
rect 142380 16000 142620 16020
rect 142880 16000 143120 16020
rect 143380 16000 143500 16020
rect 140500 15900 143500 16000
rect 16000 13700 20000 13900
rect -13500 13300 -11500 13400
rect -13500 13280 -13380 13300
rect -13120 13280 -12880 13300
rect -12620 13280 -12380 13300
rect -12120 13280 -11880 13300
rect -11620 13280 -11500 13300
rect -13500 13020 -13400 13280
rect -13100 13020 -12900 13280
rect -12600 13020 -12400 13280
rect -12100 13020 -11900 13280
rect -11600 13020 -11500 13280
rect -13500 13000 -13380 13020
rect -13120 13000 -12880 13020
rect -12620 13000 -12380 13020
rect -12120 13000 -11880 13020
rect -11620 13000 -11500 13020
rect -13500 12800 -11500 13000
rect -13500 12780 -13380 12800
rect -13120 12780 -12880 12800
rect -12620 12780 -12380 12800
rect -12120 12780 -11880 12800
rect -11620 12780 -11500 12800
rect -13500 12520 -13400 12780
rect -13100 12520 -12900 12780
rect -12600 12520 -12400 12780
rect -12100 12520 -11900 12780
rect -11600 12520 -11500 12780
rect -13500 12500 -13380 12520
rect -13120 12500 -12880 12520
rect -12620 12500 -12380 12520
rect -12120 12500 -11880 12520
rect -11620 12500 -11500 12520
rect -13500 12300 -11500 12500
rect -13500 12280 -13380 12300
rect -13120 12280 -12880 12300
rect -12620 12280 -12380 12300
rect -12120 12280 -11880 12300
rect -11620 12280 -11500 12300
rect -13500 12020 -13400 12280
rect -13100 12020 -12900 12280
rect -12600 12020 -12400 12280
rect -12100 12020 -11900 12280
rect -11600 12020 -11500 12280
rect -13500 12000 -13380 12020
rect -13120 12000 -12880 12020
rect -12620 12000 -12380 12020
rect -12120 12000 -11880 12020
rect -11620 12000 -11500 12020
rect -13500 11800 -11500 12000
rect -13500 11780 -13380 11800
rect -13120 11780 -12880 11800
rect -12620 11780 -12380 11800
rect -12120 11780 -11880 11800
rect -11620 11780 -11500 11800
rect -13500 11520 -13400 11780
rect -13100 11520 -12900 11780
rect -12600 11520 -12400 11780
rect -12100 11520 -11900 11780
rect -11600 11520 -11500 11780
rect -13500 11500 -13380 11520
rect -13120 11500 -12880 11520
rect -12620 11500 -12380 11520
rect -12120 11500 -11880 11520
rect -11620 11500 -11500 11520
rect -13500 11300 -11500 11500
rect -13500 11280 -13380 11300
rect -13120 11280 -12880 11300
rect -12620 11280 -12380 11300
rect -12120 11280 -11880 11300
rect -11620 11280 -11500 11300
rect -13500 11020 -13400 11280
rect -13100 11020 -12900 11280
rect -12600 11020 -12400 11280
rect -12100 11020 -11900 11280
rect -11600 11020 -11500 11280
rect -13500 11000 -13380 11020
rect -13120 11000 -12880 11020
rect -12620 11000 -12380 11020
rect -12120 11000 -11880 11020
rect -11620 11000 -11500 11020
rect -13500 10900 -11500 11000
rect -13500 10800 -3000 10900
rect -13500 10780 -13380 10800
rect -13120 10780 -12880 10800
rect -12620 10780 -12380 10800
rect -12120 10780 -11880 10800
rect -11620 10780 -11380 10800
rect -11120 10780 -10880 10800
rect -10620 10780 -10380 10800
rect -10120 10780 -9880 10800
rect -9620 10780 -9380 10800
rect -9120 10780 -8880 10800
rect -8620 10780 -8380 10800
rect -8120 10780 -7880 10800
rect -7620 10780 -7380 10800
rect -7120 10780 -6880 10800
rect -6620 10780 -6380 10800
rect -6120 10780 -5880 10800
rect -5620 10780 -5380 10800
rect -5120 10780 -4880 10800
rect -4620 10780 -4380 10800
rect -4120 10780 -3880 10800
rect -3620 10780 -3380 10800
rect -3120 10780 -3000 10800
rect -13500 10520 -13400 10780
rect -13100 10520 -12900 10780
rect -12600 10520 -12400 10780
rect -12100 10520 -11900 10780
rect -11600 10520 -11400 10780
rect -11100 10520 -10900 10780
rect -10600 10520 -10400 10780
rect -10100 10520 -9900 10780
rect -9600 10520 -9400 10780
rect -9100 10520 -8900 10780
rect -8600 10520 -8400 10780
rect -8100 10520 -7900 10780
rect -7600 10520 -7400 10780
rect -7100 10520 -6900 10780
rect -6600 10520 -6400 10780
rect -6100 10520 -5900 10780
rect -5600 10520 -5400 10780
rect -5100 10520 -4900 10780
rect -4600 10520 -4400 10780
rect -4100 10520 -3900 10780
rect -3600 10520 -3400 10780
rect -3100 10520 -3000 10780
rect -13500 10500 -13380 10520
rect -13120 10500 -12880 10520
rect -12620 10500 -12380 10520
rect -12120 10500 -11880 10520
rect -11620 10500 -11380 10520
rect -11120 10500 -10880 10520
rect -10620 10500 -10380 10520
rect -10120 10500 -9880 10520
rect -9620 10500 -9380 10520
rect -9120 10500 -8880 10520
rect -8620 10500 -8380 10520
rect -8120 10500 -7880 10520
rect -7620 10500 -7380 10520
rect -7120 10500 -6880 10520
rect -6620 10500 -6380 10520
rect -6120 10500 -5880 10520
rect -5620 10500 -5380 10520
rect -5120 10500 -4880 10520
rect -4620 10500 -4380 10520
rect -4120 10500 -3880 10520
rect -3620 10500 -3380 10520
rect -3120 10500 -3000 10520
rect -13500 10300 -3000 10500
rect -13500 10280 -13380 10300
rect -13120 10280 -12880 10300
rect -12620 10280 -12380 10300
rect -12120 10280 -11880 10300
rect -11620 10280 -11380 10300
rect -11120 10280 -10880 10300
rect -10620 10280 -10380 10300
rect -10120 10280 -9880 10300
rect -9620 10280 -9380 10300
rect -9120 10280 -8880 10300
rect -8620 10280 -8380 10300
rect -8120 10280 -7880 10300
rect -7620 10280 -7380 10300
rect -7120 10280 -6880 10300
rect -6620 10280 -6380 10300
rect -6120 10280 -5880 10300
rect -5620 10280 -5380 10300
rect -5120 10280 -4880 10300
rect -4620 10280 -4380 10300
rect -4120 10280 -3880 10300
rect -3620 10280 -3380 10300
rect -3120 10280 -3000 10300
rect -13500 10020 -13400 10280
rect -13100 10020 -12900 10280
rect -12600 10020 -12400 10280
rect -12100 10020 -11900 10280
rect -11600 10020 -11400 10280
rect -11100 10020 -10900 10280
rect -10600 10020 -10400 10280
rect -10100 10020 -9900 10280
rect -9600 10020 -9400 10280
rect -9100 10020 -8900 10280
rect -8600 10020 -8400 10280
rect -8100 10020 -7900 10280
rect -7600 10020 -7400 10280
rect -7100 10020 -6900 10280
rect -6600 10020 -6400 10280
rect -6100 10020 -5900 10280
rect -5600 10020 -5400 10280
rect -5100 10020 -4900 10280
rect -4600 10020 -4400 10280
rect -4100 10020 -3900 10280
rect -3600 10020 -3400 10280
rect -3100 10020 -3000 10280
rect -13500 10000 -13380 10020
rect -13120 10000 -12880 10020
rect -12620 10000 -12380 10020
rect -12120 10000 -11880 10020
rect -11620 10000 -11380 10020
rect -11120 10000 -10880 10020
rect -10620 10000 -10380 10020
rect -10120 10000 -9880 10020
rect -9620 10000 -9380 10020
rect -9120 10000 -8880 10020
rect -8620 10000 -8380 10020
rect -8120 10000 -7880 10020
rect -7620 10000 -7380 10020
rect -7120 10000 -6880 10020
rect -6620 10000 -6380 10020
rect -6120 10000 -5880 10020
rect -5620 10000 -5380 10020
rect -5120 10000 -4880 10020
rect -4620 10000 -4380 10020
rect -4120 10000 -3880 10020
rect -3620 10000 -3380 10020
rect -3120 10000 -3000 10020
rect -13500 9800 -3000 10000
rect -13500 9780 -13380 9800
rect -13120 9780 -12880 9800
rect -12620 9780 -12380 9800
rect -12120 9780 -11880 9800
rect -11620 9780 -11380 9800
rect -11120 9780 -10880 9800
rect -10620 9780 -10380 9800
rect -10120 9780 -9880 9800
rect -9620 9780 -9380 9800
rect -9120 9780 -8880 9800
rect -8620 9780 -8380 9800
rect -8120 9780 -7880 9800
rect -7620 9780 -7380 9800
rect -7120 9780 -6880 9800
rect -6620 9780 -6380 9800
rect -6120 9780 -5880 9800
rect -5620 9780 -5380 9800
rect -5120 9780 -4880 9800
rect -4620 9780 -4380 9800
rect -4120 9780 -3880 9800
rect -3620 9780 -3380 9800
rect -3120 9780 -3000 9800
rect -13500 9520 -13400 9780
rect -13100 9520 -12900 9780
rect -12600 9520 -12400 9780
rect -12100 9520 -11900 9780
rect -11600 9520 -11400 9780
rect -11100 9520 -10900 9780
rect -10600 9520 -10400 9780
rect -10100 9520 -9900 9780
rect -9600 9520 -9400 9780
rect -9100 9520 -8900 9780
rect -8600 9520 -8400 9780
rect -8100 9520 -7900 9780
rect -7600 9520 -7400 9780
rect -7100 9520 -6900 9780
rect -6600 9520 -6400 9780
rect -6100 9520 -5900 9780
rect -5600 9520 -5400 9780
rect -5100 9520 -4900 9780
rect -4600 9520 -4400 9780
rect -4100 9520 -3900 9780
rect -3600 9520 -3400 9780
rect -3100 9520 -3000 9780
rect -13500 9500 -13380 9520
rect -13120 9500 -12880 9520
rect -12620 9500 -12380 9520
rect -12120 9500 -11880 9520
rect -11620 9500 -11380 9520
rect -11120 9500 -10880 9520
rect -10620 9500 -10380 9520
rect -10120 9500 -9880 9520
rect -9620 9500 -9380 9520
rect -9120 9500 -8880 9520
rect -8620 9500 -8380 9520
rect -8120 9500 -7880 9520
rect -7620 9500 -7380 9520
rect -7120 9500 -6880 9520
rect -6620 9500 -6380 9520
rect -6120 9500 -5880 9520
rect -5620 9500 -5380 9520
rect -5120 9500 -4880 9520
rect -4620 9500 -4380 9520
rect -4120 9500 -3880 9520
rect -3620 9500 -3380 9520
rect -3120 9500 -3000 9520
rect -13500 9300 -3000 9500
rect -13500 9280 -13380 9300
rect -13120 9280 -12880 9300
rect -12620 9280 -12380 9300
rect -12120 9280 -11880 9300
rect -11620 9280 -11380 9300
rect -11120 9280 -10880 9300
rect -10620 9280 -10380 9300
rect -10120 9280 -9880 9300
rect -9620 9280 -9380 9300
rect -9120 9280 -8880 9300
rect -8620 9280 -8380 9300
rect -8120 9280 -7880 9300
rect -7620 9280 -7380 9300
rect -7120 9280 -6880 9300
rect -6620 9280 -6380 9300
rect -6120 9280 -5880 9300
rect -5620 9280 -5380 9300
rect -5120 9280 -4880 9300
rect -4620 9280 -4380 9300
rect -4120 9280 -3880 9300
rect -3620 9280 -3380 9300
rect -3120 9280 -3000 9300
rect -13500 9020 -13400 9280
rect -13100 9020 -12900 9280
rect -12600 9020 -12400 9280
rect -12100 9020 -11900 9280
rect -11600 9020 -11400 9280
rect -11100 9020 -10900 9280
rect -10600 9020 -10400 9280
rect -10100 9020 -9900 9280
rect -9600 9020 -9400 9280
rect -9100 9020 -8900 9280
rect -8600 9020 -8400 9280
rect -8100 9020 -7900 9280
rect -7600 9020 -7400 9280
rect -7100 9020 -6900 9280
rect -6600 9020 -6400 9280
rect -6100 9020 -5900 9280
rect -5600 9020 -5400 9280
rect -5100 9020 -4900 9280
rect -4600 9020 -4400 9280
rect -4100 9020 -3900 9280
rect -3600 9020 -3400 9280
rect -3100 9020 -3000 9280
rect -13500 9000 -13380 9020
rect -13120 9000 -12880 9020
rect -12620 9000 -12380 9020
rect -12120 9000 -11880 9020
rect -11620 9000 -11380 9020
rect -11120 9000 -10880 9020
rect -10620 9000 -10380 9020
rect -10120 9000 -9880 9020
rect -9620 9000 -9380 9020
rect -9120 9000 -8880 9020
rect -8620 9000 -8380 9020
rect -8120 9000 -7880 9020
rect -7620 9000 -7380 9020
rect -7120 9000 -6880 9020
rect -6620 9000 -6380 9020
rect -6120 9000 -5880 9020
rect -5620 9000 -5380 9020
rect -5120 9000 -4880 9020
rect -4620 9000 -4380 9020
rect -4120 9000 -3880 9020
rect -3620 9000 -3380 9020
rect -3120 9000 -3000 9020
rect -13500 8900 -3000 9000
rect -5500 8800 -3000 8900
rect -5500 8780 -5380 8800
rect -5120 8780 -4880 8800
rect -4620 8780 -4380 8800
rect -4120 8780 -3880 8800
rect -3620 8780 -3380 8800
rect -3120 8780 -3000 8800
rect -5500 8520 -5400 8780
rect -5100 8520 -4900 8780
rect -4600 8520 -4400 8780
rect -4100 8520 -3900 8780
rect -3600 8520 -3400 8780
rect -3100 8520 -3000 8780
rect -5500 8500 -5380 8520
rect -5120 8500 -4880 8520
rect -4620 8500 -4380 8520
rect -4120 8500 -3880 8520
rect -3620 8500 -3380 8520
rect -3120 8500 -3000 8520
rect -23000 8300 -15500 8400
rect -23000 8280 -22880 8300
rect -22620 8280 -22380 8300
rect -22120 8280 -21880 8300
rect -21620 8280 -21380 8300
rect -21120 8280 -20880 8300
rect -20620 8280 -20380 8300
rect -20120 8280 -19880 8300
rect -19620 8280 -19380 8300
rect -19120 8280 -18880 8300
rect -18620 8280 -18380 8300
rect -18120 8280 -17880 8300
rect -17620 8280 -17380 8300
rect -17120 8280 -16880 8300
rect -16620 8280 -16380 8300
rect -16120 8280 -15880 8300
rect -15620 8280 -15500 8300
rect -23000 8020 -22900 8280
rect -22600 8020 -22400 8280
rect -22100 8020 -21900 8280
rect -21600 8020 -21400 8280
rect -21100 8020 -20900 8280
rect -20600 8020 -20400 8280
rect -20100 8020 -19900 8280
rect -19600 8020 -19400 8280
rect -19100 8020 -18900 8280
rect -18600 8020 -18400 8280
rect -18100 8020 -17900 8280
rect -17600 8020 -17400 8280
rect -17100 8020 -16900 8280
rect -16600 8020 -16400 8280
rect -16100 8020 -15900 8280
rect -15600 8020 -15500 8280
rect -23000 8000 -22880 8020
rect -22620 8000 -22380 8020
rect -22120 8000 -21880 8020
rect -21620 8000 -21380 8020
rect -21120 8000 -20880 8020
rect -20620 8000 -20380 8020
rect -20120 8000 -19880 8020
rect -19620 8000 -19380 8020
rect -19120 8000 -18880 8020
rect -18620 8000 -18380 8020
rect -18120 8000 -17880 8020
rect -17620 8000 -17380 8020
rect -17120 8000 -16880 8020
rect -16620 8000 -16380 8020
rect -16120 8000 -15880 8020
rect -15620 8000 -15500 8020
rect -23000 7800 -15500 8000
rect -11500 8300 -7500 8400
rect -11500 8280 -11380 8300
rect -11120 8280 -10880 8300
rect -10620 8280 -10380 8300
rect -10120 8280 -9880 8300
rect -9620 8280 -9380 8300
rect -9120 8280 -8880 8300
rect -8620 8280 -8380 8300
rect -8120 8280 -7880 8300
rect -7620 8280 -7500 8300
rect -11500 8020 -11400 8280
rect -11100 8020 -10900 8280
rect -10600 8020 -10400 8280
rect -10100 8020 -9900 8280
rect -9600 8020 -9400 8280
rect -9100 8020 -8900 8280
rect -8600 8020 -8400 8280
rect -8100 8020 -7900 8280
rect -7600 8020 -7500 8280
rect -11500 8000 -11380 8020
rect -11120 8000 -10880 8020
rect -10620 8000 -10380 8020
rect -10120 8000 -9880 8020
rect -9620 8000 -9380 8020
rect -9120 8000 -8880 8020
rect -8620 8000 -8380 8020
rect -8120 8000 -7880 8020
rect -7620 8000 -7500 8020
rect -11500 7900 -7500 8000
rect -5500 8300 -3000 8500
rect -5500 8280 -5380 8300
rect -5120 8280 -4880 8300
rect -4620 8280 -4380 8300
rect -4120 8280 -3880 8300
rect -3620 8280 -3380 8300
rect -3120 8280 -3000 8300
rect -5500 8020 -5400 8280
rect -5100 8020 -4900 8280
rect -4600 8020 -4400 8280
rect -4100 8020 -3900 8280
rect -3600 8020 -3400 8280
rect -3100 8020 -3000 8280
rect -5500 8000 -5380 8020
rect -5120 8000 -4880 8020
rect -4620 8000 -4380 8020
rect -4120 8000 -3880 8020
rect -3620 8000 -3380 8020
rect -3120 8000 -3000 8020
rect -23000 7780 -22880 7800
rect -22620 7780 -22380 7800
rect -22120 7780 -21880 7800
rect -21620 7780 -21380 7800
rect -21120 7780 -20880 7800
rect -20620 7780 -20380 7800
rect -20120 7780 -19880 7800
rect -19620 7780 -19380 7800
rect -19120 7780 -18880 7800
rect -18620 7780 -18380 7800
rect -18120 7780 -17880 7800
rect -17620 7780 -17380 7800
rect -17120 7780 -16880 7800
rect -16620 7780 -16380 7800
rect -16120 7780 -15880 7800
rect -15620 7780 -15500 7800
rect -23000 7520 -22900 7780
rect -22600 7520 -22400 7780
rect -22100 7520 -21900 7780
rect -21600 7520 -21400 7780
rect -21100 7520 -20900 7780
rect -20600 7520 -20400 7780
rect -20100 7520 -19900 7780
rect -19600 7520 -19400 7780
rect -19100 7520 -18900 7780
rect -18600 7520 -18400 7780
rect -18100 7520 -17900 7780
rect -17600 7520 -17400 7780
rect -17100 7520 -16900 7780
rect -16600 7520 -16400 7780
rect -16100 7520 -15900 7780
rect -15600 7520 -15500 7780
rect -23000 7500 -22880 7520
rect -22620 7500 -22380 7520
rect -22120 7500 -21880 7520
rect -21620 7500 -21380 7520
rect -21120 7500 -20880 7520
rect -20620 7500 -20380 7520
rect -20120 7500 -19880 7520
rect -19620 7500 -19380 7520
rect -19120 7500 -18880 7520
rect -18620 7500 -18380 7520
rect -18120 7500 -17880 7520
rect -17620 7500 -17380 7520
rect -17120 7500 -16880 7520
rect -16620 7500 -16380 7520
rect -16120 7500 -15880 7520
rect -15620 7500 -15500 7520
rect -23000 7300 -15500 7500
rect -23000 7280 -22880 7300
rect -22620 7280 -22380 7300
rect -22120 7280 -21880 7300
rect -21620 7280 -21380 7300
rect -21120 7280 -20880 7300
rect -20620 7280 -20380 7300
rect -20120 7280 -19880 7300
rect -19620 7280 -19380 7300
rect -19120 7280 -18880 7300
rect -18620 7280 -18380 7300
rect -18120 7280 -17880 7300
rect -17620 7280 -17380 7300
rect -17120 7280 -16880 7300
rect -16620 7280 -16380 7300
rect -16120 7280 -15880 7300
rect -15620 7280 -15500 7300
rect -23000 7020 -22900 7280
rect -22600 7020 -22400 7280
rect -22100 7020 -21900 7280
rect -21600 7020 -21400 7280
rect -21100 7020 -20900 7280
rect -20600 7020 -20400 7280
rect -20100 7020 -19900 7280
rect -19600 7020 -19400 7280
rect -19100 7020 -18900 7280
rect -18600 7020 -18400 7280
rect -18100 7020 -17900 7280
rect -17600 7020 -17400 7280
rect -17100 7020 -16900 7280
rect -16600 7020 -16400 7280
rect -16100 7020 -15900 7280
rect -15600 7020 -15500 7280
rect -23000 7000 -22880 7020
rect -22620 7000 -22380 7020
rect -22120 7000 -21880 7020
rect -21620 7000 -21380 7020
rect -21120 7000 -20880 7020
rect -20620 7000 -20380 7020
rect -20120 7000 -19880 7020
rect -19620 7000 -19380 7020
rect -19120 7000 -18880 7020
rect -18620 7000 -18380 7020
rect -18120 7000 -17880 7020
rect -17620 7000 -17380 7020
rect -17120 7000 -16880 7020
rect -16620 7000 -16380 7020
rect -16120 7000 -15880 7020
rect -15620 7000 -15500 7020
rect -23000 6800 -15500 7000
rect -23000 6780 -22880 6800
rect -22620 6780 -22380 6800
rect -22120 6780 -21880 6800
rect -21620 6780 -21380 6800
rect -21120 6780 -20880 6800
rect -20620 6780 -20380 6800
rect -20120 6780 -19880 6800
rect -19620 6780 -19380 6800
rect -19120 6780 -18880 6800
rect -18620 6780 -18380 6800
rect -18120 6780 -17880 6800
rect -17620 6780 -17380 6800
rect -17120 6780 -16880 6800
rect -16620 6780 -16380 6800
rect -16120 6780 -15880 6800
rect -15620 6780 -15500 6800
rect -23000 6520 -22900 6780
rect -22600 6520 -22400 6780
rect -22100 6520 -21900 6780
rect -21600 6520 -21400 6780
rect -21100 6520 -20900 6780
rect -20600 6520 -20400 6780
rect -20100 6520 -19900 6780
rect -19600 6520 -19400 6780
rect -19100 6520 -18900 6780
rect -18600 6520 -18400 6780
rect -18100 6520 -17900 6780
rect -17600 6520 -17400 6780
rect -17100 6520 -16900 6780
rect -16600 6520 -16400 6780
rect -16100 6520 -15900 6780
rect -15600 6520 -15500 6780
rect -23000 6500 -22880 6520
rect -22620 6500 -22380 6520
rect -22120 6500 -21880 6520
rect -21620 6500 -21380 6520
rect -21120 6500 -20880 6520
rect -20620 6500 -20380 6520
rect -20120 6500 -19880 6520
rect -19620 6500 -19380 6520
rect -19120 6500 -18880 6520
rect -18620 6500 -18380 6520
rect -18120 6500 -17880 6520
rect -17620 6500 -17380 6520
rect -17120 6500 -16880 6520
rect -16620 6500 -16380 6520
rect -16120 6500 -15880 6520
rect -15620 6500 -15500 6520
rect -23000 6300 -15500 6500
rect -23000 6280 -22880 6300
rect -22620 6280 -22380 6300
rect -22120 6280 -21880 6300
rect -21620 6280 -21380 6300
rect -21120 6280 -20880 6300
rect -20620 6280 -20380 6300
rect -20120 6280 -19880 6300
rect -19620 6280 -19380 6300
rect -19120 6280 -18880 6300
rect -18620 6280 -18380 6300
rect -18120 6280 -17880 6300
rect -17620 6280 -17380 6300
rect -17120 6280 -16880 6300
rect -16620 6280 -16380 6300
rect -16120 6280 -15880 6300
rect -15620 6280 -15500 6300
rect -23000 6020 -22900 6280
rect -22600 6020 -22400 6280
rect -22100 6020 -21900 6280
rect -21600 6020 -21400 6280
rect -21100 6020 -20900 6280
rect -20600 6020 -20400 6280
rect -20100 6020 -19900 6280
rect -19600 6020 -19400 6280
rect -19100 6020 -18900 6280
rect -18600 6020 -18400 6280
rect -18100 6020 -17900 6280
rect -17600 6020 -17400 6280
rect -17100 6020 -16900 6280
rect -16600 6020 -16400 6280
rect -16100 6020 -15900 6280
rect -15600 6020 -15500 6280
rect -23000 6000 -22880 6020
rect -22620 6000 -22380 6020
rect -22120 6000 -21880 6020
rect -21620 6000 -21380 6020
rect -21120 6000 -20880 6020
rect -20620 6000 -20380 6020
rect -20120 6000 -19880 6020
rect -19620 6000 -19380 6020
rect -19120 6000 -18880 6020
rect -18620 6000 -18380 6020
rect -18120 6000 -17880 6020
rect -17620 6000 -17380 6020
rect -17120 6000 -16880 6020
rect -16620 6000 -16380 6020
rect -16120 6000 -15880 6020
rect -15620 6000 -15500 6020
rect -23000 5900 -15500 6000
rect -5500 7800 -3000 8000
rect -5500 7780 -5380 7800
rect -5120 7780 -4880 7800
rect -4620 7780 -4380 7800
rect -4120 7780 -3880 7800
rect -3620 7780 -3380 7800
rect -3120 7780 -3000 7800
rect -5500 7520 -5400 7780
rect -5100 7520 -4900 7780
rect -4600 7520 -4400 7780
rect -4100 7520 -3900 7780
rect -3600 7520 -3400 7780
rect -3100 7520 -3000 7780
rect -5500 7500 -5380 7520
rect -5120 7500 -4880 7520
rect -4620 7500 -4380 7520
rect -4120 7500 -3880 7520
rect -3620 7500 -3380 7520
rect -3120 7500 -3000 7520
rect -5500 7300 -3000 7500
rect -5500 7280 -5380 7300
rect -5120 7280 -4880 7300
rect -4620 7280 -4380 7300
rect -4120 7280 -3880 7300
rect -3620 7280 -3380 7300
rect -3120 7280 -3000 7300
rect -5500 7020 -5400 7280
rect -5100 7020 -4900 7280
rect -4600 7020 -4400 7280
rect -4100 7020 -3900 7280
rect -3600 7020 -3400 7280
rect -3100 7020 -3000 7280
rect -5500 7000 -5380 7020
rect -5120 7000 -4880 7020
rect -4620 7000 -4380 7020
rect -4120 7000 -3880 7020
rect -3620 7000 -3380 7020
rect -3120 7000 -3000 7020
rect -5500 6800 -3000 7000
rect -5500 6780 -5380 6800
rect -5120 6780 -4880 6800
rect -4620 6780 -4380 6800
rect -4120 6780 -3880 6800
rect -3620 6780 -3380 6800
rect -3120 6780 -3000 6800
rect -5500 6520 -5400 6780
rect -5100 6520 -4900 6780
rect -4600 6520 -4400 6780
rect -4100 6520 -3900 6780
rect -3600 6520 -3400 6780
rect -3100 6520 -3000 6780
rect -5500 6500 -5380 6520
rect -5120 6500 -4880 6520
rect -4620 6500 -4380 6520
rect -4120 6500 -3880 6520
rect -3620 6500 -3380 6520
rect -3120 6500 -3000 6520
rect -5500 6300 -3000 6500
rect -5500 6280 -5380 6300
rect -5120 6280 -4880 6300
rect -4620 6280 -4380 6300
rect -4120 6280 -3880 6300
rect -3620 6280 -3380 6300
rect -3120 6280 -3000 6300
rect -5500 6020 -5400 6280
rect -5100 6020 -4900 6280
rect -4600 6020 -4400 6280
rect -4100 6020 -3900 6280
rect -3600 6020 -3400 6280
rect -3100 6020 -3000 6280
rect -5500 6000 -5380 6020
rect -5120 6000 -4880 6020
rect -4620 6000 -4380 6020
rect -4120 6000 -3880 6020
rect -3620 6000 -3380 6020
rect -3120 6000 -3000 6020
rect -5500 5900 -3000 6000
rect -23000 5800 -21000 5900
rect -23000 5780 -22880 5800
rect -22620 5780 -22380 5800
rect -22120 5780 -21880 5800
rect -21620 5780 -21380 5800
rect -21120 5780 -21000 5800
rect -23000 5520 -22900 5780
rect -22600 5520 -22400 5780
rect -22100 5520 -21900 5780
rect -21600 5520 -21400 5780
rect -21100 5520 -21000 5780
rect -23000 5500 -22880 5520
rect -22620 5500 -22380 5520
rect -22120 5500 -21880 5520
rect -21620 5500 -21380 5520
rect -21120 5500 -21000 5520
rect -23000 5300 -21000 5500
rect -23000 5280 -22880 5300
rect -22620 5280 -22380 5300
rect -22120 5280 -21880 5300
rect -21620 5280 -21380 5300
rect -21120 5280 -21000 5300
rect -23000 5020 -22900 5280
rect -22600 5020 -22400 5280
rect -22100 5020 -21900 5280
rect -21600 5020 -21400 5280
rect -21100 5020 -21000 5280
rect -23000 5000 -22880 5020
rect -22620 5000 -22380 5020
rect -22120 5000 -21880 5020
rect -21620 5000 -21380 5020
rect -21120 5000 -21000 5020
rect -23000 4900 -21000 5000
rect -25000 4800 -21000 4900
rect -25000 4780 -24880 4800
rect -24620 4780 -24380 4800
rect -24120 4780 -23880 4800
rect -23620 4780 -23380 4800
rect -23120 4780 -22880 4800
rect -22620 4780 -22380 4800
rect -22120 4780 -21880 4800
rect -21620 4780 -21380 4800
rect -21120 4780 -21000 4800
rect -25000 4520 -24900 4780
rect -24600 4520 -24400 4780
rect -24100 4520 -23900 4780
rect -23600 4520 -23400 4780
rect -23100 4520 -22900 4780
rect -22600 4520 -22400 4780
rect -22100 4520 -21900 4780
rect -21600 4520 -21400 4780
rect -21100 4520 -21000 4780
rect -25000 4500 -24880 4520
rect -24620 4500 -24380 4520
rect -24120 4500 -23880 4520
rect -23620 4500 -23380 4520
rect -23120 4500 -22880 4520
rect -22620 4500 -22380 4520
rect -22120 4500 -21880 4520
rect -21620 4500 -21380 4520
rect -21120 4500 -21000 4520
rect -25000 4300 -21000 4500
rect -25000 4280 -24880 4300
rect -24620 4280 -24380 4300
rect -24120 4280 -23880 4300
rect -23620 4280 -23380 4300
rect -23120 4280 -22880 4300
rect -22620 4280 -22380 4300
rect -22120 4280 -21880 4300
rect -21620 4280 -21380 4300
rect -21120 4280 -21000 4300
rect -25000 4020 -24900 4280
rect -24600 4020 -24400 4280
rect -24100 4020 -23900 4280
rect -23600 4020 -23400 4280
rect -23100 4020 -22900 4280
rect -22600 4020 -22400 4280
rect -22100 4020 -21900 4280
rect -21600 4020 -21400 4280
rect -21100 4020 -21000 4280
rect -25000 4000 -24880 4020
rect -24620 4000 -24380 4020
rect -24120 4000 -23880 4020
rect -23620 4000 -23380 4020
rect -23120 4000 -22880 4020
rect -22620 4000 -22380 4020
rect -22120 4000 -21880 4020
rect -21620 4000 -21380 4020
rect -21120 4000 -21000 4020
rect -25000 3800 -21000 4000
rect -5000 5300 -3700 5400
rect -5000 4300 -4800 5300
rect -5000 3900 -3500 4300
rect -25000 3780 -24880 3800
rect -24620 3780 -24380 3800
rect -24120 3780 -23880 3800
rect -23620 3780 -23380 3800
rect -23120 3780 -22880 3800
rect -22620 3780 -22380 3800
rect -22120 3780 -21880 3800
rect -21620 3780 -21380 3800
rect -21120 3780 -21000 3800
rect -25000 3520 -24900 3780
rect -24600 3520 -24400 3780
rect -24100 3520 -23900 3780
rect -23600 3520 -23400 3780
rect -23100 3520 -22900 3780
rect -22600 3520 -22400 3780
rect -22100 3520 -21900 3780
rect -21600 3520 -21400 3780
rect -21100 3520 -21000 3780
rect -25000 3500 -24880 3520
rect -24620 3500 -24380 3520
rect -24120 3500 -23880 3520
rect -23620 3500 -23380 3520
rect -23120 3500 -22880 3520
rect -22620 3500 -22380 3520
rect -22120 3500 -21880 3520
rect -21620 3500 -21380 3520
rect -21120 3500 -21000 3520
rect -25000 3300 -21000 3500
rect -25000 3280 -24880 3300
rect -24620 3280 -24380 3300
rect -24120 3280 -23880 3300
rect -23620 3280 -23380 3300
rect -23120 3280 -22880 3300
rect -22620 3280 -22380 3300
rect -22120 3280 -21880 3300
rect -21620 3280 -21380 3300
rect -21120 3280 -21000 3300
rect -25000 3020 -24900 3280
rect -24600 3020 -24400 3280
rect -24100 3020 -23900 3280
rect -23600 3020 -23400 3280
rect -23100 3020 -22900 3280
rect -22600 3020 -22400 3280
rect -22100 3020 -21900 3280
rect -21600 3020 -21400 3280
rect -21100 3020 -21000 3280
rect -25000 3000 -24880 3020
rect -24620 3000 -24380 3020
rect -24120 3000 -23880 3020
rect -23620 3000 -23380 3020
rect -23120 3000 -22880 3020
rect -22620 3000 -22380 3020
rect -22120 3000 -21880 3020
rect -21620 3000 -21380 3020
rect -21120 3000 -21000 3020
rect -25000 2800 -21000 3000
rect -25000 2780 -24880 2800
rect -24620 2780 -24380 2800
rect -24120 2780 -23880 2800
rect -23620 2780 -23380 2800
rect -23120 2780 -22880 2800
rect -22620 2780 -22380 2800
rect -22120 2780 -21880 2800
rect -21620 2780 -21380 2800
rect -21120 2780 -21000 2800
rect -25000 2520 -24900 2780
rect -24600 2520 -24400 2780
rect -24100 2520 -23900 2780
rect -23600 2520 -23400 2780
rect -23100 2520 -22900 2780
rect -22600 2520 -22400 2780
rect -22100 2520 -21900 2780
rect -21600 2520 -21400 2780
rect -21100 2520 -21000 2780
rect -25000 2500 -24880 2520
rect -24620 2500 -24380 2520
rect -24120 2500 -23880 2520
rect -23620 2500 -23380 2520
rect -23120 2500 -22880 2520
rect -22620 2500 -22380 2520
rect -22120 2500 -21880 2520
rect -21620 2500 -21380 2520
rect -21120 2500 -21000 2520
rect -25000 2300 -21000 2500
rect -25000 2280 -24880 2300
rect -24620 2280 -24380 2300
rect -24120 2280 -23880 2300
rect -23620 2280 -23380 2300
rect -23120 2280 -22880 2300
rect -22620 2280 -22380 2300
rect -22120 2280 -21880 2300
rect -21620 2280 -21380 2300
rect -21120 2280 -21000 2300
rect -25000 2020 -24900 2280
rect -24600 2020 -24400 2280
rect -24100 2020 -23900 2280
rect -23600 2020 -23400 2280
rect -23100 2020 -22900 2280
rect -22600 2020 -22400 2280
rect -22100 2020 -21900 2280
rect -21600 2020 -21400 2280
rect -21100 2020 -21000 2280
rect -25000 2000 -24880 2020
rect -24620 2000 -24380 2020
rect -24120 2000 -23880 2020
rect -23620 2000 -23380 2020
rect -23120 2000 -22880 2020
rect -22620 2000 -22380 2020
rect -22120 2000 -21880 2020
rect -21620 2000 -21380 2020
rect -21120 2000 -21000 2020
rect -25000 1800 -21000 2000
rect -25000 1780 -24880 1800
rect -24620 1780 -24380 1800
rect -24120 1780 -23880 1800
rect -23620 1780 -23380 1800
rect -23120 1780 -22880 1800
rect -22620 1780 -22380 1800
rect -22120 1780 -21880 1800
rect -21620 1780 -21380 1800
rect -21120 1780 -21000 1800
rect -25000 1520 -24900 1780
rect -24600 1520 -24400 1780
rect -24100 1520 -23900 1780
rect -23600 1520 -23400 1780
rect -23100 1520 -22900 1780
rect -22600 1520 -22400 1780
rect -22100 1520 -21900 1780
rect -21600 1520 -21400 1780
rect -21100 1520 -21000 1780
rect -25000 1500 -24880 1520
rect -24620 1500 -24380 1520
rect -24120 1500 -23880 1520
rect -23620 1500 -23380 1520
rect -23120 1500 -22880 1520
rect -22620 1500 -22380 1520
rect -22120 1500 -21880 1520
rect -21620 1500 -21380 1520
rect -21120 1500 -21000 1520
rect -25000 1300 -21000 1500
rect -25000 1280 -24880 1300
rect -24620 1280 -24380 1300
rect -24120 1280 -23880 1300
rect -23620 1280 -23380 1300
rect -23120 1280 -22880 1300
rect -22620 1280 -22380 1300
rect -22120 1280 -21880 1300
rect -21620 1280 -21380 1300
rect -21120 1280 -21000 1300
rect -25000 1020 -24900 1280
rect -24600 1020 -24400 1280
rect -24100 1020 -23900 1280
rect -23600 1020 -23400 1280
rect -23100 1020 -22900 1280
rect -22600 1020 -22400 1280
rect -22100 1020 -21900 1280
rect -21600 1020 -21400 1280
rect -21100 1020 -21000 1280
rect -25000 1000 -24880 1020
rect -24620 1000 -24380 1020
rect -24120 1000 -23880 1020
rect -23620 1000 -23380 1020
rect -23120 1000 -22880 1020
rect -22620 1000 -22380 1020
rect -22120 1000 -21880 1020
rect -21620 1000 -21380 1020
rect -21120 1000 -21000 1020
rect -25000 800 -21000 1000
rect -25000 780 -24880 800
rect -24620 780 -24380 800
rect -24120 780 -23880 800
rect -23620 780 -23380 800
rect -23120 780 -22880 800
rect -22620 780 -22380 800
rect -22120 780 -21880 800
rect -21620 780 -21380 800
rect -21120 780 -21000 800
rect -25000 520 -24900 780
rect -24600 520 -24400 780
rect -24100 520 -23900 780
rect -23600 520 -23400 780
rect -23100 520 -22900 780
rect -22600 520 -22400 780
rect -22100 520 -21900 780
rect -21600 520 -21400 780
rect -21100 520 -21000 780
rect -25000 500 -24880 520
rect -24620 500 -24380 520
rect -24120 500 -23880 520
rect -23620 500 -23380 520
rect -23120 500 -22880 520
rect -22620 500 -22380 520
rect -22120 500 -21880 520
rect -21620 500 -21380 520
rect -21120 500 -21000 520
rect -25000 300 -21000 500
rect 13000 2300 15500 2400
rect 13000 2280 13120 2300
rect 13380 2280 13620 2300
rect 13880 2280 14120 2300
rect 14380 2280 14620 2300
rect 14880 2280 15120 2300
rect 15380 2280 15500 2300
rect 13000 2020 13100 2280
rect 13400 2020 13600 2280
rect 13900 2020 14100 2280
rect 14400 2020 14600 2280
rect 14900 2020 15100 2280
rect 15400 2020 15500 2280
rect 13000 2000 13120 2020
rect 13380 2000 13620 2020
rect 13880 2000 14120 2020
rect 14380 2000 14620 2020
rect 14880 2000 15120 2020
rect 15380 2000 15500 2020
rect 13000 1800 15500 2000
rect 13000 1780 13120 1800
rect 13380 1780 13620 1800
rect 13880 1780 14120 1800
rect 14380 1780 14620 1800
rect 14880 1780 15120 1800
rect 15380 1780 15500 1800
rect 13000 1520 13100 1780
rect 13400 1520 13600 1780
rect 13900 1520 14100 1780
rect 14400 1520 14600 1780
rect 14900 1520 15100 1780
rect 15400 1520 15500 1780
rect 13000 1500 13120 1520
rect 13380 1500 13620 1520
rect 13880 1500 14120 1520
rect 14380 1500 14620 1520
rect 14880 1500 15120 1520
rect 15380 1500 15500 1520
rect 13000 1300 15500 1500
rect 13000 1280 13120 1300
rect 13380 1280 13620 1300
rect 13880 1280 14120 1300
rect 14380 1280 14620 1300
rect 14880 1280 15120 1300
rect 15380 1280 15500 1300
rect 13000 1020 13100 1280
rect 13400 1020 13600 1280
rect 13900 1020 14100 1280
rect 14400 1020 14600 1280
rect 14900 1020 15100 1280
rect 15400 1020 15500 1280
rect 13000 1000 13120 1020
rect 13380 1000 13620 1020
rect 13880 1000 14120 1020
rect 14380 1000 14620 1020
rect 14880 1000 15120 1020
rect 15380 1000 15500 1020
rect 13000 800 15500 1000
rect 13000 780 13120 800
rect 13380 780 13620 800
rect 13880 780 14120 800
rect 14380 780 14620 800
rect 14880 780 15120 800
rect 15380 780 15500 800
rect 13000 520 13100 780
rect 13400 520 13600 780
rect 13900 520 14100 780
rect 14400 520 14600 780
rect 14900 520 15100 780
rect 15400 520 15500 780
rect 13000 500 13120 520
rect 13380 500 13620 520
rect 13880 500 14120 520
rect 14380 500 14620 520
rect 14880 500 15120 520
rect 15380 500 15500 520
rect 13000 400 15500 500
rect 17500 1300 19500 1400
rect 17500 1280 17620 1300
rect 17880 1280 18120 1300
rect 18380 1280 18620 1300
rect 18880 1280 19120 1300
rect 19380 1280 19500 1300
rect 17500 1020 17600 1280
rect 17900 1020 18100 1280
rect 18400 1020 18600 1280
rect 18900 1020 19100 1280
rect 19400 1020 19500 1280
rect 17500 1000 17620 1020
rect 17880 1000 18120 1020
rect 18380 1000 18620 1020
rect 18880 1000 19120 1020
rect 19380 1000 19500 1020
rect 17500 800 19500 1000
rect 17500 780 17620 800
rect 17880 780 18120 800
rect 18380 780 18620 800
rect 18880 780 19120 800
rect 19380 780 19500 800
rect 17500 520 17600 780
rect 17900 520 18100 780
rect 18400 520 18600 780
rect 18900 520 19100 780
rect 19400 520 19500 780
rect 17500 500 17620 520
rect 17880 500 18120 520
rect 18380 500 18620 520
rect 18880 500 19120 520
rect 19380 500 19500 520
rect -25000 280 -24880 300
rect -24620 280 -24380 300
rect -24120 280 -23880 300
rect -23620 280 -23380 300
rect -23120 280 -22880 300
rect -22620 280 -22380 300
rect -22120 280 -21880 300
rect -21620 280 -21380 300
rect -21120 280 -21000 300
rect -25000 20 -24900 280
rect -24600 20 -24400 280
rect -24100 20 -23900 280
rect -23600 20 -23400 280
rect -23100 20 -22900 280
rect -22600 20 -22400 280
rect -22100 20 -21900 280
rect -21600 20 -21400 280
rect -21100 20 -21000 280
rect -25000 0 -24880 20
rect -24620 0 -24380 20
rect -24120 0 -23880 20
rect -23620 0 -23380 20
rect -23120 0 -22880 20
rect -22620 0 -22380 20
rect -22120 0 -21880 20
rect -21620 0 -21380 20
rect -21120 0 -21000 20
rect -25000 -200 -21000 0
rect -25000 -220 -24880 -200
rect -24620 -220 -24380 -200
rect -24120 -220 -23880 -200
rect -23620 -220 -23380 -200
rect -23120 -220 -22880 -200
rect -22620 -220 -22380 -200
rect -22120 -220 -21880 -200
rect -21620 -220 -21380 -200
rect -21120 -220 -21000 -200
rect -25000 -480 -24900 -220
rect -24600 -480 -24400 -220
rect -24100 -480 -23900 -220
rect -23600 -480 -23400 -220
rect -23100 -480 -22900 -220
rect -22600 -480 -22400 -220
rect -22100 -480 -21900 -220
rect -21600 -480 -21400 -220
rect -21100 -480 -21000 -220
rect -25000 -500 -24880 -480
rect -24620 -500 -24380 -480
rect -24120 -500 -23880 -480
rect -23620 -500 -23380 -480
rect -23120 -500 -22880 -480
rect -22620 -500 -22380 -480
rect -22120 -500 -21880 -480
rect -21620 -500 -21380 -480
rect -21120 -500 -21000 -480
rect -25000 -700 -21000 -500
rect -25000 -720 -24880 -700
rect -24620 -720 -24380 -700
rect -24120 -720 -23880 -700
rect -23620 -720 -23380 -700
rect -23120 -720 -22880 -700
rect -22620 -720 -22380 -700
rect -22120 -720 -21880 -700
rect -21620 -720 -21380 -700
rect -21120 -720 -21000 -700
rect -25000 -980 -24900 -720
rect -24600 -980 -24400 -720
rect -24100 -980 -23900 -720
rect -23600 -980 -23400 -720
rect -23100 -980 -22900 -720
rect -22600 -980 -22400 -720
rect -22100 -980 -21900 -720
rect -21600 -980 -21400 -720
rect -21100 -980 -21000 -720
rect -25000 -1000 -24880 -980
rect -24620 -1000 -24380 -980
rect -24120 -1000 -23880 -980
rect -23620 -1000 -23380 -980
rect -23120 -1000 -22880 -980
rect -22620 -1000 -22380 -980
rect -22120 -1000 -21880 -980
rect -21620 -1000 -21380 -980
rect -21120 -1000 -21000 -980
rect -25000 -1200 -21000 -1000
rect -25000 -1220 -24880 -1200
rect -24620 -1220 -24380 -1200
rect -24120 -1220 -23880 -1200
rect -23620 -1220 -23380 -1200
rect -23120 -1220 -22880 -1200
rect -22620 -1220 -22380 -1200
rect -22120 -1220 -21880 -1200
rect -21620 -1220 -21380 -1200
rect -21120 -1220 -21000 -1200
rect -25000 -1480 -24900 -1220
rect -24600 -1480 -24400 -1220
rect -24100 -1480 -23900 -1220
rect -23600 -1480 -23400 -1220
rect -23100 -1480 -22900 -1220
rect -22600 -1480 -22400 -1220
rect -22100 -1480 -21900 -1220
rect -21600 -1480 -21400 -1220
rect -21100 -1480 -21000 -1220
rect -25000 -1500 -24880 -1480
rect -24620 -1500 -24380 -1480
rect -24120 -1500 -23880 -1480
rect -23620 -1500 -23380 -1480
rect -23120 -1500 -22880 -1480
rect -22620 -1500 -22380 -1480
rect -22120 -1500 -21880 -1480
rect -21620 -1500 -21380 -1480
rect -21120 -1500 -21000 -1480
rect -25000 -1700 -21000 -1500
rect -25000 -1720 -24880 -1700
rect -24620 -1720 -24380 -1700
rect -24120 -1720 -23880 -1700
rect -23620 -1720 -23380 -1700
rect -23120 -1720 -22880 -1700
rect -22620 -1720 -22380 -1700
rect -22120 -1720 -21880 -1700
rect -21620 -1720 -21380 -1700
rect -21120 -1720 -21000 -1700
rect -25000 -1980 -24900 -1720
rect -24600 -1980 -24400 -1720
rect -24100 -1980 -23900 -1720
rect -23600 -1980 -23400 -1720
rect -23100 -1980 -22900 -1720
rect -22600 -1980 -22400 -1720
rect -22100 -1980 -21900 -1720
rect -21600 -1980 -21400 -1720
rect -21100 -1980 -21000 -1720
rect -25000 -2000 -24880 -1980
rect -24620 -2000 -24380 -1980
rect -24120 -2000 -23880 -1980
rect -23620 -2000 -23380 -1980
rect -23120 -2000 -22880 -1980
rect -22620 -2000 -22380 -1980
rect -22120 -2000 -21880 -1980
rect -21620 -2000 -21380 -1980
rect -21120 -2000 -21000 -1980
rect -25000 -2200 -21000 -2000
rect -25000 -2220 -24880 -2200
rect -24620 -2220 -24380 -2200
rect -24120 -2220 -23880 -2200
rect -23620 -2220 -23380 -2200
rect -23120 -2220 -22880 -2200
rect -22620 -2220 -22380 -2200
rect -22120 -2220 -21880 -2200
rect -21620 -2220 -21380 -2200
rect -21120 -2220 -21000 -2200
rect -25000 -2480 -24900 -2220
rect -24600 -2480 -24400 -2220
rect -24100 -2480 -23900 -2220
rect -23600 -2480 -23400 -2220
rect -23100 -2480 -22900 -2220
rect -22600 -2480 -22400 -2220
rect -22100 -2480 -21900 -2220
rect -21600 -2480 -21400 -2220
rect -21100 -2480 -21000 -2220
rect -25000 -2500 -24880 -2480
rect -24620 -2500 -24380 -2480
rect -24120 -2500 -23880 -2480
rect -23620 -2500 -23380 -2480
rect -23120 -2500 -22880 -2480
rect -22620 -2500 -22380 -2480
rect -22120 -2500 -21880 -2480
rect -21620 -2500 -21380 -2480
rect -21120 -2500 -21000 -2480
rect -25000 -2700 -21000 -2500
rect -25000 -2720 -24880 -2700
rect -24620 -2720 -24380 -2700
rect -24120 -2720 -23880 -2700
rect -23620 -2720 -23380 -2700
rect -23120 -2720 -22880 -2700
rect -22620 -2720 -22380 -2700
rect -22120 -2720 -21880 -2700
rect -21620 -2720 -21380 -2700
rect -21120 -2720 -21000 -2700
rect -25000 -2980 -24900 -2720
rect -24600 -2980 -24400 -2720
rect -24100 -2980 -23900 -2720
rect -23600 -2980 -23400 -2720
rect -23100 -2980 -22900 -2720
rect -22600 -2980 -22400 -2720
rect -22100 -2980 -21900 -2720
rect -21600 -2980 -21400 -2720
rect -21100 -2980 -21000 -2720
rect -25000 -3000 -24880 -2980
rect -24620 -3000 -24380 -2980
rect -24120 -3000 -23880 -2980
rect -23620 -3000 -23380 -2980
rect -23120 -3000 -22880 -2980
rect -22620 -3000 -22380 -2980
rect -22120 -3000 -21880 -2980
rect -21620 -3000 -21380 -2980
rect -21120 -3000 -21000 -2980
rect -25000 -3100 -21000 -3000
rect 12000 300 17000 400
rect 12000 280 12120 300
rect 12380 280 12620 300
rect 12880 280 13120 300
rect 13380 280 13620 300
rect 13880 280 14120 300
rect 14380 280 14620 300
rect 14880 280 15120 300
rect 15380 280 15620 300
rect 15880 280 16120 300
rect 16380 280 16620 300
rect 16880 280 17000 300
rect 12000 20 12100 280
rect 12400 20 12600 280
rect 12900 20 13100 280
rect 13400 20 13600 280
rect 13900 20 14100 280
rect 14400 20 14600 280
rect 14900 20 15100 280
rect 15400 20 15600 280
rect 15900 20 16100 280
rect 16400 20 16600 280
rect 16900 20 17000 280
rect 12000 0 12120 20
rect 12380 0 12620 20
rect 12880 0 13120 20
rect 13380 0 13620 20
rect 13880 0 14120 20
rect 14380 0 14620 20
rect 14880 0 15120 20
rect 15380 0 15620 20
rect 15880 0 16120 20
rect 16380 0 16620 20
rect 16880 0 17000 20
rect 12000 -200 17000 0
rect 12000 -220 12120 -200
rect 12380 -220 12620 -200
rect 12880 -220 13120 -200
rect 13380 -220 13620 -200
rect 13880 -220 14120 -200
rect 14380 -220 14620 -200
rect 14880 -220 15120 -200
rect 15380 -220 15620 -200
rect 15880 -220 16120 -200
rect 16380 -220 16620 -200
rect 16880 -220 17000 -200
rect 12000 -480 12100 -220
rect 12400 -480 12600 -220
rect 12900 -480 13100 -220
rect 13400 -480 13600 -220
rect 13900 -480 14100 -220
rect 14400 -480 14600 -220
rect 14900 -480 15100 -220
rect 15400 -480 15600 -220
rect 15900 -480 16100 -220
rect 16400 -480 16600 -220
rect 16900 -480 17000 -220
rect 12000 -500 12120 -480
rect 12380 -500 12620 -480
rect 12880 -500 13120 -480
rect 13380 -500 13620 -480
rect 13880 -500 14120 -480
rect 14380 -500 14620 -480
rect 14880 -500 15120 -480
rect 15380 -500 15620 -480
rect 15880 -500 16120 -480
rect 16380 -500 16620 -480
rect 16880 -500 17000 -480
rect 12000 -700 17000 -500
rect 12000 -720 12120 -700
rect 12380 -720 12620 -700
rect 12880 -720 13120 -700
rect 13380 -720 13620 -700
rect 13880 -720 14120 -700
rect 14380 -720 14620 -700
rect 14880 -720 15120 -700
rect 15380 -720 15620 -700
rect 15880 -720 16120 -700
rect 16380 -720 16620 -700
rect 16880 -720 17000 -700
rect 12000 -980 12100 -720
rect 12400 -980 12600 -720
rect 12900 -980 13100 -720
rect 13400 -980 13600 -720
rect 13900 -980 14100 -720
rect 14400 -980 14600 -720
rect 14900 -980 15100 -720
rect 15400 -980 15600 -720
rect 15900 -980 16100 -720
rect 16400 -980 16600 -720
rect 16900 -980 17000 -720
rect 12000 -1000 12120 -980
rect 12380 -1000 12620 -980
rect 12880 -1000 13120 -980
rect 13380 -1000 13620 -980
rect 13880 -1000 14120 -980
rect 14380 -1000 14620 -980
rect 14880 -1000 15120 -980
rect 15380 -1000 15620 -980
rect 15880 -1000 16120 -980
rect 16380 -1000 16620 -980
rect 16880 -1000 17000 -980
rect 12000 -1200 17000 -1000
rect 12000 -1220 12120 -1200
rect 12380 -1220 12620 -1200
rect 12880 -1220 13120 -1200
rect 13380 -1220 13620 -1200
rect 13880 -1220 14120 -1200
rect 14380 -1220 14620 -1200
rect 14880 -1220 15120 -1200
rect 15380 -1220 15620 -1200
rect 15880 -1220 16120 -1200
rect 16380 -1220 16620 -1200
rect 16880 -1220 17000 -1200
rect 12000 -1480 12100 -1220
rect 12400 -1480 12600 -1220
rect 12900 -1480 13100 -1220
rect 13400 -1480 13600 -1220
rect 13900 -1480 14100 -1220
rect 14400 -1480 14600 -1220
rect 14900 -1480 15100 -1220
rect 15400 -1480 15600 -1220
rect 15900 -1480 16100 -1220
rect 16400 -1480 16600 -1220
rect 16900 -1480 17000 -1220
rect 12000 -1500 12120 -1480
rect 12380 -1500 12620 -1480
rect 12880 -1500 13120 -1480
rect 13380 -1500 13620 -1480
rect 13880 -1500 14120 -1480
rect 14380 -1500 14620 -1480
rect 14880 -1500 15120 -1480
rect 15380 -1500 15620 -1480
rect 15880 -1500 16120 -1480
rect 16380 -1500 16620 -1480
rect 16880 -1500 17000 -1480
rect 12000 -1700 17000 -1500
rect 12000 -1720 12120 -1700
rect 12380 -1720 12620 -1700
rect 12880 -1720 13120 -1700
rect 13380 -1720 13620 -1700
rect 13880 -1720 14120 -1700
rect 14380 -1720 14620 -1700
rect 14880 -1720 15120 -1700
rect 15380 -1720 15620 -1700
rect 15880 -1720 16120 -1700
rect 16380 -1720 16620 -1700
rect 16880 -1720 17000 -1700
rect 12000 -1980 12100 -1720
rect 12400 -1980 12600 -1720
rect 12900 -1980 13100 -1720
rect 13400 -1980 13600 -1720
rect 13900 -1980 14100 -1720
rect 14400 -1980 14600 -1720
rect 14900 -1980 15100 -1720
rect 15400 -1980 15600 -1720
rect 15900 -1980 16100 -1720
rect 16400 -1980 16600 -1720
rect 16900 -1980 17000 -1720
rect 12000 -2000 12120 -1980
rect 12380 -2000 12620 -1980
rect 12880 -2000 13120 -1980
rect 13380 -2000 13620 -1980
rect 13880 -2000 14120 -1980
rect 14380 -2000 14620 -1980
rect 14880 -2000 15120 -1980
rect 15380 -2000 15620 -1980
rect 15880 -2000 16120 -1980
rect 16380 -2000 16620 -1980
rect 16880 -2000 17000 -1980
rect 12000 -2200 17000 -2000
rect 12000 -2220 12120 -2200
rect 12380 -2220 12620 -2200
rect 12880 -2220 13120 -2200
rect 13380 -2220 13620 -2200
rect 13880 -2220 14120 -2200
rect 14380 -2220 14620 -2200
rect 14880 -2220 15120 -2200
rect 15380 -2220 15620 -2200
rect 15880 -2220 16120 -2200
rect 16380 -2220 16620 -2200
rect 16880 -2220 17000 -2200
rect 12000 -2480 12100 -2220
rect 12400 -2480 12600 -2220
rect 12900 -2480 13100 -2220
rect 13400 -2480 13600 -2220
rect 13900 -2480 14100 -2220
rect 14400 -2480 14600 -2220
rect 14900 -2480 15100 -2220
rect 15400 -2480 15600 -2220
rect 15900 -2480 16100 -2220
rect 16400 -2480 16600 -2220
rect 16900 -2480 17000 -2220
rect 12000 -2500 12120 -2480
rect 12380 -2500 12620 -2480
rect 12880 -2500 13120 -2480
rect 13380 -2500 13620 -2480
rect 13880 -2500 14120 -2480
rect 14380 -2500 14620 -2480
rect 14880 -2500 15120 -2480
rect 15380 -2500 15620 -2480
rect 15880 -2500 16120 -2480
rect 16380 -2500 16620 -2480
rect 16880 -2500 17000 -2480
rect 12000 -2700 17000 -2500
rect 12000 -2720 12120 -2700
rect 12380 -2720 12620 -2700
rect 12880 -2720 13120 -2700
rect 13380 -2720 13620 -2700
rect 13880 -2720 14120 -2700
rect 14380 -2720 14620 -2700
rect 14880 -2720 15120 -2700
rect 15380 -2720 15620 -2700
rect 15880 -2720 16120 -2700
rect 16380 -2720 16620 -2700
rect 16880 -2720 17000 -2700
rect 12000 -2980 12100 -2720
rect 12400 -2980 12600 -2720
rect 12900 -2980 13100 -2720
rect 13400 -2980 13600 -2720
rect 13900 -2980 14100 -2720
rect 14400 -2980 14600 -2720
rect 14900 -2980 15100 -2720
rect 15400 -2980 15600 -2720
rect 15900 -2980 16100 -2720
rect 16400 -2980 16600 -2720
rect 16900 -2980 17000 -2720
rect 12000 -3000 12120 -2980
rect 12380 -3000 12620 -2980
rect 12880 -3000 13120 -2980
rect 13380 -3000 13620 -2980
rect 13880 -3000 14120 -2980
rect 14380 -3000 14620 -2980
rect 14880 -3000 15120 -2980
rect 15380 -3000 15620 -2980
rect 15880 -3000 16120 -2980
rect 16380 -3000 16620 -2980
rect 16880 -3000 17000 -2980
rect -23500 -3200 -14500 -3100
rect -23500 -3220 -23380 -3200
rect -23120 -3220 -22880 -3200
rect -22620 -3220 -22380 -3200
rect -22120 -3220 -21880 -3200
rect -21620 -3220 -21380 -3200
rect -21120 -3220 -20880 -3200
rect -20620 -3220 -20380 -3200
rect -20120 -3220 -19880 -3200
rect -19620 -3220 -19380 -3200
rect -19120 -3220 -18880 -3200
rect -18620 -3220 -18380 -3200
rect -18120 -3220 -17880 -3200
rect -17620 -3220 -17380 -3200
rect -17120 -3220 -16880 -3200
rect -16620 -3220 -16380 -3200
rect -16120 -3220 -15880 -3200
rect -15620 -3220 -15380 -3200
rect -15120 -3220 -14880 -3200
rect -14620 -3220 -14500 -3200
rect -23500 -3480 -23400 -3220
rect -23100 -3480 -22900 -3220
rect -22600 -3480 -22400 -3220
rect -22100 -3480 -21900 -3220
rect -21600 -3480 -21400 -3220
rect -21100 -3480 -20900 -3220
rect -20600 -3480 -20400 -3220
rect -20100 -3480 -19900 -3220
rect -19600 -3480 -19400 -3220
rect -19100 -3480 -18900 -3220
rect -18600 -3480 -18400 -3220
rect -18100 -3480 -17900 -3220
rect -17600 -3480 -17400 -3220
rect -17100 -3480 -16900 -3220
rect -16600 -3480 -16400 -3220
rect -16100 -3480 -15900 -3220
rect -15600 -3480 -15400 -3220
rect -15100 -3480 -14900 -3220
rect -14600 -3480 -14500 -3220
rect -23500 -3500 -23380 -3480
rect -23120 -3500 -22880 -3480
rect -22620 -3500 -22380 -3480
rect -22120 -3500 -21880 -3480
rect -21620 -3500 -21380 -3480
rect -21120 -3500 -20880 -3480
rect -20620 -3500 -20380 -3480
rect -20120 -3500 -19880 -3480
rect -19620 -3500 -19380 -3480
rect -19120 -3500 -18880 -3480
rect -18620 -3500 -18380 -3480
rect -18120 -3500 -17880 -3480
rect -17620 -3500 -17380 -3480
rect -17120 -3500 -16880 -3480
rect -16620 -3500 -16380 -3480
rect -16120 -3500 -15880 -3480
rect -15620 -3500 -15380 -3480
rect -15120 -3500 -14880 -3480
rect -14620 -3500 -14500 -3480
rect -23500 -3600 -14500 -3500
rect 12000 -3200 17000 -3000
rect 12000 -3220 12120 -3200
rect 12380 -3220 12620 -3200
rect 12880 -3220 13120 -3200
rect 13380 -3220 13620 -3200
rect 13880 -3220 14120 -3200
rect 14380 -3220 14620 -3200
rect 14880 -3220 15120 -3200
rect 15380 -3220 15620 -3200
rect 15880 -3220 16120 -3200
rect 16380 -3220 16620 -3200
rect 16880 -3220 17000 -3200
rect 12000 -3480 12100 -3220
rect 12400 -3480 12600 -3220
rect 12900 -3480 13100 -3220
rect 13400 -3480 13600 -3220
rect 13900 -3480 14100 -3220
rect 14400 -3480 14600 -3220
rect 14900 -3480 15100 -3220
rect 15400 -3480 15600 -3220
rect 15900 -3480 16100 -3220
rect 16400 -3480 16600 -3220
rect 16900 -3480 17000 -3220
rect 12000 -3500 12120 -3480
rect 12380 -3500 12620 -3480
rect 12880 -3500 13120 -3480
rect 13380 -3500 13620 -3480
rect 13880 -3500 14120 -3480
rect 14380 -3500 14620 -3480
rect 14880 -3500 15120 -3480
rect 15380 -3500 15620 -3480
rect 15880 -3500 16120 -3480
rect 16380 -3500 16620 -3480
rect 16880 -3500 17000 -3480
rect 12000 -3600 17000 -3500
rect 17500 300 19500 500
rect 17500 280 17620 300
rect 17880 280 18120 300
rect 18380 280 18620 300
rect 18880 280 19120 300
rect 19380 280 19500 300
rect 17500 20 17600 280
rect 17900 20 18100 280
rect 18400 20 18600 280
rect 18900 20 19100 280
rect 19400 20 19500 280
rect 17500 0 17620 20
rect 17880 0 18120 20
rect 18380 0 18620 20
rect 18880 0 19120 20
rect 19380 0 19500 20
rect 17500 -200 19500 0
rect 17500 -220 17620 -200
rect 17880 -220 18120 -200
rect 18380 -220 18620 -200
rect 18880 -220 19120 -200
rect 19380 -220 19500 -200
rect 17500 -480 17600 -220
rect 17900 -480 18100 -220
rect 18400 -480 18600 -220
rect 18900 -480 19100 -220
rect 19400 -480 19500 -220
rect 17500 -500 17620 -480
rect 17880 -500 18120 -480
rect 18380 -500 18620 -480
rect 18880 -500 19120 -480
rect 19380 -500 19500 -480
rect 17500 -700 19500 -500
rect 17500 -720 17620 -700
rect 17880 -720 18120 -700
rect 18380 -720 18620 -700
rect 18880 -720 19120 -700
rect 19380 -720 19500 -700
rect 17500 -980 17600 -720
rect 17900 -980 18100 -720
rect 18400 -980 18600 -720
rect 18900 -980 19100 -720
rect 19400 -980 19500 -720
rect 17500 -1000 17620 -980
rect 17880 -1000 18120 -980
rect 18380 -1000 18620 -980
rect 18880 -1000 19120 -980
rect 19380 -1000 19500 -980
rect 17500 -1200 19500 -1000
rect 17500 -1220 17620 -1200
rect 17880 -1220 18120 -1200
rect 18380 -1220 18620 -1200
rect 18880 -1220 19120 -1200
rect 19380 -1220 19500 -1200
rect 17500 -1480 17600 -1220
rect 17900 -1480 18100 -1220
rect 18400 -1480 18600 -1220
rect 18900 -1480 19100 -1220
rect 19400 -1480 19500 -1220
rect 17500 -1500 17620 -1480
rect 17880 -1500 18120 -1480
rect 18380 -1500 18620 -1480
rect 18880 -1500 19120 -1480
rect 19380 -1500 19500 -1480
rect 17500 -1700 19500 -1500
rect 17500 -1720 17620 -1700
rect 17880 -1720 18120 -1700
rect 18380 -1720 18620 -1700
rect 18880 -1720 19120 -1700
rect 19380 -1720 19500 -1700
rect 17500 -1980 17600 -1720
rect 17900 -1980 18100 -1720
rect 18400 -1980 18600 -1720
rect 18900 -1980 19100 -1720
rect 19400 -1980 19500 -1720
rect 17500 -2000 17620 -1980
rect 17880 -2000 18120 -1980
rect 18380 -2000 18620 -1980
rect 18880 -2000 19120 -1980
rect 19380 -2000 19500 -1980
rect 17500 -2200 19500 -2000
rect 17500 -2220 17620 -2200
rect 17880 -2220 18120 -2200
rect 18380 -2220 18620 -2200
rect 18880 -2220 19120 -2200
rect 19380 -2220 19500 -2200
rect 17500 -2480 17600 -2220
rect 17900 -2480 18100 -2220
rect 18400 -2480 18600 -2220
rect 18900 -2480 19100 -2220
rect 19400 -2480 19500 -2220
rect 17500 -2500 17620 -2480
rect 17880 -2500 18120 -2480
rect 18380 -2500 18620 -2480
rect 18880 -2500 19120 -2480
rect 19380 -2500 19500 -2480
rect 17500 -2700 19500 -2500
rect 17500 -2720 17620 -2700
rect 17880 -2720 18120 -2700
rect 18380 -2720 18620 -2700
rect 18880 -2720 19120 -2700
rect 19380 -2720 19500 -2700
rect 17500 -2980 17600 -2720
rect 17900 -2980 18100 -2720
rect 18400 -2980 18600 -2720
rect 18900 -2980 19100 -2720
rect 19400 -2980 19500 -2720
rect 17500 -3000 17620 -2980
rect 17880 -3000 18120 -2980
rect 18380 -3000 18620 -2980
rect 18880 -3000 19120 -2980
rect 19380 -3000 19500 -2980
rect 17500 -3200 19500 -3000
rect 17500 -3220 17620 -3200
rect 17880 -3220 18120 -3200
rect 18380 -3220 18620 -3200
rect 18880 -3220 19120 -3200
rect 19380 -3220 19500 -3200
rect 17500 -3480 17600 -3220
rect 17900 -3480 18100 -3220
rect 18400 -3480 18600 -3220
rect 18900 -3480 19100 -3220
rect 19400 -3480 19500 -3220
rect 17500 -3500 17620 -3480
rect 17880 -3500 18120 -3480
rect 18380 -3500 18620 -3480
rect 18880 -3500 19120 -3480
rect 19380 -3500 19500 -3480
rect 17500 -3600 19500 -3500
rect 32500 1300 33500 1400
rect 32500 1280 32620 1300
rect 32880 1280 33120 1300
rect 33380 1280 33500 1300
rect 32500 1020 32600 1280
rect 32900 1020 33100 1280
rect 33400 1020 33500 1280
rect 32500 1000 32620 1020
rect 32880 1000 33120 1020
rect 33380 1000 33500 1020
rect 32500 800 33500 1000
rect 32500 780 32620 800
rect 32880 780 33120 800
rect 33380 780 33500 800
rect 32500 520 32600 780
rect 32900 520 33100 780
rect 33400 520 33500 780
rect 32500 500 32620 520
rect 32880 500 33120 520
rect 33380 500 33500 520
rect 32500 300 33500 500
rect 32500 280 32620 300
rect 32880 280 33120 300
rect 33380 280 33500 300
rect 32500 20 32600 280
rect 32900 20 33100 280
rect 33400 20 33500 280
rect 32500 0 32620 20
rect 32880 0 33120 20
rect 33380 0 33500 20
rect 32500 -200 33500 0
rect 32500 -220 32620 -200
rect 32880 -220 33120 -200
rect 33380 -220 33500 -200
rect 32500 -480 32600 -220
rect 32900 -480 33100 -220
rect 33400 -480 33500 -220
rect 32500 -500 32620 -480
rect 32880 -500 33120 -480
rect 33380 -500 33500 -480
rect 32500 -700 33500 -500
rect 32500 -720 32620 -700
rect 32880 -720 33120 -700
rect 33380 -720 33500 -700
rect 32500 -980 32600 -720
rect 32900 -980 33100 -720
rect 33400 -980 33500 -720
rect 32500 -1000 32620 -980
rect 32880 -1000 33120 -980
rect 33380 -1000 33500 -980
rect 32500 -1200 33500 -1000
rect 32500 -1220 32620 -1200
rect 32880 -1220 33120 -1200
rect 33380 -1220 33500 -1200
rect 32500 -1480 32600 -1220
rect 32900 -1480 33100 -1220
rect 33400 -1480 33500 -1220
rect 32500 -1500 32620 -1480
rect 32880 -1500 33120 -1480
rect 33380 -1500 33500 -1480
rect 32500 -1700 33500 -1500
rect 32500 -1720 32620 -1700
rect 32880 -1720 33120 -1700
rect 33380 -1720 33500 -1700
rect 32500 -1980 32600 -1720
rect 32900 -1980 33100 -1720
rect 33400 -1980 33500 -1720
rect 32500 -2000 32620 -1980
rect 32880 -2000 33120 -1980
rect 33380 -2000 33500 -1980
rect 32500 -2200 33500 -2000
rect 32500 -2220 32620 -2200
rect 32880 -2220 33120 -2200
rect 33380 -2220 33500 -2200
rect 32500 -2480 32600 -2220
rect 32900 -2480 33100 -2220
rect 33400 -2480 33500 -2220
rect 32500 -2500 32620 -2480
rect 32880 -2500 33120 -2480
rect 33380 -2500 33500 -2480
rect 32500 -2700 33500 -2500
rect 32500 -2720 32620 -2700
rect 32880 -2720 33120 -2700
rect 33380 -2720 33500 -2700
rect 32500 -2980 32600 -2720
rect 32900 -2980 33100 -2720
rect 33400 -2980 33500 -2720
rect 32500 -3000 32620 -2980
rect 32880 -3000 33120 -2980
rect 33380 -3000 33500 -2980
rect 32500 -3200 33500 -3000
rect 32500 -3220 32620 -3200
rect 32880 -3220 33120 -3200
rect 33380 -3220 33500 -3200
rect 32500 -3480 32600 -3220
rect 32900 -3480 33100 -3220
rect 33400 -3480 33500 -3220
rect 32500 -3500 32620 -3480
rect 32880 -3500 33120 -3480
rect 33380 -3500 33500 -3480
rect 32500 -3600 33500 -3500
rect -23500 -3700 -15000 -3600
rect -23500 -3720 -23380 -3700
rect -23120 -3720 -22880 -3700
rect -22620 -3720 -22380 -3700
rect -22120 -3720 -21880 -3700
rect -21620 -3720 -21380 -3700
rect -21120 -3720 -20880 -3700
rect -20620 -3720 -20380 -3700
rect -20120 -3720 -19880 -3700
rect -19620 -3720 -19380 -3700
rect -19120 -3720 -18880 -3700
rect -18620 -3720 -18380 -3700
rect -18120 -3720 -17880 -3700
rect -17620 -3720 -17380 -3700
rect -17120 -3720 -16880 -3700
rect -16620 -3720 -16380 -3700
rect -16120 -3720 -15880 -3700
rect -15620 -3720 -15380 -3700
rect -15120 -3720 -15000 -3700
rect -23500 -3980 -23400 -3720
rect -23100 -3980 -22900 -3720
rect -22600 -3980 -22400 -3720
rect -22100 -3980 -21900 -3720
rect -21600 -3980 -21400 -3720
rect -21100 -3980 -20900 -3720
rect -20600 -3980 -20400 -3720
rect -20100 -3980 -19900 -3720
rect -19600 -3980 -19400 -3720
rect -19100 -3980 -18900 -3720
rect -18600 -3980 -18400 -3720
rect -18100 -3980 -17900 -3720
rect -17600 -3980 -17400 -3720
rect -17100 -3980 -16900 -3720
rect -16600 -3980 -16400 -3720
rect -16100 -3980 -15900 -3720
rect -15600 -3980 -15400 -3720
rect -15100 -3980 -15000 -3720
rect -23500 -4000 -23380 -3980
rect -23120 -4000 -22880 -3980
rect -22620 -4000 -22380 -3980
rect -22120 -4000 -21880 -3980
rect -21620 -4000 -21380 -3980
rect -21120 -4000 -20880 -3980
rect -20620 -4000 -20380 -3980
rect -20120 -4000 -19880 -3980
rect -19620 -4000 -19380 -3980
rect -19120 -4000 -18880 -3980
rect -18620 -4000 -18380 -3980
rect -18120 -4000 -17880 -3980
rect -17620 -4000 -17380 -3980
rect -17120 -4000 -16880 -3980
rect -16620 -4000 -16380 -3980
rect -16120 -4000 -15880 -3980
rect -15620 -4000 -15380 -3980
rect -15120 -4000 -15000 -3980
rect -23500 -4200 -15000 -4000
rect -23500 -4220 -23380 -4200
rect -23120 -4220 -22880 -4200
rect -22620 -4220 -22380 -4200
rect -22120 -4220 -21880 -4200
rect -21620 -4220 -21380 -4200
rect -21120 -4220 -20880 -4200
rect -20620 -4220 -20380 -4200
rect -20120 -4220 -19880 -4200
rect -19620 -4220 -19380 -4200
rect -19120 -4220 -18880 -4200
rect -18620 -4220 -18380 -4200
rect -18120 -4220 -17880 -4200
rect -17620 -4220 -17380 -4200
rect -17120 -4220 -16880 -4200
rect -16620 -4220 -16380 -4200
rect -16120 -4220 -15880 -4200
rect -15620 -4220 -15380 -4200
rect -15120 -4220 -15000 -4200
rect -23500 -4480 -23400 -4220
rect -23100 -4480 -22900 -4220
rect -22600 -4480 -22400 -4220
rect -22100 -4480 -21900 -4220
rect -21600 -4480 -21400 -4220
rect -21100 -4480 -20900 -4220
rect -20600 -4480 -20400 -4220
rect -20100 -4480 -19900 -4220
rect -19600 -4480 -19400 -4220
rect -19100 -4480 -18900 -4220
rect -18600 -4480 -18400 -4220
rect -18100 -4480 -17900 -4220
rect -17600 -4480 -17400 -4220
rect -17100 -4480 -16900 -4220
rect -16600 -4480 -16400 -4220
rect -16100 -4480 -15900 -4220
rect -15600 -4480 -15400 -4220
rect -15100 -4480 -15000 -4220
rect -23500 -4500 -23380 -4480
rect -23120 -4500 -22880 -4480
rect -22620 -4500 -22380 -4480
rect -22120 -4500 -21880 -4480
rect -21620 -4500 -21380 -4480
rect -21120 -4500 -20880 -4480
rect -20620 -4500 -20380 -4480
rect -20120 -4500 -19880 -4480
rect -19620 -4500 -19380 -4480
rect -19120 -4500 -18880 -4480
rect -18620 -4500 -18380 -4480
rect -18120 -4500 -17880 -4480
rect -17620 -4500 -17380 -4480
rect -17120 -4500 -16880 -4480
rect -16620 -4500 -16380 -4480
rect -16120 -4500 -15880 -4480
rect -15620 -4500 -15380 -4480
rect -15120 -4500 -15000 -4480
rect -23500 -4700 -15000 -4500
rect -23500 -4720 -23380 -4700
rect -23120 -4720 -22880 -4700
rect -22620 -4720 -22380 -4700
rect -22120 -4720 -21880 -4700
rect -21620 -4720 -21380 -4700
rect -21120 -4720 -20880 -4700
rect -20620 -4720 -20380 -4700
rect -20120 -4720 -19880 -4700
rect -19620 -4720 -19380 -4700
rect -19120 -4720 -18880 -4700
rect -18620 -4720 -18380 -4700
rect -18120 -4720 -17880 -4700
rect -17620 -4720 -17380 -4700
rect -17120 -4720 -16880 -4700
rect -16620 -4720 -16380 -4700
rect -16120 -4720 -15880 -4700
rect -15620 -4720 -15380 -4700
rect -15120 -4720 -15000 -4700
rect -23500 -4980 -23400 -4720
rect -23100 -4980 -22900 -4720
rect -22600 -4980 -22400 -4720
rect -22100 -4980 -21900 -4720
rect -21600 -4980 -21400 -4720
rect -21100 -4980 -20900 -4720
rect -20600 -4980 -20400 -4720
rect -20100 -4980 -19900 -4720
rect -19600 -4980 -19400 -4720
rect -19100 -4980 -18900 -4720
rect -18600 -4980 -18400 -4720
rect -18100 -4980 -17900 -4720
rect -17600 -4980 -17400 -4720
rect -17100 -4980 -16900 -4720
rect -16600 -4980 -16400 -4720
rect -16100 -4980 -15900 -4720
rect -15600 -4980 -15400 -4720
rect -15100 -4980 -15000 -4720
rect -23500 -5000 -23380 -4980
rect -23120 -5000 -22880 -4980
rect -22620 -5000 -22380 -4980
rect -22120 -5000 -21880 -4980
rect -21620 -5000 -21380 -4980
rect -21120 -5000 -20880 -4980
rect -20620 -5000 -20380 -4980
rect -20120 -5000 -19880 -4980
rect -19620 -5000 -19380 -4980
rect -19120 -5000 -18880 -4980
rect -18620 -5000 -18380 -4980
rect -18120 -5000 -17880 -4980
rect -17620 -5000 -17380 -4980
rect -17120 -5000 -16880 -4980
rect -16620 -5000 -16380 -4980
rect -16120 -5000 -15880 -4980
rect -15620 -5000 -15380 -4980
rect -15120 -5000 -15000 -4980
rect -23500 -5200 -15000 -5000
rect -23500 -5220 -23380 -5200
rect -23120 -5220 -22880 -5200
rect -22620 -5220 -22380 -5200
rect -22120 -5220 -21880 -5200
rect -21620 -5220 -21380 -5200
rect -21120 -5220 -20880 -5200
rect -20620 -5220 -20380 -5200
rect -20120 -5220 -19880 -5200
rect -19620 -5220 -19380 -5200
rect -19120 -5220 -18880 -5200
rect -18620 -5220 -18380 -5200
rect -18120 -5220 -17880 -5200
rect -17620 -5220 -17380 -5200
rect -17120 -5220 -16880 -5200
rect -16620 -5220 -16380 -5200
rect -16120 -5220 -15880 -5200
rect -15620 -5220 -15380 -5200
rect -15120 -5220 -15000 -5200
rect -23500 -5480 -23400 -5220
rect -23100 -5480 -22900 -5220
rect -22600 -5480 -22400 -5220
rect -22100 -5480 -21900 -5220
rect -21600 -5480 -21400 -5220
rect -21100 -5480 -20900 -5220
rect -20600 -5480 -20400 -5220
rect -20100 -5480 -19900 -5220
rect -19600 -5480 -19400 -5220
rect -19100 -5480 -18900 -5220
rect -18600 -5480 -18400 -5220
rect -18100 -5480 -17900 -5220
rect -17600 -5480 -17400 -5220
rect -17100 -5480 -16900 -5220
rect -16600 -5480 -16400 -5220
rect -16100 -5480 -15900 -5220
rect -15600 -5480 -15400 -5220
rect -15100 -5480 -15000 -5220
rect -23500 -5500 -23380 -5480
rect -23120 -5500 -22880 -5480
rect -22620 -5500 -22380 -5480
rect -22120 -5500 -21880 -5480
rect -21620 -5500 -21380 -5480
rect -21120 -5500 -20880 -5480
rect -20620 -5500 -20380 -5480
rect -20120 -5500 -19880 -5480
rect -19620 -5500 -19380 -5480
rect -19120 -5500 -18880 -5480
rect -18620 -5500 -18380 -5480
rect -18120 -5500 -17880 -5480
rect -17620 -5500 -17380 -5480
rect -17120 -5500 -16880 -5480
rect -16620 -5500 -16380 -5480
rect -16120 -5500 -15880 -5480
rect -15620 -5500 -15380 -5480
rect -15120 -5500 -15000 -5480
rect -23500 -5700 -15000 -5500
rect -23500 -5720 -23380 -5700
rect -23120 -5720 -22880 -5700
rect -22620 -5720 -22380 -5700
rect -22120 -5720 -21880 -5700
rect -21620 -5720 -21380 -5700
rect -21120 -5720 -20880 -5700
rect -20620 -5720 -20380 -5700
rect -20120 -5720 -19880 -5700
rect -19620 -5720 -19380 -5700
rect -19120 -5720 -18880 -5700
rect -18620 -5720 -18380 -5700
rect -18120 -5720 -17880 -5700
rect -17620 -5720 -17380 -5700
rect -17120 -5720 -16880 -5700
rect -16620 -5720 -16380 -5700
rect -16120 -5720 -15880 -5700
rect -15620 -5720 -15380 -5700
rect -15120 -5720 -15000 -5700
rect -23500 -5980 -23400 -5720
rect -23100 -5980 -22900 -5720
rect -22600 -5980 -22400 -5720
rect -22100 -5980 -21900 -5720
rect -21600 -5980 -21400 -5720
rect -21100 -5980 -20900 -5720
rect -20600 -5980 -20400 -5720
rect -20100 -5980 -19900 -5720
rect -19600 -5980 -19400 -5720
rect -19100 -5980 -18900 -5720
rect -18600 -5980 -18400 -5720
rect -18100 -5980 -17900 -5720
rect -17600 -5980 -17400 -5720
rect -17100 -5980 -16900 -5720
rect -16600 -5980 -16400 -5720
rect -16100 -5980 -15900 -5720
rect -15600 -5980 -15400 -5720
rect -15100 -5980 -15000 -5720
rect -23500 -6000 -23380 -5980
rect -23120 -6000 -22880 -5980
rect -22620 -6000 -22380 -5980
rect -22120 -6000 -21880 -5980
rect -21620 -6000 -21380 -5980
rect -21120 -6000 -20880 -5980
rect -20620 -6000 -20380 -5980
rect -20120 -6000 -19880 -5980
rect -19620 -6000 -19380 -5980
rect -19120 -6000 -18880 -5980
rect -18620 -6000 -18380 -5980
rect -18120 -6000 -17880 -5980
rect -17620 -6000 -17380 -5980
rect -17120 -6000 -16880 -5980
rect -16620 -6000 -16380 -5980
rect -16120 -6000 -15880 -5980
rect -15620 -6000 -15380 -5980
rect -15120 -6000 -15000 -5980
rect -23500 -6200 -15000 -6000
rect -23500 -6220 -23380 -6200
rect -23120 -6220 -22880 -6200
rect -22620 -6220 -22380 -6200
rect -22120 -6220 -21880 -6200
rect -21620 -6220 -21380 -6200
rect -21120 -6220 -20880 -6200
rect -20620 -6220 -20380 -6200
rect -20120 -6220 -19880 -6200
rect -19620 -6220 -19380 -6200
rect -19120 -6220 -18880 -6200
rect -18620 -6220 -18380 -6200
rect -18120 -6220 -17880 -6200
rect -17620 -6220 -17380 -6200
rect -17120 -6220 -16880 -6200
rect -16620 -6220 -16380 -6200
rect -16120 -6220 -15880 -6200
rect -15620 -6220 -15380 -6200
rect -15120 -6220 -15000 -6200
rect -23500 -6480 -23400 -6220
rect -23100 -6480 -22900 -6220
rect -22600 -6480 -22400 -6220
rect -22100 -6480 -21900 -6220
rect -21600 -6480 -21400 -6220
rect -21100 -6480 -20900 -6220
rect -20600 -6480 -20400 -6220
rect -20100 -6480 -19900 -6220
rect -19600 -6480 -19400 -6220
rect -19100 -6480 -18900 -6220
rect -18600 -6480 -18400 -6220
rect -18100 -6480 -17900 -6220
rect -17600 -6480 -17400 -6220
rect -17100 -6480 -16900 -6220
rect -16600 -6480 -16400 -6220
rect -16100 -6480 -15900 -6220
rect -15600 -6480 -15400 -6220
rect -15100 -6480 -15000 -6220
rect -23500 -6500 -23380 -6480
rect -23120 -6500 -22880 -6480
rect -22620 -6500 -22380 -6480
rect -22120 -6500 -21880 -6480
rect -21620 -6500 -21380 -6480
rect -21120 -6500 -20880 -6480
rect -20620 -6500 -20380 -6480
rect -20120 -6500 -19880 -6480
rect -19620 -6500 -19380 -6480
rect -19120 -6500 -18880 -6480
rect -18620 -6500 -18380 -6480
rect -18120 -6500 -17880 -6480
rect -17620 -6500 -17380 -6480
rect -17120 -6500 -16880 -6480
rect -16620 -6500 -16380 -6480
rect -16120 -6500 -15880 -6480
rect -15620 -6500 -15380 -6480
rect -15120 -6500 -15000 -6480
rect -23500 -6700 -15000 -6500
rect -23500 -6720 -23380 -6700
rect -23120 -6720 -22880 -6700
rect -22620 -6720 -22380 -6700
rect -22120 -6720 -21880 -6700
rect -21620 -6720 -21380 -6700
rect -21120 -6720 -20880 -6700
rect -20620 -6720 -20380 -6700
rect -20120 -6720 -19880 -6700
rect -19620 -6720 -19380 -6700
rect -19120 -6720 -18880 -6700
rect -18620 -6720 -18380 -6700
rect -18120 -6720 -17880 -6700
rect -17620 -6720 -17380 -6700
rect -17120 -6720 -16880 -6700
rect -16620 -6720 -16380 -6700
rect -16120 -6720 -15880 -6700
rect -15620 -6720 -15380 -6700
rect -15120 -6720 -15000 -6700
rect -23500 -6980 -23400 -6720
rect -23100 -6980 -22900 -6720
rect -22600 -6980 -22400 -6720
rect -22100 -6980 -21900 -6720
rect -21600 -6980 -21400 -6720
rect -21100 -6980 -20900 -6720
rect -20600 -6980 -20400 -6720
rect -20100 -6980 -19900 -6720
rect -19600 -6980 -19400 -6720
rect -19100 -6980 -18900 -6720
rect -18600 -6980 -18400 -6720
rect -18100 -6980 -17900 -6720
rect -17600 -6980 -17400 -6720
rect -17100 -6980 -16900 -6720
rect -16600 -6980 -16400 -6720
rect -16100 -6980 -15900 -6720
rect -15600 -6980 -15400 -6720
rect -15100 -6980 -15000 -6720
rect -23500 -7000 -23380 -6980
rect -23120 -7000 -22880 -6980
rect -22620 -7000 -22380 -6980
rect -22120 -7000 -21880 -6980
rect -21620 -7000 -21380 -6980
rect -21120 -7000 -20880 -6980
rect -20620 -7000 -20380 -6980
rect -20120 -7000 -19880 -6980
rect -19620 -7000 -19380 -6980
rect -19120 -7000 -18880 -6980
rect -18620 -7000 -18380 -6980
rect -18120 -7000 -17880 -6980
rect -17620 -7000 -17380 -6980
rect -17120 -7000 -16880 -6980
rect -16620 -7000 -16380 -6980
rect -16120 -7000 -15880 -6980
rect -15620 -7000 -15380 -6980
rect -15120 -7000 -15000 -6980
rect -23500 -7200 -15000 -7000
rect -23500 -7220 -23380 -7200
rect -23120 -7220 -22880 -7200
rect -22620 -7220 -22380 -7200
rect -22120 -7220 -21880 -7200
rect -21620 -7220 -21380 -7200
rect -21120 -7220 -20880 -7200
rect -20620 -7220 -20380 -7200
rect -20120 -7220 -19880 -7200
rect -19620 -7220 -19380 -7200
rect -19120 -7220 -18880 -7200
rect -18620 -7220 -18380 -7200
rect -18120 -7220 -17880 -7200
rect -17620 -7220 -17380 -7200
rect -17120 -7220 -16880 -7200
rect -16620 -7220 -16380 -7200
rect -16120 -7220 -15880 -7200
rect -15620 -7220 -15380 -7200
rect -15120 -7220 -15000 -7200
rect -23500 -7480 -23400 -7220
rect -23100 -7480 -22900 -7220
rect -22600 -7480 -22400 -7220
rect -22100 -7480 -21900 -7220
rect -21600 -7480 -21400 -7220
rect -21100 -7480 -20900 -7220
rect -20600 -7480 -20400 -7220
rect -20100 -7480 -19900 -7220
rect -19600 -7480 -19400 -7220
rect -19100 -7480 -18900 -7220
rect -18600 -7480 -18400 -7220
rect -18100 -7480 -17900 -7220
rect -17600 -7480 -17400 -7220
rect -17100 -7480 -16900 -7220
rect -16600 -7480 -16400 -7220
rect -16100 -7480 -15900 -7220
rect -15600 -7480 -15400 -7220
rect -15100 -7480 -15000 -7220
rect -23500 -7500 -23380 -7480
rect -23120 -7500 -22880 -7480
rect -22620 -7500 -22380 -7480
rect -22120 -7500 -21880 -7480
rect -21620 -7500 -21380 -7480
rect -21120 -7500 -20880 -7480
rect -20620 -7500 -20380 -7480
rect -20120 -7500 -19880 -7480
rect -19620 -7500 -19380 -7480
rect -19120 -7500 -18880 -7480
rect -18620 -7500 -18380 -7480
rect -18120 -7500 -17880 -7480
rect -17620 -7500 -17380 -7480
rect -17120 -7500 -16880 -7480
rect -16620 -7500 -16380 -7480
rect -16120 -7500 -15880 -7480
rect -15620 -7500 -15380 -7480
rect -15120 -7500 -15000 -7480
rect -28000 -8100 -27500 -7600
rect -23500 -7700 -15000 -7500
rect -23500 -7720 -23380 -7700
rect -23120 -7720 -22880 -7700
rect -22620 -7720 -22380 -7700
rect -22120 -7720 -21880 -7700
rect -21620 -7720 -21380 -7700
rect -21120 -7720 -20880 -7700
rect -20620 -7720 -20380 -7700
rect -20120 -7720 -19880 -7700
rect -19620 -7720 -19380 -7700
rect -19120 -7720 -18880 -7700
rect -18620 -7720 -18380 -7700
rect -18120 -7720 -17880 -7700
rect -17620 -7720 -17380 -7700
rect -17120 -7720 -16880 -7700
rect -16620 -7720 -16380 -7700
rect -16120 -7720 -15880 -7700
rect -15620 -7720 -15380 -7700
rect -15120 -7720 -15000 -7700
rect -23500 -7980 -23400 -7720
rect -23100 -7980 -22900 -7720
rect -22600 -7980 -22400 -7720
rect -22100 -7980 -21900 -7720
rect -21600 -7980 -21400 -7720
rect -21100 -7980 -20900 -7720
rect -20600 -7980 -20400 -7720
rect -20100 -7980 -19900 -7720
rect -19600 -7980 -19400 -7720
rect -19100 -7980 -18900 -7720
rect -18600 -7980 -18400 -7720
rect -18100 -7980 -17900 -7720
rect -17600 -7980 -17400 -7720
rect -17100 -7980 -16900 -7720
rect -16600 -7980 -16400 -7720
rect -16100 -7980 -15900 -7720
rect -15600 -7980 -15400 -7720
rect -15100 -7980 -15000 -7720
rect -23500 -8000 -23380 -7980
rect -23120 -8000 -22880 -7980
rect -22620 -8000 -22380 -7980
rect -22120 -8000 -21880 -7980
rect -21620 -8000 -21380 -7980
rect -21120 -8000 -20880 -7980
rect -20620 -8000 -20380 -7980
rect -20120 -8000 -19880 -7980
rect -19620 -8000 -19380 -7980
rect -19120 -8000 -18880 -7980
rect -18620 -8000 -18380 -7980
rect -18120 -8000 -17880 -7980
rect -17620 -8000 -17380 -7980
rect -17120 -8000 -16880 -7980
rect -16620 -8000 -16380 -7980
rect -16120 -8000 -15880 -7980
rect -15620 -8000 -15380 -7980
rect -15120 -8000 -15000 -7980
rect -23500 -8100 -15000 -8000
rect -27500 -8200 -15000 -8100
rect -27500 -8220 -27380 -8200
rect -27120 -8220 -26880 -8200
rect -26620 -8220 -26380 -8200
rect -26120 -8220 -25880 -8200
rect -25620 -8220 -25380 -8200
rect -25120 -8220 -24880 -8200
rect -24620 -8220 -24380 -8200
rect -24120 -8220 -23880 -8200
rect -23620 -8220 -23380 -8200
rect -23120 -8220 -22880 -8200
rect -22620 -8220 -22380 -8200
rect -22120 -8220 -21880 -8200
rect -21620 -8220 -21380 -8200
rect -21120 -8220 -20880 -8200
rect -20620 -8220 -20380 -8200
rect -20120 -8220 -19880 -8200
rect -19620 -8220 -19380 -8200
rect -19120 -8220 -18880 -8200
rect -18620 -8220 -18380 -8200
rect -18120 -8220 -17880 -8200
rect -17620 -8220 -17380 -8200
rect -17120 -8220 -16880 -8200
rect -16620 -8220 -16380 -8200
rect -16120 -8220 -15880 -8200
rect -15620 -8220 -15380 -8200
rect -15120 -8220 -15000 -8200
rect -27500 -8480 -27400 -8220
rect -27100 -8480 -26900 -8220
rect -26600 -8480 -26400 -8220
rect -26100 -8480 -25900 -8220
rect -25600 -8480 -25400 -8220
rect -25100 -8480 -24900 -8220
rect -24600 -8480 -24400 -8220
rect -24100 -8480 -23900 -8220
rect -23600 -8480 -23400 -8220
rect -23100 -8480 -22900 -8220
rect -22600 -8480 -22400 -8220
rect -22100 -8480 -21900 -8220
rect -21600 -8480 -21400 -8220
rect -21100 -8480 -20900 -8220
rect -20600 -8480 -20400 -8220
rect -20100 -8480 -19900 -8220
rect -19600 -8480 -19400 -8220
rect -19100 -8480 -18900 -8220
rect -18600 -8480 -18400 -8220
rect -18100 -8480 -17900 -8220
rect -17600 -8480 -17400 -8220
rect -17100 -8480 -16900 -8220
rect -16600 -8480 -16400 -8220
rect -16100 -8480 -15900 -8220
rect -15600 -8480 -15400 -8220
rect -15100 -8480 -15000 -8220
rect -27500 -8500 -27380 -8480
rect -27120 -8500 -26880 -8480
rect -26620 -8500 -26380 -8480
rect -26120 -8500 -25880 -8480
rect -25620 -8500 -25380 -8480
rect -25120 -8500 -24880 -8480
rect -24620 -8500 -24380 -8480
rect -24120 -8500 -23880 -8480
rect -23620 -8500 -23380 -8480
rect -23120 -8500 -22880 -8480
rect -22620 -8500 -22380 -8480
rect -22120 -8500 -21880 -8480
rect -21620 -8500 -21380 -8480
rect -21120 -8500 -20880 -8480
rect -20620 -8500 -20380 -8480
rect -20120 -8500 -19880 -8480
rect -19620 -8500 -19380 -8480
rect -19120 -8500 -18880 -8480
rect -18620 -8500 -18380 -8480
rect -18120 -8500 -17880 -8480
rect -17620 -8500 -17380 -8480
rect -17120 -8500 -16880 -8480
rect -16620 -8500 -16380 -8480
rect -16120 -8500 -15880 -8480
rect -15620 -8500 -15380 -8480
rect -15120 -8500 -15000 -8480
rect -27500 -8700 -15000 -8500
rect -27500 -8720 -27380 -8700
rect -27120 -8720 -26880 -8700
rect -26620 -8720 -26380 -8700
rect -26120 -8720 -25880 -8700
rect -25620 -8720 -25380 -8700
rect -25120 -8720 -24880 -8700
rect -24620 -8720 -24380 -8700
rect -24120 -8720 -23880 -8700
rect -23620 -8720 -23380 -8700
rect -23120 -8720 -22880 -8700
rect -22620 -8720 -22380 -8700
rect -22120 -8720 -21880 -8700
rect -21620 -8720 -21380 -8700
rect -21120 -8720 -20880 -8700
rect -20620 -8720 -20380 -8700
rect -20120 -8720 -19880 -8700
rect -19620 -8720 -19380 -8700
rect -19120 -8720 -18880 -8700
rect -18620 -8720 -18380 -8700
rect -18120 -8720 -17880 -8700
rect -17620 -8720 -17380 -8700
rect -17120 -8720 -16880 -8700
rect -16620 -8720 -16380 -8700
rect -16120 -8720 -15880 -8700
rect -15620 -8720 -15380 -8700
rect -15120 -8720 -15000 -8700
rect -27500 -8980 -27400 -8720
rect -27100 -8980 -26900 -8720
rect -26600 -8980 -26400 -8720
rect -26100 -8980 -25900 -8720
rect -25600 -8980 -25400 -8720
rect -25100 -8980 -24900 -8720
rect -24600 -8980 -24400 -8720
rect -24100 -8980 -23900 -8720
rect -23600 -8980 -23400 -8720
rect -23100 -8980 -22900 -8720
rect -22600 -8980 -22400 -8720
rect -22100 -8980 -21900 -8720
rect -21600 -8980 -21400 -8720
rect -21100 -8980 -20900 -8720
rect -20600 -8980 -20400 -8720
rect -20100 -8980 -19900 -8720
rect -19600 -8980 -19400 -8720
rect -19100 -8980 -18900 -8720
rect -18600 -8980 -18400 -8720
rect -18100 -8980 -17900 -8720
rect -17600 -8980 -17400 -8720
rect -17100 -8980 -16900 -8720
rect -16600 -8980 -16400 -8720
rect -16100 -8980 -15900 -8720
rect -15600 -8980 -15400 -8720
rect -15100 -8980 -15000 -8720
rect -27500 -9000 -27380 -8980
rect -27120 -9000 -26880 -8980
rect -26620 -9000 -26380 -8980
rect -26120 -9000 -25880 -8980
rect -25620 -9000 -25380 -8980
rect -25120 -9000 -24880 -8980
rect -24620 -9000 -24380 -8980
rect -24120 -9000 -23880 -8980
rect -23620 -9000 -23380 -8980
rect -23120 -9000 -22880 -8980
rect -22620 -9000 -22380 -8980
rect -22120 -9000 -21880 -8980
rect -21620 -9000 -21380 -8980
rect -21120 -9000 -20880 -8980
rect -20620 -9000 -20380 -8980
rect -20120 -9000 -19880 -8980
rect -19620 -9000 -19380 -8980
rect -19120 -9000 -18880 -8980
rect -18620 -9000 -18380 -8980
rect -18120 -9000 -17880 -8980
rect -17620 -9000 -17380 -8980
rect -17120 -9000 -16880 -8980
rect -16620 -9000 -16380 -8980
rect -16120 -9000 -15880 -8980
rect -15620 -9000 -15380 -8980
rect -15120 -9000 -15000 -8980
rect -27500 -9200 -15000 -9000
rect -27500 -9220 -27380 -9200
rect -27120 -9220 -26880 -9200
rect -26620 -9220 -26380 -9200
rect -26120 -9220 -25880 -9200
rect -25620 -9220 -25380 -9200
rect -25120 -9220 -24880 -9200
rect -24620 -9220 -24380 -9200
rect -24120 -9220 -23880 -9200
rect -23620 -9220 -23380 -9200
rect -23120 -9220 -22880 -9200
rect -22620 -9220 -22380 -9200
rect -22120 -9220 -21880 -9200
rect -21620 -9220 -21380 -9200
rect -21120 -9220 -20880 -9200
rect -20620 -9220 -20380 -9200
rect -20120 -9220 -19880 -9200
rect -19620 -9220 -19380 -9200
rect -19120 -9220 -18880 -9200
rect -18620 -9220 -18380 -9200
rect -18120 -9220 -17880 -9200
rect -17620 -9220 -17380 -9200
rect -17120 -9220 -16880 -9200
rect -16620 -9220 -16380 -9200
rect -16120 -9220 -15880 -9200
rect -15620 -9220 -15380 -9200
rect -15120 -9220 -15000 -9200
rect -27500 -9480 -27400 -9220
rect -27100 -9480 -26900 -9220
rect -26600 -9480 -26400 -9220
rect -26100 -9480 -25900 -9220
rect -25600 -9480 -25400 -9220
rect -25100 -9480 -24900 -9220
rect -24600 -9480 -24400 -9220
rect -24100 -9480 -23900 -9220
rect -23600 -9480 -23400 -9220
rect -23100 -9480 -22900 -9220
rect -22600 -9480 -22400 -9220
rect -22100 -9480 -21900 -9220
rect -21600 -9480 -21400 -9220
rect -21100 -9480 -20900 -9220
rect -20600 -9480 -20400 -9220
rect -20100 -9480 -19900 -9220
rect -19600 -9480 -19400 -9220
rect -19100 -9480 -18900 -9220
rect -18600 -9480 -18400 -9220
rect -18100 -9480 -17900 -9220
rect -17600 -9480 -17400 -9220
rect -17100 -9480 -16900 -9220
rect -16600 -9480 -16400 -9220
rect -16100 -9480 -15900 -9220
rect -15600 -9480 -15400 -9220
rect -15100 -9480 -15000 -9220
rect -27500 -9500 -27380 -9480
rect -27120 -9500 -26880 -9480
rect -26620 -9500 -26380 -9480
rect -26120 -9500 -25880 -9480
rect -25620 -9500 -25380 -9480
rect -25120 -9500 -24880 -9480
rect -24620 -9500 -24380 -9480
rect -24120 -9500 -23880 -9480
rect -23620 -9500 -23380 -9480
rect -23120 -9500 -22880 -9480
rect -22620 -9500 -22380 -9480
rect -22120 -9500 -21880 -9480
rect -21620 -9500 -21380 -9480
rect -21120 -9500 -20880 -9480
rect -20620 -9500 -20380 -9480
rect -20120 -9500 -19880 -9480
rect -19620 -9500 -19380 -9480
rect -19120 -9500 -18880 -9480
rect -18620 -9500 -18380 -9480
rect -18120 -9500 -17880 -9480
rect -17620 -9500 -17380 -9480
rect -17120 -9500 -16880 -9480
rect -16620 -9500 -16380 -9480
rect -16120 -9500 -15880 -9480
rect -15620 -9500 -15380 -9480
rect -15120 -9500 -15000 -9480
rect -27500 -9700 -15000 -9500
rect -27500 -9720 -27380 -9700
rect -27120 -9720 -26880 -9700
rect -26620 -9720 -26380 -9700
rect -26120 -9720 -25880 -9700
rect -25620 -9720 -25380 -9700
rect -25120 -9720 -24880 -9700
rect -24620 -9720 -24380 -9700
rect -24120 -9720 -23880 -9700
rect -23620 -9720 -23380 -9700
rect -23120 -9720 -22880 -9700
rect -22620 -9720 -22380 -9700
rect -22120 -9720 -21880 -9700
rect -21620 -9720 -21380 -9700
rect -21120 -9720 -20880 -9700
rect -20620 -9720 -20380 -9700
rect -20120 -9720 -19880 -9700
rect -19620 -9720 -19380 -9700
rect -19120 -9720 -18880 -9700
rect -18620 -9720 -18380 -9700
rect -18120 -9720 -17880 -9700
rect -17620 -9720 -17380 -9700
rect -17120 -9720 -16880 -9700
rect -16620 -9720 -16380 -9700
rect -16120 -9720 -15880 -9700
rect -15620 -9720 -15380 -9700
rect -15120 -9720 -15000 -9700
rect -27500 -9980 -27400 -9720
rect -27100 -9980 -26900 -9720
rect -26600 -9980 -26400 -9720
rect -26100 -9980 -25900 -9720
rect -25600 -9980 -25400 -9720
rect -25100 -9980 -24900 -9720
rect -24600 -9980 -24400 -9720
rect -24100 -9980 -23900 -9720
rect -23600 -9980 -23400 -9720
rect -23100 -9980 -22900 -9720
rect -22600 -9980 -22400 -9720
rect -22100 -9980 -21900 -9720
rect -21600 -9980 -21400 -9720
rect -21100 -9980 -20900 -9720
rect -20600 -9980 -20400 -9720
rect -20100 -9980 -19900 -9720
rect -19600 -9980 -19400 -9720
rect -19100 -9980 -18900 -9720
rect -18600 -9980 -18400 -9720
rect -18100 -9980 -17900 -9720
rect -17600 -9980 -17400 -9720
rect -17100 -9980 -16900 -9720
rect -16600 -9980 -16400 -9720
rect -16100 -9980 -15900 -9720
rect -15600 -9980 -15400 -9720
rect -15100 -9980 -15000 -9720
rect -27500 -10000 -27380 -9980
rect -27120 -10000 -26880 -9980
rect -26620 -10000 -26380 -9980
rect -26120 -10000 -25880 -9980
rect -25620 -10000 -25380 -9980
rect -25120 -10000 -24880 -9980
rect -24620 -10000 -24380 -9980
rect -24120 -10000 -23880 -9980
rect -23620 -10000 -23380 -9980
rect -23120 -10000 -22880 -9980
rect -22620 -10000 -22380 -9980
rect -22120 -10000 -21880 -9980
rect -21620 -10000 -21380 -9980
rect -21120 -10000 -20880 -9980
rect -20620 -10000 -20380 -9980
rect -20120 -10000 -19880 -9980
rect -19620 -10000 -19380 -9980
rect -19120 -10000 -18880 -9980
rect -18620 -10000 -18380 -9980
rect -18120 -10000 -17880 -9980
rect -17620 -10000 -17380 -9980
rect -17120 -10000 -16880 -9980
rect -16620 -10000 -16380 -9980
rect -16120 -10000 -15880 -9980
rect -15620 -10000 -15380 -9980
rect -15120 -10000 -15000 -9980
rect -27500 -10200 -15000 -10000
rect -27500 -10220 -27380 -10200
rect -27120 -10220 -26880 -10200
rect -26620 -10220 -26380 -10200
rect -26120 -10220 -25880 -10200
rect -25620 -10220 -25380 -10200
rect -25120 -10220 -24880 -10200
rect -24620 -10220 -24380 -10200
rect -24120 -10220 -23880 -10200
rect -23620 -10220 -23380 -10200
rect -23120 -10220 -22880 -10200
rect -22620 -10220 -22380 -10200
rect -22120 -10220 -21880 -10200
rect -21620 -10220 -21380 -10200
rect -21120 -10220 -20880 -10200
rect -20620 -10220 -20380 -10200
rect -20120 -10220 -19880 -10200
rect -19620 -10220 -19380 -10200
rect -19120 -10220 -18880 -10200
rect -18620 -10220 -18380 -10200
rect -18120 -10220 -17880 -10200
rect -17620 -10220 -17380 -10200
rect -17120 -10220 -16880 -10200
rect -16620 -10220 -16380 -10200
rect -16120 -10220 -15880 -10200
rect -15620 -10220 -15380 -10200
rect -15120 -10220 -15000 -10200
rect -27500 -10480 -27400 -10220
rect -27100 -10480 -26900 -10220
rect -26600 -10480 -26400 -10220
rect -26100 -10480 -25900 -10220
rect -25600 -10480 -25400 -10220
rect -25100 -10480 -24900 -10220
rect -24600 -10480 -24400 -10220
rect -24100 -10480 -23900 -10220
rect -23600 -10480 -23400 -10220
rect -23100 -10480 -22900 -10220
rect -22600 -10480 -22400 -10220
rect -22100 -10480 -21900 -10220
rect -21600 -10480 -21400 -10220
rect -21100 -10480 -20900 -10220
rect -20600 -10480 -20400 -10220
rect -20100 -10480 -19900 -10220
rect -19600 -10480 -19400 -10220
rect -19100 -10480 -18900 -10220
rect -18600 -10480 -18400 -10220
rect -18100 -10480 -17900 -10220
rect -17600 -10480 -17400 -10220
rect -17100 -10480 -16900 -10220
rect -16600 -10480 -16400 -10220
rect -16100 -10480 -15900 -10220
rect -15600 -10480 -15400 -10220
rect -15100 -10480 -15000 -10220
rect -27500 -10500 -27380 -10480
rect -27120 -10500 -26880 -10480
rect -26620 -10500 -26380 -10480
rect -26120 -10500 -25880 -10480
rect -25620 -10500 -25380 -10480
rect -25120 -10500 -24880 -10480
rect -24620 -10500 -24380 -10480
rect -24120 -10500 -23880 -10480
rect -23620 -10500 -23380 -10480
rect -23120 -10500 -22880 -10480
rect -22620 -10500 -22380 -10480
rect -22120 -10500 -21880 -10480
rect -21620 -10500 -21380 -10480
rect -21120 -10500 -20880 -10480
rect -20620 -10500 -20380 -10480
rect -20120 -10500 -19880 -10480
rect -19620 -10500 -19380 -10480
rect -19120 -10500 -18880 -10480
rect -18620 -10500 -18380 -10480
rect -18120 -10500 -17880 -10480
rect -17620 -10500 -17380 -10480
rect -17120 -10500 -16880 -10480
rect -16620 -10500 -16380 -10480
rect -16120 -10500 -15880 -10480
rect -15620 -10500 -15380 -10480
rect -15120 -10500 -15000 -10480
rect -27500 -10700 -15000 -10500
rect -27500 -10720 -27380 -10700
rect -27120 -10720 -26880 -10700
rect -26620 -10720 -26380 -10700
rect -26120 -10720 -25880 -10700
rect -25620 -10720 -25380 -10700
rect -25120 -10720 -24880 -10700
rect -24620 -10720 -24380 -10700
rect -24120 -10720 -23880 -10700
rect -23620 -10720 -23380 -10700
rect -23120 -10720 -22880 -10700
rect -22620 -10720 -22380 -10700
rect -22120 -10720 -21880 -10700
rect -21620 -10720 -21380 -10700
rect -21120 -10720 -20880 -10700
rect -20620 -10720 -20380 -10700
rect -20120 -10720 -19880 -10700
rect -19620 -10720 -19380 -10700
rect -19120 -10720 -18880 -10700
rect -18620 -10720 -18380 -10700
rect -18120 -10720 -17880 -10700
rect -17620 -10720 -17380 -10700
rect -17120 -10720 -16880 -10700
rect -16620 -10720 -16380 -10700
rect -16120 -10720 -15880 -10700
rect -15620 -10720 -15380 -10700
rect -15120 -10720 -15000 -10700
rect -27500 -10980 -27400 -10720
rect -27100 -10980 -26900 -10720
rect -26600 -10980 -26400 -10720
rect -26100 -10980 -25900 -10720
rect -25600 -10980 -25400 -10720
rect -25100 -10980 -24900 -10720
rect -24600 -10980 -24400 -10720
rect -24100 -10980 -23900 -10720
rect -23600 -10980 -23400 -10720
rect -23100 -10980 -22900 -10720
rect -22600 -10980 -22400 -10720
rect -22100 -10980 -21900 -10720
rect -21600 -10980 -21400 -10720
rect -21100 -10980 -20900 -10720
rect -20600 -10980 -20400 -10720
rect -20100 -10980 -19900 -10720
rect -19600 -10980 -19400 -10720
rect -19100 -10980 -18900 -10720
rect -18600 -10980 -18400 -10720
rect -18100 -10980 -17900 -10720
rect -17600 -10980 -17400 -10720
rect -17100 -10980 -16900 -10720
rect -16600 -10980 -16400 -10720
rect -16100 -10980 -15900 -10720
rect -15600 -10980 -15400 -10720
rect -15100 -10980 -15000 -10720
rect -27500 -11000 -27380 -10980
rect -27120 -11000 -26880 -10980
rect -26620 -11000 -26380 -10980
rect -26120 -11000 -25880 -10980
rect -25620 -11000 -25380 -10980
rect -25120 -11000 -24880 -10980
rect -24620 -11000 -24380 -10980
rect -24120 -11000 -23880 -10980
rect -23620 -11000 -23380 -10980
rect -23120 -11000 -22880 -10980
rect -22620 -11000 -22380 -10980
rect -22120 -11000 -21880 -10980
rect -21620 -11000 -21380 -10980
rect -21120 -11000 -20880 -10980
rect -20620 -11000 -20380 -10980
rect -20120 -11000 -19880 -10980
rect -19620 -11000 -19380 -10980
rect -19120 -11000 -18880 -10980
rect -18620 -11000 -18380 -10980
rect -18120 -11000 -17880 -10980
rect -17620 -11000 -17380 -10980
rect -17120 -11000 -16880 -10980
rect -16620 -11000 -16380 -10980
rect -16120 -11000 -15880 -10980
rect -15620 -11000 -15380 -10980
rect -15120 -11000 -15000 -10980
rect -27500 -11200 -15000 -11000
rect -27500 -11220 -27380 -11200
rect -27120 -11220 -26880 -11200
rect -26620 -11220 -26380 -11200
rect -26120 -11220 -25880 -11200
rect -25620 -11220 -25380 -11200
rect -25120 -11220 -24880 -11200
rect -24620 -11220 -24380 -11200
rect -24120 -11220 -23880 -11200
rect -23620 -11220 -23380 -11200
rect -23120 -11220 -22880 -11200
rect -22620 -11220 -22380 -11200
rect -22120 -11220 -21880 -11200
rect -21620 -11220 -21380 -11200
rect -21120 -11220 -20880 -11200
rect -20620 -11220 -20380 -11200
rect -20120 -11220 -19880 -11200
rect -19620 -11220 -19380 -11200
rect -19120 -11220 -18880 -11200
rect -18620 -11220 -18380 -11200
rect -18120 -11220 -17880 -11200
rect -17620 -11220 -17380 -11200
rect -17120 -11220 -16880 -11200
rect -16620 -11220 -16380 -11200
rect -16120 -11220 -15880 -11200
rect -15620 -11220 -15380 -11200
rect -15120 -11220 -15000 -11200
rect -27500 -11480 -27400 -11220
rect -27100 -11480 -26900 -11220
rect -26600 -11480 -26400 -11220
rect -26100 -11480 -25900 -11220
rect -25600 -11480 -25400 -11220
rect -25100 -11480 -24900 -11220
rect -24600 -11480 -24400 -11220
rect -24100 -11480 -23900 -11220
rect -23600 -11480 -23400 -11220
rect -23100 -11480 -22900 -11220
rect -22600 -11480 -22400 -11220
rect -22100 -11480 -21900 -11220
rect -21600 -11480 -21400 -11220
rect -21100 -11480 -20900 -11220
rect -20600 -11480 -20400 -11220
rect -20100 -11480 -19900 -11220
rect -19600 -11480 -19400 -11220
rect -19100 -11480 -18900 -11220
rect -18600 -11480 -18400 -11220
rect -18100 -11480 -17900 -11220
rect -17600 -11480 -17400 -11220
rect -17100 -11480 -16900 -11220
rect -16600 -11480 -16400 -11220
rect -16100 -11480 -15900 -11220
rect -15600 -11480 -15400 -11220
rect -15100 -11480 -15000 -11220
rect -27500 -11500 -27380 -11480
rect -27120 -11500 -26880 -11480
rect -26620 -11500 -26380 -11480
rect -26120 -11500 -25880 -11480
rect -25620 -11500 -25380 -11480
rect -25120 -11500 -24880 -11480
rect -24620 -11500 -24380 -11480
rect -24120 -11500 -23880 -11480
rect -23620 -11500 -23380 -11480
rect -23120 -11500 -22880 -11480
rect -22620 -11500 -22380 -11480
rect -22120 -11500 -21880 -11480
rect -21620 -11500 -21380 -11480
rect -21120 -11500 -20880 -11480
rect -20620 -11500 -20380 -11480
rect -20120 -11500 -19880 -11480
rect -19620 -11500 -19380 -11480
rect -19120 -11500 -18880 -11480
rect -18620 -11500 -18380 -11480
rect -18120 -11500 -17880 -11480
rect -17620 -11500 -17380 -11480
rect -17120 -11500 -16880 -11480
rect -16620 -11500 -16380 -11480
rect -16120 -11500 -15880 -11480
rect -15620 -11500 -15380 -11480
rect -15120 -11500 -15000 -11480
rect -27500 -11600 -15000 -11500
rect -27500 -11700 -18200 -11600
rect -18000 -11700 -15000 -11600
rect -27500 -11720 -27380 -11700
rect -27120 -11720 -26880 -11700
rect -26620 -11720 -26380 -11700
rect -26120 -11720 -25880 -11700
rect -25620 -11720 -25380 -11700
rect -25120 -11720 -24880 -11700
rect -24620 -11720 -24380 -11700
rect -24120 -11720 -23880 -11700
rect -23620 -11720 -23380 -11700
rect -23120 -11720 -22880 -11700
rect -22620 -11720 -22380 -11700
rect -22120 -11720 -21880 -11700
rect -21620 -11720 -21380 -11700
rect -21120 -11720 -20880 -11700
rect -20620 -11720 -20380 -11700
rect -20120 -11720 -19880 -11700
rect -19620 -11720 -19380 -11700
rect -19120 -11720 -18880 -11700
rect -18620 -11720 -18380 -11700
rect -18000 -11720 -17880 -11700
rect -17620 -11720 -17380 -11700
rect -17120 -11720 -16880 -11700
rect -16620 -11720 -16380 -11700
rect -16120 -11720 -15880 -11700
rect -15620 -11720 -15380 -11700
rect -15120 -11720 -15000 -11700
rect -27500 -11980 -27400 -11720
rect -27100 -11980 -26900 -11720
rect -26600 -11980 -26400 -11720
rect -26100 -11980 -25900 -11720
rect -25600 -11980 -25400 -11720
rect -25100 -11980 -24900 -11720
rect -24600 -11980 -24400 -11720
rect -24100 -11980 -23900 -11720
rect -23600 -11980 -23400 -11720
rect -23100 -11980 -22900 -11720
rect -22600 -11980 -22400 -11720
rect -22100 -11980 -21900 -11720
rect -21600 -11980 -21400 -11720
rect -21100 -11980 -20900 -11720
rect -20600 -11980 -20400 -11720
rect -20100 -11980 -19900 -11720
rect -19600 -11980 -19400 -11720
rect -19100 -11980 -18900 -11720
rect -18600 -11980 -18400 -11720
rect -18000 -11900 -17900 -11720
rect -18100 -11980 -17900 -11900
rect -17600 -11980 -17400 -11720
rect -17100 -11980 -16900 -11720
rect -16600 -11980 -16400 -11720
rect -16100 -11980 -15900 -11720
rect -15600 -11980 -15400 -11720
rect -15100 -11980 -15000 -11720
rect -27500 -12000 -27380 -11980
rect -27120 -12000 -26880 -11980
rect -26620 -12000 -26380 -11980
rect -26120 -12000 -25880 -11980
rect -25620 -12000 -25380 -11980
rect -25120 -12000 -24880 -11980
rect -24620 -12000 -24380 -11980
rect -24120 -12000 -23880 -11980
rect -23620 -12000 -23380 -11980
rect -23120 -12000 -22880 -11980
rect -22620 -12000 -22380 -11980
rect -22120 -12000 -21880 -11980
rect -21620 -12000 -21380 -11980
rect -21120 -12000 -20880 -11980
rect -20620 -12000 -20380 -11980
rect -20120 -12000 -19880 -11980
rect -19620 -12000 -19380 -11980
rect -19120 -12000 -18880 -11980
rect -18620 -12000 -18380 -11980
rect -18120 -12000 -17880 -11980
rect -17620 -12000 -17380 -11980
rect -17120 -12000 -16880 -11980
rect -16620 -12000 -16380 -11980
rect -16120 -12000 -15880 -11980
rect -15620 -12000 -15380 -11980
rect -15120 -12000 -15000 -11980
rect -27500 -12200 -15000 -12000
rect -27500 -12220 -27380 -12200
rect -27120 -12220 -26880 -12200
rect -26620 -12220 -26380 -12200
rect -26120 -12220 -25880 -12200
rect -25620 -12220 -25380 -12200
rect -25120 -12220 -24880 -12200
rect -24620 -12220 -24380 -12200
rect -24120 -12220 -23880 -12200
rect -23620 -12220 -23380 -12200
rect -23120 -12220 -22880 -12200
rect -22620 -12220 -22380 -12200
rect -22120 -12220 -21880 -12200
rect -21620 -12220 -21380 -12200
rect -21120 -12220 -20880 -12200
rect -20620 -12220 -20380 -12200
rect -20120 -12220 -19880 -12200
rect -19620 -12220 -19380 -12200
rect -19120 -12220 -18880 -12200
rect -18620 -12220 -18380 -12200
rect -18120 -12220 -17880 -12200
rect -17620 -12220 -17380 -12200
rect -17120 -12220 -16880 -12200
rect -16620 -12220 -16380 -12200
rect -16120 -12220 -15880 -12200
rect -15620 -12220 -15380 -12200
rect -15120 -12220 -15000 -12200
rect -27500 -12480 -27400 -12220
rect -27100 -12480 -26900 -12220
rect -26600 -12480 -26400 -12220
rect -26100 -12480 -25900 -12220
rect -25600 -12480 -25400 -12220
rect -25100 -12480 -24900 -12220
rect -24600 -12480 -24400 -12220
rect -24100 -12480 -23900 -12220
rect -23600 -12480 -23400 -12220
rect -23100 -12480 -22900 -12220
rect -22600 -12480 -22400 -12220
rect -22100 -12480 -21900 -12220
rect -21600 -12480 -21400 -12220
rect -21100 -12480 -20900 -12220
rect -20600 -12480 -20400 -12220
rect -20100 -12480 -19900 -12220
rect -19600 -12480 -19400 -12220
rect -19100 -12480 -18900 -12220
rect -18600 -12480 -18400 -12220
rect -18100 -12480 -17900 -12220
rect -17600 -12480 -17400 -12220
rect -17100 -12480 -16900 -12220
rect -16600 -12480 -16400 -12220
rect -16100 -12480 -15900 -12220
rect -15600 -12480 -15400 -12220
rect -15100 -12480 -15000 -12220
rect -27500 -12500 -27380 -12480
rect -27120 -12500 -26880 -12480
rect -26620 -12500 -26380 -12480
rect -26120 -12500 -25880 -12480
rect -25620 -12500 -25380 -12480
rect -25120 -12500 -24880 -12480
rect -24620 -12500 -24380 -12480
rect -24120 -12500 -23880 -12480
rect -23620 -12500 -23380 -12480
rect -23120 -12500 -22880 -12480
rect -22620 -12500 -22380 -12480
rect -22120 -12500 -21880 -12480
rect -21620 -12500 -21380 -12480
rect -21120 -12500 -20880 -12480
rect -20620 -12500 -20380 -12480
rect -20120 -12500 -19880 -12480
rect -19620 -12500 -19380 -12480
rect -19120 -12500 -18880 -12480
rect -18620 -12500 -18380 -12480
rect -18120 -12500 -17880 -12480
rect -17620 -12500 -17380 -12480
rect -17120 -12500 -16880 -12480
rect -16620 -12500 -16380 -12480
rect -16120 -12500 -15880 -12480
rect -15620 -12500 -15380 -12480
rect -15120 -12500 -15000 -12480
rect -27500 -12700 -15000 -12500
rect -27500 -12720 -27380 -12700
rect -27120 -12720 -26880 -12700
rect -26620 -12720 -26380 -12700
rect -26120 -12720 -25880 -12700
rect -25620 -12720 -25380 -12700
rect -25120 -12720 -24880 -12700
rect -24620 -12720 -24380 -12700
rect -24120 -12720 -23880 -12700
rect -23620 -12720 -23380 -12700
rect -23120 -12720 -22880 -12700
rect -22620 -12720 -22380 -12700
rect -22120 -12720 -21880 -12700
rect -21620 -12720 -21380 -12700
rect -21120 -12720 -20880 -12700
rect -20620 -12720 -20380 -12700
rect -20120 -12720 -19880 -12700
rect -19620 -12720 -19380 -12700
rect -19120 -12720 -18880 -12700
rect -18620 -12720 -18380 -12700
rect -18120 -12720 -17880 -12700
rect -17620 -12720 -17380 -12700
rect -17120 -12720 -16880 -12700
rect -16620 -12720 -16380 -12700
rect -16120 -12720 -15880 -12700
rect -15620 -12720 -15380 -12700
rect -15120 -12720 -15000 -12700
rect -27500 -12980 -27400 -12720
rect -27100 -12980 -26900 -12720
rect -26600 -12980 -26400 -12720
rect -26100 -12980 -25900 -12720
rect -25600 -12980 -25400 -12720
rect -25100 -12980 -24900 -12720
rect -24600 -12980 -24400 -12720
rect -24100 -12980 -23900 -12720
rect -23600 -12980 -23400 -12720
rect -23100 -12980 -22900 -12720
rect -22600 -12980 -22400 -12720
rect -22100 -12980 -21900 -12720
rect -21600 -12980 -21400 -12720
rect -21100 -12980 -20900 -12720
rect -20600 -12980 -20400 -12720
rect -20100 -12980 -19900 -12720
rect -19600 -12980 -19400 -12720
rect -19100 -12980 -18900 -12720
rect -18600 -12980 -18400 -12720
rect -18100 -12980 -17900 -12720
rect -17600 -12980 -17400 -12720
rect -17100 -12980 -16900 -12720
rect -16600 -12980 -16400 -12720
rect -16100 -12980 -15900 -12720
rect -15600 -12980 -15400 -12720
rect -15100 -12980 -15000 -12720
rect -27500 -13000 -27380 -12980
rect -27120 -13000 -26880 -12980
rect -26620 -13000 -26380 -12980
rect -26120 -13000 -25880 -12980
rect -25620 -13000 -25380 -12980
rect -25120 -13000 -24880 -12980
rect -24620 -13000 -24380 -12980
rect -24120 -13000 -23880 -12980
rect -23620 -13000 -23380 -12980
rect -23120 -13000 -22880 -12980
rect -22620 -13000 -22380 -12980
rect -22120 -13000 -21880 -12980
rect -21620 -13000 -21380 -12980
rect -21120 -13000 -20880 -12980
rect -20620 -13000 -20380 -12980
rect -20120 -13000 -19880 -12980
rect -19620 -13000 -19380 -12980
rect -19120 -13000 -18880 -12980
rect -18620 -13000 -18380 -12980
rect -18120 -13000 -17880 -12980
rect -17620 -13000 -17380 -12980
rect -17120 -13000 -16880 -12980
rect -16620 -13000 -16380 -12980
rect -16120 -13000 -15880 -12980
rect -15620 -13000 -15380 -12980
rect -15120 -13000 -15000 -12980
rect -27500 -13200 -15000 -13000
rect 14500 -3700 33500 -3600
rect 14500 -3720 14620 -3700
rect 14880 -3720 15120 -3700
rect 15380 -3720 15620 -3700
rect 15880 -3720 16120 -3700
rect 16380 -3720 16620 -3700
rect 16880 -3720 17120 -3700
rect 17380 -3720 17620 -3700
rect 17880 -3720 18120 -3700
rect 18380 -3720 18620 -3700
rect 18880 -3720 19120 -3700
rect 19380 -3720 19620 -3700
rect 19880 -3720 20120 -3700
rect 20380 -3720 20620 -3700
rect 20880 -3720 21120 -3700
rect 21380 -3720 21620 -3700
rect 21880 -3720 22120 -3700
rect 22380 -3720 22620 -3700
rect 22880 -3720 23120 -3700
rect 23380 -3720 23620 -3700
rect 23880 -3720 24120 -3700
rect 24380 -3720 24620 -3700
rect 24880 -3720 25120 -3700
rect 25380 -3720 25620 -3700
rect 25880 -3720 26120 -3700
rect 26380 -3720 26620 -3700
rect 26880 -3720 27120 -3700
rect 27380 -3720 27620 -3700
rect 27880 -3720 28120 -3700
rect 28380 -3720 28620 -3700
rect 28880 -3720 29120 -3700
rect 29380 -3720 29620 -3700
rect 29880 -3720 30120 -3700
rect 30380 -3720 30620 -3700
rect 30880 -3720 31120 -3700
rect 31380 -3720 31620 -3700
rect 31880 -3720 32120 -3700
rect 32380 -3720 32620 -3700
rect 32880 -3720 33120 -3700
rect 33380 -3720 33500 -3700
rect 14500 -3980 14600 -3720
rect 14900 -3980 15100 -3720
rect 15400 -3980 15600 -3720
rect 15900 -3980 16100 -3720
rect 16400 -3980 16600 -3720
rect 16900 -3980 17100 -3720
rect 17400 -3980 17600 -3720
rect 17900 -3980 18100 -3720
rect 18400 -3980 18600 -3720
rect 18900 -3980 19100 -3720
rect 19400 -3980 19600 -3720
rect 19900 -3980 20100 -3720
rect 20400 -3980 20600 -3720
rect 20900 -3980 21100 -3720
rect 21400 -3980 21600 -3720
rect 21900 -3980 22100 -3720
rect 22400 -3980 22600 -3720
rect 22900 -3980 23100 -3720
rect 23400 -3980 23600 -3720
rect 23900 -3980 24100 -3720
rect 24400 -3980 24600 -3720
rect 24900 -3980 25100 -3720
rect 25400 -3980 25600 -3720
rect 25900 -3980 26100 -3720
rect 26400 -3980 26600 -3720
rect 26900 -3980 27100 -3720
rect 27400 -3980 27600 -3720
rect 27900 -3980 28100 -3720
rect 28400 -3980 28600 -3720
rect 28900 -3980 29100 -3720
rect 29400 -3980 29600 -3720
rect 29900 -3980 30100 -3720
rect 30400 -3980 30600 -3720
rect 30900 -3980 31100 -3720
rect 31400 -3980 31600 -3720
rect 31900 -3980 32100 -3720
rect 32400 -3980 32600 -3720
rect 32900 -3980 33100 -3720
rect 33400 -3980 33500 -3720
rect 14500 -4000 14620 -3980
rect 14880 -4000 15120 -3980
rect 15380 -4000 15620 -3980
rect 15880 -4000 16120 -3980
rect 16380 -4000 16620 -3980
rect 16880 -4000 17120 -3980
rect 17380 -4000 17620 -3980
rect 17880 -4000 18120 -3980
rect 18380 -4000 18620 -3980
rect 18880 -4000 19120 -3980
rect 19380 -4000 19620 -3980
rect 19880 -4000 20120 -3980
rect 20380 -4000 20620 -3980
rect 20880 -4000 21120 -3980
rect 21380 -4000 21620 -3980
rect 21880 -4000 22120 -3980
rect 22380 -4000 22620 -3980
rect 22880 -4000 23120 -3980
rect 23380 -4000 23620 -3980
rect 23880 -4000 24120 -3980
rect 24380 -4000 24620 -3980
rect 24880 -4000 25120 -3980
rect 25380 -4000 25620 -3980
rect 25880 -4000 26120 -3980
rect 26380 -4000 26620 -3980
rect 26880 -4000 27120 -3980
rect 27380 -4000 27620 -3980
rect 27880 -4000 28120 -3980
rect 28380 -4000 28620 -3980
rect 28880 -4000 29120 -3980
rect 29380 -4000 29620 -3980
rect 29880 -4000 30120 -3980
rect 30380 -4000 30620 -3980
rect 30880 -4000 31120 -3980
rect 31380 -4000 31620 -3980
rect 31880 -4000 32120 -3980
rect 32380 -4000 32620 -3980
rect 32880 -4000 33120 -3980
rect 33380 -4000 33500 -3980
rect 14500 -4200 33500 -4000
rect 14500 -4220 14620 -4200
rect 14880 -4220 15120 -4200
rect 15380 -4220 15620 -4200
rect 15880 -4220 16120 -4200
rect 16380 -4220 16620 -4200
rect 16880 -4220 17120 -4200
rect 17380 -4220 17620 -4200
rect 17880 -4220 18120 -4200
rect 18380 -4220 18620 -4200
rect 18880 -4220 19120 -4200
rect 19380 -4220 19620 -4200
rect 19880 -4220 20120 -4200
rect 20380 -4220 20620 -4200
rect 20880 -4220 21120 -4200
rect 21380 -4220 21620 -4200
rect 21880 -4220 22120 -4200
rect 22380 -4220 22620 -4200
rect 22880 -4220 23120 -4200
rect 23380 -4220 23620 -4200
rect 23880 -4220 24120 -4200
rect 24380 -4220 24620 -4200
rect 24880 -4220 25120 -4200
rect 25380 -4220 25620 -4200
rect 25880 -4220 26120 -4200
rect 26380 -4220 26620 -4200
rect 26880 -4220 27120 -4200
rect 27380 -4220 27620 -4200
rect 27880 -4220 28120 -4200
rect 28380 -4220 28620 -4200
rect 28880 -4220 29120 -4200
rect 29380 -4220 29620 -4200
rect 29880 -4220 30120 -4200
rect 30380 -4220 30620 -4200
rect 30880 -4220 31120 -4200
rect 31380 -4220 31620 -4200
rect 31880 -4220 32120 -4200
rect 32380 -4220 32620 -4200
rect 32880 -4220 33120 -4200
rect 33380 -4220 33500 -4200
rect 14500 -4480 14600 -4220
rect 14900 -4480 15100 -4220
rect 15400 -4480 15600 -4220
rect 15900 -4480 16100 -4220
rect 16400 -4480 16600 -4220
rect 16900 -4480 17100 -4220
rect 17400 -4480 17600 -4220
rect 17900 -4480 18100 -4220
rect 18400 -4480 18600 -4220
rect 18900 -4480 19100 -4220
rect 19400 -4480 19600 -4220
rect 19900 -4480 20100 -4220
rect 20400 -4480 20600 -4220
rect 20900 -4480 21100 -4220
rect 21400 -4480 21600 -4220
rect 21900 -4480 22100 -4220
rect 22400 -4480 22600 -4220
rect 22900 -4480 23100 -4220
rect 23400 -4480 23600 -4220
rect 23900 -4480 24100 -4220
rect 24400 -4480 24600 -4220
rect 24900 -4480 25100 -4220
rect 25400 -4480 25600 -4220
rect 25900 -4480 26100 -4220
rect 26400 -4480 26600 -4220
rect 26900 -4480 27100 -4220
rect 27400 -4480 27600 -4220
rect 27900 -4480 28100 -4220
rect 28400 -4480 28600 -4220
rect 28900 -4480 29100 -4220
rect 29400 -4480 29600 -4220
rect 29900 -4480 30100 -4220
rect 30400 -4480 30600 -4220
rect 30900 -4480 31100 -4220
rect 31400 -4480 31600 -4220
rect 31900 -4480 32100 -4220
rect 32400 -4480 32600 -4220
rect 32900 -4480 33100 -4220
rect 33400 -4480 33500 -4220
rect 14500 -4500 14620 -4480
rect 14880 -4500 15120 -4480
rect 15380 -4500 15620 -4480
rect 15880 -4500 16120 -4480
rect 16380 -4500 16620 -4480
rect 16880 -4500 17120 -4480
rect 17380 -4500 17620 -4480
rect 17880 -4500 18120 -4480
rect 18380 -4500 18620 -4480
rect 18880 -4500 19120 -4480
rect 19380 -4500 19620 -4480
rect 19880 -4500 20120 -4480
rect 20380 -4500 20620 -4480
rect 20880 -4500 21120 -4480
rect 21380 -4500 21620 -4480
rect 21880 -4500 22120 -4480
rect 22380 -4500 22620 -4480
rect 22880 -4500 23120 -4480
rect 23380 -4500 23620 -4480
rect 23880 -4500 24120 -4480
rect 24380 -4500 24620 -4480
rect 24880 -4500 25120 -4480
rect 25380 -4500 25620 -4480
rect 25880 -4500 26120 -4480
rect 26380 -4500 26620 -4480
rect 26880 -4500 27120 -4480
rect 27380 -4500 27620 -4480
rect 27880 -4500 28120 -4480
rect 28380 -4500 28620 -4480
rect 28880 -4500 29120 -4480
rect 29380 -4500 29620 -4480
rect 29880 -4500 30120 -4480
rect 30380 -4500 30620 -4480
rect 30880 -4500 31120 -4480
rect 31380 -4500 31620 -4480
rect 31880 -4500 32120 -4480
rect 32380 -4500 32620 -4480
rect 32880 -4500 33120 -4480
rect 33380 -4500 33500 -4480
rect 14500 -4700 33500 -4500
rect 14500 -4720 14620 -4700
rect 14880 -4720 15120 -4700
rect 15380 -4720 15620 -4700
rect 15880 -4720 16120 -4700
rect 16380 -4720 16620 -4700
rect 16880 -4720 17120 -4700
rect 17380 -4720 17620 -4700
rect 17880 -4720 18120 -4700
rect 18380 -4720 18620 -4700
rect 18880 -4720 19120 -4700
rect 19380 -4720 19620 -4700
rect 19880 -4720 20120 -4700
rect 20380 -4720 20620 -4700
rect 20880 -4720 21120 -4700
rect 21380 -4720 21620 -4700
rect 21880 -4720 22120 -4700
rect 22380 -4720 22620 -4700
rect 22880 -4720 23120 -4700
rect 23380 -4720 23620 -4700
rect 23880 -4720 24120 -4700
rect 24380 -4720 24620 -4700
rect 24880 -4720 25120 -4700
rect 25380 -4720 25620 -4700
rect 25880 -4720 26120 -4700
rect 26380 -4720 26620 -4700
rect 26880 -4720 27120 -4700
rect 27380 -4720 27620 -4700
rect 27880 -4720 28120 -4700
rect 28380 -4720 28620 -4700
rect 28880 -4720 29120 -4700
rect 29380 -4720 29620 -4700
rect 29880 -4720 30120 -4700
rect 30380 -4720 30620 -4700
rect 30880 -4720 31120 -4700
rect 31380 -4720 31620 -4700
rect 31880 -4720 32120 -4700
rect 32380 -4720 32620 -4700
rect 32880 -4720 33120 -4700
rect 33380 -4720 33500 -4700
rect 14500 -4980 14600 -4720
rect 14900 -4980 15100 -4720
rect 15400 -4980 15600 -4720
rect 15900 -4980 16100 -4720
rect 16400 -4980 16600 -4720
rect 16900 -4980 17100 -4720
rect 17400 -4980 17600 -4720
rect 17900 -4980 18100 -4720
rect 18400 -4980 18600 -4720
rect 18900 -4980 19100 -4720
rect 19400 -4980 19600 -4720
rect 19900 -4980 20100 -4720
rect 20400 -4980 20600 -4720
rect 20900 -4980 21100 -4720
rect 21400 -4980 21600 -4720
rect 21900 -4980 22100 -4720
rect 22400 -4980 22600 -4720
rect 22900 -4980 23100 -4720
rect 23400 -4980 23600 -4720
rect 23900 -4980 24100 -4720
rect 24400 -4980 24600 -4720
rect 24900 -4980 25100 -4720
rect 25400 -4980 25600 -4720
rect 25900 -4980 26100 -4720
rect 26400 -4980 26600 -4720
rect 26900 -4980 27100 -4720
rect 27400 -4980 27600 -4720
rect 27900 -4980 28100 -4720
rect 28400 -4980 28600 -4720
rect 28900 -4980 29100 -4720
rect 29400 -4980 29600 -4720
rect 29900 -4980 30100 -4720
rect 30400 -4980 30600 -4720
rect 30900 -4980 31100 -4720
rect 31400 -4980 31600 -4720
rect 31900 -4980 32100 -4720
rect 32400 -4980 32600 -4720
rect 32900 -4980 33100 -4720
rect 33400 -4980 33500 -4720
rect 14500 -5000 14620 -4980
rect 14880 -5000 15120 -4980
rect 15380 -5000 15620 -4980
rect 15880 -5000 16120 -4980
rect 16380 -5000 16620 -4980
rect 16880 -5000 17120 -4980
rect 17380 -5000 17620 -4980
rect 17880 -5000 18120 -4980
rect 18380 -5000 18620 -4980
rect 18880 -5000 19120 -4980
rect 19380 -5000 19620 -4980
rect 19880 -5000 20120 -4980
rect 20380 -5000 20620 -4980
rect 20880 -5000 21120 -4980
rect 21380 -5000 21620 -4980
rect 21880 -5000 22120 -4980
rect 22380 -5000 22620 -4980
rect 22880 -5000 23120 -4980
rect 23380 -5000 23620 -4980
rect 23880 -5000 24120 -4980
rect 24380 -5000 24620 -4980
rect 24880 -5000 25120 -4980
rect 25380 -5000 25620 -4980
rect 25880 -5000 26120 -4980
rect 26380 -5000 26620 -4980
rect 26880 -5000 27120 -4980
rect 27380 -5000 27620 -4980
rect 27880 -5000 28120 -4980
rect 28380 -5000 28620 -4980
rect 28880 -5000 29120 -4980
rect 29380 -5000 29620 -4980
rect 29880 -5000 30120 -4980
rect 30380 -5000 30620 -4980
rect 30880 -5000 31120 -4980
rect 31380 -5000 31620 -4980
rect 31880 -5000 32120 -4980
rect 32380 -5000 32620 -4980
rect 32880 -5000 33120 -4980
rect 33380 -5000 33500 -4980
rect 14500 -5200 33500 -5000
rect 14500 -5220 14620 -5200
rect 14880 -5220 15120 -5200
rect 15380 -5220 15620 -5200
rect 15880 -5220 16120 -5200
rect 16380 -5220 16620 -5200
rect 16880 -5220 17120 -5200
rect 17380 -5220 17620 -5200
rect 17880 -5220 18120 -5200
rect 18380 -5220 18620 -5200
rect 18880 -5220 19120 -5200
rect 19380 -5220 19620 -5200
rect 19880 -5220 20120 -5200
rect 20380 -5220 20620 -5200
rect 20880 -5220 21120 -5200
rect 21380 -5220 21620 -5200
rect 21880 -5220 22120 -5200
rect 22380 -5220 22620 -5200
rect 22880 -5220 23120 -5200
rect 23380 -5220 23620 -5200
rect 23880 -5220 24120 -5200
rect 24380 -5220 24620 -5200
rect 24880 -5220 25120 -5200
rect 25380 -5220 25620 -5200
rect 25880 -5220 26120 -5200
rect 26380 -5220 26620 -5200
rect 26880 -5220 27120 -5200
rect 27380 -5220 27620 -5200
rect 27880 -5220 28120 -5200
rect 28380 -5220 28620 -5200
rect 28880 -5220 29120 -5200
rect 29380 -5220 29620 -5200
rect 29880 -5220 30120 -5200
rect 30380 -5220 30620 -5200
rect 30880 -5220 31120 -5200
rect 31380 -5220 31620 -5200
rect 31880 -5220 32120 -5200
rect 32380 -5220 32620 -5200
rect 32880 -5220 33120 -5200
rect 33380 -5220 33500 -5200
rect 14500 -5480 14600 -5220
rect 14900 -5480 15100 -5220
rect 15400 -5480 15600 -5220
rect 15900 -5480 16100 -5220
rect 16400 -5480 16600 -5220
rect 16900 -5480 17100 -5220
rect 17400 -5480 17600 -5220
rect 17900 -5480 18100 -5220
rect 18400 -5480 18600 -5220
rect 18900 -5480 19100 -5220
rect 19400 -5480 19600 -5220
rect 19900 -5480 20100 -5220
rect 20400 -5480 20600 -5220
rect 20900 -5480 21100 -5220
rect 21400 -5480 21600 -5220
rect 21900 -5480 22100 -5220
rect 22400 -5480 22600 -5220
rect 22900 -5480 23100 -5220
rect 23400 -5480 23600 -5220
rect 23900 -5480 24100 -5220
rect 24400 -5480 24600 -5220
rect 24900 -5480 25100 -5220
rect 25400 -5480 25600 -5220
rect 25900 -5480 26100 -5220
rect 26400 -5480 26600 -5220
rect 26900 -5480 27100 -5220
rect 27400 -5480 27600 -5220
rect 27900 -5480 28100 -5220
rect 28400 -5480 28600 -5220
rect 28900 -5480 29100 -5220
rect 29400 -5480 29600 -5220
rect 29900 -5480 30100 -5220
rect 30400 -5480 30600 -5220
rect 30900 -5480 31100 -5220
rect 31400 -5480 31600 -5220
rect 31900 -5480 32100 -5220
rect 32400 -5480 32600 -5220
rect 32900 -5480 33100 -5220
rect 33400 -5480 33500 -5220
rect 14500 -5500 14620 -5480
rect 14880 -5500 15120 -5480
rect 15380 -5500 15620 -5480
rect 15880 -5500 16120 -5480
rect 16380 -5500 16620 -5480
rect 16880 -5500 17120 -5480
rect 17380 -5500 17620 -5480
rect 17880 -5500 18120 -5480
rect 18380 -5500 18620 -5480
rect 18880 -5500 19120 -5480
rect 19380 -5500 19620 -5480
rect 19880 -5500 20120 -5480
rect 20380 -5500 20620 -5480
rect 20880 -5500 21120 -5480
rect 21380 -5500 21620 -5480
rect 21880 -5500 22120 -5480
rect 22380 -5500 22620 -5480
rect 22880 -5500 23120 -5480
rect 23380 -5500 23620 -5480
rect 23880 -5500 24120 -5480
rect 24380 -5500 24620 -5480
rect 24880 -5500 25120 -5480
rect 25380 -5500 25620 -5480
rect 25880 -5500 26120 -5480
rect 26380 -5500 26620 -5480
rect 26880 -5500 27120 -5480
rect 27380 -5500 27620 -5480
rect 27880 -5500 28120 -5480
rect 28380 -5500 28620 -5480
rect 28880 -5500 29120 -5480
rect 29380 -5500 29620 -5480
rect 29880 -5500 30120 -5480
rect 30380 -5500 30620 -5480
rect 30880 -5500 31120 -5480
rect 31380 -5500 31620 -5480
rect 31880 -5500 32120 -5480
rect 32380 -5500 32620 -5480
rect 32880 -5500 33120 -5480
rect 33380 -5500 33500 -5480
rect 14500 -5600 33500 -5500
rect 14500 -5700 24000 -5600
rect 14500 -5720 14620 -5700
rect 14880 -5720 15120 -5700
rect 15380 -5720 15620 -5700
rect 15880 -5720 16120 -5700
rect 16380 -5720 16620 -5700
rect 16880 -5720 17120 -5700
rect 17380 -5720 17620 -5700
rect 17880 -5720 18120 -5700
rect 18380 -5720 18620 -5700
rect 18880 -5720 19120 -5700
rect 19380 -5720 19620 -5700
rect 19880 -5720 20120 -5700
rect 20380 -5720 20620 -5700
rect 20880 -5720 21120 -5700
rect 21380 -5720 21620 -5700
rect 21880 -5720 22120 -5700
rect 22380 -5720 22620 -5700
rect 22880 -5720 23120 -5700
rect 23380 -5720 23620 -5700
rect 23880 -5720 24000 -5700
rect 14500 -5980 14600 -5720
rect 14900 -5980 15100 -5720
rect 15400 -5980 15600 -5720
rect 15900 -5980 16100 -5720
rect 16400 -5980 16600 -5720
rect 16900 -5980 17100 -5720
rect 17400 -5980 17600 -5720
rect 17900 -5980 18100 -5720
rect 18400 -5980 18600 -5720
rect 18900 -5980 19100 -5720
rect 19400 -5980 19600 -5720
rect 19900 -5980 20100 -5720
rect 20400 -5980 20600 -5720
rect 20900 -5980 21100 -5720
rect 21400 -5980 21600 -5720
rect 21900 -5980 22100 -5720
rect 22400 -5980 22600 -5720
rect 22900 -5980 23100 -5720
rect 23400 -5980 23600 -5720
rect 23900 -5980 24000 -5720
rect 14500 -6000 14620 -5980
rect 14880 -6000 15120 -5980
rect 15380 -6000 15620 -5980
rect 15880 -6000 16120 -5980
rect 16380 -6000 16620 -5980
rect 16880 -6000 17120 -5980
rect 17380 -6000 17620 -5980
rect 17880 -6000 18120 -5980
rect 18380 -6000 18620 -5980
rect 18880 -6000 19120 -5980
rect 19380 -6000 19620 -5980
rect 19880 -6000 20120 -5980
rect 20380 -6000 20620 -5980
rect 20880 -6000 21120 -5980
rect 21380 -6000 21620 -5980
rect 21880 -6000 22120 -5980
rect 22380 -6000 22620 -5980
rect 22880 -6000 23120 -5980
rect 23380 -6000 23620 -5980
rect 23880 -6000 24000 -5980
rect 14500 -6200 24000 -6000
rect 14500 -6220 14620 -6200
rect 14880 -6220 15120 -6200
rect 15380 -6220 15620 -6200
rect 15880 -6220 16120 -6200
rect 16380 -6220 16620 -6200
rect 16880 -6220 17120 -6200
rect 17380 -6220 17620 -6200
rect 17880 -6220 18120 -6200
rect 18380 -6220 18620 -6200
rect 18880 -6220 19120 -6200
rect 19380 -6220 19620 -6200
rect 19880 -6220 20120 -6200
rect 20380 -6220 20620 -6200
rect 20880 -6220 21120 -6200
rect 21380 -6220 21620 -6200
rect 21880 -6220 22120 -6200
rect 22380 -6220 22620 -6200
rect 22880 -6220 23120 -6200
rect 23380 -6220 23620 -6200
rect 23880 -6220 24000 -6200
rect 14500 -6480 14600 -6220
rect 14900 -6480 15100 -6220
rect 15400 -6480 15600 -6220
rect 15900 -6480 16100 -6220
rect 16400 -6480 16600 -6220
rect 16900 -6480 17100 -6220
rect 17400 -6480 17600 -6220
rect 17900 -6480 18100 -6220
rect 18400 -6480 18600 -6220
rect 18900 -6480 19100 -6220
rect 19400 -6480 19600 -6220
rect 19900 -6480 20100 -6220
rect 20400 -6480 20600 -6220
rect 20900 -6480 21100 -6220
rect 21400 -6480 21600 -6220
rect 21900 -6480 22100 -6220
rect 22400 -6480 22600 -6220
rect 22900 -6480 23100 -6220
rect 23400 -6480 23600 -6220
rect 23900 -6480 24000 -6220
rect 14500 -6500 14620 -6480
rect 14880 -6500 15120 -6480
rect 15380 -6500 15620 -6480
rect 15880 -6500 16120 -6480
rect 16380 -6500 16620 -6480
rect 16880 -6500 17120 -6480
rect 17380 -6500 17620 -6480
rect 17880 -6500 18120 -6480
rect 18380 -6500 18620 -6480
rect 18880 -6500 19120 -6480
rect 19380 -6500 19620 -6480
rect 19880 -6500 20120 -6480
rect 20380 -6500 20620 -6480
rect 20880 -6500 21120 -6480
rect 21380 -6500 21620 -6480
rect 21880 -6500 22120 -6480
rect 22380 -6500 22620 -6480
rect 22880 -6500 23120 -6480
rect 23380 -6500 23620 -6480
rect 23880 -6500 24000 -6480
rect 14500 -6700 24000 -6500
rect 14500 -6720 14620 -6700
rect 14880 -6720 15120 -6700
rect 15380 -6720 15620 -6700
rect 15880 -6720 16120 -6700
rect 16380 -6720 16620 -6700
rect 16880 -6720 17120 -6700
rect 17380 -6720 17620 -6700
rect 17880 -6720 18120 -6700
rect 18380 -6720 18620 -6700
rect 18880 -6720 19120 -6700
rect 19380 -6720 19620 -6700
rect 19880 -6720 20120 -6700
rect 20380 -6720 20620 -6700
rect 20880 -6720 21120 -6700
rect 21380 -6720 21620 -6700
rect 21880 -6720 22120 -6700
rect 22380 -6720 22620 -6700
rect 22880 -6720 23120 -6700
rect 23380 -6720 23620 -6700
rect 23880 -6720 24000 -6700
rect 14500 -6980 14600 -6720
rect 14900 -6980 15100 -6720
rect 15400 -6980 15600 -6720
rect 15900 -6980 16100 -6720
rect 16400 -6980 16600 -6720
rect 16900 -6980 17100 -6720
rect 17400 -6980 17600 -6720
rect 17900 -6980 18100 -6720
rect 18400 -6980 18600 -6720
rect 18900 -6980 19100 -6720
rect 19400 -6980 19600 -6720
rect 19900 -6980 20100 -6720
rect 20400 -6980 20600 -6720
rect 20900 -6980 21100 -6720
rect 21400 -6980 21600 -6720
rect 21900 -6980 22100 -6720
rect 22400 -6980 22600 -6720
rect 22900 -6980 23100 -6720
rect 23400 -6980 23600 -6720
rect 23900 -6980 24000 -6720
rect 14500 -7000 14620 -6980
rect 14880 -7000 15120 -6980
rect 15380 -7000 15620 -6980
rect 15880 -7000 16120 -6980
rect 16380 -7000 16620 -6980
rect 16880 -7000 17120 -6980
rect 17380 -7000 17620 -6980
rect 17880 -7000 18120 -6980
rect 18380 -7000 18620 -6980
rect 18880 -7000 19120 -6980
rect 19380 -7000 19620 -6980
rect 19880 -7000 20120 -6980
rect 20380 -7000 20620 -6980
rect 20880 -7000 21120 -6980
rect 21380 -7000 21620 -6980
rect 21880 -7000 22120 -6980
rect 22380 -7000 22620 -6980
rect 22880 -7000 23120 -6980
rect 23380 -7000 23620 -6980
rect 23880 -7000 24000 -6980
rect 14500 -7200 24000 -7000
rect 14500 -7220 14620 -7200
rect 14880 -7220 15120 -7200
rect 15380 -7220 15620 -7200
rect 15880 -7220 16120 -7200
rect 16380 -7220 16620 -7200
rect 16880 -7220 17120 -7200
rect 17380 -7220 17620 -7200
rect 17880 -7220 18120 -7200
rect 18380 -7220 18620 -7200
rect 18880 -7220 19120 -7200
rect 19380 -7220 19620 -7200
rect 19880 -7220 20120 -7200
rect 20380 -7220 20620 -7200
rect 20880 -7220 21120 -7200
rect 21380 -7220 21620 -7200
rect 21880 -7220 22120 -7200
rect 22380 -7220 22620 -7200
rect 22880 -7220 23120 -7200
rect 23380 -7220 23620 -7200
rect 23880 -7220 24000 -7200
rect 14500 -7480 14600 -7220
rect 14900 -7480 15100 -7220
rect 15400 -7480 15600 -7220
rect 15900 -7480 16100 -7220
rect 16400 -7480 16600 -7220
rect 16900 -7480 17100 -7220
rect 17400 -7480 17600 -7220
rect 17900 -7480 18100 -7220
rect 18400 -7480 18600 -7220
rect 18900 -7480 19100 -7220
rect 19400 -7480 19600 -7220
rect 19900 -7480 20100 -7220
rect 20400 -7480 20600 -7220
rect 20900 -7480 21100 -7220
rect 21400 -7480 21600 -7220
rect 21900 -7480 22100 -7220
rect 22400 -7480 22600 -7220
rect 22900 -7480 23100 -7220
rect 23400 -7480 23600 -7220
rect 23900 -7480 24000 -7220
rect 14500 -7500 14620 -7480
rect 14880 -7500 15120 -7480
rect 15380 -7500 15620 -7480
rect 15880 -7500 16120 -7480
rect 16380 -7500 16620 -7480
rect 16880 -7500 17120 -7480
rect 17380 -7500 17620 -7480
rect 17880 -7500 18120 -7480
rect 18380 -7500 18620 -7480
rect 18880 -7500 19120 -7480
rect 19380 -7500 19620 -7480
rect 19880 -7500 20120 -7480
rect 20380 -7500 20620 -7480
rect 20880 -7500 21120 -7480
rect 21380 -7500 21620 -7480
rect 21880 -7500 22120 -7480
rect 22380 -7500 22620 -7480
rect 22880 -7500 23120 -7480
rect 23380 -7500 23620 -7480
rect 23880 -7500 24000 -7480
rect 14500 -7700 24000 -7500
rect 14500 -7720 14620 -7700
rect 14880 -7720 15120 -7700
rect 15380 -7720 15620 -7700
rect 15880 -7720 16120 -7700
rect 16380 -7720 16620 -7700
rect 16880 -7720 17120 -7700
rect 17380 -7720 17620 -7700
rect 17880 -7720 18120 -7700
rect 18380 -7720 18620 -7700
rect 18880 -7720 19120 -7700
rect 19380 -7720 19620 -7700
rect 19880 -7720 20120 -7700
rect 20380 -7720 20620 -7700
rect 20880 -7720 21120 -7700
rect 21380 -7720 21620 -7700
rect 21880 -7720 22120 -7700
rect 22380 -7720 22620 -7700
rect 22880 -7720 23120 -7700
rect 23380 -7720 23620 -7700
rect 23880 -7720 24000 -7700
rect 14500 -7980 14600 -7720
rect 14900 -7980 15100 -7720
rect 15400 -7980 15600 -7720
rect 15900 -7980 16100 -7720
rect 16400 -7980 16600 -7720
rect 16900 -7980 17100 -7720
rect 17400 -7980 17600 -7720
rect 17900 -7980 18100 -7720
rect 18400 -7980 18600 -7720
rect 18900 -7980 19100 -7720
rect 19400 -7980 19600 -7720
rect 19900 -7980 20100 -7720
rect 20400 -7980 20600 -7720
rect 20900 -7980 21100 -7720
rect 21400 -7980 21600 -7720
rect 21900 -7980 22100 -7720
rect 22400 -7980 22600 -7720
rect 22900 -7980 23100 -7720
rect 23400 -7980 23600 -7720
rect 23900 -7980 24000 -7720
rect 14500 -8000 14620 -7980
rect 14880 -8000 15120 -7980
rect 15380 -8000 15620 -7980
rect 15880 -8000 16120 -7980
rect 16380 -8000 16620 -7980
rect 16880 -8000 17120 -7980
rect 17380 -8000 17620 -7980
rect 17880 -8000 18120 -7980
rect 18380 -8000 18620 -7980
rect 18880 -8000 19120 -7980
rect 19380 -8000 19620 -7980
rect 19880 -8000 20120 -7980
rect 20380 -8000 20620 -7980
rect 20880 -8000 21120 -7980
rect 21380 -8000 21620 -7980
rect 21880 -8000 22120 -7980
rect 22380 -8000 22620 -7980
rect 22880 -8000 23120 -7980
rect 23380 -8000 23620 -7980
rect 23880 -8000 24000 -7980
rect 14500 -8200 24000 -8000
rect 14500 -8220 14620 -8200
rect 14880 -8220 15120 -8200
rect 15380 -8220 15620 -8200
rect 15880 -8220 16120 -8200
rect 16380 -8220 16620 -8200
rect 16880 -8220 17120 -8200
rect 17380 -8220 17620 -8200
rect 17880 -8220 18120 -8200
rect 18380 -8220 18620 -8200
rect 18880 -8220 19120 -8200
rect 19380 -8220 19620 -8200
rect 19880 -8220 20120 -8200
rect 20380 -8220 20620 -8200
rect 20880 -8220 21120 -8200
rect 21380 -8220 21620 -8200
rect 21880 -8220 22120 -8200
rect 22380 -8220 22620 -8200
rect 22880 -8220 23120 -8200
rect 23380 -8220 23620 -8200
rect 23880 -8220 24000 -8200
rect 14500 -8480 14600 -8220
rect 14900 -8480 15100 -8220
rect 15400 -8480 15600 -8220
rect 15900 -8480 16100 -8220
rect 16400 -8480 16600 -8220
rect 16900 -8480 17100 -8220
rect 17400 -8480 17600 -8220
rect 17900 -8480 18100 -8220
rect 18400 -8480 18600 -8220
rect 18900 -8480 19100 -8220
rect 19400 -8480 19600 -8220
rect 19900 -8480 20100 -8220
rect 20400 -8480 20600 -8220
rect 20900 -8480 21100 -8220
rect 21400 -8480 21600 -8220
rect 21900 -8480 22100 -8220
rect 22400 -8480 22600 -8220
rect 22900 -8480 23100 -8220
rect 23400 -8480 23600 -8220
rect 23900 -8480 24000 -8220
rect 14500 -8500 14620 -8480
rect 14880 -8500 15120 -8480
rect 15380 -8500 15620 -8480
rect 15880 -8500 16120 -8480
rect 16380 -8500 16620 -8480
rect 16880 -8500 17120 -8480
rect 17380 -8500 17620 -8480
rect 17880 -8500 18120 -8480
rect 18380 -8500 18620 -8480
rect 18880 -8500 19120 -8480
rect 19380 -8500 19620 -8480
rect 19880 -8500 20120 -8480
rect 20380 -8500 20620 -8480
rect 20880 -8500 21120 -8480
rect 21380 -8500 21620 -8480
rect 21880 -8500 22120 -8480
rect 22380 -8500 22620 -8480
rect 22880 -8500 23120 -8480
rect 23380 -8500 23620 -8480
rect 23880 -8500 24000 -8480
rect 14500 -8600 24000 -8500
rect 14500 -8700 17000 -8600
rect 14500 -8720 14620 -8700
rect 14880 -8720 15120 -8700
rect 15380 -8720 15620 -8700
rect 15880 -8720 16120 -8700
rect 16380 -8720 16620 -8700
rect 16880 -8720 17000 -8700
rect 14500 -8980 14600 -8720
rect 14900 -8980 15100 -8720
rect 15400 -8980 15600 -8720
rect 15900 -8980 16100 -8720
rect 16400 -8980 16600 -8720
rect 16900 -8980 17000 -8720
rect 14500 -9000 14620 -8980
rect 14880 -9000 15120 -8980
rect 15380 -9000 15620 -8980
rect 15880 -9000 16120 -8980
rect 16380 -9000 16620 -8980
rect 16880 -9000 17000 -8980
rect 14500 -9200 17000 -9000
rect 14500 -9220 14620 -9200
rect 14880 -9220 15120 -9200
rect 15380 -9220 15620 -9200
rect 15880 -9220 16120 -9200
rect 16380 -9220 16620 -9200
rect 16880 -9220 17000 -9200
rect 14500 -9480 14600 -9220
rect 14900 -9480 15100 -9220
rect 15400 -9480 15600 -9220
rect 15900 -9480 16100 -9220
rect 16400 -9480 16600 -9220
rect 16900 -9480 17000 -9220
rect 14500 -9500 14620 -9480
rect 14880 -9500 15120 -9480
rect 15380 -9500 15620 -9480
rect 15880 -9500 16120 -9480
rect 16380 -9500 16620 -9480
rect 16880 -9500 17000 -9480
rect 14500 -9700 17000 -9500
rect 14500 -9720 14620 -9700
rect 14880 -9720 15120 -9700
rect 15380 -9720 15620 -9700
rect 15880 -9720 16120 -9700
rect 16380 -9720 16620 -9700
rect 16880 -9720 17000 -9700
rect 14500 -9980 14600 -9720
rect 14900 -9980 15100 -9720
rect 15400 -9980 15600 -9720
rect 15900 -9980 16100 -9720
rect 16400 -9980 16600 -9720
rect 16900 -9980 17000 -9720
rect 14500 -10000 14620 -9980
rect 14880 -10000 15120 -9980
rect 15380 -10000 15620 -9980
rect 15880 -10000 16120 -9980
rect 16380 -10000 16620 -9980
rect 16880 -10000 17000 -9980
rect 14500 -10200 17000 -10000
rect 14500 -10220 14620 -10200
rect 14880 -10220 15120 -10200
rect 15380 -10220 15620 -10200
rect 15880 -10220 16120 -10200
rect 16380 -10220 16620 -10200
rect 16880 -10220 17000 -10200
rect 14500 -10480 14600 -10220
rect 14900 -10480 15100 -10220
rect 15400 -10480 15600 -10220
rect 15900 -10480 16100 -10220
rect 16400 -10480 16600 -10220
rect 16900 -10480 17000 -10220
rect 14500 -10500 14620 -10480
rect 14880 -10500 15120 -10480
rect 15380 -10500 15620 -10480
rect 15880 -10500 16120 -10480
rect 16380 -10500 16620 -10480
rect 16880 -10500 17000 -10480
rect 14500 -10700 17000 -10500
rect 14500 -10720 14620 -10700
rect 14880 -10720 15120 -10700
rect 15380 -10720 15620 -10700
rect 15880 -10720 16120 -10700
rect 16380 -10720 16620 -10700
rect 16880 -10720 17000 -10700
rect 14500 -10980 14600 -10720
rect 14900 -10980 15100 -10720
rect 15400 -10980 15600 -10720
rect 15900 -10980 16100 -10720
rect 16400 -10980 16600 -10720
rect 16900 -10980 17000 -10720
rect 14500 -11000 14620 -10980
rect 14880 -11000 15120 -10980
rect 15380 -11000 15620 -10980
rect 15880 -11000 16120 -10980
rect 16380 -11000 16620 -10980
rect 16880 -11000 17000 -10980
rect 14500 -11200 17000 -11000
rect 14500 -11220 14620 -11200
rect 14880 -11220 15120 -11200
rect 15380 -11220 15620 -11200
rect 15880 -11220 16120 -11200
rect 16380 -11220 16620 -11200
rect 16880 -11220 17000 -11200
rect 14500 -11480 14600 -11220
rect 14900 -11480 15100 -11220
rect 15400 -11480 15600 -11220
rect 15900 -11480 16100 -11220
rect 16400 -11480 16600 -11220
rect 16900 -11480 17000 -11220
rect 14500 -11500 14620 -11480
rect 14880 -11500 15120 -11480
rect 15380 -11500 15620 -11480
rect 15880 -11500 16120 -11480
rect 16380 -11500 16620 -11480
rect 16880 -11500 17000 -11480
rect 14500 -11700 17000 -11500
rect 14500 -11720 14620 -11700
rect 14880 -11720 15120 -11700
rect 15380 -11720 15620 -11700
rect 15880 -11720 16120 -11700
rect 16380 -11720 16620 -11700
rect 16880 -11720 17000 -11700
rect 14500 -11980 14600 -11720
rect 14900 -11980 15100 -11720
rect 15400 -11980 15600 -11720
rect 15900 -11980 16100 -11720
rect 16400 -11980 16600 -11720
rect 16900 -11980 17000 -11720
rect 14500 -12000 14620 -11980
rect 14880 -12000 15120 -11980
rect 15380 -12000 15620 -11980
rect 15880 -12000 16120 -11980
rect 16380 -12000 16620 -11980
rect 16880 -12000 17000 -11980
rect 14500 -12100 17000 -12000
rect 23500 -8700 24000 -8600
rect 23500 -8720 23620 -8700
rect 23880 -8720 24000 -8700
rect 23500 -8980 23600 -8720
rect 23900 -8980 24000 -8720
rect 23500 -9000 23620 -8980
rect 23880 -9000 24000 -8980
rect 23500 -9200 24000 -9000
rect 23500 -9220 23620 -9200
rect 23880 -9220 24000 -9200
rect 23500 -9480 23600 -9220
rect 23900 -9480 24000 -9220
rect 23500 -9500 23620 -9480
rect 23880 -9500 24000 -9480
rect 23500 -9700 24000 -9500
rect 23500 -9720 23620 -9700
rect 23880 -9720 24000 -9700
rect 23500 -9980 23600 -9720
rect 23900 -9980 24000 -9720
rect 23500 -10000 23620 -9980
rect 23880 -10000 24000 -9980
rect 23500 -10200 24000 -10000
rect 23500 -10220 23620 -10200
rect 23880 -10220 24000 -10200
rect 23500 -10480 23600 -10220
rect 23900 -10480 24000 -10220
rect 23500 -10500 23620 -10480
rect 23880 -10500 24000 -10480
rect 23500 -10700 24000 -10500
rect 23500 -10720 23620 -10700
rect 23880 -10720 24000 -10700
rect 23500 -10980 23600 -10720
rect 23900 -10980 24000 -10720
rect 23500 -11000 23620 -10980
rect 23880 -11000 24000 -10980
rect 23500 -11200 24000 -11000
rect 23500 -11220 23620 -11200
rect 23880 -11220 24000 -11200
rect 23500 -11480 23600 -11220
rect 23900 -11480 24000 -11220
rect 23500 -11500 23620 -11480
rect 23880 -11500 24000 -11480
rect 23500 -11700 24000 -11500
rect 23500 -11720 23620 -11700
rect 23880 -11720 24000 -11700
rect 23500 -11980 23600 -11720
rect 23900 -11980 24000 -11720
rect 23500 -12000 23620 -11980
rect 23880 -12000 24000 -11980
rect 14500 -12200 18500 -12100
rect 14500 -12220 14620 -12200
rect 14880 -12220 15120 -12200
rect 15380 -12220 15620 -12200
rect 15880 -12220 16120 -12200
rect 16380 -12220 16620 -12200
rect 16880 -12220 17120 -12200
rect 17380 -12220 17620 -12200
rect 17880 -12220 18120 -12200
rect 18380 -12220 18500 -12200
rect 14500 -12480 14600 -12220
rect 14900 -12480 15100 -12220
rect 15400 -12480 15600 -12220
rect 15900 -12480 16100 -12220
rect 16400 -12480 16600 -12220
rect 16900 -12480 17100 -12220
rect 17400 -12480 17600 -12220
rect 17900 -12480 18100 -12220
rect 18400 -12480 18500 -12220
rect 14500 -12500 14620 -12480
rect 14880 -12500 15120 -12480
rect 15380 -12500 15620 -12480
rect 15880 -12500 16120 -12480
rect 16380 -12500 16620 -12480
rect 16880 -12500 17120 -12480
rect 17380 -12500 17620 -12480
rect 17880 -12500 18120 -12480
rect 18380 -12500 18500 -12480
rect 14500 -12700 18500 -12500
rect 14500 -12720 14620 -12700
rect 14880 -12720 15120 -12700
rect 15380 -12720 15620 -12700
rect 15880 -12720 16120 -12700
rect 16380 -12720 16620 -12700
rect 16880 -12720 17120 -12700
rect 17380 -12720 17620 -12700
rect 17880 -12720 18120 -12700
rect 18380 -12720 18500 -12700
rect 14500 -12980 14600 -12720
rect 14900 -12980 15100 -12720
rect 15400 -12980 15600 -12720
rect 15900 -12980 16100 -12720
rect 16400 -12980 16600 -12720
rect 16900 -12980 17100 -12720
rect 17400 -12980 17600 -12720
rect 17900 -12980 18100 -12720
rect 18400 -12980 18500 -12720
rect 14500 -13000 14620 -12980
rect 14880 -13000 15120 -12980
rect 15380 -13000 15620 -12980
rect 15880 -13000 16120 -12980
rect 16380 -13000 16620 -12980
rect 16880 -13000 17120 -12980
rect 17380 -13000 17620 -12980
rect 17880 -13000 18120 -12980
rect 18380 -13000 18500 -12980
rect 14500 -13100 18500 -13000
rect -27500 -13220 -27380 -13200
rect -27120 -13220 -26880 -13200
rect -26620 -13220 -26380 -13200
rect -26120 -13220 -25880 -13200
rect -25620 -13220 -25380 -13200
rect -25120 -13220 -24880 -13200
rect -24620 -13220 -24380 -13200
rect -24120 -13220 -23880 -13200
rect -23620 -13220 -23380 -13200
rect -23120 -13220 -22880 -13200
rect -22620 -13220 -22380 -13200
rect -22120 -13220 -21880 -13200
rect -21620 -13220 -21380 -13200
rect -21120 -13220 -20880 -13200
rect -20620 -13220 -20380 -13200
rect -20120 -13220 -19880 -13200
rect -19620 -13220 -19380 -13200
rect -19120 -13220 -18880 -13200
rect -18620 -13220 -18380 -13200
rect -18120 -13220 -17880 -13200
rect -17620 -13220 -17380 -13200
rect -17120 -13220 -16880 -13200
rect -16620 -13220 -16380 -13200
rect -16120 -13220 -15880 -13200
rect -15620 -13220 -15380 -13200
rect -15120 -13220 -15000 -13200
rect -27500 -13480 -27400 -13220
rect -27100 -13480 -26900 -13220
rect -26600 -13480 -26400 -13220
rect -26100 -13480 -25900 -13220
rect -25600 -13480 -25400 -13220
rect -25100 -13480 -24900 -13220
rect -24600 -13480 -24400 -13220
rect -24100 -13480 -23900 -13220
rect -23600 -13480 -23400 -13220
rect -23100 -13480 -22900 -13220
rect -22600 -13480 -22400 -13220
rect -22100 -13480 -21900 -13220
rect -21600 -13480 -21400 -13220
rect -21100 -13480 -20900 -13220
rect -20600 -13480 -20400 -13220
rect -20100 -13480 -19900 -13220
rect -19600 -13480 -19400 -13220
rect -19100 -13480 -18900 -13220
rect -18600 -13480 -18400 -13220
rect -18100 -13480 -17900 -13220
rect -17600 -13480 -17400 -13220
rect -17100 -13480 -16900 -13220
rect -16600 -13480 -16400 -13220
rect -16100 -13480 -15900 -13220
rect -15600 -13480 -15400 -13220
rect -15100 -13480 -15000 -13220
rect -27500 -13500 -27380 -13480
rect -27120 -13500 -26880 -13480
rect -26620 -13500 -26380 -13480
rect -26120 -13500 -25880 -13480
rect -25620 -13500 -25380 -13480
rect -25120 -13500 -24880 -13480
rect -24620 -13500 -24380 -13480
rect -24120 -13500 -23880 -13480
rect -23620 -13500 -23380 -13480
rect -23120 -13500 -22880 -13480
rect -22620 -13500 -22380 -13480
rect -22120 -13500 -21880 -13480
rect -21620 -13500 -21380 -13480
rect -21120 -13500 -20880 -13480
rect -20620 -13500 -20380 -13480
rect -20120 -13500 -19880 -13480
rect -19620 -13500 -19380 -13480
rect -19120 -13500 -18880 -13480
rect -18620 -13500 -18380 -13480
rect -18120 -13500 -17880 -13480
rect -17620 -13500 -17380 -13480
rect -17120 -13500 -16880 -13480
rect -16620 -13500 -16380 -13480
rect -16120 -13500 -15880 -13480
rect -15620 -13500 -15380 -13480
rect -15120 -13500 -15000 -13480
rect -27500 -13600 -15000 -13500
rect -29500 -13700 -15000 -13600
rect -29500 -13720 -29380 -13700
rect -29120 -13720 -28880 -13700
rect -28620 -13720 -28380 -13700
rect -28120 -13720 -27880 -13700
rect -27620 -13720 -27380 -13700
rect -27120 -13720 -26880 -13700
rect -26620 -13720 -26380 -13700
rect -26120 -13720 -25880 -13700
rect -25620 -13720 -25380 -13700
rect -25120 -13720 -24880 -13700
rect -24620 -13720 -24380 -13700
rect -24120 -13720 -23880 -13700
rect -23620 -13720 -23380 -13700
rect -23120 -13720 -22880 -13700
rect -22620 -13720 -22380 -13700
rect -22120 -13720 -21880 -13700
rect -21620 -13720 -21380 -13700
rect -21120 -13720 -20880 -13700
rect -20620 -13720 -20380 -13700
rect -20120 -13720 -19880 -13700
rect -19620 -13720 -19380 -13700
rect -19120 -13720 -18880 -13700
rect -18620 -13720 -18380 -13700
rect -18120 -13720 -17880 -13700
rect -17620 -13720 -17380 -13700
rect -17120 -13720 -16880 -13700
rect -16620 -13720 -16380 -13700
rect -16120 -13720 -15880 -13700
rect -15620 -13720 -15380 -13700
rect -15120 -13720 -15000 -13700
rect -29500 -13980 -29400 -13720
rect -29100 -13980 -28900 -13720
rect -28600 -13980 -28400 -13720
rect -28100 -13980 -27900 -13720
rect -27600 -13980 -27400 -13720
rect -27100 -13980 -26900 -13720
rect -26600 -13980 -26400 -13720
rect -26100 -13980 -25900 -13720
rect -25600 -13980 -25400 -13720
rect -25100 -13980 -24900 -13720
rect -24600 -13980 -24400 -13720
rect -24100 -13980 -23900 -13720
rect -23600 -13980 -23400 -13720
rect -23100 -13980 -22900 -13720
rect -22600 -13980 -22400 -13720
rect -22100 -13980 -21900 -13720
rect -21600 -13980 -21400 -13720
rect -21100 -13980 -20900 -13720
rect -20600 -13980 -20400 -13720
rect -20100 -13980 -19900 -13720
rect -19600 -13980 -19400 -13720
rect -19100 -13980 -18900 -13720
rect -18600 -13980 -18400 -13720
rect -18100 -13980 -17900 -13720
rect -17600 -13980 -17400 -13720
rect -17100 -13980 -16900 -13720
rect -16600 -13980 -16400 -13720
rect -16100 -13980 -15900 -13720
rect -15600 -13980 -15400 -13720
rect -15100 -13980 -15000 -13720
rect -29500 -14000 -29380 -13980
rect -29120 -14000 -28880 -13980
rect -28620 -14000 -28380 -13980
rect -28120 -14000 -27880 -13980
rect -27620 -14000 -27380 -13980
rect -27120 -14000 -26880 -13980
rect -26620 -14000 -26380 -13980
rect -26120 -14000 -25880 -13980
rect -25620 -14000 -25380 -13980
rect -25120 -14000 -24880 -13980
rect -24620 -14000 -24380 -13980
rect -24120 -14000 -23880 -13980
rect -23620 -14000 -23380 -13980
rect -23120 -14000 -22880 -13980
rect -22620 -14000 -22380 -13980
rect -22120 -14000 -21880 -13980
rect -21620 -14000 -21380 -13980
rect -21120 -14000 -20880 -13980
rect -20620 -14000 -20380 -13980
rect -20120 -14000 -19880 -13980
rect -19620 -14000 -19380 -13980
rect -19120 -14000 -18880 -13980
rect -18620 -14000 -18380 -13980
rect -18120 -14000 -17880 -13980
rect -17620 -14000 -17380 -13980
rect -17120 -14000 -16880 -13980
rect -16620 -14000 -16380 -13980
rect -16120 -14000 -15880 -13980
rect -15620 -14000 -15380 -13980
rect -15120 -14000 -15000 -13980
rect -29500 -14200 -15000 -14000
rect -29500 -14220 -29380 -14200
rect -29120 -14220 -28880 -14200
rect -28620 -14220 -28380 -14200
rect -28120 -14220 -27880 -14200
rect -27620 -14220 -27380 -14200
rect -27120 -14220 -26880 -14200
rect -26620 -14220 -26380 -14200
rect -26120 -14220 -25880 -14200
rect -25620 -14220 -25380 -14200
rect -25120 -14220 -24880 -14200
rect -24620 -14220 -24380 -14200
rect -24120 -14220 -23880 -14200
rect -23620 -14220 -23380 -14200
rect -23120 -14220 -22880 -14200
rect -22620 -14220 -22380 -14200
rect -22120 -14220 -21880 -14200
rect -21620 -14220 -21380 -14200
rect -21120 -14220 -20880 -14200
rect -20620 -14220 -20380 -14200
rect -20120 -14220 -19880 -14200
rect -19620 -14220 -19380 -14200
rect -19120 -14220 -18880 -14200
rect -18620 -14220 -18380 -14200
rect -18120 -14220 -17880 -14200
rect -17620 -14220 -17380 -14200
rect -17120 -14220 -16880 -14200
rect -16620 -14220 -16380 -14200
rect -16120 -14220 -15880 -14200
rect -15620 -14220 -15380 -14200
rect -15120 -14220 -15000 -14200
rect -29500 -14480 -29400 -14220
rect -29100 -14480 -28900 -14220
rect -28600 -14480 -28400 -14220
rect -28100 -14480 -27900 -14220
rect -27600 -14480 -27400 -14220
rect -27100 -14480 -26900 -14220
rect -26600 -14480 -26400 -14220
rect -26100 -14480 -25900 -14220
rect -25600 -14480 -25400 -14220
rect -25100 -14480 -24900 -14220
rect -24600 -14480 -24400 -14220
rect -24100 -14480 -23900 -14220
rect -23600 -14480 -23400 -14220
rect -23100 -14480 -22900 -14220
rect -22600 -14480 -22400 -14220
rect -22100 -14480 -21900 -14220
rect -21600 -14480 -21400 -14220
rect -21100 -14480 -20900 -14220
rect -20600 -14480 -20400 -14220
rect -20100 -14480 -19900 -14220
rect -19600 -14480 -19400 -14220
rect -19100 -14480 -18900 -14220
rect -18600 -14480 -18400 -14220
rect -18100 -14480 -17900 -14220
rect -17600 -14480 -17400 -14220
rect -17100 -14480 -16900 -14220
rect -16600 -14480 -16400 -14220
rect -16100 -14480 -15900 -14220
rect -15600 -14480 -15400 -14220
rect -15100 -14480 -15000 -14220
rect -29500 -14500 -29380 -14480
rect -29120 -14500 -28880 -14480
rect -28620 -14500 -28380 -14480
rect -28120 -14500 -27880 -14480
rect -27620 -14500 -27380 -14480
rect -27120 -14500 -26880 -14480
rect -26620 -14500 -26380 -14480
rect -26120 -14500 -25880 -14480
rect -25620 -14500 -25380 -14480
rect -25120 -14500 -24880 -14480
rect -24620 -14500 -24380 -14480
rect -24120 -14500 -23880 -14480
rect -23620 -14500 -23380 -14480
rect -23120 -14500 -22880 -14480
rect -22620 -14500 -22380 -14480
rect -22120 -14500 -21880 -14480
rect -21620 -14500 -21380 -14480
rect -21120 -14500 -20880 -14480
rect -20620 -14500 -20380 -14480
rect -20120 -14500 -19880 -14480
rect -19620 -14500 -19380 -14480
rect -19120 -14500 -18880 -14480
rect -18620 -14500 -18380 -14480
rect -18120 -14500 -17880 -14480
rect -17620 -14500 -17380 -14480
rect -17120 -14500 -16880 -14480
rect -16620 -14500 -16380 -14480
rect -16120 -14500 -15880 -14480
rect -15620 -14500 -15380 -14480
rect -15120 -14500 -15000 -14480
rect -29500 -14700 -15000 -14500
rect -29500 -14720 -29380 -14700
rect -29120 -14720 -28880 -14700
rect -28620 -14720 -28380 -14700
rect -28120 -14720 -27880 -14700
rect -27620 -14720 -27380 -14700
rect -27120 -14720 -26880 -14700
rect -26620 -14720 -26380 -14700
rect -26120 -14720 -25880 -14700
rect -25620 -14720 -25380 -14700
rect -25120 -14720 -24880 -14700
rect -24620 -14720 -24380 -14700
rect -24120 -14720 -23880 -14700
rect -23620 -14720 -23380 -14700
rect -23120 -14720 -22880 -14700
rect -22620 -14720 -22380 -14700
rect -22120 -14720 -21880 -14700
rect -21620 -14720 -21380 -14700
rect -21120 -14720 -20880 -14700
rect -20620 -14720 -20380 -14700
rect -20120 -14720 -19880 -14700
rect -19620 -14720 -19380 -14700
rect -19120 -14720 -18880 -14700
rect -18620 -14720 -18380 -14700
rect -18120 -14720 -17880 -14700
rect -17620 -14720 -17380 -14700
rect -17120 -14720 -16880 -14700
rect -16620 -14720 -16380 -14700
rect -16120 -14720 -15880 -14700
rect -15620 -14720 -15380 -14700
rect -15120 -14720 -15000 -14700
rect -29500 -14980 -29400 -14720
rect -29100 -14980 -28900 -14720
rect -28600 -14980 -28400 -14720
rect -28100 -14980 -27900 -14720
rect -27600 -14980 -27400 -14720
rect -27100 -14980 -26900 -14720
rect -26600 -14980 -26400 -14720
rect -26100 -14980 -25900 -14720
rect -25600 -14980 -25400 -14720
rect -25100 -14980 -24900 -14720
rect -24600 -14980 -24400 -14720
rect -24100 -14980 -23900 -14720
rect -23600 -14980 -23400 -14720
rect -23100 -14980 -22900 -14720
rect -22600 -14980 -22400 -14720
rect -22100 -14980 -21900 -14720
rect -21600 -14980 -21400 -14720
rect -21100 -14980 -20900 -14720
rect -20600 -14980 -20400 -14720
rect -20100 -14980 -19900 -14720
rect -19600 -14980 -19400 -14720
rect -19100 -14980 -18900 -14720
rect -18600 -14980 -18400 -14720
rect -18100 -14980 -17900 -14720
rect -17600 -14980 -17400 -14720
rect -17100 -14980 -16900 -14720
rect -16600 -14980 -16400 -14720
rect -16100 -14980 -15900 -14720
rect -15600 -14980 -15400 -14720
rect -15100 -14980 -15000 -14720
rect -29500 -15000 -29380 -14980
rect -29120 -15000 -28880 -14980
rect -28620 -15000 -28380 -14980
rect -28120 -15000 -27880 -14980
rect -27620 -15000 -27380 -14980
rect -27120 -15000 -26880 -14980
rect -26620 -15000 -26380 -14980
rect -26120 -15000 -25880 -14980
rect -25620 -15000 -25380 -14980
rect -25120 -15000 -24880 -14980
rect -24620 -15000 -24380 -14980
rect -24120 -15000 -23880 -14980
rect -23620 -15000 -23380 -14980
rect -23120 -15000 -22880 -14980
rect -22620 -15000 -22380 -14980
rect -22120 -15000 -21880 -14980
rect -21620 -15000 -21380 -14980
rect -21120 -15000 -20880 -14980
rect -20620 -15000 -20380 -14980
rect -20120 -15000 -19880 -14980
rect -19620 -15000 -19380 -14980
rect -19120 -15000 -18880 -14980
rect -18620 -15000 -18380 -14980
rect -18120 -15000 -17880 -14980
rect -17620 -15000 -17380 -14980
rect -17120 -15000 -16880 -14980
rect -16620 -15000 -16380 -14980
rect -16120 -15000 -15880 -14980
rect -15620 -15000 -15380 -14980
rect -15120 -15000 -15000 -14980
rect -29500 -15200 -15000 -15000
rect -29500 -15220 -29380 -15200
rect -29120 -15220 -28880 -15200
rect -28620 -15220 -28380 -15200
rect -28120 -15220 -27880 -15200
rect -27620 -15220 -27380 -15200
rect -27120 -15220 -26880 -15200
rect -26620 -15220 -26380 -15200
rect -26120 -15220 -25880 -15200
rect -25620 -15220 -25380 -15200
rect -25120 -15220 -24880 -15200
rect -24620 -15220 -24380 -15200
rect -24120 -15220 -23880 -15200
rect -23620 -15220 -23380 -15200
rect -23120 -15220 -22880 -15200
rect -22620 -15220 -22380 -15200
rect -22120 -15220 -21880 -15200
rect -21620 -15220 -21380 -15200
rect -21120 -15220 -20880 -15200
rect -20620 -15220 -20380 -15200
rect -20120 -15220 -19880 -15200
rect -19620 -15220 -19380 -15200
rect -19120 -15220 -18880 -15200
rect -18620 -15220 -18380 -15200
rect -18120 -15220 -17880 -15200
rect -17620 -15220 -17380 -15200
rect -17120 -15220 -16880 -15200
rect -16620 -15220 -16380 -15200
rect -16120 -15220 -15880 -15200
rect -15620 -15220 -15380 -15200
rect -15120 -15220 -15000 -15200
rect -29500 -15480 -29400 -15220
rect -29100 -15480 -28900 -15220
rect -28600 -15480 -28400 -15220
rect -28100 -15480 -27900 -15220
rect -27600 -15480 -27400 -15220
rect -27100 -15480 -26900 -15220
rect -26600 -15480 -26400 -15220
rect -26100 -15480 -25900 -15220
rect -25600 -15480 -25400 -15220
rect -25100 -15480 -24900 -15220
rect -24600 -15480 -24400 -15220
rect -24100 -15480 -23900 -15220
rect -23600 -15480 -23400 -15220
rect -23100 -15480 -22900 -15220
rect -22600 -15480 -22400 -15220
rect -22100 -15480 -21900 -15220
rect -21600 -15480 -21400 -15220
rect -21100 -15480 -20900 -15220
rect -20600 -15480 -20400 -15220
rect -20100 -15480 -19900 -15220
rect -19600 -15480 -19400 -15220
rect -19100 -15480 -18900 -15220
rect -18600 -15480 -18400 -15220
rect -18100 -15480 -17900 -15220
rect -17600 -15480 -17400 -15220
rect -17100 -15480 -16900 -15220
rect -16600 -15480 -16400 -15220
rect -16100 -15480 -15900 -15220
rect -15600 -15480 -15400 -15220
rect -15100 -15480 -15000 -15220
rect -29500 -15500 -29380 -15480
rect -29120 -15500 -28880 -15480
rect -28620 -15500 -28380 -15480
rect -28120 -15500 -27880 -15480
rect -27620 -15500 -27380 -15480
rect -27120 -15500 -26880 -15480
rect -26620 -15500 -26380 -15480
rect -26120 -15500 -25880 -15480
rect -25620 -15500 -25380 -15480
rect -25120 -15500 -24880 -15480
rect -24620 -15500 -24380 -15480
rect -24120 -15500 -23880 -15480
rect -23620 -15500 -23380 -15480
rect -23120 -15500 -22880 -15480
rect -22620 -15500 -22380 -15480
rect -22120 -15500 -21880 -15480
rect -21620 -15500 -21380 -15480
rect -21120 -15500 -20880 -15480
rect -20620 -15500 -20380 -15480
rect -20120 -15500 -19880 -15480
rect -19620 -15500 -19380 -15480
rect -19120 -15500 -18880 -15480
rect -18620 -15500 -18380 -15480
rect -18120 -15500 -17880 -15480
rect -17620 -15500 -17380 -15480
rect -17120 -15500 -16880 -15480
rect -16620 -15500 -16380 -15480
rect -16120 -15500 -15880 -15480
rect -15620 -15500 -15380 -15480
rect -15120 -15500 -15000 -15480
rect -29500 -15700 -15000 -15500
rect -29500 -15720 -29380 -15700
rect -29120 -15720 -28880 -15700
rect -28620 -15720 -28380 -15700
rect -28120 -15720 -27880 -15700
rect -27620 -15720 -27380 -15700
rect -27120 -15720 -26880 -15700
rect -26620 -15720 -26380 -15700
rect -26120 -15720 -25880 -15700
rect -25620 -15720 -25380 -15700
rect -25120 -15720 -24880 -15700
rect -24620 -15720 -24380 -15700
rect -24120 -15720 -23880 -15700
rect -23620 -15720 -23380 -15700
rect -23120 -15720 -22880 -15700
rect -22620 -15720 -22380 -15700
rect -22120 -15720 -21880 -15700
rect -21620 -15720 -21380 -15700
rect -21120 -15720 -20880 -15700
rect -20620 -15720 -20380 -15700
rect -20120 -15720 -19880 -15700
rect -19620 -15720 -19380 -15700
rect -19120 -15720 -18880 -15700
rect -18620 -15720 -18380 -15700
rect -18120 -15720 -17880 -15700
rect -17620 -15720 -17380 -15700
rect -17120 -15720 -16880 -15700
rect -16620 -15720 -16380 -15700
rect -16120 -15720 -15880 -15700
rect -15620 -15720 -15380 -15700
rect -15120 -15720 -15000 -15700
rect -29500 -15980 -29400 -15720
rect -29100 -15980 -28900 -15720
rect -28600 -15980 -28400 -15720
rect -28100 -15980 -27900 -15720
rect -27600 -15980 -27400 -15720
rect -27100 -15980 -26900 -15720
rect -26600 -15980 -26400 -15720
rect -26100 -15980 -25900 -15720
rect -25600 -15980 -25400 -15720
rect -25100 -15980 -24900 -15720
rect -24600 -15980 -24400 -15720
rect -24100 -15980 -23900 -15720
rect -23600 -15980 -23400 -15720
rect -23100 -15980 -22900 -15720
rect -22600 -15980 -22400 -15720
rect -22100 -15980 -21900 -15720
rect -21600 -15980 -21400 -15720
rect -21100 -15980 -20900 -15720
rect -20600 -15980 -20400 -15720
rect -20100 -15980 -19900 -15720
rect -19600 -15980 -19400 -15720
rect -19100 -15980 -18900 -15720
rect -18600 -15980 -18400 -15720
rect -18100 -15980 -17900 -15720
rect -17600 -15980 -17400 -15720
rect -17100 -15980 -16900 -15720
rect -16600 -15980 -16400 -15720
rect -16100 -15980 -15900 -15720
rect -15600 -15980 -15400 -15720
rect -15100 -15980 -15000 -15720
rect -29500 -16000 -29380 -15980
rect -29120 -16000 -28880 -15980
rect -28620 -16000 -28380 -15980
rect -28120 -16000 -27880 -15980
rect -27620 -16000 -27380 -15980
rect -27120 -16000 -26880 -15980
rect -26620 -16000 -26380 -15980
rect -26120 -16000 -25880 -15980
rect -25620 -16000 -25380 -15980
rect -25120 -16000 -24880 -15980
rect -24620 -16000 -24380 -15980
rect -24120 -16000 -23880 -15980
rect -23620 -16000 -23380 -15980
rect -23120 -16000 -22880 -15980
rect -22620 -16000 -22380 -15980
rect -22120 -16000 -21880 -15980
rect -21620 -16000 -21380 -15980
rect -21120 -16000 -20880 -15980
rect -20620 -16000 -20380 -15980
rect -20120 -16000 -19880 -15980
rect -19620 -16000 -19380 -15980
rect -19120 -16000 -18880 -15980
rect -18620 -16000 -18380 -15980
rect -18120 -16000 -17880 -15980
rect -17620 -16000 -17380 -15980
rect -17120 -16000 -16880 -15980
rect -16620 -16000 -16380 -15980
rect -16120 -16000 -15880 -15980
rect -15620 -16000 -15380 -15980
rect -15120 -16000 -15000 -15980
rect -29500 -16100 -15000 -16000
rect -31500 -16200 -15000 -16100
rect -31500 -16220 -31380 -16200
rect -31120 -16220 -30880 -16200
rect -30620 -16220 -30380 -16200
rect -30120 -16220 -29880 -16200
rect -29620 -16220 -29380 -16200
rect -29120 -16220 -28880 -16200
rect -28620 -16220 -28380 -16200
rect -28120 -16220 -27880 -16200
rect -27620 -16220 -27380 -16200
rect -27120 -16220 -26880 -16200
rect -26620 -16220 -26380 -16200
rect -26120 -16220 -25880 -16200
rect -25620 -16220 -25380 -16200
rect -25120 -16220 -24880 -16200
rect -24620 -16220 -24380 -16200
rect -24120 -16220 -23880 -16200
rect -23620 -16220 -23380 -16200
rect -23120 -16220 -22880 -16200
rect -22620 -16220 -22380 -16200
rect -22120 -16220 -21880 -16200
rect -21620 -16220 -21380 -16200
rect -21120 -16220 -20880 -16200
rect -20620 -16220 -20380 -16200
rect -20120 -16220 -19880 -16200
rect -19620 -16220 -19380 -16200
rect -19120 -16220 -18880 -16200
rect -18620 -16220 -18380 -16200
rect -18120 -16220 -17880 -16200
rect -17620 -16220 -17380 -16200
rect -17120 -16220 -16880 -16200
rect -16620 -16220 -16380 -16200
rect -16120 -16220 -15880 -16200
rect -15620 -16220 -15380 -16200
rect -15120 -16220 -15000 -16200
rect -31500 -16480 -31400 -16220
rect -31100 -16480 -30900 -16220
rect -30600 -16480 -30400 -16220
rect -30100 -16480 -29900 -16220
rect -29600 -16480 -29400 -16220
rect -29100 -16480 -28900 -16220
rect -28600 -16480 -28400 -16220
rect -28100 -16480 -27900 -16220
rect -27600 -16480 -27400 -16220
rect -27100 -16480 -26900 -16220
rect -26600 -16480 -26400 -16220
rect -26100 -16480 -25900 -16220
rect -25600 -16480 -25400 -16220
rect -25100 -16480 -24900 -16220
rect -24600 -16480 -24400 -16220
rect -24100 -16480 -23900 -16220
rect -23600 -16480 -23400 -16220
rect -23100 -16480 -22900 -16220
rect -22600 -16480 -22400 -16220
rect -22100 -16480 -21900 -16220
rect -21600 -16480 -21400 -16220
rect -21100 -16480 -20900 -16220
rect -20600 -16480 -20400 -16220
rect -20100 -16480 -19900 -16220
rect -19600 -16480 -19400 -16220
rect -19100 -16480 -18900 -16220
rect -18600 -16480 -18400 -16220
rect -18100 -16480 -17900 -16220
rect -17600 -16480 -17400 -16220
rect -17100 -16480 -16900 -16220
rect -16600 -16480 -16400 -16220
rect -16100 -16480 -15900 -16220
rect -15600 -16480 -15400 -16220
rect -15100 -16480 -15000 -16220
rect -31500 -16500 -31380 -16480
rect -31120 -16500 -30880 -16480
rect -30620 -16500 -30380 -16480
rect -30120 -16500 -29880 -16480
rect -29620 -16500 -29380 -16480
rect -29120 -16500 -28880 -16480
rect -28620 -16500 -28380 -16480
rect -28120 -16500 -27880 -16480
rect -27620 -16500 -27380 -16480
rect -27120 -16500 -26880 -16480
rect -26620 -16500 -26380 -16480
rect -26120 -16500 -25880 -16480
rect -25620 -16500 -25380 -16480
rect -25120 -16500 -24880 -16480
rect -24620 -16500 -24380 -16480
rect -24120 -16500 -23880 -16480
rect -23620 -16500 -23380 -16480
rect -23120 -16500 -22880 -16480
rect -22620 -16500 -22380 -16480
rect -22120 -16500 -21880 -16480
rect -21620 -16500 -21380 -16480
rect -21120 -16500 -20880 -16480
rect -20620 -16500 -20380 -16480
rect -20120 -16500 -19880 -16480
rect -19620 -16500 -19380 -16480
rect -19120 -16500 -18880 -16480
rect -18620 -16500 -18380 -16480
rect -18120 -16500 -17880 -16480
rect -17620 -16500 -17380 -16480
rect -17120 -16500 -16880 -16480
rect -16620 -16500 -16380 -16480
rect -16120 -16500 -15880 -16480
rect -15620 -16500 -15380 -16480
rect -15120 -16500 -15000 -16480
rect -31500 -16700 -15000 -16500
rect -31500 -16720 -31380 -16700
rect -31120 -16720 -30880 -16700
rect -30620 -16720 -30380 -16700
rect -30120 -16720 -29880 -16700
rect -29620 -16720 -29380 -16700
rect -29120 -16720 -28880 -16700
rect -28620 -16720 -28380 -16700
rect -28120 -16720 -27880 -16700
rect -27620 -16720 -27380 -16700
rect -27120 -16720 -26880 -16700
rect -26620 -16720 -26380 -16700
rect -26120 -16720 -25880 -16700
rect -25620 -16720 -25380 -16700
rect -25120 -16720 -24880 -16700
rect -24620 -16720 -24380 -16700
rect -24120 -16720 -23880 -16700
rect -23620 -16720 -23380 -16700
rect -23120 -16720 -22880 -16700
rect -22620 -16720 -22380 -16700
rect -22120 -16720 -21880 -16700
rect -21620 -16720 -21380 -16700
rect -21120 -16720 -20880 -16700
rect -20620 -16720 -20380 -16700
rect -20120 -16720 -19880 -16700
rect -19620 -16720 -19380 -16700
rect -19120 -16720 -18880 -16700
rect -18620 -16720 -18380 -16700
rect -18120 -16720 -17880 -16700
rect -17620 -16720 -17380 -16700
rect -17120 -16720 -16880 -16700
rect -16620 -16720 -16380 -16700
rect -16120 -16720 -15880 -16700
rect -15620 -16720 -15380 -16700
rect -15120 -16720 -15000 -16700
rect -31500 -16980 -31400 -16720
rect -31100 -16980 -30900 -16720
rect -30600 -16980 -30400 -16720
rect -30100 -16980 -29900 -16720
rect -29600 -16980 -29400 -16720
rect -29100 -16980 -28900 -16720
rect -28600 -16980 -28400 -16720
rect -28100 -16980 -27900 -16720
rect -27600 -16980 -27400 -16720
rect -27100 -16980 -26900 -16720
rect -26600 -16980 -26400 -16720
rect -26100 -16980 -25900 -16720
rect -25600 -16980 -25400 -16720
rect -25100 -16980 -24900 -16720
rect -24600 -16980 -24400 -16720
rect -24100 -16980 -23900 -16720
rect -23600 -16980 -23400 -16720
rect -23100 -16980 -22900 -16720
rect -22600 -16980 -22400 -16720
rect -22100 -16980 -21900 -16720
rect -21600 -16980 -21400 -16720
rect -21100 -16980 -20900 -16720
rect -20600 -16980 -20400 -16720
rect -20100 -16980 -19900 -16720
rect -19600 -16980 -19400 -16720
rect -19100 -16980 -18900 -16720
rect -18600 -16980 -18400 -16720
rect -18100 -16980 -17900 -16720
rect -17600 -16980 -17400 -16720
rect -17100 -16980 -16900 -16720
rect -16600 -16980 -16400 -16720
rect -16100 -16980 -15900 -16720
rect -15600 -16980 -15400 -16720
rect -15100 -16980 -15000 -16720
rect -31500 -17000 -31380 -16980
rect -31120 -17000 -30880 -16980
rect -30620 -17000 -30380 -16980
rect -30120 -17000 -29880 -16980
rect -29620 -17000 -29380 -16980
rect -29120 -17000 -28880 -16980
rect -28620 -17000 -28380 -16980
rect -28120 -17000 -27880 -16980
rect -27620 -17000 -27380 -16980
rect -27120 -17000 -26880 -16980
rect -26620 -17000 -26380 -16980
rect -26120 -17000 -25880 -16980
rect -25620 -17000 -25380 -16980
rect -25120 -17000 -24880 -16980
rect -24620 -17000 -24380 -16980
rect -24120 -17000 -23880 -16980
rect -23620 -17000 -23380 -16980
rect -23120 -17000 -22880 -16980
rect -22620 -17000 -22380 -16980
rect -22120 -17000 -21880 -16980
rect -21620 -17000 -21380 -16980
rect -21120 -17000 -20880 -16980
rect -20620 -17000 -20380 -16980
rect -20120 -17000 -19880 -16980
rect -19620 -17000 -19380 -16980
rect -19120 -17000 -18880 -16980
rect -18620 -17000 -18380 -16980
rect -18120 -17000 -17880 -16980
rect -17620 -17000 -17380 -16980
rect -17120 -17000 -16880 -16980
rect -16620 -17000 -16380 -16980
rect -16120 -17000 -15880 -16980
rect -15620 -17000 -15380 -16980
rect -15120 -17000 -15000 -16980
rect -31500 -17200 -15000 -17000
rect -31500 -17220 -31380 -17200
rect -31120 -17220 -30880 -17200
rect -30620 -17220 -30380 -17200
rect -30120 -17220 -29880 -17200
rect -29620 -17220 -29380 -17200
rect -29120 -17220 -28880 -17200
rect -28620 -17220 -28380 -17200
rect -28120 -17220 -27880 -17200
rect -27620 -17220 -27380 -17200
rect -27120 -17220 -26880 -17200
rect -26620 -17220 -26380 -17200
rect -26120 -17220 -25880 -17200
rect -25620 -17220 -25380 -17200
rect -25120 -17220 -24880 -17200
rect -24620 -17220 -24380 -17200
rect -24120 -17220 -23880 -17200
rect -23620 -17220 -23380 -17200
rect -23120 -17220 -22880 -17200
rect -22620 -17220 -22380 -17200
rect -22120 -17220 -21880 -17200
rect -21620 -17220 -21380 -17200
rect -21120 -17220 -20880 -17200
rect -20620 -17220 -20380 -17200
rect -20120 -17220 -19880 -17200
rect -19620 -17220 -19380 -17200
rect -19120 -17220 -18880 -17200
rect -18620 -17220 -18380 -17200
rect -18120 -17220 -17880 -17200
rect -17620 -17220 -17380 -17200
rect -17120 -17220 -16880 -17200
rect -16620 -17220 -16380 -17200
rect -16120 -17220 -15880 -17200
rect -15620 -17220 -15380 -17200
rect -15120 -17220 -15000 -17200
rect -31500 -17480 -31400 -17220
rect -31100 -17480 -30900 -17220
rect -30600 -17480 -30400 -17220
rect -30100 -17480 -29900 -17220
rect -29600 -17480 -29400 -17220
rect -29100 -17480 -28900 -17220
rect -28600 -17480 -28400 -17220
rect -28100 -17480 -27900 -17220
rect -27600 -17480 -27400 -17220
rect -27100 -17480 -26900 -17220
rect -26600 -17480 -26400 -17220
rect -26100 -17480 -25900 -17220
rect -25600 -17480 -25400 -17220
rect -25100 -17480 -24900 -17220
rect -24600 -17480 -24400 -17220
rect -24100 -17480 -23900 -17220
rect -23600 -17480 -23400 -17220
rect -23100 -17480 -22900 -17220
rect -22600 -17480 -22400 -17220
rect -22100 -17480 -21900 -17220
rect -21600 -17480 -21400 -17220
rect -21100 -17480 -20900 -17220
rect -20600 -17480 -20400 -17220
rect -20100 -17480 -19900 -17220
rect -19600 -17480 -19400 -17220
rect -19100 -17480 -18900 -17220
rect -18600 -17480 -18400 -17220
rect -18100 -17480 -17900 -17220
rect -17600 -17480 -17400 -17220
rect -17100 -17480 -16900 -17220
rect -16600 -17480 -16400 -17220
rect -16100 -17480 -15900 -17220
rect -15600 -17480 -15400 -17220
rect -15100 -17480 -15000 -17220
rect -31500 -17500 -31380 -17480
rect -31120 -17500 -30880 -17480
rect -30620 -17500 -30380 -17480
rect -30120 -17500 -29880 -17480
rect -29620 -17500 -29380 -17480
rect -29120 -17500 -28880 -17480
rect -28620 -17500 -28380 -17480
rect -28120 -17500 -27880 -17480
rect -27620 -17500 -27380 -17480
rect -27120 -17500 -26880 -17480
rect -26620 -17500 -26380 -17480
rect -26120 -17500 -25880 -17480
rect -25620 -17500 -25380 -17480
rect -25120 -17500 -24880 -17480
rect -24620 -17500 -24380 -17480
rect -24120 -17500 -23880 -17480
rect -23620 -17500 -23380 -17480
rect -23120 -17500 -22880 -17480
rect -22620 -17500 -22380 -17480
rect -22120 -17500 -21880 -17480
rect -21620 -17500 -21380 -17480
rect -21120 -17500 -20880 -17480
rect -20620 -17500 -20380 -17480
rect -20120 -17500 -19880 -17480
rect -19620 -17500 -19380 -17480
rect -19120 -17500 -18880 -17480
rect -18620 -17500 -18380 -17480
rect -18120 -17500 -17880 -17480
rect -17620 -17500 -17380 -17480
rect -17120 -17500 -16880 -17480
rect -16620 -17500 -16380 -17480
rect -16120 -17500 -15880 -17480
rect -15620 -17500 -15380 -17480
rect -15120 -17500 -15000 -17480
rect -31500 -17600 -15000 -17500
rect -31500 -17700 -27500 -17600
rect -31500 -17720 -31380 -17700
rect -31120 -17720 -30880 -17700
rect -30620 -17720 -30380 -17700
rect -30120 -17720 -29880 -17700
rect -29620 -17720 -29380 -17700
rect -29120 -17720 -28880 -17700
rect -28620 -17720 -28380 -17700
rect -28120 -17720 -27880 -17700
rect -27620 -17720 -27500 -17700
rect -31500 -17980 -31400 -17720
rect -31100 -17980 -30900 -17720
rect -30600 -17980 -30400 -17720
rect -30100 -17980 -29900 -17720
rect -29600 -17980 -29400 -17720
rect -29100 -17980 -28900 -17720
rect -28600 -17980 -28400 -17720
rect -28100 -17980 -27900 -17720
rect -27600 -17980 -27500 -17720
rect -31500 -18000 -31380 -17980
rect -31120 -18000 -30880 -17980
rect -30620 -18000 -30380 -17980
rect -30120 -18000 -29880 -17980
rect -29620 -18000 -29380 -17980
rect -29120 -18000 -28880 -17980
rect -28620 -18000 -28380 -17980
rect -28120 -18000 -27880 -17980
rect -27620 -18000 -27500 -17980
rect -31500 -18100 -27500 -18000
rect -26500 -17700 -15000 -17600
rect -26500 -17720 -26380 -17700
rect -26120 -17720 -25880 -17700
rect -25620 -17720 -25380 -17700
rect -25120 -17720 -24880 -17700
rect -24620 -17720 -24380 -17700
rect -24120 -17720 -23880 -17700
rect -23620 -17720 -23380 -17700
rect -23120 -17720 -22880 -17700
rect -22620 -17720 -22380 -17700
rect -22120 -17720 -21880 -17700
rect -21620 -17720 -21380 -17700
rect -21120 -17720 -20880 -17700
rect -20620 -17720 -20380 -17700
rect -20120 -17720 -19880 -17700
rect -19620 -17720 -19380 -17700
rect -19120 -17720 -18880 -17700
rect -18620 -17720 -18380 -17700
rect -18120 -17720 -17880 -17700
rect -17620 -17720 -17380 -17700
rect -17120 -17720 -16880 -17700
rect -16620 -17720 -16380 -17700
rect -16120 -17720 -15880 -17700
rect -15620 -17720 -15380 -17700
rect -15120 -17720 -15000 -17700
rect -26500 -17980 -26400 -17720
rect -26100 -17980 -25900 -17720
rect -25600 -17980 -25400 -17720
rect -25100 -17980 -24900 -17720
rect -24600 -17980 -24400 -17720
rect -24100 -17980 -23900 -17720
rect -23600 -17980 -23400 -17720
rect -23100 -17980 -22900 -17720
rect -22600 -17980 -22400 -17720
rect -22100 -17980 -21900 -17720
rect -21600 -17980 -21400 -17720
rect -21100 -17980 -20900 -17720
rect -20600 -17980 -20400 -17720
rect -20100 -17980 -19900 -17720
rect -19600 -17980 -19400 -17720
rect -19100 -17980 -18900 -17720
rect -18600 -17980 -18400 -17720
rect -18100 -17980 -17900 -17720
rect -17600 -17980 -17400 -17720
rect -17100 -17980 -16900 -17720
rect -16600 -17980 -16400 -17720
rect -16100 -17980 -15900 -17720
rect -15600 -17980 -15400 -17720
rect -15100 -17980 -15000 -17720
rect -26500 -18000 -26380 -17980
rect -26120 -18000 -25880 -17980
rect -25620 -18000 -25380 -17980
rect -25120 -18000 -24880 -17980
rect -24620 -18000 -24380 -17980
rect -24120 -18000 -23880 -17980
rect -23620 -18000 -23380 -17980
rect -23120 -18000 -22880 -17980
rect -22620 -18000 -22380 -17980
rect -22120 -18000 -21880 -17980
rect -21620 -18000 -21380 -17980
rect -21120 -18000 -20880 -17980
rect -20620 -18000 -20380 -17980
rect -20120 -18000 -19880 -17980
rect -19620 -18000 -19380 -17980
rect -19120 -18000 -18880 -17980
rect -18620 -18000 -18380 -17980
rect -18120 -18000 -17880 -17980
rect -17620 -18000 -17380 -17980
rect -17120 -18000 -16880 -17980
rect -16620 -18000 -16380 -17980
rect -16120 -18000 -15880 -17980
rect -15620 -18000 -15380 -17980
rect -15120 -18000 -15000 -17980
rect -31500 -18200 -29500 -18100
rect -31500 -18220 -31380 -18200
rect -31120 -18220 -30880 -18200
rect -30620 -18220 -30380 -18200
rect -30120 -18220 -29880 -18200
rect -29620 -18220 -29500 -18200
rect -31500 -18480 -31400 -18220
rect -31100 -18480 -30900 -18220
rect -30600 -18480 -30400 -18220
rect -30100 -18480 -29900 -18220
rect -29600 -18480 -29500 -18220
rect -31500 -18500 -31380 -18480
rect -31120 -18500 -30880 -18480
rect -30620 -18500 -30380 -18480
rect -30120 -18500 -29880 -18480
rect -29620 -18500 -29500 -18480
rect -31500 -18700 -29500 -18500
rect -31500 -18720 -31380 -18700
rect -31120 -18720 -30880 -18700
rect -30620 -18720 -30380 -18700
rect -30120 -18720 -29880 -18700
rect -29620 -18720 -29500 -18700
rect -31500 -18980 -31400 -18720
rect -31100 -18980 -30900 -18720
rect -30600 -18980 -30400 -18720
rect -30100 -18980 -29900 -18720
rect -29600 -18980 -29500 -18720
rect -31500 -19000 -31380 -18980
rect -31120 -19000 -30880 -18980
rect -30620 -19000 -30380 -18980
rect -30120 -19000 -29880 -18980
rect -29620 -19000 -29500 -18980
rect -31500 -19200 -29500 -19000
rect -31500 -19220 -31380 -19200
rect -31120 -19220 -30880 -19200
rect -30620 -19220 -30380 -19200
rect -30120 -19220 -29880 -19200
rect -29620 -19220 -29500 -19200
rect -31500 -19480 -31400 -19220
rect -31100 -19480 -30900 -19220
rect -30600 -19480 -30400 -19220
rect -30100 -19480 -29900 -19220
rect -29600 -19480 -29500 -19220
rect -31500 -19500 -31380 -19480
rect -31120 -19500 -30880 -19480
rect -30620 -19500 -30380 -19480
rect -30120 -19500 -29880 -19480
rect -29620 -19500 -29500 -19480
rect -31500 -19700 -29500 -19500
rect -31500 -19720 -31380 -19700
rect -31120 -19720 -30880 -19700
rect -30620 -19720 -30380 -19700
rect -30120 -19720 -29880 -19700
rect -29620 -19720 -29500 -19700
rect -31500 -19980 -31400 -19720
rect -31100 -19980 -30900 -19720
rect -30600 -19980 -30400 -19720
rect -30100 -19980 -29900 -19720
rect -29600 -19980 -29500 -19720
rect -31500 -20000 -31380 -19980
rect -31120 -20000 -30880 -19980
rect -30620 -20000 -30380 -19980
rect -30120 -20000 -29880 -19980
rect -29620 -20000 -29500 -19980
rect -31500 -20200 -29500 -20000
rect -31500 -20220 -31380 -20200
rect -31120 -20220 -30880 -20200
rect -30620 -20220 -30380 -20200
rect -30120 -20220 -29880 -20200
rect -29620 -20220 -29500 -20200
rect -31500 -20480 -31400 -20220
rect -31100 -20480 -30900 -20220
rect -30600 -20480 -30400 -20220
rect -30100 -20480 -29900 -20220
rect -29600 -20480 -29500 -20220
rect -31500 -20500 -31380 -20480
rect -31120 -20500 -30880 -20480
rect -30620 -20500 -30380 -20480
rect -30120 -20500 -29880 -20480
rect -29620 -20500 -29500 -20480
rect -31500 -20700 -29500 -20500
rect -31500 -20720 -31380 -20700
rect -31120 -20720 -30880 -20700
rect -30620 -20720 -30380 -20700
rect -30120 -20720 -29880 -20700
rect -29620 -20720 -29500 -20700
rect -31500 -20980 -31400 -20720
rect -31100 -20980 -30900 -20720
rect -30600 -20980 -30400 -20720
rect -30100 -20980 -29900 -20720
rect -29600 -20980 -29500 -20720
rect -31500 -21000 -31380 -20980
rect -31120 -21000 -30880 -20980
rect -30620 -21000 -30380 -20980
rect -30120 -21000 -29880 -20980
rect -29620 -21000 -29500 -20980
rect -31500 -21200 -29500 -21000
rect -31500 -21220 -31380 -21200
rect -31120 -21220 -30880 -21200
rect -30620 -21220 -30380 -21200
rect -30120 -21220 -29880 -21200
rect -29620 -21220 -29500 -21200
rect -31500 -21480 -31400 -21220
rect -31100 -21480 -30900 -21220
rect -30600 -21480 -30400 -21220
rect -30100 -21480 -29900 -21220
rect -29600 -21480 -29500 -21220
rect -31500 -21500 -31380 -21480
rect -31120 -21500 -30880 -21480
rect -30620 -21500 -30380 -21480
rect -30120 -21500 -29880 -21480
rect -29620 -21500 -29500 -21480
rect -31500 -21700 -29500 -21500
rect -31500 -21720 -31380 -21700
rect -31120 -21720 -30880 -21700
rect -30620 -21720 -30380 -21700
rect -30120 -21720 -29880 -21700
rect -29620 -21720 -29500 -21700
rect -31500 -21980 -31400 -21720
rect -31100 -21980 -30900 -21720
rect -30600 -21980 -30400 -21720
rect -30100 -21980 -29900 -21720
rect -29600 -21980 -29500 -21720
rect -31500 -22000 -31380 -21980
rect -31120 -22000 -30880 -21980
rect -30620 -22000 -30380 -21980
rect -30120 -22000 -29880 -21980
rect -29620 -22000 -29500 -21980
rect -31500 -22200 -29500 -22000
rect -31500 -22220 -31380 -22200
rect -31120 -22220 -30880 -22200
rect -30620 -22220 -30380 -22200
rect -30120 -22220 -29880 -22200
rect -29620 -22220 -29500 -22200
rect -31500 -22480 -31400 -22220
rect -31100 -22480 -30900 -22220
rect -30600 -22480 -30400 -22220
rect -30100 -22480 -29900 -22220
rect -29600 -22480 -29500 -22220
rect -31500 -22500 -31380 -22480
rect -31120 -22500 -30880 -22480
rect -30620 -22500 -30380 -22480
rect -30120 -22500 -29880 -22480
rect -29620 -22500 -29500 -22480
rect -31500 -22700 -29500 -22500
rect -31500 -22720 -31380 -22700
rect -31120 -22720 -30880 -22700
rect -30620 -22720 -30380 -22700
rect -30120 -22720 -29880 -22700
rect -29620 -22720 -29500 -22700
rect -31500 -22980 -31400 -22720
rect -31100 -22980 -30900 -22720
rect -30600 -22980 -30400 -22720
rect -30100 -22980 -29900 -22720
rect -29600 -22980 -29500 -22720
rect -31500 -23000 -31380 -22980
rect -31120 -23000 -30880 -22980
rect -30620 -23000 -30380 -22980
rect -30120 -23000 -29880 -22980
rect -29620 -23000 -29500 -22980
rect -31500 -23200 -29500 -23000
rect -31500 -23220 -31380 -23200
rect -31120 -23220 -30880 -23200
rect -30620 -23220 -30380 -23200
rect -30120 -23220 -29880 -23200
rect -29620 -23220 -29500 -23200
rect -31500 -23480 -31400 -23220
rect -31100 -23480 -30900 -23220
rect -30600 -23480 -30400 -23220
rect -30100 -23480 -29900 -23220
rect -29600 -23480 -29500 -23220
rect -31500 -23500 -31380 -23480
rect -31120 -23500 -30880 -23480
rect -30620 -23500 -30380 -23480
rect -30120 -23500 -29880 -23480
rect -29620 -23500 -29500 -23480
rect -31500 -23700 -29500 -23500
rect -31500 -23720 -31380 -23700
rect -31120 -23720 -30880 -23700
rect -30620 -23720 -30380 -23700
rect -30120 -23720 -29880 -23700
rect -29620 -23720 -29500 -23700
rect -31500 -23980 -31400 -23720
rect -31100 -23980 -30900 -23720
rect -30600 -23980 -30400 -23720
rect -30100 -23980 -29900 -23720
rect -29600 -23980 -29500 -23720
rect -31500 -24000 -31380 -23980
rect -31120 -24000 -30880 -23980
rect -30620 -24000 -30380 -23980
rect -30120 -24000 -29880 -23980
rect -29620 -24000 -29500 -23980
rect -31500 -24200 -29500 -24000
rect -31500 -24220 -31380 -24200
rect -31120 -24220 -30880 -24200
rect -30620 -24220 -30380 -24200
rect -30120 -24220 -29880 -24200
rect -29620 -24220 -29500 -24200
rect -31500 -24480 -31400 -24220
rect -31100 -24480 -30900 -24220
rect -30600 -24480 -30400 -24220
rect -30100 -24480 -29900 -24220
rect -29600 -24480 -29500 -24220
rect -31500 -24500 -31380 -24480
rect -31120 -24500 -30880 -24480
rect -30620 -24500 -30380 -24480
rect -30120 -24500 -29880 -24480
rect -29620 -24500 -29500 -24480
rect -31500 -24700 -29500 -24500
rect -31500 -24720 -31380 -24700
rect -31120 -24720 -30880 -24700
rect -30620 -24720 -30380 -24700
rect -30120 -24720 -29880 -24700
rect -29620 -24720 -29500 -24700
rect -31500 -24980 -31400 -24720
rect -31100 -24980 -30900 -24720
rect -30600 -24980 -30400 -24720
rect -30100 -24980 -29900 -24720
rect -29600 -24980 -29500 -24720
rect -31500 -25000 -31380 -24980
rect -31120 -25000 -30880 -24980
rect -30620 -25000 -30380 -24980
rect -30120 -25000 -29880 -24980
rect -29620 -25000 -29500 -24980
rect -31500 -25200 -29500 -25000
rect -31500 -25220 -31380 -25200
rect -31120 -25220 -30880 -25200
rect -30620 -25220 -30380 -25200
rect -30120 -25220 -29880 -25200
rect -29620 -25220 -29500 -25200
rect -31500 -25480 -31400 -25220
rect -31100 -25480 -30900 -25220
rect -30600 -25480 -30400 -25220
rect -30100 -25480 -29900 -25220
rect -29600 -25480 -29500 -25220
rect -31500 -25500 -31380 -25480
rect -31120 -25500 -30880 -25480
rect -30620 -25500 -30380 -25480
rect -30120 -25500 -29880 -25480
rect -29620 -25500 -29500 -25480
rect -31500 -25700 -29500 -25500
rect -31500 -25720 -31380 -25700
rect -31120 -25720 -30880 -25700
rect -30620 -25720 -30380 -25700
rect -30120 -25720 -29880 -25700
rect -29620 -25720 -29500 -25700
rect -31500 -25980 -31400 -25720
rect -31100 -25980 -30900 -25720
rect -30600 -25980 -30400 -25720
rect -30100 -25980 -29900 -25720
rect -29600 -25980 -29500 -25720
rect -31500 -26000 -31380 -25980
rect -31120 -26000 -30880 -25980
rect -30620 -26000 -30380 -25980
rect -30120 -26000 -29880 -25980
rect -29620 -26000 -29500 -25980
rect -31500 -26200 -29500 -26000
rect -31500 -26220 -31380 -26200
rect -31120 -26220 -30880 -26200
rect -30620 -26220 -30380 -26200
rect -30120 -26220 -29880 -26200
rect -29620 -26220 -29500 -26200
rect -31500 -26480 -31400 -26220
rect -31100 -26480 -30900 -26220
rect -30600 -26480 -30400 -26220
rect -30100 -26480 -29900 -26220
rect -29600 -26480 -29500 -26220
rect -31500 -26500 -31380 -26480
rect -31120 -26500 -30880 -26480
rect -30620 -26500 -30380 -26480
rect -30120 -26500 -29880 -26480
rect -29620 -26500 -29500 -26480
rect -31500 -26700 -29500 -26500
rect -31500 -26720 -31380 -26700
rect -31120 -26720 -30880 -26700
rect -30620 -26720 -30380 -26700
rect -30120 -26720 -29880 -26700
rect -29620 -26720 -29500 -26700
rect -31500 -26980 -31400 -26720
rect -31100 -26980 -30900 -26720
rect -30600 -26980 -30400 -26720
rect -30100 -26980 -29900 -26720
rect -29600 -26980 -29500 -26720
rect -31500 -27000 -31380 -26980
rect -31120 -27000 -30880 -26980
rect -30620 -27000 -30380 -26980
rect -30120 -27000 -29880 -26980
rect -29620 -27000 -29500 -26980
rect -31500 -27200 -29500 -27000
rect -31500 -27220 -31380 -27200
rect -31120 -27220 -30880 -27200
rect -30620 -27220 -30380 -27200
rect -30120 -27220 -29880 -27200
rect -29620 -27220 -29500 -27200
rect -31500 -27480 -31400 -27220
rect -31100 -27480 -30900 -27220
rect -30600 -27480 -30400 -27220
rect -30100 -27480 -29900 -27220
rect -29600 -27480 -29500 -27220
rect -31500 -27500 -31380 -27480
rect -31120 -27500 -30880 -27480
rect -30620 -27500 -30380 -27480
rect -30120 -27500 -29880 -27480
rect -29620 -27500 -29500 -27480
rect -31500 -27700 -29500 -27500
rect -31500 -27720 -31380 -27700
rect -31120 -27720 -30880 -27700
rect -30620 -27720 -30380 -27700
rect -30120 -27720 -29880 -27700
rect -29620 -27720 -29500 -27700
rect -31500 -27980 -31400 -27720
rect -31100 -27980 -30900 -27720
rect -30600 -27980 -30400 -27720
rect -30100 -27980 -29900 -27720
rect -29600 -27980 -29500 -27720
rect -31500 -28000 -31380 -27980
rect -31120 -28000 -30880 -27980
rect -30620 -28000 -30380 -27980
rect -30120 -28000 -29880 -27980
rect -29620 -28000 -29500 -27980
rect -31500 -28200 -29500 -28000
rect -31500 -28220 -31380 -28200
rect -31120 -28220 -30880 -28200
rect -30620 -28220 -30380 -28200
rect -30120 -28220 -29880 -28200
rect -29620 -28220 -29500 -28200
rect -31500 -28480 -31400 -28220
rect -31100 -28480 -30900 -28220
rect -30600 -28480 -30400 -28220
rect -30100 -28480 -29900 -28220
rect -29600 -28480 -29500 -28220
rect -31500 -28500 -31380 -28480
rect -31120 -28500 -30880 -28480
rect -30620 -28500 -30380 -28480
rect -30120 -28500 -29880 -28480
rect -29620 -28500 -29500 -28480
rect -31500 -28700 -29500 -28500
rect -31500 -28720 -31380 -28700
rect -31120 -28720 -30880 -28700
rect -30620 -28720 -30380 -28700
rect -30120 -28720 -29880 -28700
rect -29620 -28720 -29500 -28700
rect -31500 -28980 -31400 -28720
rect -31100 -28980 -30900 -28720
rect -30600 -28980 -30400 -28720
rect -30100 -28980 -29900 -28720
rect -29600 -28980 -29500 -28720
rect -31500 -29000 -31380 -28980
rect -31120 -29000 -30880 -28980
rect -30620 -29000 -30380 -28980
rect -30120 -29000 -29880 -28980
rect -29620 -29000 -29500 -28980
rect -31500 -29200 -29500 -29000
rect -31500 -29220 -31380 -29200
rect -31120 -29220 -30880 -29200
rect -30620 -29220 -30380 -29200
rect -30120 -29220 -29880 -29200
rect -29620 -29220 -29500 -29200
rect -31500 -29480 -31400 -29220
rect -31100 -29480 -30900 -29220
rect -30600 -29480 -30400 -29220
rect -30100 -29480 -29900 -29220
rect -29600 -29480 -29500 -29220
rect -31500 -29500 -31380 -29480
rect -31120 -29500 -30880 -29480
rect -30620 -29500 -30380 -29480
rect -30120 -29500 -29880 -29480
rect -29620 -29500 -29500 -29480
rect -31500 -29600 -29500 -29500
rect -26500 -18200 -15000 -18000
rect -26500 -18220 -26380 -18200
rect -26120 -18220 -25880 -18200
rect -25620 -18220 -25380 -18200
rect -25120 -18220 -24880 -18200
rect -24620 -18220 -24380 -18200
rect -24120 -18220 -23880 -18200
rect -23620 -18220 -23380 -18200
rect -23120 -18220 -22880 -18200
rect -22620 -18220 -22380 -18200
rect -22120 -18220 -21880 -18200
rect -21620 -18220 -21380 -18200
rect -21120 -18220 -20880 -18200
rect -20620 -18220 -20380 -18200
rect -20120 -18220 -19880 -18200
rect -19620 -18220 -19380 -18200
rect -19120 -18220 -18880 -18200
rect -18620 -18220 -18380 -18200
rect -18120 -18220 -17880 -18200
rect -17620 -18220 -17380 -18200
rect -17120 -18220 -16880 -18200
rect -16620 -18220 -16380 -18200
rect -16120 -18220 -15880 -18200
rect -15620 -18220 -15380 -18200
rect -15120 -18220 -15000 -18200
rect -26500 -18480 -26400 -18220
rect -26100 -18480 -25900 -18220
rect -25600 -18480 -25400 -18220
rect -25100 -18480 -24900 -18220
rect -24600 -18480 -24400 -18220
rect -24100 -18480 -23900 -18220
rect -23600 -18480 -23400 -18220
rect -23100 -18480 -22900 -18220
rect -22600 -18480 -22400 -18220
rect -22100 -18480 -21900 -18220
rect -21600 -18480 -21400 -18220
rect -21100 -18480 -20900 -18220
rect -20600 -18480 -20400 -18220
rect -20100 -18480 -19900 -18220
rect -19600 -18480 -19400 -18220
rect -19100 -18480 -18900 -18220
rect -18600 -18480 -18400 -18220
rect -18100 -18480 -17900 -18220
rect -17600 -18480 -17400 -18220
rect -17100 -18480 -16900 -18220
rect -16600 -18480 -16400 -18220
rect -16100 -18480 -15900 -18220
rect -15600 -18480 -15400 -18220
rect -15100 -18480 -15000 -18220
rect -26500 -18500 -26380 -18480
rect -26120 -18500 -25880 -18480
rect -25620 -18500 -25380 -18480
rect -25120 -18500 -24880 -18480
rect -24620 -18500 -24380 -18480
rect -24120 -18500 -23880 -18480
rect -23620 -18500 -23380 -18480
rect -23120 -18500 -22880 -18480
rect -22620 -18500 -22380 -18480
rect -22120 -18500 -21880 -18480
rect -21620 -18500 -21380 -18480
rect -21120 -18500 -20880 -18480
rect -20620 -18500 -20380 -18480
rect -20120 -18500 -19880 -18480
rect -19620 -18500 -19380 -18480
rect -19120 -18500 -18880 -18480
rect -18620 -18500 -18380 -18480
rect -18120 -18500 -17880 -18480
rect -17620 -18500 -17380 -18480
rect -17120 -18500 -16880 -18480
rect -16620 -18500 -16380 -18480
rect -16120 -18500 -15880 -18480
rect -15620 -18500 -15380 -18480
rect -15120 -18500 -15000 -18480
rect -26500 -18700 -15000 -18500
rect -26500 -18720 -26380 -18700
rect -26120 -18720 -25880 -18700
rect -25620 -18720 -25380 -18700
rect -25120 -18720 -24880 -18700
rect -24620 -18720 -24380 -18700
rect -24120 -18720 -23880 -18700
rect -23620 -18720 -23380 -18700
rect -23120 -18720 -22880 -18700
rect -22620 -18720 -22380 -18700
rect -22120 -18720 -21880 -18700
rect -21620 -18720 -21380 -18700
rect -21120 -18720 -20880 -18700
rect -20620 -18720 -20380 -18700
rect -20120 -18720 -19880 -18700
rect -19620 -18720 -19380 -18700
rect -19120 -18720 -18880 -18700
rect -18620 -18720 -18380 -18700
rect -18120 -18720 -17880 -18700
rect -17620 -18720 -17380 -18700
rect -17120 -18720 -16880 -18700
rect -16620 -18720 -16380 -18700
rect -16120 -18720 -15880 -18700
rect -15620 -18720 -15380 -18700
rect -15120 -18720 -15000 -18700
rect -26500 -18980 -26400 -18720
rect -26100 -18980 -25900 -18720
rect -25600 -18980 -25400 -18720
rect -25100 -18980 -24900 -18720
rect -24600 -18980 -24400 -18720
rect -24100 -18980 -23900 -18720
rect -23600 -18980 -23400 -18720
rect -23100 -18980 -22900 -18720
rect -22600 -18980 -22400 -18720
rect -22100 -18980 -21900 -18720
rect -21600 -18980 -21400 -18720
rect -21100 -18980 -20900 -18720
rect -20600 -18980 -20400 -18720
rect -20100 -18980 -19900 -18720
rect -19600 -18980 -19400 -18720
rect -19100 -18980 -18900 -18720
rect -18600 -18980 -18400 -18720
rect -18100 -18980 -17900 -18720
rect -17600 -18980 -17400 -18720
rect -17100 -18980 -16900 -18720
rect -16600 -18980 -16400 -18720
rect -16100 -18980 -15900 -18720
rect -15600 -18980 -15400 -18720
rect -15100 -18980 -15000 -18720
rect -26500 -19000 -26380 -18980
rect -26120 -19000 -25880 -18980
rect -25620 -19000 -25380 -18980
rect -25120 -19000 -24880 -18980
rect -24620 -19000 -24380 -18980
rect -24120 -19000 -23880 -18980
rect -23620 -19000 -23380 -18980
rect -23120 -19000 -22880 -18980
rect -22620 -19000 -22380 -18980
rect -22120 -19000 -21880 -18980
rect -21620 -19000 -21380 -18980
rect -21120 -19000 -20880 -18980
rect -20620 -19000 -20380 -18980
rect -20120 -19000 -19880 -18980
rect -19620 -19000 -19380 -18980
rect -19120 -19000 -18880 -18980
rect -18620 -19000 -18380 -18980
rect -18120 -19000 -17880 -18980
rect -17620 -19000 -17380 -18980
rect -17120 -19000 -16880 -18980
rect -16620 -19000 -16380 -18980
rect -16120 -19000 -15880 -18980
rect -15620 -19000 -15380 -18980
rect -15120 -19000 -15000 -18980
rect -26500 -19200 -15000 -19000
rect -26500 -19220 -26380 -19200
rect -26120 -19220 -25880 -19200
rect -25620 -19220 -25380 -19200
rect -25120 -19220 -24880 -19200
rect -24620 -19220 -24380 -19200
rect -24120 -19220 -23880 -19200
rect -23620 -19220 -23380 -19200
rect -23120 -19220 -22880 -19200
rect -22620 -19220 -22380 -19200
rect -22120 -19220 -21880 -19200
rect -21620 -19220 -21380 -19200
rect -21120 -19220 -20880 -19200
rect -20620 -19220 -20380 -19200
rect -20120 -19220 -19880 -19200
rect -19620 -19220 -19380 -19200
rect -19120 -19220 -18880 -19200
rect -18620 -19220 -18380 -19200
rect -18120 -19220 -17880 -19200
rect -17620 -19220 -17380 -19200
rect -17120 -19220 -16880 -19200
rect -16620 -19220 -16380 -19200
rect -16120 -19220 -15880 -19200
rect -15620 -19220 -15380 -19200
rect -15120 -19220 -15000 -19200
rect -26500 -19480 -26400 -19220
rect -26100 -19480 -25900 -19220
rect -25600 -19480 -25400 -19220
rect -25100 -19480 -24900 -19220
rect -24600 -19480 -24400 -19220
rect -24100 -19480 -23900 -19220
rect -23600 -19480 -23400 -19220
rect -23100 -19480 -22900 -19220
rect -22600 -19480 -22400 -19220
rect -22100 -19480 -21900 -19220
rect -21600 -19480 -21400 -19220
rect -21100 -19480 -20900 -19220
rect -20600 -19480 -20400 -19220
rect -20100 -19480 -19900 -19220
rect -19600 -19480 -19400 -19220
rect -19100 -19480 -18900 -19220
rect -18600 -19480 -18400 -19220
rect -18100 -19480 -17900 -19220
rect -17600 -19480 -17400 -19220
rect -17100 -19480 -16900 -19220
rect -16600 -19480 -16400 -19220
rect -16100 -19480 -15900 -19220
rect -15600 -19480 -15400 -19220
rect -15100 -19480 -15000 -19220
rect -26500 -19500 -26380 -19480
rect -26120 -19500 -25880 -19480
rect -25620 -19500 -25380 -19480
rect -25120 -19500 -24880 -19480
rect -24620 -19500 -24380 -19480
rect -24120 -19500 -23880 -19480
rect -23620 -19500 -23380 -19480
rect -23120 -19500 -22880 -19480
rect -22620 -19500 -22380 -19480
rect -22120 -19500 -21880 -19480
rect -21620 -19500 -21380 -19480
rect -21120 -19500 -20880 -19480
rect -20620 -19500 -20380 -19480
rect -20120 -19500 -19880 -19480
rect -19620 -19500 -19380 -19480
rect -19120 -19500 -18880 -19480
rect -18620 -19500 -18380 -19480
rect -18120 -19500 -17880 -19480
rect -17620 -19500 -17380 -19480
rect -17120 -19500 -16880 -19480
rect -16620 -19500 -16380 -19480
rect -16120 -19500 -15880 -19480
rect -15620 -19500 -15380 -19480
rect -15120 -19500 -15000 -19480
rect -26500 -19700 -15000 -19500
rect -26500 -19720 -26380 -19700
rect -26120 -19720 -25880 -19700
rect -25620 -19720 -25380 -19700
rect -25120 -19720 -24880 -19700
rect -24620 -19720 -24380 -19700
rect -24120 -19720 -23880 -19700
rect -23620 -19720 -23380 -19700
rect -23120 -19720 -22880 -19700
rect -22620 -19720 -22380 -19700
rect -22120 -19720 -21880 -19700
rect -21620 -19720 -21380 -19700
rect -21120 -19720 -20880 -19700
rect -20620 -19720 -20380 -19700
rect -20120 -19720 -19880 -19700
rect -19620 -19720 -19380 -19700
rect -19120 -19720 -18880 -19700
rect -18620 -19720 -18380 -19700
rect -18120 -19720 -17880 -19700
rect -17620 -19720 -17380 -19700
rect -17120 -19720 -16880 -19700
rect -16620 -19720 -16380 -19700
rect -16120 -19720 -15880 -19700
rect -15620 -19720 -15380 -19700
rect -15120 -19720 -15000 -19700
rect -26500 -19980 -26400 -19720
rect -26100 -19980 -25900 -19720
rect -25600 -19980 -25400 -19720
rect -25100 -19980 -24900 -19720
rect -24600 -19980 -24400 -19720
rect -24100 -19980 -23900 -19720
rect -23600 -19980 -23400 -19720
rect -23100 -19980 -22900 -19720
rect -22600 -19980 -22400 -19720
rect -22100 -19980 -21900 -19720
rect -21600 -19980 -21400 -19720
rect -21100 -19980 -20900 -19720
rect -20600 -19980 -20400 -19720
rect -20100 -19980 -19900 -19720
rect -19600 -19980 -19400 -19720
rect -19100 -19980 -18900 -19720
rect -18600 -19980 -18400 -19720
rect -18100 -19980 -17900 -19720
rect -17600 -19980 -17400 -19720
rect -17100 -19980 -16900 -19720
rect -16600 -19980 -16400 -19720
rect -16100 -19980 -15900 -19720
rect -15600 -19980 -15400 -19720
rect -15100 -19980 -15000 -19720
rect -26500 -20000 -26380 -19980
rect -26120 -20000 -25880 -19980
rect -25620 -20000 -25380 -19980
rect -25120 -20000 -24880 -19980
rect -24620 -20000 -24380 -19980
rect -24120 -20000 -23880 -19980
rect -23620 -20000 -23380 -19980
rect -23120 -20000 -22880 -19980
rect -22620 -20000 -22380 -19980
rect -22120 -20000 -21880 -19980
rect -21620 -20000 -21380 -19980
rect -21120 -20000 -20880 -19980
rect -20620 -20000 -20380 -19980
rect -20120 -20000 -19880 -19980
rect -19620 -20000 -19380 -19980
rect -19120 -20000 -18880 -19980
rect -18620 -20000 -18380 -19980
rect -18120 -20000 -17880 -19980
rect -17620 -20000 -17380 -19980
rect -17120 -20000 -16880 -19980
rect -16620 -20000 -16380 -19980
rect -16120 -20000 -15880 -19980
rect -15620 -20000 -15380 -19980
rect -15120 -20000 -15000 -19980
rect -26500 -20200 -15000 -20000
rect -26500 -20220 -26380 -20200
rect -26120 -20220 -25880 -20200
rect -25620 -20220 -25380 -20200
rect -25120 -20220 -24880 -20200
rect -24620 -20220 -24380 -20200
rect -24120 -20220 -23880 -20200
rect -23620 -20220 -23380 -20200
rect -23120 -20220 -22880 -20200
rect -22620 -20220 -22380 -20200
rect -22120 -20220 -21880 -20200
rect -21620 -20220 -21380 -20200
rect -21120 -20220 -20880 -20200
rect -20620 -20220 -20380 -20200
rect -20120 -20220 -19880 -20200
rect -19620 -20220 -19380 -20200
rect -19120 -20220 -18880 -20200
rect -18620 -20220 -18380 -20200
rect -18120 -20220 -17880 -20200
rect -17620 -20220 -17380 -20200
rect -17120 -20220 -16880 -20200
rect -16620 -20220 -16380 -20200
rect -16120 -20220 -15880 -20200
rect -15620 -20220 -15380 -20200
rect -15120 -20220 -15000 -20200
rect -26500 -20480 -26400 -20220
rect -26100 -20480 -25900 -20220
rect -25600 -20480 -25400 -20220
rect -25100 -20480 -24900 -20220
rect -24600 -20480 -24400 -20220
rect -24100 -20480 -23900 -20220
rect -23600 -20480 -23400 -20220
rect -23100 -20480 -22900 -20220
rect -22600 -20480 -22400 -20220
rect -22100 -20480 -21900 -20220
rect -21600 -20480 -21400 -20220
rect -21100 -20480 -20900 -20220
rect -20600 -20480 -20400 -20220
rect -20100 -20480 -19900 -20220
rect -19600 -20480 -19400 -20220
rect -19100 -20480 -18900 -20220
rect -18600 -20480 -18400 -20220
rect -18100 -20480 -17900 -20220
rect -17600 -20480 -17400 -20220
rect -17100 -20480 -16900 -20220
rect -16600 -20480 -16400 -20220
rect -16100 -20480 -15900 -20220
rect -15600 -20480 -15400 -20220
rect -15100 -20480 -15000 -20220
rect -26500 -20500 -26380 -20480
rect -26120 -20500 -25880 -20480
rect -25620 -20500 -25380 -20480
rect -25120 -20500 -24880 -20480
rect -24620 -20500 -24380 -20480
rect -24120 -20500 -23880 -20480
rect -23620 -20500 -23380 -20480
rect -23120 -20500 -22880 -20480
rect -22620 -20500 -22380 -20480
rect -22120 -20500 -21880 -20480
rect -21620 -20500 -21380 -20480
rect -21120 -20500 -20880 -20480
rect -20620 -20500 -20380 -20480
rect -20120 -20500 -19880 -20480
rect -19620 -20500 -19380 -20480
rect -19120 -20500 -18880 -20480
rect -18620 -20500 -18380 -20480
rect -18120 -20500 -17880 -20480
rect -17620 -20500 -17380 -20480
rect -17120 -20500 -16880 -20480
rect -16620 -20500 -16380 -20480
rect -16120 -20500 -15880 -20480
rect -15620 -20500 -15380 -20480
rect -15120 -20500 -15000 -20480
rect -26500 -20700 -15000 -20500
rect -26500 -20720 -26380 -20700
rect -26120 -20720 -25880 -20700
rect -25620 -20720 -25380 -20700
rect -25120 -20720 -24880 -20700
rect -24620 -20720 -24380 -20700
rect -24120 -20720 -23880 -20700
rect -23620 -20720 -23380 -20700
rect -23120 -20720 -22880 -20700
rect -22620 -20720 -22380 -20700
rect -22120 -20720 -21880 -20700
rect -21620 -20720 -21380 -20700
rect -21120 -20720 -20880 -20700
rect -20620 -20720 -20380 -20700
rect -20120 -20720 -19880 -20700
rect -19620 -20720 -19380 -20700
rect -19120 -20720 -18880 -20700
rect -18620 -20720 -18380 -20700
rect -18120 -20720 -17880 -20700
rect -17620 -20720 -17380 -20700
rect -17120 -20720 -16880 -20700
rect -16620 -20720 -16380 -20700
rect -16120 -20720 -15880 -20700
rect -15620 -20720 -15380 -20700
rect -15120 -20720 -15000 -20700
rect -26500 -20980 -26400 -20720
rect -26100 -20980 -25900 -20720
rect -25600 -20980 -25400 -20720
rect -25100 -20980 -24900 -20720
rect -24600 -20980 -24400 -20720
rect -24100 -20980 -23900 -20720
rect -23600 -20980 -23400 -20720
rect -23100 -20980 -22900 -20720
rect -22600 -20980 -22400 -20720
rect -22100 -20980 -21900 -20720
rect -21600 -20980 -21400 -20720
rect -21100 -20980 -20900 -20720
rect -20600 -20980 -20400 -20720
rect -20100 -20980 -19900 -20720
rect -19600 -20980 -19400 -20720
rect -19100 -20980 -18900 -20720
rect -18600 -20980 -18400 -20720
rect -18100 -20980 -17900 -20720
rect -17600 -20980 -17400 -20720
rect -17100 -20980 -16900 -20720
rect -16600 -20980 -16400 -20720
rect -16100 -20980 -15900 -20720
rect -15600 -20980 -15400 -20720
rect -15100 -20980 -15000 -20720
rect -26500 -21000 -26380 -20980
rect -26120 -21000 -25880 -20980
rect -25620 -21000 -25380 -20980
rect -25120 -21000 -24880 -20980
rect -24620 -21000 -24380 -20980
rect -24120 -21000 -23880 -20980
rect -23620 -21000 -23380 -20980
rect -23120 -21000 -22880 -20980
rect -22620 -21000 -22380 -20980
rect -22120 -21000 -21880 -20980
rect -21620 -21000 -21380 -20980
rect -21120 -21000 -20880 -20980
rect -20620 -21000 -20380 -20980
rect -20120 -21000 -19880 -20980
rect -19620 -21000 -19380 -20980
rect -19120 -21000 -18880 -20980
rect -18620 -21000 -18380 -20980
rect -18120 -21000 -17880 -20980
rect -17620 -21000 -17380 -20980
rect -17120 -21000 -16880 -20980
rect -16620 -21000 -16380 -20980
rect -16120 -21000 -15880 -20980
rect -15620 -21000 -15380 -20980
rect -15120 -21000 -15000 -20980
rect -26500 -21200 -15000 -21000
rect 17500 -13200 18500 -13100
rect 17500 -13220 17620 -13200
rect 17880 -13220 18120 -13200
rect 18380 -13220 18500 -13200
rect 17500 -13480 17600 -13220
rect 17900 -13480 18100 -13220
rect 18400 -13480 18500 -13220
rect 17500 -13500 17620 -13480
rect 17880 -13500 18120 -13480
rect 18380 -13500 18500 -13480
rect 17500 -13700 18500 -13500
rect 17500 -13720 17620 -13700
rect 17880 -13720 18120 -13700
rect 18380 -13720 18500 -13700
rect 17500 -13980 17600 -13720
rect 17900 -13980 18100 -13720
rect 18400 -13980 18500 -13720
rect 17500 -14000 17620 -13980
rect 17880 -14000 18120 -13980
rect 18380 -14000 18500 -13980
rect 17500 -14200 18500 -14000
rect 17500 -14220 17620 -14200
rect 17880 -14220 18120 -14200
rect 18380 -14220 18500 -14200
rect 17500 -14480 17600 -14220
rect 17900 -14480 18100 -14220
rect 18400 -14480 18500 -14220
rect 17500 -14500 17620 -14480
rect 17880 -14500 18120 -14480
rect 18380 -14500 18500 -14480
rect 17500 -14700 18500 -14500
rect 17500 -14720 17620 -14700
rect 17880 -14720 18120 -14700
rect 18380 -14720 18500 -14700
rect 17500 -14980 17600 -14720
rect 17900 -14980 18100 -14720
rect 18400 -14980 18500 -14720
rect 17500 -15000 17620 -14980
rect 17880 -15000 18120 -14980
rect 18380 -15000 18500 -14980
rect 17500 -15200 18500 -15000
rect 17500 -15220 17620 -15200
rect 17880 -15220 18120 -15200
rect 18380 -15220 18500 -15200
rect 17500 -15480 17600 -15220
rect 17900 -15480 18100 -15220
rect 18400 -15480 18500 -15220
rect 17500 -15500 17620 -15480
rect 17880 -15500 18120 -15480
rect 18380 -15500 18500 -15480
rect 17500 -15700 18500 -15500
rect 17500 -15720 17620 -15700
rect 17880 -15720 18120 -15700
rect 18380 -15720 18500 -15700
rect 17500 -15980 17600 -15720
rect 17900 -15980 18100 -15720
rect 18400 -15980 18500 -15720
rect 17500 -16000 17620 -15980
rect 17880 -16000 18120 -15980
rect 18380 -16000 18500 -15980
rect 17500 -16200 18500 -16000
rect 17500 -16220 17620 -16200
rect 17880 -16220 18120 -16200
rect 18380 -16220 18500 -16200
rect 17500 -16480 17600 -16220
rect 17900 -16480 18100 -16220
rect 18400 -16480 18500 -16220
rect 17500 -16500 17620 -16480
rect 17880 -16500 18120 -16480
rect 18380 -16500 18500 -16480
rect 17500 -16700 18500 -16500
rect 17500 -16720 17620 -16700
rect 17880 -16720 18120 -16700
rect 18380 -16720 18500 -16700
rect 17500 -16980 17600 -16720
rect 17900 -16980 18100 -16720
rect 18400 -16980 18500 -16720
rect 17500 -17000 17620 -16980
rect 17880 -17000 18120 -16980
rect 18380 -17000 18500 -16980
rect 17500 -17200 18500 -17000
rect 17500 -17220 17620 -17200
rect 17880 -17220 18120 -17200
rect 18380 -17220 18500 -17200
rect 17500 -17480 17600 -17220
rect 17900 -17480 18100 -17220
rect 18400 -17480 18500 -17220
rect 17500 -17500 17620 -17480
rect 17880 -17500 18120 -17480
rect 18380 -17500 18500 -17480
rect 17500 -17700 18500 -17500
rect 17500 -17720 17620 -17700
rect 17880 -17720 18120 -17700
rect 18380 -17720 18500 -17700
rect 17500 -17980 17600 -17720
rect 17900 -17980 18100 -17720
rect 18400 -17980 18500 -17720
rect 17500 -18000 17620 -17980
rect 17880 -18000 18120 -17980
rect 18380 -18000 18500 -17980
rect 17500 -18200 18500 -18000
rect 17500 -18220 17620 -18200
rect 17880 -18220 18120 -18200
rect 18380 -18220 18500 -18200
rect 17500 -18480 17600 -18220
rect 17900 -18480 18100 -18220
rect 18400 -18480 18500 -18220
rect 17500 -18500 17620 -18480
rect 17880 -18500 18120 -18480
rect 18380 -18500 18500 -18480
rect 17500 -18700 18500 -18500
rect 17500 -18720 17620 -18700
rect 17880 -18720 18120 -18700
rect 18380 -18720 18500 -18700
rect 17500 -18980 17600 -18720
rect 17900 -18980 18100 -18720
rect 18400 -18980 18500 -18720
rect 17500 -19000 17620 -18980
rect 17880 -19000 18120 -18980
rect 18380 -19000 18500 -18980
rect 17500 -19200 18500 -19000
rect 17500 -19220 17620 -19200
rect 17880 -19220 18120 -19200
rect 18380 -19220 18500 -19200
rect 17500 -19480 17600 -19220
rect 17900 -19480 18100 -19220
rect 18400 -19480 18500 -19220
rect 17500 -19500 17620 -19480
rect 17880 -19500 18120 -19480
rect 18380 -19500 18500 -19480
rect 17500 -19700 18500 -19500
rect 17500 -19720 17620 -19700
rect 17880 -19720 18120 -19700
rect 18380 -19720 18500 -19700
rect 17500 -19980 17600 -19720
rect 17900 -19980 18100 -19720
rect 18400 -19980 18500 -19720
rect 17500 -20000 17620 -19980
rect 17880 -20000 18120 -19980
rect 18380 -20000 18500 -19980
rect 17500 -20100 18500 -20000
rect 23500 -12200 24000 -12000
rect 23500 -12220 23620 -12200
rect 23880 -12220 24000 -12200
rect 23500 -12480 23600 -12220
rect 23900 -12480 24000 -12220
rect 23500 -12500 23620 -12480
rect 23880 -12500 24000 -12480
rect 23500 -12700 24000 -12500
rect 23500 -12720 23620 -12700
rect 23880 -12720 24000 -12700
rect 23500 -12980 23600 -12720
rect 23900 -12980 24000 -12720
rect 23500 -13000 23620 -12980
rect 23880 -13000 24000 -12980
rect 23500 -13200 24000 -13000
rect 23500 -13220 23620 -13200
rect 23880 -13220 24000 -13200
rect 23500 -13480 23600 -13220
rect 23900 -13480 24000 -13220
rect 23500 -13500 23620 -13480
rect 23880 -13500 24000 -13480
rect 23500 -13700 24000 -13500
rect 23500 -13720 23620 -13700
rect 23880 -13720 24000 -13700
rect 23500 -13980 23600 -13720
rect 23900 -13980 24000 -13720
rect 23500 -14000 23620 -13980
rect 23880 -14000 24000 -13980
rect 23500 -14200 24000 -14000
rect 23500 -14220 23620 -14200
rect 23880 -14220 24000 -14200
rect 23500 -14480 23600 -14220
rect 23900 -14480 24000 -14220
rect 23500 -14500 23620 -14480
rect 23880 -14500 24000 -14480
rect 23500 -14700 24000 -14500
rect 23500 -14720 23620 -14700
rect 23880 -14720 24000 -14700
rect 23500 -14980 23600 -14720
rect 23900 -14980 24000 -14720
rect 23500 -15000 23620 -14980
rect 23880 -15000 24000 -14980
rect 23500 -15200 24000 -15000
rect 23500 -15220 23620 -15200
rect 23880 -15220 24000 -15200
rect 23500 -15480 23600 -15220
rect 23900 -15480 24000 -15220
rect 23500 -15500 23620 -15480
rect 23880 -15500 24000 -15480
rect 23500 -15700 24000 -15500
rect 23500 -15720 23620 -15700
rect 23880 -15720 24000 -15700
rect 23500 -15980 23600 -15720
rect 23900 -15980 24000 -15720
rect 23500 -16000 23620 -15980
rect 23880 -16000 24000 -15980
rect 23500 -16200 24000 -16000
rect 23500 -16220 23620 -16200
rect 23880 -16220 24000 -16200
rect 23500 -16480 23600 -16220
rect 23900 -16480 24000 -16220
rect 23500 -16500 23620 -16480
rect 23880 -16500 24000 -16480
rect 23500 -16700 24000 -16500
rect 23500 -16720 23620 -16700
rect 23880 -16720 24000 -16700
rect 23500 -16980 23600 -16720
rect 23900 -16980 24000 -16720
rect 23500 -17000 23620 -16980
rect 23880 -17000 24000 -16980
rect 23500 -17200 24000 -17000
rect 23500 -17220 23620 -17200
rect 23880 -17220 24000 -17200
rect 23500 -17480 23600 -17220
rect 23900 -17480 24000 -17220
rect 23500 -17500 23620 -17480
rect 23880 -17500 24000 -17480
rect 23500 -17700 24000 -17500
rect 23500 -17720 23620 -17700
rect 23880 -17720 24000 -17700
rect 23500 -17980 23600 -17720
rect 23900 -17980 24000 -17720
rect 23500 -18000 23620 -17980
rect 23880 -18000 24000 -17980
rect 23500 -18200 24000 -18000
rect 23500 -18220 23620 -18200
rect 23880 -18220 24000 -18200
rect 23500 -18480 23600 -18220
rect 23900 -18480 24000 -18220
rect 23500 -18500 23620 -18480
rect 23880 -18500 24000 -18480
rect 23500 -18700 24000 -18500
rect 23500 -18720 23620 -18700
rect 23880 -18720 24000 -18700
rect 23500 -18980 23600 -18720
rect 23900 -18980 24000 -18720
rect 23500 -19000 23620 -18980
rect 23880 -19000 24000 -18980
rect 23500 -19200 24000 -19000
rect 23500 -19220 23620 -19200
rect 23880 -19220 24000 -19200
rect 23500 -19480 23600 -19220
rect 23900 -19480 24000 -19220
rect 23500 -19500 23620 -19480
rect 23880 -19500 24000 -19480
rect 23500 -19700 24000 -19500
rect 23500 -19720 23620 -19700
rect 23880 -19720 24000 -19700
rect 23500 -19980 23600 -19720
rect 23900 -19980 24000 -19720
rect 23500 -20000 23620 -19980
rect 23880 -20000 24000 -19980
rect 17500 -20200 20500 -20100
rect 17500 -20220 17620 -20200
rect 17880 -20220 18120 -20200
rect 18380 -20220 18620 -20200
rect 18880 -20220 19120 -20200
rect 19380 -20220 19620 -20200
rect 19880 -20220 20120 -20200
rect 20380 -20220 20500 -20200
rect 17500 -20480 17600 -20220
rect 17900 -20480 18100 -20220
rect 18400 -20480 18600 -20220
rect 18900 -20480 19100 -20220
rect 19400 -20480 19600 -20220
rect 19900 -20480 20100 -20220
rect 20400 -20480 20500 -20220
rect 17500 -20500 17620 -20480
rect 17880 -20500 18120 -20480
rect 18380 -20500 18620 -20480
rect 18880 -20500 19120 -20480
rect 19380 -20500 19620 -20480
rect 19880 -20500 20120 -20480
rect 20380 -20500 20500 -20480
rect 17500 -20700 20500 -20500
rect 17500 -20720 17620 -20700
rect 17880 -20720 18120 -20700
rect 18380 -20720 18620 -20700
rect 18880 -20720 19120 -20700
rect 19380 -20720 19620 -20700
rect 19880 -20720 20120 -20700
rect 20380 -20720 20500 -20700
rect 17500 -20980 17600 -20720
rect 17900 -20980 18100 -20720
rect 18400 -20980 18600 -20720
rect 18900 -20980 19100 -20720
rect 19400 -20980 19600 -20720
rect 19900 -20980 20100 -20720
rect 20400 -20980 20500 -20720
rect 17500 -21000 17620 -20980
rect 17880 -21000 18120 -20980
rect 18380 -21000 18620 -20980
rect 18880 -21000 19120 -20980
rect 19380 -21000 19620 -20980
rect 19880 -21000 20120 -20980
rect 20380 -21000 20500 -20980
rect 17500 -21100 20500 -21000
rect -26500 -21220 -26380 -21200
rect -26120 -21220 -25880 -21200
rect -25620 -21220 -25380 -21200
rect -25120 -21220 -24880 -21200
rect -24620 -21220 -24380 -21200
rect -24120 -21220 -23880 -21200
rect -23620 -21220 -23380 -21200
rect -23120 -21220 -22880 -21200
rect -22620 -21220 -22380 -21200
rect -22120 -21220 -21880 -21200
rect -21620 -21220 -21380 -21200
rect -21120 -21220 -20880 -21200
rect -20620 -21220 -20380 -21200
rect -20120 -21220 -19880 -21200
rect -19620 -21220 -19380 -21200
rect -19120 -21220 -18880 -21200
rect -18620 -21220 -18380 -21200
rect -18120 -21220 -17880 -21200
rect -17620 -21220 -17380 -21200
rect -17120 -21220 -16880 -21200
rect -16620 -21220 -16380 -21200
rect -16120 -21220 -15880 -21200
rect -15620 -21220 -15380 -21200
rect -15120 -21220 -15000 -21200
rect -26500 -21480 -26400 -21220
rect -26100 -21480 -25900 -21220
rect -25600 -21480 -25400 -21220
rect -25100 -21480 -24900 -21220
rect -24600 -21480 -24400 -21220
rect -24100 -21480 -23900 -21220
rect -23600 -21480 -23400 -21220
rect -23100 -21480 -22900 -21220
rect -22600 -21480 -22400 -21220
rect -22100 -21480 -21900 -21220
rect -21600 -21480 -21400 -21220
rect -21100 -21480 -20900 -21220
rect -20600 -21480 -20400 -21220
rect -20100 -21480 -19900 -21220
rect -19600 -21480 -19400 -21220
rect -19100 -21480 -18900 -21220
rect -18600 -21480 -18400 -21220
rect -18100 -21480 -17900 -21220
rect -17600 -21480 -17400 -21220
rect -17100 -21480 -16900 -21220
rect -16600 -21480 -16400 -21220
rect -16100 -21480 -15900 -21220
rect -15600 -21480 -15400 -21220
rect -15100 -21480 -15000 -21220
rect -26500 -21500 -26380 -21480
rect -26120 -21500 -25880 -21480
rect -25620 -21500 -25380 -21480
rect -25120 -21500 -24880 -21480
rect -24620 -21500 -24380 -21480
rect -24120 -21500 -23880 -21480
rect -23620 -21500 -23380 -21480
rect -23120 -21500 -22880 -21480
rect -22620 -21500 -22380 -21480
rect -22120 -21500 -21880 -21480
rect -21620 -21500 -21380 -21480
rect -21120 -21500 -20880 -21480
rect -20620 -21500 -20380 -21480
rect -20120 -21500 -19880 -21480
rect -19620 -21500 -19380 -21480
rect -19120 -21500 -18880 -21480
rect -18620 -21500 -18380 -21480
rect -18120 -21500 -17880 -21480
rect -17620 -21500 -17380 -21480
rect -17120 -21500 -16880 -21480
rect -16620 -21500 -16380 -21480
rect -16120 -21500 -15880 -21480
rect -15620 -21500 -15380 -21480
rect -15120 -21500 -15000 -21480
rect -26500 -21700 -15000 -21500
rect -26500 -21720 -26380 -21700
rect -26120 -21720 -25880 -21700
rect -25620 -21720 -25380 -21700
rect -25120 -21720 -24880 -21700
rect -24620 -21720 -24380 -21700
rect -24120 -21720 -23880 -21700
rect -23620 -21720 -23380 -21700
rect -23120 -21720 -22880 -21700
rect -22620 -21720 -22380 -21700
rect -22120 -21720 -21880 -21700
rect -21620 -21720 -21380 -21700
rect -21120 -21720 -20880 -21700
rect -20620 -21720 -20380 -21700
rect -20120 -21720 -19880 -21700
rect -19620 -21720 -19380 -21700
rect -19120 -21720 -18880 -21700
rect -18620 -21720 -18380 -21700
rect -18120 -21720 -17880 -21700
rect -17620 -21720 -17380 -21700
rect -17120 -21720 -16880 -21700
rect -16620 -21720 -16380 -21700
rect -16120 -21720 -15880 -21700
rect -15620 -21720 -15380 -21700
rect -15120 -21720 -15000 -21700
rect -26500 -21980 -26400 -21720
rect -26100 -21980 -25900 -21720
rect -25600 -21980 -25400 -21720
rect -25100 -21980 -24900 -21720
rect -24600 -21980 -24400 -21720
rect -24100 -21980 -23900 -21720
rect -23600 -21980 -23400 -21720
rect -23100 -21980 -22900 -21720
rect -22600 -21980 -22400 -21720
rect -22100 -21980 -21900 -21720
rect -21600 -21980 -21400 -21720
rect -21100 -21980 -20900 -21720
rect -20600 -21980 -20400 -21720
rect -20100 -21980 -19900 -21720
rect -19600 -21980 -19400 -21720
rect -19100 -21980 -18900 -21720
rect -18600 -21980 -18400 -21720
rect -18100 -21980 -17900 -21720
rect -17600 -21980 -17400 -21720
rect -17100 -21980 -16900 -21720
rect -16600 -21980 -16400 -21720
rect -16100 -21980 -15900 -21720
rect -15600 -21980 -15400 -21720
rect -15100 -21980 -15000 -21720
rect -26500 -22000 -26380 -21980
rect -26120 -22000 -25880 -21980
rect -25620 -22000 -25380 -21980
rect -25120 -22000 -24880 -21980
rect -24620 -22000 -24380 -21980
rect -24120 -22000 -23880 -21980
rect -23620 -22000 -23380 -21980
rect -23120 -22000 -22880 -21980
rect -22620 -22000 -22380 -21980
rect -22120 -22000 -21880 -21980
rect -21620 -22000 -21380 -21980
rect -21120 -22000 -20880 -21980
rect -20620 -22000 -20380 -21980
rect -20120 -22000 -19880 -21980
rect -19620 -22000 -19380 -21980
rect -19120 -22000 -18880 -21980
rect -18620 -22000 -18380 -21980
rect -18120 -22000 -17880 -21980
rect -17620 -22000 -17380 -21980
rect -17120 -22000 -16880 -21980
rect -16620 -22000 -16380 -21980
rect -16120 -22000 -15880 -21980
rect -15620 -22000 -15380 -21980
rect -15120 -22000 -15000 -21980
rect -26500 -22200 -15000 -22000
rect -26500 -22220 -26380 -22200
rect -26120 -22220 -25880 -22200
rect -25620 -22220 -25380 -22200
rect -25120 -22220 -24880 -22200
rect -24620 -22220 -24380 -22200
rect -24120 -22220 -23880 -22200
rect -23620 -22220 -23380 -22200
rect -23120 -22220 -22880 -22200
rect -22620 -22220 -22380 -22200
rect -22120 -22220 -21880 -22200
rect -21620 -22220 -21380 -22200
rect -21120 -22220 -20880 -22200
rect -20620 -22220 -20380 -22200
rect -20120 -22220 -19880 -22200
rect -19620 -22220 -19380 -22200
rect -19120 -22220 -18880 -22200
rect -18620 -22220 -18380 -22200
rect -18120 -22220 -17880 -22200
rect -17620 -22220 -17380 -22200
rect -17120 -22220 -16880 -22200
rect -16620 -22220 -16380 -22200
rect -16120 -22220 -15880 -22200
rect -15620 -22220 -15380 -22200
rect -15120 -22220 -15000 -22200
rect -26500 -22480 -26400 -22220
rect -26100 -22480 -25900 -22220
rect -25600 -22480 -25400 -22220
rect -25100 -22480 -24900 -22220
rect -24600 -22480 -24400 -22220
rect -24100 -22480 -23900 -22220
rect -23600 -22480 -23400 -22220
rect -23100 -22480 -22900 -22220
rect -22600 -22480 -22400 -22220
rect -22100 -22480 -21900 -22220
rect -21600 -22480 -21400 -22220
rect -21100 -22480 -20900 -22220
rect -20600 -22480 -20400 -22220
rect -20100 -22480 -19900 -22220
rect -19600 -22480 -19400 -22220
rect -19100 -22480 -18900 -22220
rect -18600 -22480 -18400 -22220
rect -18100 -22480 -17900 -22220
rect -17600 -22480 -17400 -22220
rect -17100 -22480 -16900 -22220
rect -16600 -22480 -16400 -22220
rect -16100 -22480 -15900 -22220
rect -15600 -22480 -15400 -22220
rect -15100 -22480 -15000 -22220
rect -26500 -22500 -26380 -22480
rect -26120 -22500 -25880 -22480
rect -25620 -22500 -25380 -22480
rect -25120 -22500 -24880 -22480
rect -24620 -22500 -24380 -22480
rect -24120 -22500 -23880 -22480
rect -23620 -22500 -23380 -22480
rect -23120 -22500 -22880 -22480
rect -22620 -22500 -22380 -22480
rect -22120 -22500 -21880 -22480
rect -21620 -22500 -21380 -22480
rect -21120 -22500 -20880 -22480
rect -20620 -22500 -20380 -22480
rect -20120 -22500 -19880 -22480
rect -19620 -22500 -19380 -22480
rect -19120 -22500 -18880 -22480
rect -18620 -22500 -18380 -22480
rect -18120 -22500 -17880 -22480
rect -17620 -22500 -17380 -22480
rect -17120 -22500 -16880 -22480
rect -16620 -22500 -16380 -22480
rect -16120 -22500 -15880 -22480
rect -15620 -22500 -15380 -22480
rect -15120 -22500 -15000 -22480
rect -26500 -22700 -15000 -22500
rect -26500 -22720 -26380 -22700
rect -26120 -22720 -25880 -22700
rect -25620 -22720 -25380 -22700
rect -25120 -22720 -24880 -22700
rect -24620 -22720 -24380 -22700
rect -24120 -22720 -23880 -22700
rect -23620 -22720 -23380 -22700
rect -23120 -22720 -22880 -22700
rect -22620 -22720 -22380 -22700
rect -22120 -22720 -21880 -22700
rect -21620 -22720 -21380 -22700
rect -21120 -22720 -20880 -22700
rect -20620 -22720 -20380 -22700
rect -20120 -22720 -19880 -22700
rect -19620 -22720 -19380 -22700
rect -19120 -22720 -18880 -22700
rect -18620 -22720 -18380 -22700
rect -18120 -22720 -17880 -22700
rect -17620 -22720 -17380 -22700
rect -17120 -22720 -16880 -22700
rect -16620 -22720 -16380 -22700
rect -16120 -22720 -15880 -22700
rect -15620 -22720 -15380 -22700
rect -15120 -22720 -15000 -22700
rect -26500 -22980 -26400 -22720
rect -26100 -22980 -25900 -22720
rect -25600 -22980 -25400 -22720
rect -25100 -22980 -24900 -22720
rect -24600 -22980 -24400 -22720
rect -24100 -22980 -23900 -22720
rect -23600 -22980 -23400 -22720
rect -23100 -22980 -22900 -22720
rect -22600 -22980 -22400 -22720
rect -22100 -22980 -21900 -22720
rect -21600 -22980 -21400 -22720
rect -21100 -22980 -20900 -22720
rect -20600 -22980 -20400 -22720
rect -20100 -22980 -19900 -22720
rect -19600 -22980 -19400 -22720
rect -19100 -22980 -18900 -22720
rect -18600 -22980 -18400 -22720
rect -18100 -22980 -17900 -22720
rect -17600 -22980 -17400 -22720
rect -17100 -22980 -16900 -22720
rect -16600 -22980 -16400 -22720
rect -16100 -22980 -15900 -22720
rect -15600 -22980 -15400 -22720
rect -15100 -22980 -15000 -22720
rect -26500 -23000 -26380 -22980
rect -26120 -23000 -25880 -22980
rect -25620 -23000 -25380 -22980
rect -25120 -23000 -24880 -22980
rect -24620 -23000 -24380 -22980
rect -24120 -23000 -23880 -22980
rect -23620 -23000 -23380 -22980
rect -23120 -23000 -22880 -22980
rect -22620 -23000 -22380 -22980
rect -22120 -23000 -21880 -22980
rect -21620 -23000 -21380 -22980
rect -21120 -23000 -20880 -22980
rect -20620 -23000 -20380 -22980
rect -20120 -23000 -19880 -22980
rect -19620 -23000 -19380 -22980
rect -19120 -23000 -18880 -22980
rect -18620 -23000 -18380 -22980
rect -18120 -23000 -17880 -22980
rect -17620 -23000 -17380 -22980
rect -17120 -23000 -16880 -22980
rect -16620 -23000 -16380 -22980
rect -16120 -23000 -15880 -22980
rect -15620 -23000 -15380 -22980
rect -15120 -23000 -15000 -22980
rect -26500 -23200 -15000 -23000
rect -26500 -23220 -26380 -23200
rect -26120 -23220 -25880 -23200
rect -25620 -23220 -25380 -23200
rect -25120 -23220 -24880 -23200
rect -24620 -23220 -24380 -23200
rect -24120 -23220 -23880 -23200
rect -23620 -23220 -23380 -23200
rect -23120 -23220 -22880 -23200
rect -22620 -23220 -22380 -23200
rect -22120 -23220 -21880 -23200
rect -21620 -23220 -21380 -23200
rect -21120 -23220 -20880 -23200
rect -20620 -23220 -20380 -23200
rect -20120 -23220 -19880 -23200
rect -19620 -23220 -19380 -23200
rect -19120 -23220 -18880 -23200
rect -18620 -23220 -18380 -23200
rect -18120 -23220 -17880 -23200
rect -17620 -23220 -17380 -23200
rect -17120 -23220 -16880 -23200
rect -16620 -23220 -16380 -23200
rect -16120 -23220 -15880 -23200
rect -15620 -23220 -15380 -23200
rect -15120 -23220 -15000 -23200
rect -26500 -23480 -26400 -23220
rect -26100 -23480 -25900 -23220
rect -25600 -23480 -25400 -23220
rect -25100 -23480 -24900 -23220
rect -24600 -23480 -24400 -23220
rect -24100 -23480 -23900 -23220
rect -23600 -23480 -23400 -23220
rect -23100 -23480 -22900 -23220
rect -22600 -23480 -22400 -23220
rect -22100 -23480 -21900 -23220
rect -21600 -23480 -21400 -23220
rect -21100 -23480 -20900 -23220
rect -20600 -23480 -20400 -23220
rect -20100 -23480 -19900 -23220
rect -19600 -23480 -19400 -23220
rect -19100 -23480 -18900 -23220
rect -18600 -23480 -18400 -23220
rect -18100 -23480 -17900 -23220
rect -17600 -23480 -17400 -23220
rect -17100 -23480 -16900 -23220
rect -16600 -23480 -16400 -23220
rect -16100 -23480 -15900 -23220
rect -15600 -23480 -15400 -23220
rect -15100 -23480 -15000 -23220
rect -26500 -23500 -26380 -23480
rect -26120 -23500 -25880 -23480
rect -25620 -23500 -25380 -23480
rect -25120 -23500 -24880 -23480
rect -24620 -23500 -24380 -23480
rect -24120 -23500 -23880 -23480
rect -23620 -23500 -23380 -23480
rect -23120 -23500 -22880 -23480
rect -22620 -23500 -22380 -23480
rect -22120 -23500 -21880 -23480
rect -21620 -23500 -21380 -23480
rect -21120 -23500 -20880 -23480
rect -20620 -23500 -20380 -23480
rect -20120 -23500 -19880 -23480
rect -19620 -23500 -19380 -23480
rect -19120 -23500 -18880 -23480
rect -18620 -23500 -18380 -23480
rect -18120 -23500 -17880 -23480
rect -17620 -23500 -17380 -23480
rect -17120 -23500 -16880 -23480
rect -16620 -23500 -16380 -23480
rect -16120 -23500 -15880 -23480
rect -15620 -23500 -15380 -23480
rect -15120 -23500 -15000 -23480
rect -26500 -23700 -15000 -23500
rect -26500 -23720 -26380 -23700
rect -26120 -23720 -25880 -23700
rect -25620 -23720 -25380 -23700
rect -25120 -23720 -24880 -23700
rect -24620 -23720 -24380 -23700
rect -24120 -23720 -23880 -23700
rect -23620 -23720 -23380 -23700
rect -23120 -23720 -22880 -23700
rect -22620 -23720 -22380 -23700
rect -22120 -23720 -21880 -23700
rect -21620 -23720 -21380 -23700
rect -21120 -23720 -20880 -23700
rect -20620 -23720 -20380 -23700
rect -20120 -23720 -19880 -23700
rect -19620 -23720 -19380 -23700
rect -19120 -23720 -18880 -23700
rect -18620 -23720 -18380 -23700
rect -18120 -23720 -17880 -23700
rect -17620 -23720 -17380 -23700
rect -17120 -23720 -16880 -23700
rect -16620 -23720 -16380 -23700
rect -16120 -23720 -15880 -23700
rect -15620 -23720 -15380 -23700
rect -15120 -23720 -15000 -23700
rect -26500 -23980 -26400 -23720
rect -26100 -23980 -25900 -23720
rect -25600 -23980 -25400 -23720
rect -25100 -23980 -24900 -23720
rect -24600 -23980 -24400 -23720
rect -24100 -23980 -23900 -23720
rect -23600 -23980 -23400 -23720
rect -23100 -23980 -22900 -23720
rect -22600 -23980 -22400 -23720
rect -22100 -23980 -21900 -23720
rect -21600 -23980 -21400 -23720
rect -21100 -23980 -20900 -23720
rect -20600 -23980 -20400 -23720
rect -20100 -23980 -19900 -23720
rect -19600 -23980 -19400 -23720
rect -19100 -23980 -18900 -23720
rect -18600 -23980 -18400 -23720
rect -18100 -23980 -17900 -23720
rect -17600 -23980 -17400 -23720
rect -17100 -23980 -16900 -23720
rect -16600 -23980 -16400 -23720
rect -16100 -23980 -15900 -23720
rect -15600 -23980 -15400 -23720
rect -15100 -23980 -15000 -23720
rect -26500 -24000 -26380 -23980
rect -26120 -24000 -25880 -23980
rect -25620 -24000 -25380 -23980
rect -25120 -24000 -24880 -23980
rect -24620 -24000 -24380 -23980
rect -24120 -24000 -23880 -23980
rect -23620 -24000 -23380 -23980
rect -23120 -24000 -22880 -23980
rect -22620 -24000 -22380 -23980
rect -22120 -24000 -21880 -23980
rect -21620 -24000 -21380 -23980
rect -21120 -24000 -20880 -23980
rect -20620 -24000 -20380 -23980
rect -20120 -24000 -19880 -23980
rect -19620 -24000 -19380 -23980
rect -19120 -24000 -18880 -23980
rect -18620 -24000 -18380 -23980
rect -18120 -24000 -17880 -23980
rect -17620 -24000 -17380 -23980
rect -17120 -24000 -16880 -23980
rect -16620 -24000 -16380 -23980
rect -16120 -24000 -15880 -23980
rect -15620 -24000 -15380 -23980
rect -15120 -24000 -15000 -23980
rect -26500 -24100 -15000 -24000
rect 19500 -21200 20500 -21100
rect 19500 -21220 19620 -21200
rect 19880 -21220 20120 -21200
rect 20380 -21220 20500 -21200
rect 19500 -21480 19600 -21220
rect 19900 -21480 20100 -21220
rect 20400 -21480 20500 -21220
rect 19500 -21500 19620 -21480
rect 19880 -21500 20120 -21480
rect 20380 -21500 20500 -21480
rect 19500 -21700 20500 -21500
rect 19500 -21720 19620 -21700
rect 19880 -21720 20120 -21700
rect 20380 -21720 20500 -21700
rect 19500 -21980 19600 -21720
rect 19900 -21980 20100 -21720
rect 20400 -21980 20500 -21720
rect 19500 -22000 19620 -21980
rect 19880 -22000 20120 -21980
rect 20380 -22000 20500 -21980
rect 19500 -22200 20500 -22000
rect 19500 -22220 19620 -22200
rect 19880 -22220 20120 -22200
rect 20380 -22220 20500 -22200
rect 19500 -22480 19600 -22220
rect 19900 -22480 20100 -22220
rect 20400 -22480 20500 -22220
rect 19500 -22500 19620 -22480
rect 19880 -22500 20120 -22480
rect 20380 -22500 20500 -22480
rect 19500 -22700 20500 -22500
rect 19500 -22720 19620 -22700
rect 19880 -22720 20120 -22700
rect 20380 -22720 20500 -22700
rect 19500 -22980 19600 -22720
rect 19900 -22980 20100 -22720
rect 20400 -22980 20500 -22720
rect 19500 -23000 19620 -22980
rect 19880 -23000 20120 -22980
rect 20380 -23000 20500 -22980
rect 19500 -23200 20500 -23000
rect 19500 -23220 19620 -23200
rect 19880 -23220 20120 -23200
rect 20380 -23220 20500 -23200
rect 19500 -23480 19600 -23220
rect 19900 -23480 20100 -23220
rect 20400 -23480 20500 -23220
rect 19500 -23500 19620 -23480
rect 19880 -23500 20120 -23480
rect 20380 -23500 20500 -23480
rect 19500 -23700 20500 -23500
rect 19500 -23720 19620 -23700
rect 19880 -23720 20120 -23700
rect 20380 -23720 20500 -23700
rect 19500 -23980 19600 -23720
rect 19900 -23980 20100 -23720
rect 20400 -23980 20500 -23720
rect 19500 -24000 19620 -23980
rect 19880 -24000 20120 -23980
rect 20380 -24000 20500 -23980
rect -26500 -24200 -17000 -24100
rect -26500 -24220 -26380 -24200
rect -26120 -24220 -25880 -24200
rect -25620 -24220 -25380 -24200
rect -25120 -24220 -24880 -24200
rect -24620 -24220 -24380 -24200
rect -24120 -24220 -23880 -24200
rect -23620 -24220 -23380 -24200
rect -23120 -24220 -22880 -24200
rect -22620 -24220 -22380 -24200
rect -22120 -24220 -21880 -24200
rect -21620 -24220 -21380 -24200
rect -21120 -24220 -20880 -24200
rect -20620 -24220 -20380 -24200
rect -20120 -24220 -19880 -24200
rect -19620 -24220 -19380 -24200
rect -19120 -24220 -18880 -24200
rect -18620 -24220 -18380 -24200
rect -18120 -24220 -17880 -24200
rect -17620 -24220 -17380 -24200
rect -17120 -24220 -17000 -24200
rect -26500 -24480 -26400 -24220
rect -26100 -24480 -25900 -24220
rect -25600 -24480 -25400 -24220
rect -25100 -24480 -24900 -24220
rect -24600 -24480 -24400 -24220
rect -24100 -24480 -23900 -24220
rect -23600 -24480 -23400 -24220
rect -23100 -24480 -22900 -24220
rect -22600 -24480 -22400 -24220
rect -22100 -24480 -21900 -24220
rect -21600 -24480 -21400 -24220
rect -21100 -24480 -20900 -24220
rect -20600 -24480 -20400 -24220
rect -20100 -24480 -19900 -24220
rect -19600 -24480 -19400 -24220
rect -19100 -24480 -18900 -24220
rect -18600 -24480 -18400 -24220
rect -18100 -24480 -17900 -24220
rect -17600 -24480 -17400 -24220
rect -17100 -24480 -17000 -24220
rect -26500 -24500 -26380 -24480
rect -26120 -24500 -25880 -24480
rect -25620 -24500 -25380 -24480
rect -25120 -24500 -24880 -24480
rect -24620 -24500 -24380 -24480
rect -24120 -24500 -23880 -24480
rect -23620 -24500 -23380 -24480
rect -23120 -24500 -22880 -24480
rect -22620 -24500 -22380 -24480
rect -22120 -24500 -21880 -24480
rect -21620 -24500 -21380 -24480
rect -21120 -24500 -20880 -24480
rect -20620 -24500 -20380 -24480
rect -20120 -24500 -19880 -24480
rect -19620 -24500 -19380 -24480
rect -19120 -24500 -18880 -24480
rect -18620 -24500 -18380 -24480
rect -18120 -24500 -17880 -24480
rect -17620 -24500 -17380 -24480
rect -17120 -24500 -17000 -24480
rect -26500 -24600 -17000 -24500
rect 19500 -24200 20500 -24000
rect 19500 -24220 19620 -24200
rect 19880 -24220 20120 -24200
rect 20380 -24220 20500 -24200
rect 19500 -24480 19600 -24220
rect 19900 -24480 20100 -24220
rect 20400 -24480 20500 -24220
rect 19500 -24500 19620 -24480
rect 19880 -24500 20120 -24480
rect 20380 -24500 20500 -24480
rect -26500 -24700 -19000 -24600
rect -26500 -24720 -26380 -24700
rect -26120 -24720 -25880 -24700
rect -25620 -24720 -25380 -24700
rect -25120 -24720 -24880 -24700
rect -24620 -24720 -24380 -24700
rect -24120 -24720 -23880 -24700
rect -23620 -24720 -23380 -24700
rect -23120 -24720 -22880 -24700
rect -22620 -24720 -22380 -24700
rect -22120 -24720 -21880 -24700
rect -21620 -24720 -21380 -24700
rect -21120 -24720 -20880 -24700
rect -20620 -24720 -20380 -24700
rect -20120 -24720 -19880 -24700
rect -19620 -24720 -19380 -24700
rect -19120 -24720 -19000 -24700
rect -26500 -24980 -26400 -24720
rect -26100 -24980 -25900 -24720
rect -25600 -24980 -25400 -24720
rect -25100 -24980 -24900 -24720
rect -24600 -24980 -24400 -24720
rect -24100 -24980 -23900 -24720
rect -23600 -24980 -23400 -24720
rect -23100 -24980 -22900 -24720
rect -22600 -24980 -22400 -24720
rect -22100 -24980 -21900 -24720
rect -21600 -24980 -21400 -24720
rect -21100 -24980 -20900 -24720
rect -20600 -24980 -20400 -24720
rect -20100 -24980 -19900 -24720
rect -19600 -24980 -19400 -24720
rect -19100 -24980 -19000 -24720
rect -26500 -25000 -26380 -24980
rect -26120 -25000 -25880 -24980
rect -25620 -25000 -25380 -24980
rect -25120 -25000 -24880 -24980
rect -24620 -25000 -24380 -24980
rect -24120 -25000 -23880 -24980
rect -23620 -25000 -23380 -24980
rect -23120 -25000 -22880 -24980
rect -22620 -25000 -22380 -24980
rect -22120 -25000 -21880 -24980
rect -21620 -25000 -21380 -24980
rect -21120 -25000 -20880 -24980
rect -20620 -25000 -20380 -24980
rect -20120 -25000 -19880 -24980
rect -19620 -25000 -19380 -24980
rect -19120 -25000 -19000 -24980
rect -26500 -25100 -19000 -25000
rect 19500 -24700 20500 -24500
rect 19500 -24720 19620 -24700
rect 19880 -24720 20120 -24700
rect 20380 -24720 20500 -24700
rect 19500 -24980 19600 -24720
rect 19900 -24980 20100 -24720
rect 20400 -24980 20500 -24720
rect 19500 -25000 19620 -24980
rect 19880 -25000 20120 -24980
rect 20380 -25000 20500 -24980
rect -26500 -25200 -21500 -25100
rect -26500 -25220 -26380 -25200
rect -26120 -25220 -25880 -25200
rect -25620 -25220 -25380 -25200
rect -25120 -25220 -24880 -25200
rect -24620 -25220 -24380 -25200
rect -24120 -25220 -23880 -25200
rect -23620 -25220 -23380 -25200
rect -23120 -25220 -22880 -25200
rect -22620 -25220 -22380 -25200
rect -22120 -25220 -21880 -25200
rect -21620 -25220 -21500 -25200
rect -26500 -25480 -26400 -25220
rect -26100 -25480 -25900 -25220
rect -25600 -25480 -25400 -25220
rect -25100 -25480 -24900 -25220
rect -24600 -25480 -24400 -25220
rect -24100 -25480 -23900 -25220
rect -23600 -25480 -23400 -25220
rect -23100 -25480 -22900 -25220
rect -22600 -25480 -22400 -25220
rect -22100 -25480 -21900 -25220
rect -21600 -25480 -21500 -25220
rect -26500 -25500 -26380 -25480
rect -26120 -25500 -25880 -25480
rect -25620 -25500 -25380 -25480
rect -25120 -25500 -24880 -25480
rect -24620 -25500 -24380 -25480
rect -24120 -25500 -23880 -25480
rect -23620 -25500 -23380 -25480
rect -23120 -25500 -22880 -25480
rect -22620 -25500 -22380 -25480
rect -22120 -25500 -21880 -25480
rect -21620 -25500 -21500 -25480
rect -26500 -25700 -21500 -25500
rect -26500 -25720 -26380 -25700
rect -26120 -25720 -25880 -25700
rect -25620 -25720 -25380 -25700
rect -25120 -25720 -24880 -25700
rect -24620 -25720 -24380 -25700
rect -24120 -25720 -23880 -25700
rect -23620 -25720 -23380 -25700
rect -23120 -25720 -22880 -25700
rect -22620 -25720 -22380 -25700
rect -22120 -25720 -21880 -25700
rect -21620 -25720 -21500 -25700
rect -26500 -25980 -26400 -25720
rect -26100 -25980 -25900 -25720
rect -25600 -25980 -25400 -25720
rect -25100 -25980 -24900 -25720
rect -24600 -25980 -24400 -25720
rect -24100 -25980 -23900 -25720
rect -23600 -25980 -23400 -25720
rect -23100 -25980 -22900 -25720
rect -22600 -25980 -22400 -25720
rect -22100 -25980 -21900 -25720
rect -21600 -25980 -21500 -25720
rect -26500 -26000 -26380 -25980
rect -26120 -26000 -25880 -25980
rect -25620 -26000 -25380 -25980
rect -25120 -26000 -24880 -25980
rect -24620 -26000 -24380 -25980
rect -24120 -26000 -23880 -25980
rect -23620 -26000 -23380 -25980
rect -23120 -26000 -22880 -25980
rect -22620 -26000 -22380 -25980
rect -22120 -26000 -21880 -25980
rect -21620 -26000 -21500 -25980
rect -26500 -26200 -21500 -26000
rect -26500 -26220 -26380 -26200
rect -26120 -26220 -25880 -26200
rect -25620 -26220 -25380 -26200
rect -25120 -26220 -24880 -26200
rect -24620 -26220 -24380 -26200
rect -24120 -26220 -23880 -26200
rect -23620 -26220 -23380 -26200
rect -23120 -26220 -22880 -26200
rect -22620 -26220 -22380 -26200
rect -22120 -26220 -21880 -26200
rect -21620 -26220 -21500 -26200
rect -26500 -26480 -26400 -26220
rect -26100 -26480 -25900 -26220
rect -25600 -26480 -25400 -26220
rect -25100 -26480 -24900 -26220
rect -24600 -26480 -24400 -26220
rect -24100 -26480 -23900 -26220
rect -23600 -26480 -23400 -26220
rect -23100 -26480 -22900 -26220
rect -22600 -26480 -22400 -26220
rect -22100 -26480 -21900 -26220
rect -21600 -26480 -21500 -26220
rect -26500 -26500 -26380 -26480
rect -26120 -26500 -25880 -26480
rect -25620 -26500 -25380 -26480
rect -25120 -26500 -24880 -26480
rect -24620 -26500 -24380 -26480
rect -24120 -26500 -23880 -26480
rect -23620 -26500 -23380 -26480
rect -23120 -26500 -22880 -26480
rect -22620 -26500 -22380 -26480
rect -22120 -26500 -21880 -26480
rect -21620 -26500 -21500 -26480
rect -26500 -26700 -21500 -26500
rect -26500 -26720 -26380 -26700
rect -26120 -26720 -25880 -26700
rect -25620 -26720 -25380 -26700
rect -25120 -26720 -24880 -26700
rect -24620 -26720 -24380 -26700
rect -24120 -26720 -23880 -26700
rect -23620 -26720 -23380 -26700
rect -23120 -26720 -22880 -26700
rect -22620 -26720 -22380 -26700
rect -22120 -26720 -21880 -26700
rect -21620 -26720 -21500 -26700
rect -26500 -26980 -26400 -26720
rect -26100 -26980 -25900 -26720
rect -25600 -26980 -25400 -26720
rect -25100 -26980 -24900 -26720
rect -24600 -26980 -24400 -26720
rect -24100 -26980 -23900 -26720
rect -23600 -26980 -23400 -26720
rect -23100 -26980 -22900 -26720
rect -22600 -26980 -22400 -26720
rect -22100 -26980 -21900 -26720
rect -21600 -26980 -21500 -26720
rect -26500 -27000 -26380 -26980
rect -26120 -27000 -25880 -26980
rect -25620 -27000 -25380 -26980
rect -25120 -27000 -24880 -26980
rect -24620 -27000 -24380 -26980
rect -24120 -27000 -23880 -26980
rect -23620 -27000 -23380 -26980
rect -23120 -27000 -22880 -26980
rect -22620 -27000 -22380 -26980
rect -22120 -27000 -21880 -26980
rect -21620 -27000 -21500 -26980
rect -26500 -27200 -21500 -27000
rect -26500 -27220 -26380 -27200
rect -26120 -27220 -25880 -27200
rect -25620 -27220 -25380 -27200
rect -25120 -27220 -24880 -27200
rect -24620 -27220 -24380 -27200
rect -24120 -27220 -23880 -27200
rect -23620 -27220 -23380 -27200
rect -23120 -27220 -22880 -27200
rect -22620 -27220 -22380 -27200
rect -22120 -27220 -21880 -27200
rect -21620 -27220 -21500 -27200
rect -26500 -27480 -26400 -27220
rect -26100 -27480 -25900 -27220
rect -25600 -27480 -25400 -27220
rect -25100 -27480 -24900 -27220
rect -24600 -27480 -24400 -27220
rect -24100 -27480 -23900 -27220
rect -23600 -27480 -23400 -27220
rect -23100 -27480 -22900 -27220
rect -22600 -27480 -22400 -27220
rect -22100 -27480 -21900 -27220
rect -21600 -27480 -21500 -27220
rect -26500 -27500 -26380 -27480
rect -26120 -27500 -25880 -27480
rect -25620 -27500 -25380 -27480
rect -25120 -27500 -24880 -27480
rect -24620 -27500 -24380 -27480
rect -24120 -27500 -23880 -27480
rect -23620 -27500 -23380 -27480
rect -23120 -27500 -22880 -27480
rect -22620 -27500 -22380 -27480
rect -22120 -27500 -21880 -27480
rect -21620 -27500 -21500 -27480
rect -26500 -27700 -21500 -27500
rect -26500 -27720 -26380 -27700
rect -26120 -27720 -25880 -27700
rect -25620 -27720 -25380 -27700
rect -25120 -27720 -24880 -27700
rect -24620 -27720 -24380 -27700
rect -24120 -27720 -23880 -27700
rect -23620 -27720 -23380 -27700
rect -23120 -27720 -22880 -27700
rect -22620 -27720 -22380 -27700
rect -22120 -27720 -21880 -27700
rect -21620 -27720 -21500 -27700
rect -26500 -27980 -26400 -27720
rect -26100 -27980 -25900 -27720
rect -25600 -27980 -25400 -27720
rect -25100 -27980 -24900 -27720
rect -24600 -27980 -24400 -27720
rect -24100 -27980 -23900 -27720
rect -23600 -27980 -23400 -27720
rect -23100 -27980 -22900 -27720
rect -22600 -27980 -22400 -27720
rect -22100 -27980 -21900 -27720
rect -21600 -27980 -21500 -27720
rect -26500 -28000 -26380 -27980
rect -26120 -28000 -25880 -27980
rect -25620 -28000 -25380 -27980
rect -25120 -28000 -24880 -27980
rect -24620 -28000 -24380 -27980
rect -24120 -28000 -23880 -27980
rect -23620 -28000 -23380 -27980
rect -23120 -28000 -22880 -27980
rect -22620 -28000 -22380 -27980
rect -22120 -28000 -21880 -27980
rect -21620 -28000 -21500 -27980
rect -26500 -28200 -21500 -28000
rect -26500 -28220 -26380 -28200
rect -26120 -28220 -25880 -28200
rect -25620 -28220 -25380 -28200
rect -25120 -28220 -24880 -28200
rect -24620 -28220 -24380 -28200
rect -24120 -28220 -23880 -28200
rect -23620 -28220 -23380 -28200
rect -23120 -28220 -22880 -28200
rect -22620 -28220 -22380 -28200
rect -22120 -28220 -21880 -28200
rect -21620 -28220 -21500 -28200
rect -26500 -28480 -26400 -28220
rect -26100 -28480 -25900 -28220
rect -25600 -28480 -25400 -28220
rect -25100 -28480 -24900 -28220
rect -24600 -28480 -24400 -28220
rect -24100 -28480 -23900 -28220
rect -23600 -28480 -23400 -28220
rect -23100 -28480 -22900 -28220
rect -22600 -28480 -22400 -28220
rect -22100 -28480 -21900 -28220
rect -21600 -28480 -21500 -28220
rect -26500 -28500 -26380 -28480
rect -26120 -28500 -25880 -28480
rect -25620 -28500 -25380 -28480
rect -25120 -28500 -24880 -28480
rect -24620 -28500 -24380 -28480
rect -24120 -28500 -23880 -28480
rect -23620 -28500 -23380 -28480
rect -23120 -28500 -22880 -28480
rect -22620 -28500 -22380 -28480
rect -22120 -28500 -21880 -28480
rect -21620 -28500 -21500 -28480
rect -26500 -28700 -21500 -28500
rect -26500 -28720 -26380 -28700
rect -26120 -28720 -25880 -28700
rect -25620 -28720 -25380 -28700
rect -25120 -28720 -24880 -28700
rect -24620 -28720 -24380 -28700
rect -24120 -28720 -23880 -28700
rect -23620 -28720 -23380 -28700
rect -23120 -28720 -22880 -28700
rect -22620 -28720 -22380 -28700
rect -22120 -28720 -21880 -28700
rect -21620 -28720 -21500 -28700
rect -26500 -28980 -26400 -28720
rect -26100 -28980 -25900 -28720
rect -25600 -28980 -25400 -28720
rect -25100 -28980 -24900 -28720
rect -24600 -28980 -24400 -28720
rect -24100 -28980 -23900 -28720
rect -23600 -28980 -23400 -28720
rect -23100 -28980 -22900 -28720
rect -22600 -28980 -22400 -28720
rect -22100 -28980 -21900 -28720
rect -21600 -28980 -21500 -28720
rect -26500 -29000 -26380 -28980
rect -26120 -29000 -25880 -28980
rect -25620 -29000 -25380 -28980
rect -25120 -29000 -24880 -28980
rect -24620 -29000 -24380 -28980
rect -24120 -29000 -23880 -28980
rect -23620 -29000 -23380 -28980
rect -23120 -29000 -22880 -28980
rect -22620 -29000 -22380 -28980
rect -22120 -29000 -21880 -28980
rect -21620 -29000 -21500 -28980
rect -26500 -29200 -21500 -29000
rect 19500 -25200 20500 -25000
rect 19500 -25220 19620 -25200
rect 19880 -25220 20120 -25200
rect 20380 -25220 20500 -25200
rect 19500 -25480 19600 -25220
rect 19900 -25480 20100 -25220
rect 20400 -25480 20500 -25220
rect 19500 -25500 19620 -25480
rect 19880 -25500 20120 -25480
rect 20380 -25500 20500 -25480
rect 19500 -25700 20500 -25500
rect 19500 -25720 19620 -25700
rect 19880 -25720 20120 -25700
rect 20380 -25720 20500 -25700
rect 19500 -25980 19600 -25720
rect 19900 -25980 20100 -25720
rect 20400 -25980 20500 -25720
rect 19500 -26000 19620 -25980
rect 19880 -26000 20120 -25980
rect 20380 -26000 20500 -25980
rect 19500 -26200 20500 -26000
rect 19500 -26220 19620 -26200
rect 19880 -26220 20120 -26200
rect 20380 -26220 20500 -26200
rect 19500 -26480 19600 -26220
rect 19900 -26480 20100 -26220
rect 20400 -26480 20500 -26220
rect 19500 -26500 19620 -26480
rect 19880 -26500 20120 -26480
rect 20380 -26500 20500 -26480
rect 19500 -26700 20500 -26500
rect 19500 -26720 19620 -26700
rect 19880 -26720 20120 -26700
rect 20380 -26720 20500 -26700
rect 19500 -26980 19600 -26720
rect 19900 -26980 20100 -26720
rect 20400 -26980 20500 -26720
rect 19500 -27000 19620 -26980
rect 19880 -27000 20120 -26980
rect 20380 -27000 20500 -26980
rect 19500 -27200 20500 -27000
rect 19500 -27220 19620 -27200
rect 19880 -27220 20120 -27200
rect 20380 -27220 20500 -27200
rect 19500 -27480 19600 -27220
rect 19900 -27480 20100 -27220
rect 20400 -27480 20500 -27220
rect 19500 -27500 19620 -27480
rect 19880 -27500 20120 -27480
rect 20380 -27500 20500 -27480
rect 19500 -27700 20500 -27500
rect 19500 -27720 19620 -27700
rect 19880 -27720 20120 -27700
rect 20380 -27720 20500 -27700
rect 19500 -27980 19600 -27720
rect 19900 -27980 20100 -27720
rect 20400 -27980 20500 -27720
rect 19500 -28000 19620 -27980
rect 19880 -28000 20120 -27980
rect 20380 -28000 20500 -27980
rect 19500 -28100 20500 -28000
rect 23500 -20200 24000 -20000
rect 23500 -20220 23620 -20200
rect 23880 -20220 24000 -20200
rect 23500 -20480 23600 -20220
rect 23900 -20480 24000 -20220
rect 23500 -20500 23620 -20480
rect 23880 -20500 24000 -20480
rect 23500 -20700 24000 -20500
rect 23500 -20720 23620 -20700
rect 23880 -20720 24000 -20700
rect 23500 -20980 23600 -20720
rect 23900 -20980 24000 -20720
rect 23500 -21000 23620 -20980
rect 23880 -21000 24000 -20980
rect 23500 -21200 24000 -21000
rect 23500 -21220 23620 -21200
rect 23880 -21220 24000 -21200
rect 23500 -21480 23600 -21220
rect 23900 -21480 24000 -21220
rect 23500 -21500 23620 -21480
rect 23880 -21500 24000 -21480
rect 23500 -21700 24000 -21500
rect 23500 -21720 23620 -21700
rect 23880 -21720 24000 -21700
rect 23500 -21980 23600 -21720
rect 23900 -21980 24000 -21720
rect 23500 -22000 23620 -21980
rect 23880 -22000 24000 -21980
rect 23500 -22200 24000 -22000
rect 23500 -22220 23620 -22200
rect 23880 -22220 24000 -22200
rect 23500 -22480 23600 -22220
rect 23900 -22480 24000 -22220
rect 23500 -22500 23620 -22480
rect 23880 -22500 24000 -22480
rect 23500 -22700 24000 -22500
rect 23500 -22720 23620 -22700
rect 23880 -22720 24000 -22700
rect 23500 -22980 23600 -22720
rect 23900 -22980 24000 -22720
rect 23500 -23000 23620 -22980
rect 23880 -23000 24000 -22980
rect 23500 -23200 24000 -23000
rect 23500 -23220 23620 -23200
rect 23880 -23220 24000 -23200
rect 23500 -23480 23600 -23220
rect 23900 -23480 24000 -23220
rect 23500 -23500 23620 -23480
rect 23880 -23500 24000 -23480
rect 23500 -23700 24000 -23500
rect 23500 -23720 23620 -23700
rect 23880 -23720 24000 -23700
rect 23500 -23980 23600 -23720
rect 23900 -23980 24000 -23720
rect 23500 -24000 23620 -23980
rect 23880 -24000 24000 -23980
rect 23500 -24200 24000 -24000
rect 23500 -24220 23620 -24200
rect 23880 -24220 24000 -24200
rect 23500 -24480 23600 -24220
rect 23900 -24480 24000 -24220
rect 23500 -24500 23620 -24480
rect 23880 -24500 24000 -24480
rect 23500 -24700 24000 -24500
rect 23500 -24720 23620 -24700
rect 23880 -24720 24000 -24700
rect 23500 -24980 23600 -24720
rect 23900 -24980 24000 -24720
rect 23500 -25000 23620 -24980
rect 23880 -25000 24000 -24980
rect 23500 -25200 24000 -25000
rect 23500 -25220 23620 -25200
rect 23880 -25220 24000 -25200
rect 23500 -25480 23600 -25220
rect 23900 -25480 24000 -25220
rect 23500 -25500 23620 -25480
rect 23880 -25500 24000 -25480
rect 23500 -25700 24000 -25500
rect 23500 -25720 23620 -25700
rect 23880 -25720 24000 -25700
rect 23500 -25980 23600 -25720
rect 23900 -25980 24000 -25720
rect 23500 -26000 23620 -25980
rect 23880 -26000 24000 -25980
rect 23500 -26200 24000 -26000
rect 23500 -26220 23620 -26200
rect 23880 -26220 24000 -26200
rect 23500 -26480 23600 -26220
rect 23900 -26480 24000 -26220
rect 23500 -26500 23620 -26480
rect 23880 -26500 24000 -26480
rect 23500 -26700 24000 -26500
rect 23500 -26720 23620 -26700
rect 23880 -26720 24000 -26700
rect 23500 -26980 23600 -26720
rect 23900 -26980 24000 -26720
rect 23500 -27000 23620 -26980
rect 23880 -27000 24000 -26980
rect 23500 -27200 24000 -27000
rect 23500 -27220 23620 -27200
rect 23880 -27220 24000 -27200
rect 23500 -27480 23600 -27220
rect 23900 -27480 24000 -27220
rect 23500 -27500 23620 -27480
rect 23880 -27500 24000 -27480
rect 23500 -27700 24000 -27500
rect 23500 -27720 23620 -27700
rect 23880 -27720 24000 -27700
rect 23500 -27980 23600 -27720
rect 23900 -27980 24000 -27720
rect 23500 -28000 23620 -27980
rect 23880 -28000 24000 -27980
rect 19500 -28200 22500 -28100
rect 19500 -28220 19620 -28200
rect 19880 -28220 20120 -28200
rect 20380 -28220 20620 -28200
rect 20880 -28220 21120 -28200
rect 21380 -28220 21620 -28200
rect 21880 -28220 22120 -28200
rect 22380 -28220 22500 -28200
rect 19500 -28480 19600 -28220
rect 19900 -28480 20100 -28220
rect 20400 -28480 20600 -28220
rect 20900 -28480 21100 -28220
rect 21400 -28480 21600 -28220
rect 21900 -28480 22100 -28220
rect 22400 -28480 22500 -28220
rect 19500 -28500 19620 -28480
rect 19880 -28500 20120 -28480
rect 20380 -28500 20620 -28480
rect 20880 -28500 21120 -28480
rect 21380 -28500 21620 -28480
rect 21880 -28500 22120 -28480
rect 22380 -28500 22500 -28480
rect 19500 -28600 22500 -28500
rect 23500 -28200 24000 -28000
rect 32800 -5700 33500 -5600
rect 32800 -5720 33120 -5700
rect 33380 -5720 33500 -5700
rect 32800 -5980 33100 -5720
rect 33400 -5980 33500 -5720
rect 32800 -6000 33120 -5980
rect 33380 -6000 33500 -5980
rect 32800 -6200 33500 -6000
rect 32800 -6220 33120 -6200
rect 33380 -6220 33500 -6200
rect 32800 -6480 33100 -6220
rect 33400 -6480 33500 -6220
rect 32800 -6500 33120 -6480
rect 33380 -6500 33500 -6480
rect 32800 -6700 33500 -6500
rect 32800 -6720 33120 -6700
rect 33380 -6720 33500 -6700
rect 32800 -6980 33100 -6720
rect 33400 -6980 33500 -6720
rect 32800 -7000 33120 -6980
rect 33380 -7000 33500 -6980
rect 32800 -7200 33500 -7000
rect 32800 -7220 33120 -7200
rect 33380 -7220 33500 -7200
rect 32800 -7480 33100 -7220
rect 33400 -7480 33500 -7220
rect 32800 -7500 33120 -7480
rect 33380 -7500 33500 -7480
rect 32800 -7700 33500 -7500
rect 32800 -7720 33120 -7700
rect 33380 -7720 33500 -7700
rect 32800 -7980 33100 -7720
rect 33400 -7980 33500 -7720
rect 32800 -8000 33120 -7980
rect 33380 -8000 33500 -7980
rect 32800 -8200 33500 -8000
rect 32800 -8220 33120 -8200
rect 33380 -8220 33500 -8200
rect 32800 -8480 33100 -8220
rect 33400 -8480 33500 -8220
rect 32800 -8500 33120 -8480
rect 33380 -8500 33500 -8480
rect 32800 -8700 33500 -8500
rect 32800 -8720 33120 -8700
rect 33380 -8720 33500 -8700
rect 32800 -8980 33100 -8720
rect 33400 -8980 33500 -8720
rect 32800 -9000 33120 -8980
rect 33380 -9000 33500 -8980
rect 32800 -9200 33500 -9000
rect 32800 -9220 33120 -9200
rect 33380 -9220 33500 -9200
rect 32800 -9480 33100 -9220
rect 33400 -9480 33500 -9220
rect 32800 -9500 33120 -9480
rect 33380 -9500 33500 -9480
rect 32800 -9700 33500 -9500
rect 32800 -9720 33120 -9700
rect 33380 -9720 33500 -9700
rect 32800 -9980 33100 -9720
rect 33400 -9980 33500 -9720
rect 32800 -10000 33120 -9980
rect 33380 -10000 33500 -9980
rect 32800 -10200 33500 -10000
rect 32800 -10220 33120 -10200
rect 33380 -10220 33500 -10200
rect 32800 -10480 33100 -10220
rect 33400 -10480 33500 -10220
rect 32800 -10500 33120 -10480
rect 33380 -10500 33500 -10480
rect 32800 -10700 33500 -10500
rect 32800 -10720 33120 -10700
rect 33380 -10720 33500 -10700
rect 32800 -10980 33100 -10720
rect 33400 -10980 33500 -10720
rect 32800 -11000 33120 -10980
rect 33380 -11000 33500 -10980
rect 32800 -11200 33500 -11000
rect 32800 -11220 33120 -11200
rect 33380 -11220 33500 -11200
rect 32800 -11480 33100 -11220
rect 33400 -11480 33500 -11220
rect 32800 -11500 33120 -11480
rect 33380 -11500 33500 -11480
rect 32800 -11700 33500 -11500
rect 32800 -11720 33120 -11700
rect 33380 -11720 33500 -11700
rect 32800 -11980 33100 -11720
rect 33400 -11980 33500 -11720
rect 32800 -12000 33120 -11980
rect 33380 -12000 33500 -11980
rect 32800 -12200 33500 -12000
rect 32800 -12220 33120 -12200
rect 33380 -12220 33500 -12200
rect 32800 -12480 33100 -12220
rect 33400 -12480 33500 -12220
rect 32800 -12500 33120 -12480
rect 33380 -12500 33500 -12480
rect 32800 -12700 33500 -12500
rect 32800 -12720 33120 -12700
rect 33380 -12720 33500 -12700
rect 32800 -12980 33100 -12720
rect 33400 -12980 33500 -12720
rect 32800 -13000 33120 -12980
rect 33380 -13000 33500 -12980
rect 32800 -13200 33500 -13000
rect 32800 -13220 33120 -13200
rect 33380 -13220 33500 -13200
rect 32800 -13480 33100 -13220
rect 33400 -13480 33500 -13220
rect 32800 -13500 33120 -13480
rect 33380 -13500 33500 -13480
rect 32800 -13700 33500 -13500
rect 32800 -13720 33120 -13700
rect 33380 -13720 33500 -13700
rect 32800 -13980 33100 -13720
rect 33400 -13980 33500 -13720
rect 32800 -14000 33120 -13980
rect 33380 -14000 33500 -13980
rect 32800 -14200 33500 -14000
rect 32800 -14220 33120 -14200
rect 33380 -14220 33500 -14200
rect 32800 -14480 33100 -14220
rect 33400 -14480 33500 -14220
rect 32800 -14500 33120 -14480
rect 33380 -14500 33500 -14480
rect 32800 -14700 33500 -14500
rect 32800 -14720 33120 -14700
rect 33380 -14720 33500 -14700
rect 32800 -14980 33100 -14720
rect 33400 -14980 33500 -14720
rect 32800 -15000 33120 -14980
rect 33380 -15000 33500 -14980
rect 32800 -15200 33500 -15000
rect 32800 -15220 33120 -15200
rect 33380 -15220 33500 -15200
rect 32800 -15480 33100 -15220
rect 33400 -15480 33500 -15220
rect 32800 -15500 33120 -15480
rect 33380 -15500 33500 -15480
rect 32800 -15700 33500 -15500
rect 32800 -15720 33120 -15700
rect 33380 -15720 33500 -15700
rect 32800 -15980 33100 -15720
rect 33400 -15980 33500 -15720
rect 32800 -16000 33120 -15980
rect 33380 -16000 33500 -15980
rect 32800 -16200 33500 -16000
rect 32800 -16220 33120 -16200
rect 33380 -16220 33500 -16200
rect 32800 -16480 33100 -16220
rect 33400 -16480 33500 -16220
rect 32800 -16500 33120 -16480
rect 33380 -16500 33500 -16480
rect 32800 -16700 33500 -16500
rect 32800 -16720 33120 -16700
rect 33380 -16720 33500 -16700
rect 32800 -16980 33100 -16720
rect 33400 -16980 33500 -16720
rect 32800 -17000 33120 -16980
rect 33380 -17000 33500 -16980
rect 32800 -17200 33500 -17000
rect 32800 -17220 33120 -17200
rect 33380 -17220 33500 -17200
rect 32800 -17480 33100 -17220
rect 33400 -17480 33500 -17220
rect 32800 -17500 33120 -17480
rect 33380 -17500 33500 -17480
rect 32800 -17700 33500 -17500
rect 32800 -17720 33120 -17700
rect 33380 -17720 33500 -17700
rect 32800 -17980 33100 -17720
rect 33400 -17980 33500 -17720
rect 32800 -18000 33120 -17980
rect 33380 -18000 33500 -17980
rect 32800 -18200 33500 -18000
rect 32800 -18220 33120 -18200
rect 33380 -18220 33500 -18200
rect 32800 -18480 33100 -18220
rect 33400 -18480 33500 -18220
rect 32800 -18500 33120 -18480
rect 33380 -18500 33500 -18480
rect 32800 -18700 33500 -18500
rect 32800 -18720 33120 -18700
rect 33380 -18720 33500 -18700
rect 32800 -18980 33100 -18720
rect 33400 -18980 33500 -18720
rect 32800 -19000 33120 -18980
rect 33380 -19000 33500 -18980
rect 32800 -19200 33500 -19000
rect 32800 -19220 33120 -19200
rect 33380 -19220 33500 -19200
rect 32800 -19480 33100 -19220
rect 33400 -19480 33500 -19220
rect 32800 -19500 33120 -19480
rect 33380 -19500 33500 -19480
rect 32800 -19700 33500 -19500
rect 32800 -19720 33120 -19700
rect 33380 -19720 33500 -19700
rect 32800 -19980 33100 -19720
rect 33400 -19980 33500 -19720
rect 32800 -20000 33120 -19980
rect 33380 -20000 33500 -19980
rect 32800 -20100 33500 -20000
rect 140500 -12200 143500 -12100
rect 140500 -12220 140620 -12200
rect 140880 -12220 141120 -12200
rect 141380 -12220 141620 -12200
rect 141880 -12220 142120 -12200
rect 142380 -12220 142620 -12200
rect 142880 -12220 143120 -12200
rect 143380 -12220 143500 -12200
rect 140500 -12480 140600 -12220
rect 140900 -12480 141100 -12220
rect 141400 -12480 141600 -12220
rect 141900 -12480 142100 -12220
rect 142400 -12480 142600 -12220
rect 142900 -12480 143100 -12220
rect 143400 -12480 143500 -12220
rect 140500 -12500 140620 -12480
rect 140880 -12500 141120 -12480
rect 141380 -12500 141620 -12480
rect 141880 -12500 142120 -12480
rect 142380 -12500 142620 -12480
rect 142880 -12500 143120 -12480
rect 143380 -12500 143500 -12480
rect 140500 -12700 143500 -12500
rect 140500 -12720 140620 -12700
rect 140880 -12720 141120 -12700
rect 141380 -12720 141620 -12700
rect 141880 -12720 142120 -12700
rect 142380 -12720 142620 -12700
rect 142880 -12720 143120 -12700
rect 143380 -12720 143500 -12700
rect 140500 -12980 140600 -12720
rect 140900 -12980 141100 -12720
rect 141400 -12980 141600 -12720
rect 141900 -12980 142100 -12720
rect 142400 -12980 142600 -12720
rect 142900 -12980 143100 -12720
rect 143400 -12980 143500 -12720
rect 140500 -13000 140620 -12980
rect 140880 -13000 141120 -12980
rect 141380 -13000 141620 -12980
rect 141880 -13000 142120 -12980
rect 142380 -13000 142620 -12980
rect 142880 -13000 143120 -12980
rect 143380 -13000 143500 -12980
rect 140500 -13200 143500 -13000
rect 140500 -13220 140620 -13200
rect 140880 -13220 141120 -13200
rect 141380 -13220 141620 -13200
rect 141880 -13220 142120 -13200
rect 142380 -13220 142620 -13200
rect 142880 -13220 143120 -13200
rect 143380 -13220 143500 -13200
rect 140500 -13480 140600 -13220
rect 140900 -13480 141100 -13220
rect 141400 -13480 141600 -13220
rect 141900 -13480 142100 -13220
rect 142400 -13480 142600 -13220
rect 142900 -13480 143100 -13220
rect 143400 -13480 143500 -13220
rect 140500 -13500 140620 -13480
rect 140880 -13500 141120 -13480
rect 141380 -13500 141620 -13480
rect 141880 -13500 142120 -13480
rect 142380 -13500 142620 -13480
rect 142880 -13500 143120 -13480
rect 143380 -13500 143500 -13480
rect 140500 -13700 143500 -13500
rect 140500 -13720 140620 -13700
rect 140880 -13720 141120 -13700
rect 141380 -13720 141620 -13700
rect 141880 -13720 142120 -13700
rect 142380 -13720 142620 -13700
rect 142880 -13720 143120 -13700
rect 143380 -13720 143500 -13700
rect 140500 -13980 140600 -13720
rect 140900 -13980 141100 -13720
rect 141400 -13980 141600 -13720
rect 141900 -13980 142100 -13720
rect 142400 -13980 142600 -13720
rect 142900 -13980 143100 -13720
rect 143400 -13980 143500 -13720
rect 140500 -14000 140620 -13980
rect 140880 -14000 141120 -13980
rect 141380 -14000 141620 -13980
rect 141880 -14000 142120 -13980
rect 142380 -14000 142620 -13980
rect 142880 -14000 143120 -13980
rect 143380 -14000 143500 -13980
rect 140500 -14200 143500 -14000
rect 140500 -14220 140620 -14200
rect 140880 -14220 141120 -14200
rect 141380 -14220 141620 -14200
rect 141880 -14220 142120 -14200
rect 142380 -14220 142620 -14200
rect 142880 -14220 143120 -14200
rect 143380 -14220 143500 -14200
rect 140500 -14480 140600 -14220
rect 140900 -14480 141100 -14220
rect 141400 -14480 141600 -14220
rect 141900 -14480 142100 -14220
rect 142400 -14480 142600 -14220
rect 142900 -14480 143100 -14220
rect 143400 -14480 143500 -14220
rect 140500 -14500 140620 -14480
rect 140880 -14500 141120 -14480
rect 141380 -14500 141620 -14480
rect 141880 -14500 142120 -14480
rect 142380 -14500 142620 -14480
rect 142880 -14500 143120 -14480
rect 143380 -14500 143500 -14480
rect 140500 -14700 143500 -14500
rect 140500 -14720 140620 -14700
rect 140880 -14720 141120 -14700
rect 141380 -14720 141620 -14700
rect 141880 -14720 142120 -14700
rect 142380 -14720 142620 -14700
rect 142880 -14720 143120 -14700
rect 143380 -14720 143500 -14700
rect 140500 -14980 140600 -14720
rect 140900 -14980 141100 -14720
rect 141400 -14980 141600 -14720
rect 141900 -14980 142100 -14720
rect 142400 -14980 142600 -14720
rect 142900 -14980 143100 -14720
rect 143400 -14980 143500 -14720
rect 140500 -15000 140620 -14980
rect 140880 -15000 141120 -14980
rect 141380 -15000 141620 -14980
rect 141880 -15000 142120 -14980
rect 142380 -15000 142620 -14980
rect 142880 -15000 143120 -14980
rect 143380 -15000 143500 -14980
rect 140500 -15200 143500 -15000
rect 140500 -15220 140620 -15200
rect 140880 -15220 141120 -15200
rect 141380 -15220 141620 -15200
rect 141880 -15220 142120 -15200
rect 142380 -15220 142620 -15200
rect 142880 -15220 143120 -15200
rect 143380 -15220 143500 -15200
rect 140500 -15480 140600 -15220
rect 140900 -15480 141100 -15220
rect 141400 -15480 141600 -15220
rect 141900 -15480 142100 -15220
rect 142400 -15480 142600 -15220
rect 142900 -15480 143100 -15220
rect 143400 -15480 143500 -15220
rect 140500 -15500 140620 -15480
rect 140880 -15500 141120 -15480
rect 141380 -15500 141620 -15480
rect 141880 -15500 142120 -15480
rect 142380 -15500 142620 -15480
rect 142880 -15500 143120 -15480
rect 143380 -15500 143500 -15480
rect 140500 -15700 143500 -15500
rect 140500 -15720 140620 -15700
rect 140880 -15720 141120 -15700
rect 141380 -15720 141620 -15700
rect 141880 -15720 142120 -15700
rect 142380 -15720 142620 -15700
rect 142880 -15720 143120 -15700
rect 143380 -15720 143500 -15700
rect 140500 -15980 140600 -15720
rect 140900 -15980 141100 -15720
rect 141400 -15980 141600 -15720
rect 141900 -15980 142100 -15720
rect 142400 -15980 142600 -15720
rect 142900 -15980 143100 -15720
rect 143400 -15980 143500 -15720
rect 140500 -16000 140620 -15980
rect 140880 -16000 141120 -15980
rect 141380 -16000 141620 -15980
rect 141880 -16000 142120 -15980
rect 142380 -16000 142620 -15980
rect 142880 -16000 143120 -15980
rect 143380 -16000 143500 -15980
rect 140500 -16200 143500 -16000
rect 140500 -16220 140620 -16200
rect 140880 -16220 141120 -16200
rect 141380 -16220 141620 -16200
rect 141880 -16220 142120 -16200
rect 142380 -16220 142620 -16200
rect 142880 -16220 143120 -16200
rect 143380 -16220 143500 -16200
rect 140500 -16480 140600 -16220
rect 140900 -16480 141100 -16220
rect 141400 -16480 141600 -16220
rect 141900 -16480 142100 -16220
rect 142400 -16480 142600 -16220
rect 142900 -16480 143100 -16220
rect 143400 -16480 143500 -16220
rect 140500 -16500 140620 -16480
rect 140880 -16500 141120 -16480
rect 141380 -16500 141620 -16480
rect 141880 -16500 142120 -16480
rect 142380 -16500 142620 -16480
rect 142880 -16500 143120 -16480
rect 143380 -16500 143500 -16480
rect 140500 -16700 143500 -16500
rect 140500 -16720 140620 -16700
rect 140880 -16720 141120 -16700
rect 141380 -16720 141620 -16700
rect 141880 -16720 142120 -16700
rect 142380 -16720 142620 -16700
rect 142880 -16720 143120 -16700
rect 143380 -16720 143500 -16700
rect 140500 -16980 140600 -16720
rect 140900 -16980 141100 -16720
rect 141400 -16980 141600 -16720
rect 141900 -16980 142100 -16720
rect 142400 -16980 142600 -16720
rect 142900 -16980 143100 -16720
rect 143400 -16980 143500 -16720
rect 140500 -17000 140620 -16980
rect 140880 -17000 141120 -16980
rect 141380 -17000 141620 -16980
rect 141880 -17000 142120 -16980
rect 142380 -17000 142620 -16980
rect 142880 -17000 143120 -16980
rect 143380 -17000 143500 -16980
rect 140500 -17200 143500 -17000
rect 140500 -17220 140620 -17200
rect 140880 -17220 141120 -17200
rect 141380 -17220 141620 -17200
rect 141880 -17220 142120 -17200
rect 142380 -17220 142620 -17200
rect 142880 -17220 143120 -17200
rect 143380 -17220 143500 -17200
rect 140500 -17480 140600 -17220
rect 140900 -17480 141100 -17220
rect 141400 -17480 141600 -17220
rect 141900 -17480 142100 -17220
rect 142400 -17480 142600 -17220
rect 142900 -17480 143100 -17220
rect 143400 -17480 143500 -17220
rect 140500 -17500 140620 -17480
rect 140880 -17500 141120 -17480
rect 141380 -17500 141620 -17480
rect 141880 -17500 142120 -17480
rect 142380 -17500 142620 -17480
rect 142880 -17500 143120 -17480
rect 143380 -17500 143500 -17480
rect 140500 -17700 143500 -17500
rect 140500 -17720 140620 -17700
rect 140880 -17720 141120 -17700
rect 141380 -17720 141620 -17700
rect 141880 -17720 142120 -17700
rect 142380 -17720 142620 -17700
rect 142880 -17720 143120 -17700
rect 143380 -17720 143500 -17700
rect 140500 -17980 140600 -17720
rect 140900 -17980 141100 -17720
rect 141400 -17980 141600 -17720
rect 141900 -17980 142100 -17720
rect 142400 -17980 142600 -17720
rect 142900 -17980 143100 -17720
rect 143400 -17980 143500 -17720
rect 140500 -18000 140620 -17980
rect 140880 -18000 141120 -17980
rect 141380 -18000 141620 -17980
rect 141880 -18000 142120 -17980
rect 142380 -18000 142620 -17980
rect 142880 -18000 143120 -17980
rect 143380 -18000 143500 -17980
rect 140500 -18200 143500 -18000
rect 140500 -18220 140620 -18200
rect 140880 -18220 141120 -18200
rect 141380 -18220 141620 -18200
rect 141880 -18220 142120 -18200
rect 142380 -18220 142620 -18200
rect 142880 -18220 143120 -18200
rect 143380 -18220 143500 -18200
rect 140500 -18480 140600 -18220
rect 140900 -18480 141100 -18220
rect 141400 -18480 141600 -18220
rect 141900 -18480 142100 -18220
rect 142400 -18480 142600 -18220
rect 142900 -18480 143100 -18220
rect 143400 -18480 143500 -18220
rect 140500 -18500 140620 -18480
rect 140880 -18500 141120 -18480
rect 141380 -18500 141620 -18480
rect 141880 -18500 142120 -18480
rect 142380 -18500 142620 -18480
rect 142880 -18500 143120 -18480
rect 143380 -18500 143500 -18480
rect 140500 -18700 143500 -18500
rect 140500 -18720 140620 -18700
rect 140880 -18720 141120 -18700
rect 141380 -18720 141620 -18700
rect 141880 -18720 142120 -18700
rect 142380 -18720 142620 -18700
rect 142880 -18720 143120 -18700
rect 143380 -18720 143500 -18700
rect 140500 -18980 140600 -18720
rect 140900 -18980 141100 -18720
rect 141400 -18980 141600 -18720
rect 141900 -18980 142100 -18720
rect 142400 -18980 142600 -18720
rect 142900 -18980 143100 -18720
rect 143400 -18980 143500 -18720
rect 140500 -19000 140620 -18980
rect 140880 -19000 141120 -18980
rect 141380 -19000 141620 -18980
rect 141880 -19000 142120 -18980
rect 142380 -19000 142620 -18980
rect 142880 -19000 143120 -18980
rect 143380 -19000 143500 -18980
rect 140500 -19200 143500 -19000
rect 140500 -19220 140620 -19200
rect 140880 -19220 141120 -19200
rect 141380 -19220 141620 -19200
rect 141880 -19220 142120 -19200
rect 142380 -19220 142620 -19200
rect 142880 -19220 143120 -19200
rect 143380 -19220 143500 -19200
rect 140500 -19480 140600 -19220
rect 140900 -19480 141100 -19220
rect 141400 -19480 141600 -19220
rect 141900 -19480 142100 -19220
rect 142400 -19480 142600 -19220
rect 142900 -19480 143100 -19220
rect 143400 -19480 143500 -19220
rect 140500 -19500 140620 -19480
rect 140880 -19500 141120 -19480
rect 141380 -19500 141620 -19480
rect 141880 -19500 142120 -19480
rect 142380 -19500 142620 -19480
rect 142880 -19500 143120 -19480
rect 143380 -19500 143500 -19480
rect 140500 -19700 143500 -19500
rect 140500 -19720 140620 -19700
rect 140880 -19720 141120 -19700
rect 141380 -19720 141620 -19700
rect 141880 -19720 142120 -19700
rect 142380 -19720 142620 -19700
rect 142880 -19720 143120 -19700
rect 143380 -19720 143500 -19700
rect 140500 -19980 140600 -19720
rect 140900 -19980 141100 -19720
rect 141400 -19980 141600 -19720
rect 141900 -19980 142100 -19720
rect 142400 -19980 142600 -19720
rect 142900 -19980 143100 -19720
rect 143400 -19980 143500 -19720
rect 140500 -20000 140620 -19980
rect 140880 -20000 141120 -19980
rect 141380 -20000 141620 -19980
rect 141880 -20000 142120 -19980
rect 142380 -20000 142620 -19980
rect 142880 -20000 143120 -19980
rect 143380 -20000 143500 -19980
rect 140500 -20100 143500 -20000
rect 32800 -20200 34500 -20100
rect 32800 -20220 33120 -20200
rect 33380 -20220 33620 -20200
rect 33880 -20220 34120 -20200
rect 34380 -20220 34500 -20200
rect 32800 -20480 33100 -20220
rect 33400 -20480 33600 -20220
rect 33900 -20480 34100 -20220
rect 34400 -20480 34500 -20220
rect 32800 -20500 33120 -20480
rect 33380 -20500 33620 -20480
rect 33880 -20500 34120 -20480
rect 34380 -20500 34500 -20480
rect 32800 -20700 34500 -20500
rect 32800 -20720 33120 -20700
rect 33380 -20720 33620 -20700
rect 33880 -20720 34120 -20700
rect 34380 -20720 34500 -20700
rect 32800 -20980 33100 -20720
rect 33400 -20980 33600 -20720
rect 33900 -20980 34100 -20720
rect 34400 -20980 34500 -20720
rect 32800 -21000 33120 -20980
rect 33380 -21000 33620 -20980
rect 33880 -21000 34120 -20980
rect 34380 -21000 34500 -20980
rect 32800 -21200 34500 -21000
rect 32800 -21220 33120 -21200
rect 33380 -21220 33620 -21200
rect 33880 -21220 34120 -21200
rect 34380 -21220 34500 -21200
rect 32800 -21480 33100 -21220
rect 33400 -21480 33600 -21220
rect 33900 -21480 34100 -21220
rect 34400 -21480 34500 -21220
rect 32800 -21500 33120 -21480
rect 33380 -21500 33620 -21480
rect 33880 -21500 34120 -21480
rect 34380 -21500 34500 -21480
rect 32800 -21700 34500 -21500
rect 32800 -21720 33120 -21700
rect 33380 -21720 33620 -21700
rect 33880 -21720 34120 -21700
rect 34380 -21720 34500 -21700
rect 32800 -21980 33100 -21720
rect 33400 -21980 33600 -21720
rect 33900 -21980 34100 -21720
rect 34400 -21980 34500 -21720
rect 32800 -22000 33120 -21980
rect 33380 -22000 33620 -21980
rect 33880 -22000 34120 -21980
rect 34380 -22000 34500 -21980
rect 32800 -22200 34500 -22000
rect 32800 -22220 33120 -22200
rect 33380 -22220 33620 -22200
rect 33880 -22220 34120 -22200
rect 34380 -22220 34500 -22200
rect 32800 -22480 33100 -22220
rect 33400 -22480 33600 -22220
rect 33900 -22480 34100 -22220
rect 34400 -22480 34500 -22220
rect 32800 -22500 33120 -22480
rect 33380 -22500 33620 -22480
rect 33880 -22500 34120 -22480
rect 34380 -22500 34500 -22480
rect 32800 -22700 34500 -22500
rect 32800 -22720 33120 -22700
rect 33380 -22720 33620 -22700
rect 33880 -22720 34120 -22700
rect 34380 -22720 34500 -22700
rect 32800 -22980 33100 -22720
rect 33400 -22980 33600 -22720
rect 33900 -22980 34100 -22720
rect 34400 -22980 34500 -22720
rect 32800 -23000 33120 -22980
rect 33380 -23000 33620 -22980
rect 33880 -23000 34120 -22980
rect 34380 -23000 34500 -22980
rect 32800 -23200 34500 -23000
rect 32800 -23220 33120 -23200
rect 33380 -23220 33620 -23200
rect 33880 -23220 34120 -23200
rect 34380 -23220 34500 -23200
rect 32800 -23480 33100 -23220
rect 33400 -23480 33600 -23220
rect 33900 -23480 34100 -23220
rect 34400 -23480 34500 -23220
rect 32800 -23500 33120 -23480
rect 33380 -23500 33620 -23480
rect 33880 -23500 34120 -23480
rect 34380 -23500 34500 -23480
rect 32800 -23700 34500 -23500
rect 32800 -23720 33120 -23700
rect 33380 -23720 33620 -23700
rect 33880 -23720 34120 -23700
rect 34380 -23720 34500 -23700
rect 32800 -23980 33100 -23720
rect 33400 -23980 33600 -23720
rect 33900 -23980 34100 -23720
rect 34400 -23980 34500 -23720
rect 32800 -24000 33120 -23980
rect 33380 -24000 33620 -23980
rect 33880 -24000 34120 -23980
rect 34380 -24000 34500 -23980
rect 32800 -24200 34500 -24000
rect 32800 -24220 33120 -24200
rect 33380 -24220 33620 -24200
rect 33880 -24220 34120 -24200
rect 34380 -24220 34500 -24200
rect 32800 -24480 33100 -24220
rect 33400 -24480 33600 -24220
rect 33900 -24480 34100 -24220
rect 34400 -24480 34500 -24220
rect 32800 -24500 33120 -24480
rect 33380 -24500 33620 -24480
rect 33880 -24500 34120 -24480
rect 34380 -24500 34500 -24480
rect 32800 -24700 34500 -24500
rect 32800 -24720 33120 -24700
rect 33380 -24720 33620 -24700
rect 33880 -24720 34120 -24700
rect 34380 -24720 34500 -24700
rect 32800 -24980 33100 -24720
rect 33400 -24980 33600 -24720
rect 33900 -24980 34100 -24720
rect 34400 -24980 34500 -24720
rect 32800 -25000 33120 -24980
rect 33380 -25000 33620 -24980
rect 33880 -25000 34120 -24980
rect 34380 -25000 34500 -24980
rect 32800 -25200 34500 -25000
rect 32800 -25220 33120 -25200
rect 33380 -25220 33620 -25200
rect 33880 -25220 34120 -25200
rect 34380 -25220 34500 -25200
rect 32800 -25480 33100 -25220
rect 33400 -25480 33600 -25220
rect 33900 -25480 34100 -25220
rect 34400 -25480 34500 -25220
rect 32800 -25500 33120 -25480
rect 33380 -25500 33620 -25480
rect 33880 -25500 34120 -25480
rect 34380 -25500 34500 -25480
rect 32800 -25700 34500 -25500
rect 32800 -25720 33120 -25700
rect 33380 -25720 33620 -25700
rect 33880 -25720 34120 -25700
rect 34380 -25720 34500 -25700
rect 32800 -25980 33100 -25720
rect 33400 -25980 33600 -25720
rect 33900 -25980 34100 -25720
rect 34400 -25980 34500 -25720
rect 32800 -26000 33120 -25980
rect 33380 -26000 33620 -25980
rect 33880 -26000 34120 -25980
rect 34380 -26000 34500 -25980
rect 32800 -26200 34500 -26000
rect 32800 -26220 33120 -26200
rect 33380 -26220 33620 -26200
rect 33880 -26220 34120 -26200
rect 34380 -26220 34500 -26200
rect 32800 -26480 33100 -26220
rect 33400 -26480 33600 -26220
rect 33900 -26480 34100 -26220
rect 34400 -26480 34500 -26220
rect 32800 -26500 33120 -26480
rect 33380 -26500 33620 -26480
rect 33880 -26500 34120 -26480
rect 34380 -26500 34500 -26480
rect 32800 -26700 34500 -26500
rect 32800 -26720 33120 -26700
rect 33380 -26720 33620 -26700
rect 33880 -26720 34120 -26700
rect 34380 -26720 34500 -26700
rect 32800 -26980 33100 -26720
rect 33400 -26980 33600 -26720
rect 33900 -26980 34100 -26720
rect 34400 -26980 34500 -26720
rect 32800 -27000 33120 -26980
rect 33380 -27000 33620 -26980
rect 33880 -27000 34120 -26980
rect 34380 -27000 34500 -26980
rect 32800 -27200 34500 -27000
rect 32800 -27220 33120 -27200
rect 33380 -27220 33620 -27200
rect 33880 -27220 34120 -27200
rect 34380 -27220 34500 -27200
rect 32800 -27480 33100 -27220
rect 33400 -27480 33600 -27220
rect 33900 -27480 34100 -27220
rect 34400 -27480 34500 -27220
rect 32800 -27500 33120 -27480
rect 33380 -27500 33620 -27480
rect 33880 -27500 34120 -27480
rect 34380 -27500 34500 -27480
rect 32800 -27700 34500 -27500
rect 32800 -27720 33120 -27700
rect 33380 -27720 33620 -27700
rect 33880 -27720 34120 -27700
rect 34380 -27720 34500 -27700
rect 32800 -27980 33100 -27720
rect 33400 -27980 33600 -27720
rect 33900 -27980 34100 -27720
rect 34400 -27980 34500 -27720
rect 32800 -28000 33120 -27980
rect 33380 -28000 33620 -27980
rect 33880 -28000 34120 -27980
rect 34380 -28000 34500 -27980
rect 32800 -28100 34500 -28000
rect 32800 -28200 36500 -28100
rect 23500 -28220 23620 -28200
rect 23880 -28220 26000 -28200
rect 23500 -28480 23600 -28220
rect 23900 -28480 26000 -28220
rect 23500 -28500 23620 -28480
rect 23880 -28500 26000 -28480
rect 23500 -28600 26000 -28500
rect 19500 -28700 26000 -28600
rect 19500 -28720 19620 -28700
rect 19880 -28720 20120 -28700
rect 20380 -28720 20620 -28700
rect 20880 -28720 21120 -28700
rect 21380 -28720 21620 -28700
rect 21880 -28720 22120 -28700
rect 22380 -28720 22620 -28700
rect 22880 -28720 23120 -28700
rect 23380 -28720 23620 -28700
rect 23880 -28720 26000 -28700
rect 19500 -28980 19600 -28720
rect 19900 -28980 20100 -28720
rect 20400 -28980 20600 -28720
rect 20900 -28980 21100 -28720
rect 21400 -28980 21600 -28720
rect 21900 -28980 22100 -28720
rect 22400 -28980 22600 -28720
rect 22900 -28980 23100 -28720
rect 23400 -28980 23600 -28720
rect 23900 -28980 26000 -28720
rect 19500 -29000 19620 -28980
rect 19880 -29000 20120 -28980
rect 20380 -29000 20620 -28980
rect 20880 -29000 21120 -28980
rect 21380 -29000 21620 -28980
rect 21880 -29000 22120 -28980
rect 22380 -29000 22620 -28980
rect 22880 -29000 23120 -28980
rect 23380 -29000 23620 -28980
rect 23880 -29000 26000 -28980
rect 19500 -29100 26000 -29000
rect -26500 -29220 -26380 -29200
rect -26120 -29220 -25880 -29200
rect -25620 -29220 -25380 -29200
rect -25120 -29220 -24880 -29200
rect -24620 -29220 -24380 -29200
rect -24120 -29220 -23880 -29200
rect -23620 -29220 -23380 -29200
rect -23120 -29220 -22880 -29200
rect -22620 -29220 -22380 -29200
rect -22120 -29220 -21880 -29200
rect -21620 -29220 -21500 -29200
rect -26500 -29480 -26400 -29220
rect -26100 -29480 -25900 -29220
rect -25600 -29480 -25400 -29220
rect -25100 -29480 -24900 -29220
rect -24600 -29480 -24400 -29220
rect -24100 -29480 -23900 -29220
rect -23600 -29480 -23400 -29220
rect -23100 -29480 -22900 -29220
rect -22600 -29480 -22400 -29220
rect -22100 -29480 -21900 -29220
rect -21600 -29480 -21500 -29220
rect -26500 -29500 -26380 -29480
rect -26120 -29500 -25880 -29480
rect -25620 -29500 -25380 -29480
rect -25120 -29500 -24880 -29480
rect -24620 -29500 -24380 -29480
rect -24120 -29500 -23880 -29480
rect -23620 -29500 -23380 -29480
rect -23120 -29500 -22880 -29480
rect -22620 -29500 -22380 -29480
rect -22120 -29500 -21880 -29480
rect -21620 -29500 -21500 -29480
rect -26500 -29600 -21500 -29500
rect 22500 -29120 26000 -29100
rect 22500 -29190 22650 -29120
rect 22850 -29190 23150 -29120
rect 23350 -29190 26000 -29120
rect 22500 -29200 26000 -29190
rect 22500 -29220 22620 -29200
rect 22880 -29220 23120 -29200
rect 23380 -29220 23620 -29200
rect 23880 -29220 26000 -29200
rect 22500 -29250 22600 -29220
rect 22500 -29450 22520 -29250
rect 22590 -29450 22600 -29250
rect 22500 -29480 22600 -29450
rect 22900 -29250 23100 -29220
rect 22900 -29450 22910 -29250
rect 22980 -29450 23020 -29250
rect 23090 -29450 23100 -29250
rect 22900 -29480 23100 -29450
rect 23400 -29250 23600 -29220
rect 23400 -29450 23410 -29250
rect 23480 -29450 23600 -29250
rect 23400 -29480 23600 -29450
rect 23900 -29480 26000 -29220
rect 22500 -29500 22620 -29480
rect 22880 -29500 23120 -29480
rect 23380 -29500 23620 -29480
rect 23880 -29500 26000 -29480
rect 22500 -29510 26000 -29500
rect 22500 -29580 22650 -29510
rect 22850 -29580 23150 -29510
rect 23350 -29580 26000 -29510
rect 22500 -29600 26000 -29580
rect 23500 -29700 26000 -29600
rect 23500 -29720 23620 -29700
rect 23880 -29720 26000 -29700
rect 23500 -29980 23600 -29720
rect 23900 -29980 26000 -29720
rect 23500 -30000 23620 -29980
rect 23880 -30000 26000 -29980
rect 23500 -30200 26000 -30000
rect 23500 -30220 23620 -30200
rect 23880 -30220 26000 -30200
rect 23500 -30480 23600 -30220
rect 23900 -30480 26000 -30220
rect 23500 -30500 23620 -30480
rect 23880 -30500 26000 -30480
rect 23500 -30700 26000 -30500
rect 23500 -30720 23620 -30700
rect 23880 -30720 24200 -30700
rect 23500 -30980 23600 -30720
rect 23900 -30980 24200 -30720
rect 23500 -31000 23620 -30980
rect 23880 -31000 24200 -30980
rect 23500 -31200 24200 -31000
rect 23500 -31220 23620 -31200
rect 23880 -31220 24200 -31200
rect 23500 -31480 23600 -31220
rect 23900 -31480 24200 -31220
rect 23500 -31500 23620 -31480
rect 23880 -31500 24200 -31480
rect 23500 -31700 24200 -31500
rect 23500 -31720 23620 -31700
rect 23880 -31720 24200 -31700
rect 23500 -31980 23600 -31720
rect 23900 -31980 24200 -31720
rect 23500 -32000 23620 -31980
rect 23880 -32000 24200 -31980
rect 23500 -32200 24200 -32000
rect 23500 -32220 23620 -32200
rect 23880 -32220 24200 -32200
rect 23500 -32480 23600 -32220
rect 23900 -32480 24200 -32220
rect 23500 -32500 23620 -32480
rect 23880 -32500 24200 -32480
rect 23500 -32700 24200 -32500
rect 23500 -32720 23620 -32700
rect 23880 -32720 24200 -32700
rect 23500 -32980 23600 -32720
rect 23900 -32980 24200 -32720
rect 23500 -33000 23620 -32980
rect 23880 -33000 24200 -32980
rect 23500 -33200 24200 -33000
rect 25800 -31000 26000 -30700
rect 30800 -28220 33120 -28200
rect 33380 -28220 33620 -28200
rect 33880 -28220 34120 -28200
rect 34380 -28220 34620 -28200
rect 34880 -28220 35120 -28200
rect 35380 -28220 35620 -28200
rect 35880 -28220 36120 -28200
rect 36380 -28220 36500 -28200
rect 30800 -28480 33100 -28220
rect 33400 -28480 33600 -28220
rect 33900 -28480 34100 -28220
rect 34400 -28480 34600 -28220
rect 34900 -28480 35100 -28220
rect 35400 -28480 35600 -28220
rect 35900 -28480 36100 -28220
rect 36400 -28480 36500 -28220
rect 30800 -28500 33120 -28480
rect 33380 -28500 33620 -28480
rect 33880 -28500 34120 -28480
rect 34380 -28500 34620 -28480
rect 34880 -28500 35120 -28480
rect 35380 -28500 35620 -28480
rect 35880 -28500 36120 -28480
rect 36380 -28500 36500 -28480
rect 30800 -28700 36500 -28500
rect 30800 -28720 33120 -28700
rect 33380 -28720 33620 -28700
rect 33880 -28720 34120 -28700
rect 34380 -28720 34620 -28700
rect 34880 -28720 35120 -28700
rect 35380 -28720 35620 -28700
rect 35880 -28720 36120 -28700
rect 36380 -28720 36500 -28700
rect 30800 -28980 33100 -28720
rect 33400 -28980 33600 -28720
rect 33900 -28980 34100 -28720
rect 34400 -28980 34600 -28720
rect 34900 -28980 35100 -28720
rect 35400 -28980 35600 -28720
rect 35900 -28980 36100 -28720
rect 36400 -28980 36500 -28720
rect 30800 -29000 33120 -28980
rect 33380 -29000 33620 -28980
rect 33880 -29000 34120 -28980
rect 34380 -29000 34620 -28980
rect 34880 -29000 35120 -28980
rect 35380 -29000 35620 -28980
rect 35880 -29000 36120 -28980
rect 36380 -29000 36500 -28980
rect 30800 -29100 36500 -29000
rect 30800 -29200 34500 -29100
rect 30800 -29220 33120 -29200
rect 33380 -29220 33620 -29200
rect 33880 -29220 34120 -29200
rect 34380 -29220 34500 -29200
rect 30800 -29480 33100 -29220
rect 33400 -29480 33600 -29220
rect 33900 -29480 34100 -29220
rect 34400 -29480 34500 -29220
rect 30800 -29500 33120 -29480
rect 33380 -29500 33620 -29480
rect 33880 -29500 34120 -29480
rect 34380 -29500 34500 -29480
rect 30800 -29700 34500 -29500
rect 30800 -29720 33120 -29700
rect 33380 -29720 33620 -29700
rect 33880 -29720 34120 -29700
rect 34380 -29720 34500 -29700
rect 30800 -29980 33100 -29720
rect 33400 -29980 33600 -29720
rect 33900 -29980 34100 -29720
rect 34400 -29980 34500 -29720
rect 30800 -30000 33120 -29980
rect 33380 -30000 33620 -29980
rect 33880 -30000 34120 -29980
rect 34380 -30000 34500 -29980
rect 30800 -30200 34500 -30000
rect 30800 -30220 33120 -30200
rect 33380 -30220 33620 -30200
rect 33880 -30220 34120 -30200
rect 34380 -30220 34500 -30200
rect 30800 -30480 33100 -30220
rect 33400 -30480 33600 -30220
rect 33900 -30480 34100 -30220
rect 34400 -30480 34500 -30220
rect 30800 -30500 33120 -30480
rect 33380 -30500 33620 -30480
rect 33880 -30500 34120 -30480
rect 34380 -30500 34500 -30480
rect 30800 -30700 34500 -30500
rect 30800 -31000 31000 -30700
rect 25800 -33200 31000 -31000
rect 32600 -30720 33120 -30700
rect 33380 -30720 33620 -30700
rect 33880 -30720 34120 -30700
rect 34380 -30720 34500 -30700
rect 32600 -30980 33100 -30720
rect 33400 -30980 33600 -30720
rect 33900 -30980 34100 -30720
rect 34400 -30980 34500 -30720
rect 32600 -31000 33120 -30980
rect 33380 -31000 33620 -30980
rect 33880 -31000 34120 -30980
rect 34380 -31000 34500 -30980
rect 32600 -31200 34500 -31000
rect 32600 -31220 33120 -31200
rect 33380 -31220 33620 -31200
rect 33880 -31220 34120 -31200
rect 34380 -31220 34500 -31200
rect 32600 -31480 33100 -31220
rect 33400 -31480 33600 -31220
rect 33900 -31480 34100 -31220
rect 34400 -31480 34500 -31220
rect 32600 -31500 33120 -31480
rect 33380 -31500 33620 -31480
rect 33880 -31500 34120 -31480
rect 34380 -31500 34500 -31480
rect 32600 -31700 34500 -31500
rect 32600 -31720 33120 -31700
rect 33380 -31720 33620 -31700
rect 33880 -31720 34120 -31700
rect 34380 -31720 34500 -31700
rect 32600 -31980 33100 -31720
rect 33400 -31980 33600 -31720
rect 33900 -31980 34100 -31720
rect 34400 -31980 34500 -31720
rect 32600 -32000 33120 -31980
rect 33380 -32000 33620 -31980
rect 33880 -32000 34120 -31980
rect 34380 -32000 34500 -31980
rect 32600 -32200 34500 -32000
rect 32600 -32220 33120 -32200
rect 33380 -32220 33620 -32200
rect 33880 -32220 34120 -32200
rect 34380 -32220 34500 -32200
rect 32600 -32480 33100 -32220
rect 33400 -32480 33600 -32220
rect 33900 -32480 34100 -32220
rect 34400 -32480 34500 -32220
rect 32600 -32500 33120 -32480
rect 33380 -32500 33620 -32480
rect 33880 -32500 34120 -32480
rect 34380 -32500 34500 -32480
rect 32600 -32700 34500 -32500
rect 32600 -32720 33120 -32700
rect 33380 -32720 33620 -32700
rect 33880 -32720 34120 -32700
rect 34380 -32720 34500 -32700
rect 32600 -32980 33100 -32720
rect 33400 -32980 33600 -32720
rect 33900 -32980 34100 -32720
rect 34400 -32980 34500 -32720
rect 32600 -33000 33120 -32980
rect 33380 -33000 33620 -32980
rect 33880 -33000 34120 -32980
rect 34380 -33000 34500 -32980
rect 32600 -33200 34500 -33000
rect 23500 -33220 23620 -33200
rect 23880 -33220 33120 -33200
rect 33380 -33220 33620 -33200
rect 33880 -33220 34120 -33200
rect 34380 -33220 34500 -33200
rect 23500 -33480 23600 -33220
rect 23900 -33480 33100 -33220
rect 33400 -33480 33600 -33220
rect 33900 -33480 34100 -33220
rect 34400 -33480 34500 -33220
rect 23500 -33500 23620 -33480
rect 23880 -33500 33120 -33480
rect 33380 -33500 33620 -33480
rect 33880 -33500 34120 -33480
rect 34380 -33500 34500 -33480
rect 23500 -33600 34500 -33500
rect -27500 -34800 -25500 -34700
rect -27500 -34820 -27380 -34800
rect -27120 -34820 -26880 -34800
rect -26620 -34820 -26380 -34800
rect -26120 -34820 -25880 -34800
rect -25620 -34820 -25500 -34800
rect -27500 -35080 -27400 -34820
rect -27100 -35080 -26900 -34820
rect -26600 -35080 -26400 -34820
rect -26100 -35080 -25900 -34820
rect -25600 -35080 -25500 -34820
rect -27500 -35100 -27380 -35080
rect -27120 -35100 -26880 -35080
rect -26620 -35100 -26380 -35080
rect -26120 -35100 -25880 -35080
rect -25620 -35100 -25500 -35080
rect -27500 -35300 -25500 -35100
rect -27500 -35320 -27380 -35300
rect -27120 -35320 -26880 -35300
rect -26620 -35320 -26380 -35300
rect -26120 -35320 -25880 -35300
rect -25620 -35320 -25500 -35300
rect -27500 -35580 -27400 -35320
rect -27100 -35580 -26900 -35320
rect -26600 -35580 -26400 -35320
rect -26100 -35580 -25900 -35320
rect -25600 -35580 -25500 -35320
rect -27500 -35600 -27380 -35580
rect -27120 -35600 -26880 -35580
rect -26620 -35600 -26380 -35580
rect -26120 -35600 -25880 -35580
rect -25620 -35600 -25500 -35580
rect -27500 -35800 -25500 -35600
rect -27500 -35820 -27380 -35800
rect -27120 -35820 -26880 -35800
rect -26620 -35820 -26380 -35800
rect -26120 -35820 -25880 -35800
rect -25620 -35820 -25500 -35800
rect -27500 -36080 -27400 -35820
rect -27100 -36080 -26900 -35820
rect -26600 -36080 -26400 -35820
rect -26100 -36080 -25900 -35820
rect -25600 -36080 -25500 -35820
rect -27500 -36100 -27380 -36080
rect -27120 -36100 -26880 -36080
rect -26620 -36100 -26380 -36080
rect -26120 -36100 -25880 -36080
rect -25620 -36100 -25500 -36080
rect -27500 -36300 -25500 -36100
rect -27500 -36320 -27380 -36300
rect -27120 -36320 -26880 -36300
rect -26620 -36320 -26380 -36300
rect -26120 -36320 -25880 -36300
rect -25620 -36320 -25500 -36300
rect -27500 -36580 -27400 -36320
rect -27100 -36580 -26900 -36320
rect -26600 -36580 -26400 -36320
rect -26100 -36580 -25900 -36320
rect -25600 -36580 -25500 -36320
rect -27500 -36600 -27380 -36580
rect -27120 -36600 -26880 -36580
rect -26620 -36600 -26380 -36580
rect -26120 -36600 -25880 -36580
rect -25620 -36600 -25500 -36580
rect -27500 -36700 -25500 -36600
rect 124500 -38200 136500 -38100
rect 124500 -38220 124620 -38200
rect 124880 -38220 125120 -38200
rect 125380 -38220 125620 -38200
rect 125880 -38220 126120 -38200
rect 126380 -38220 126620 -38200
rect 126880 -38220 127120 -38200
rect 127380 -38220 127620 -38200
rect 127880 -38220 128120 -38200
rect 128380 -38220 128620 -38200
rect 128880 -38220 129120 -38200
rect 129380 -38220 129620 -38200
rect 129880 -38220 130120 -38200
rect 130380 -38220 130620 -38200
rect 130880 -38220 131120 -38200
rect 131380 -38220 131620 -38200
rect 131880 -38220 132120 -38200
rect 132380 -38220 132620 -38200
rect 132880 -38220 133120 -38200
rect 133380 -38220 133620 -38200
rect 133880 -38220 134120 -38200
rect 134380 -38220 134620 -38200
rect 134880 -38220 135120 -38200
rect 135380 -38220 135620 -38200
rect 135880 -38220 136120 -38200
rect 136380 -38220 136500 -38200
rect 124500 -38480 124600 -38220
rect 124900 -38480 125100 -38220
rect 125400 -38480 125600 -38220
rect 125900 -38480 126100 -38220
rect 126400 -38480 126600 -38220
rect 126900 -38480 127100 -38220
rect 127400 -38480 127600 -38220
rect 127900 -38480 128100 -38220
rect 128400 -38480 128600 -38220
rect 128900 -38480 129100 -38220
rect 129400 -38480 129600 -38220
rect 129900 -38480 130100 -38220
rect 130400 -38480 130600 -38220
rect 130900 -38480 131100 -38220
rect 131400 -38480 131600 -38220
rect 131900 -38480 132100 -38220
rect 132400 -38480 132600 -38220
rect 132900 -38480 133100 -38220
rect 133400 -38480 133600 -38220
rect 133900 -38480 134100 -38220
rect 134400 -38480 134600 -38220
rect 134900 -38480 135100 -38220
rect 135400 -38480 135600 -38220
rect 135900 -38480 136100 -38220
rect 136400 -38480 136500 -38220
rect 124500 -38500 124620 -38480
rect 124880 -38500 125120 -38480
rect 125380 -38500 125620 -38480
rect 125880 -38500 126120 -38480
rect 126380 -38500 126620 -38480
rect 126880 -38500 127120 -38480
rect 127380 -38500 127620 -38480
rect 127880 -38500 128120 -38480
rect 128380 -38500 128620 -38480
rect 128880 -38500 129120 -38480
rect 129380 -38500 129620 -38480
rect 129880 -38500 130120 -38480
rect 130380 -38500 130620 -38480
rect 130880 -38500 131120 -38480
rect 131380 -38500 131620 -38480
rect 131880 -38500 132120 -38480
rect 132380 -38500 132620 -38480
rect 132880 -38500 133120 -38480
rect 133380 -38500 133620 -38480
rect 133880 -38500 134120 -38480
rect 134380 -38500 134620 -38480
rect 134880 -38500 135120 -38480
rect 135380 -38500 135620 -38480
rect 135880 -38500 136120 -38480
rect 136380 -38500 136500 -38480
rect 124500 -38700 136500 -38500
rect 124500 -38720 124620 -38700
rect 124880 -38720 125120 -38700
rect 125380 -38720 125620 -38700
rect 125880 -38720 126120 -38700
rect 126380 -38720 126620 -38700
rect 126880 -38720 127120 -38700
rect 127380 -38720 127620 -38700
rect 127880 -38720 128120 -38700
rect 128380 -38720 128620 -38700
rect 128880 -38720 129120 -38700
rect 129380 -38720 129620 -38700
rect 129880 -38720 130120 -38700
rect 130380 -38720 130620 -38700
rect 130880 -38720 131120 -38700
rect 131380 -38720 131620 -38700
rect 131880 -38720 132120 -38700
rect 132380 -38720 132620 -38700
rect 132880 -38720 133120 -38700
rect 133380 -38720 133620 -38700
rect 133880 -38720 134120 -38700
rect 134380 -38720 134620 -38700
rect 134880 -38720 135120 -38700
rect 135380 -38720 135620 -38700
rect 135880 -38720 136120 -38700
rect 136380 -38720 136500 -38700
rect 124500 -38980 124600 -38720
rect 124900 -38980 125100 -38720
rect 125400 -38980 125600 -38720
rect 125900 -38980 126100 -38720
rect 126400 -38980 126600 -38720
rect 126900 -38980 127100 -38720
rect 127400 -38980 127600 -38720
rect 127900 -38980 128100 -38720
rect 128400 -38980 128600 -38720
rect 128900 -38980 129100 -38720
rect 129400 -38980 129600 -38720
rect 129900 -38980 130100 -38720
rect 130400 -38980 130600 -38720
rect 130900 -38980 131100 -38720
rect 131400 -38980 131600 -38720
rect 131900 -38980 132100 -38720
rect 132400 -38980 132600 -38720
rect 132900 -38980 133100 -38720
rect 133400 -38980 133600 -38720
rect 133900 -38980 134100 -38720
rect 134400 -38980 134600 -38720
rect 134900 -38980 135100 -38720
rect 135400 -38980 135600 -38720
rect 135900 -38980 136100 -38720
rect 136400 -38980 136500 -38720
rect 124500 -39000 124620 -38980
rect 124880 -39000 125120 -38980
rect 125380 -39000 125620 -38980
rect 125880 -39000 126120 -38980
rect 126380 -39000 126620 -38980
rect 126880 -39000 127120 -38980
rect 127380 -39000 127620 -38980
rect 127880 -39000 128120 -38980
rect 128380 -39000 128620 -38980
rect 128880 -39000 129120 -38980
rect 129380 -39000 129620 -38980
rect 129880 -39000 130120 -38980
rect 130380 -39000 130620 -38980
rect 130880 -39000 131120 -38980
rect 131380 -39000 131620 -38980
rect 131880 -39000 132120 -38980
rect 132380 -39000 132620 -38980
rect 132880 -39000 133120 -38980
rect 133380 -39000 133620 -38980
rect 133880 -39000 134120 -38980
rect 134380 -39000 134620 -38980
rect 134880 -39000 135120 -38980
rect 135380 -39000 135620 -38980
rect 135880 -39000 136120 -38980
rect 136380 -39000 136500 -38980
rect 124500 -39100 136500 -39000
<< via1 >>
rect -83350 82810 -83150 82880
rect -82850 82810 -82650 82880
rect -82350 82810 -82150 82880
rect -81850 82810 -81650 82880
rect -81350 82810 -81150 82880
rect -80850 82810 -80650 82880
rect -80350 82810 -80150 82880
rect -79850 82810 -79650 82880
rect -79350 82810 -79150 82880
rect -78850 82810 -78650 82880
rect -78350 82810 -78150 82880
rect -77850 82810 -77650 82880
rect -77350 82810 -77150 82880
rect -76850 82810 -76650 82880
rect -76350 82810 -76150 82880
rect -75850 82810 -75650 82880
rect -75350 82810 -75150 82880
rect -74850 82810 -74650 82880
rect -74350 82810 -74150 82880
rect -73850 82810 -73650 82880
rect -73350 82810 -73150 82880
rect -72850 82810 -72650 82880
rect -72350 82810 -72150 82880
rect -71850 82810 -71650 82880
rect -71350 82810 -71150 82880
rect -70850 82810 -70650 82880
rect -70350 82810 -70150 82880
rect -69850 82810 -69650 82880
rect -69350 82810 -69150 82880
rect -68850 82810 -68650 82880
rect -68350 82810 -68150 82880
rect -67850 82810 -67650 82880
rect -67350 82810 -67150 82880
rect -66850 82810 -66650 82880
rect -66350 82810 -66150 82880
rect -65850 82810 -65650 82880
rect -65350 82810 -65150 82880
rect -64850 82810 -64650 82880
rect -64350 82810 -64150 82880
rect -63850 82810 -63650 82880
rect -63350 82810 -63150 82880
rect -62850 82810 -62650 82880
rect -62350 82810 -62150 82880
rect -61850 82810 -61650 82880
rect -61350 82810 -61150 82880
rect -60850 82810 -60650 82880
rect -60350 82810 -60150 82880
rect -59850 82810 -59650 82880
rect -59350 82810 -59150 82880
rect -58850 82810 -58650 82880
rect -58350 82810 -58150 82880
rect -57850 82810 -57650 82880
rect -57350 82810 -57150 82880
rect -56850 82810 -56650 82880
rect -56350 82810 -56150 82880
rect -55850 82810 -55650 82880
rect -55350 82810 -55150 82880
rect -54850 82810 -54650 82880
rect -54350 82810 -54150 82880
rect -53850 82810 -53650 82880
rect -53350 82810 -53150 82880
rect -52850 82810 -52650 82880
rect -52350 82810 -52150 82880
rect -51850 82810 -51650 82880
rect -51350 82810 -51150 82880
rect -50850 82810 -50650 82880
rect -50350 82810 -50150 82880
rect -49850 82810 -49650 82880
rect -49350 82810 -49150 82880
rect -48850 82810 -48650 82880
rect -48350 82810 -48150 82880
rect -47850 82810 -47650 82880
rect -47350 82810 -47150 82880
rect -46850 82810 -46650 82880
rect -46350 82810 -46150 82880
rect -45850 82810 -45650 82880
rect -45350 82810 -45150 82880
rect -44850 82810 -44650 82880
rect -44350 82810 -44150 82880
rect -43850 82810 -43650 82880
rect -43350 82810 -43150 82880
rect -42850 82810 -42650 82880
rect -42350 82810 -42150 82880
rect -41850 82810 -41650 82880
rect -41350 82810 -41150 82880
rect -40850 82810 -40650 82880
rect -40350 82810 -40150 82880
rect -39850 82810 -39650 82880
rect -39350 82810 -39150 82880
rect -38850 82810 -38650 82880
rect -38350 82810 -38150 82880
rect -37850 82810 -37650 82880
rect -37350 82810 -37150 82880
rect -36850 82810 -36650 82880
rect -36350 82810 -36150 82880
rect -35850 82810 -35650 82880
rect -35350 82810 -35150 82880
rect -34850 82810 -34650 82880
rect -34350 82810 -34150 82880
rect -33850 82810 -33650 82880
rect -33350 82810 -33150 82880
rect -32850 82810 -32650 82880
rect -32350 82810 -32150 82880
rect -31850 82810 -31650 82880
rect -31350 82810 -31150 82880
rect -30850 82810 -30650 82880
rect -30350 82810 -30150 82880
rect -29850 82810 -29650 82880
rect -29350 82810 -29150 82880
rect -28850 82810 -28650 82880
rect -28350 82810 -28150 82880
rect -27850 82810 -27650 82880
rect -27350 82810 -27150 82880
rect -26850 82810 -26650 82880
rect -26350 82810 -26150 82880
rect -25850 82810 -25650 82880
rect -25350 82810 -25150 82880
rect -24850 82810 -24650 82880
rect -24350 82810 -24150 82880
rect -23850 82810 -23650 82880
rect -23350 82810 -23150 82880
rect -22850 82810 -22650 82880
rect -22350 82810 -22150 82880
rect -21850 82810 -21650 82880
rect -21350 82810 -21150 82880
rect -20850 82810 -20650 82880
rect -20350 82810 -20150 82880
rect -19850 82810 -19650 82880
rect -19350 82810 -19150 82880
rect -18850 82810 -18650 82880
rect -18350 82810 -18150 82880
rect -17850 82810 -17650 82880
rect -17350 82810 -17150 82880
rect -16850 82810 -16650 82880
rect -16350 82810 -16150 82880
rect -15850 82810 -15650 82880
rect -15350 82810 -15150 82880
rect -14850 82810 -14650 82880
rect -14350 82810 -14150 82880
rect -13850 82810 -13650 82880
rect -13350 82810 -13150 82880
rect -12850 82810 -12650 82880
rect -12350 82810 -12150 82880
rect -11850 82810 -11650 82880
rect -11350 82810 -11150 82880
rect -10850 82810 -10650 82880
rect -10350 82810 -10150 82880
rect -9850 82810 -9650 82880
rect -9350 82810 -9150 82880
rect -8850 82810 -8650 82880
rect -8350 82810 -8150 82880
rect -7850 82810 -7650 82880
rect -7350 82810 -7150 82880
rect -6850 82810 -6650 82880
rect -6350 82810 -6150 82880
rect -5850 82810 -5650 82880
rect -5350 82810 -5150 82880
rect -4850 82810 -4650 82880
rect -4350 82810 -4150 82880
rect -3850 82810 -3650 82880
rect -3350 82810 -3150 82880
rect -2850 82810 -2650 82880
rect -2350 82810 -2150 82880
rect -1850 82810 -1650 82880
rect -1350 82810 -1150 82880
rect -850 82810 -650 82880
rect -350 82810 -150 82880
rect 150 82810 350 82880
rect 650 82810 850 82880
rect 1150 82810 1350 82880
rect 1650 82810 1850 82880
rect 2150 82810 2350 82880
rect 2650 82810 2850 82880
rect 3150 82810 3350 82880
rect 3650 82810 3850 82880
rect 4150 82810 4350 82880
rect 4650 82810 4850 82880
rect 5150 82810 5350 82880
rect 5650 82810 5850 82880
rect 6150 82810 6350 82880
rect 6650 82810 6850 82880
rect 7150 82810 7350 82880
rect 7650 82810 7850 82880
rect 8150 82810 8350 82880
rect 8650 82810 8850 82880
rect 9150 82810 9350 82880
rect 9650 82810 9850 82880
rect 10150 82810 10350 82880
rect 10650 82810 10850 82880
rect 11150 82810 11350 82880
rect 11650 82810 11850 82880
rect 12150 82810 12350 82880
rect 12650 82810 12850 82880
rect 13150 82810 13350 82880
rect 13650 82810 13850 82880
rect 14150 82810 14350 82880
rect 14650 82810 14850 82880
rect 15150 82810 15350 82880
rect 15650 82810 15850 82880
rect 16150 82810 16350 82880
rect 16650 82810 16850 82880
rect 17150 82810 17350 82880
rect 17650 82810 17850 82880
rect 18150 82810 18350 82880
rect 18650 82810 18850 82880
rect 19150 82810 19350 82880
rect 19650 82810 19850 82880
rect 20150 82810 20350 82880
rect 20650 82810 20850 82880
rect 21150 82810 21350 82880
rect 21650 82810 21850 82880
rect 22150 82810 22350 82880
rect 22650 82810 22850 82880
rect 23150 82810 23350 82880
rect 23650 82810 23850 82880
rect 24150 82810 24350 82880
rect 24650 82810 24850 82880
rect 25150 82810 25350 82880
rect 25650 82810 25850 82880
rect 26150 82810 26350 82880
rect 26650 82810 26850 82880
rect 27150 82810 27350 82880
rect 27650 82810 27850 82880
rect 28150 82810 28350 82880
rect 28650 82810 28850 82880
rect 29150 82810 29350 82880
rect 29650 82810 29850 82880
rect 30150 82810 30350 82880
rect 30650 82810 30850 82880
rect 31150 82810 31350 82880
rect 31650 82810 31850 82880
rect 32150 82810 32350 82880
rect 32650 82810 32850 82880
rect 33150 82810 33350 82880
rect 33650 82810 33850 82880
rect 34150 82810 34350 82880
rect 34650 82810 34850 82880
rect 35150 82810 35350 82880
rect 35650 82810 35850 82880
rect 36150 82810 36350 82880
rect 36650 82810 36850 82880
rect 37150 82810 37350 82880
rect 37650 82810 37850 82880
rect 38150 82810 38350 82880
rect 38650 82810 38850 82880
rect 39150 82810 39350 82880
rect 39650 82810 39850 82880
rect 40150 82810 40350 82880
rect 40650 82810 40850 82880
rect 41150 82810 41350 82880
rect 41650 82810 41850 82880
rect 42150 82810 42350 82880
rect 42650 82810 42850 82880
rect 43150 82810 43350 82880
rect 43650 82810 43850 82880
rect 44150 82810 44350 82880
rect 44650 82810 44850 82880
rect 45150 82810 45350 82880
rect 45650 82810 45850 82880
rect 46150 82810 46350 82880
rect 46650 82810 46850 82880
rect 47150 82810 47350 82880
rect 47650 82810 47850 82880
rect 48150 82810 48350 82880
rect 48650 82810 48850 82880
rect 49150 82810 49350 82880
rect 49650 82810 49850 82880
rect 50150 82810 50350 82880
rect 50650 82810 50850 82880
rect 51150 82810 51350 82880
rect 51650 82810 51850 82880
rect 52150 82810 52350 82880
rect 52650 82810 52850 82880
rect 53150 82810 53350 82880
rect 53650 82810 53850 82880
rect 54150 82810 54350 82880
rect 54650 82810 54850 82880
rect 55150 82810 55350 82880
rect 55650 82810 55850 82880
rect 56150 82810 56350 82880
rect 56650 82810 56850 82880
rect 57150 82810 57350 82880
rect 57650 82810 57850 82880
rect 58150 82810 58350 82880
rect 58650 82810 58850 82880
rect 59150 82810 59350 82880
rect 59650 82810 59850 82880
rect 60150 82810 60350 82880
rect 60650 82810 60850 82880
rect 61150 82810 61350 82880
rect 61650 82810 61850 82880
rect 62150 82810 62350 82880
rect 62650 82810 62850 82880
rect 63150 82810 63350 82880
rect 63650 82810 63850 82880
rect 64150 82810 64350 82880
rect 64650 82810 64850 82880
rect 65150 82810 65350 82880
rect 65650 82810 65850 82880
rect 66150 82810 66350 82880
rect 66650 82810 66850 82880
rect 67150 82810 67350 82880
rect 67650 82810 67850 82880
rect 68150 82810 68350 82880
rect 68650 82810 68850 82880
rect 69150 82810 69350 82880
rect 69650 82810 69850 82880
rect 70150 82810 70350 82880
rect 70650 82810 70850 82880
rect 71150 82810 71350 82880
rect 71650 82810 71850 82880
rect 72150 82810 72350 82880
rect 72650 82810 72850 82880
rect 73150 82810 73350 82880
rect 73650 82810 73850 82880
rect 74150 82810 74350 82880
rect 74650 82810 74850 82880
rect 75150 82810 75350 82880
rect 75650 82810 75850 82880
rect 76150 82810 76350 82880
rect 76650 82810 76850 82880
rect 77150 82810 77350 82880
rect 77650 82810 77850 82880
rect 78150 82810 78350 82880
rect 78650 82810 78850 82880
rect 79150 82810 79350 82880
rect 79650 82810 79850 82880
rect 80150 82810 80350 82880
rect 80650 82810 80850 82880
rect 81150 82810 81350 82880
rect 81650 82810 81850 82880
rect 82150 82810 82350 82880
rect 82650 82810 82850 82880
rect 83150 82810 83350 82880
rect 83650 82810 83850 82880
rect 84150 82810 84350 82880
rect 84650 82810 84850 82880
rect 85150 82810 85350 82880
rect 85650 82810 85850 82880
rect 86150 82810 86350 82880
rect 86650 82810 86850 82880
rect 87150 82810 87350 82880
rect 87650 82810 87850 82880
rect 88150 82810 88350 82880
rect 88650 82810 88850 82880
rect 89150 82810 89350 82880
rect 89650 82810 89850 82880
rect 90150 82810 90350 82880
rect 90650 82810 90850 82880
rect 91150 82810 91350 82880
rect 91650 82810 91850 82880
rect 92150 82810 92350 82880
rect 92650 82810 92850 82880
rect 93150 82810 93350 82880
rect 93650 82810 93850 82880
rect 94150 82810 94350 82880
rect 94650 82810 94850 82880
rect 95150 82810 95350 82880
rect 95650 82810 95850 82880
rect 96150 82810 96350 82880
rect 96650 82810 96850 82880
rect 97150 82810 97350 82880
rect 97650 82810 97850 82880
rect 98150 82810 98350 82880
rect 98650 82810 98850 82880
rect 99150 82810 99350 82880
rect 99650 82810 99850 82880
rect 100150 82810 100350 82880
rect -83480 82550 -83410 82750
rect -83090 82550 -83020 82750
rect -82980 82550 -82910 82750
rect -82590 82550 -82520 82750
rect -82480 82550 -82410 82750
rect -82090 82550 -82020 82750
rect -81980 82550 -81910 82750
rect -81590 82550 -81520 82750
rect -81480 82550 -81410 82750
rect -81090 82550 -81020 82750
rect -80980 82550 -80910 82750
rect -80590 82550 -80520 82750
rect -80480 82550 -80410 82750
rect -80090 82550 -80020 82750
rect -79980 82550 -79910 82750
rect -79590 82550 -79520 82750
rect -79480 82550 -79410 82750
rect -79090 82550 -79020 82750
rect -78980 82550 -78910 82750
rect -78590 82550 -78520 82750
rect -78480 82550 -78410 82750
rect -78090 82550 -78020 82750
rect -77980 82550 -77910 82750
rect -77590 82550 -77520 82750
rect -77480 82550 -77410 82750
rect -77090 82550 -77020 82750
rect -76980 82550 -76910 82750
rect -76590 82550 -76520 82750
rect -76480 82550 -76410 82750
rect -76090 82550 -76020 82750
rect -75980 82550 -75910 82750
rect -75590 82550 -75520 82750
rect -75480 82550 -75410 82750
rect -75090 82550 -75020 82750
rect -74980 82550 -74910 82750
rect -74590 82550 -74520 82750
rect -74480 82550 -74410 82750
rect -74090 82550 -74020 82750
rect -73980 82550 -73910 82750
rect -73590 82550 -73520 82750
rect -73480 82550 -73410 82750
rect -73090 82550 -73020 82750
rect -72980 82550 -72910 82750
rect -72590 82550 -72520 82750
rect -72480 82550 -72410 82750
rect -72090 82550 -72020 82750
rect -71980 82550 -71910 82750
rect -71590 82550 -71520 82750
rect -71480 82550 -71410 82750
rect -71090 82550 -71020 82750
rect -70980 82550 -70910 82750
rect -70590 82550 -70520 82750
rect -70480 82550 -70410 82750
rect -70090 82550 -70020 82750
rect -69980 82550 -69910 82750
rect -69590 82550 -69520 82750
rect -69480 82550 -69410 82750
rect -69090 82550 -69020 82750
rect -68980 82550 -68910 82750
rect -68590 82550 -68520 82750
rect -68480 82550 -68410 82750
rect -68090 82550 -68020 82750
rect -67980 82550 -67910 82750
rect -67590 82550 -67520 82750
rect -67480 82550 -67410 82750
rect -67090 82550 -67020 82750
rect -66980 82550 -66910 82750
rect -66590 82550 -66520 82750
rect -66480 82550 -66410 82750
rect -66090 82550 -66020 82750
rect -65980 82550 -65910 82750
rect -65590 82550 -65520 82750
rect -65480 82550 -65410 82750
rect -65090 82550 -65020 82750
rect -64980 82550 -64910 82750
rect -64590 82550 -64520 82750
rect -64480 82550 -64410 82750
rect -64090 82550 -64020 82750
rect -63980 82550 -63910 82750
rect -63590 82550 -63520 82750
rect -63480 82550 -63410 82750
rect -63090 82550 -63020 82750
rect -62980 82550 -62910 82750
rect -62590 82550 -62520 82750
rect -62480 82550 -62410 82750
rect -62090 82550 -62020 82750
rect -61980 82550 -61910 82750
rect -61590 82550 -61520 82750
rect -61480 82550 -61410 82750
rect -61090 82550 -61020 82750
rect -60980 82550 -60910 82750
rect -60590 82550 -60520 82750
rect -60480 82550 -60410 82750
rect -60090 82550 -60020 82750
rect -59980 82550 -59910 82750
rect -59590 82550 -59520 82750
rect -59480 82550 -59410 82750
rect -59090 82550 -59020 82750
rect -58980 82550 -58910 82750
rect -58590 82550 -58520 82750
rect -58480 82550 -58410 82750
rect -58090 82550 -58020 82750
rect -57980 82550 -57910 82750
rect -57590 82550 -57520 82750
rect -57480 82550 -57410 82750
rect -57090 82550 -57020 82750
rect -56980 82550 -56910 82750
rect -56590 82550 -56520 82750
rect -56480 82550 -56410 82750
rect -56090 82550 -56020 82750
rect -55980 82550 -55910 82750
rect -55590 82550 -55520 82750
rect -55480 82550 -55410 82750
rect -55090 82550 -55020 82750
rect -54980 82550 -54910 82750
rect -54590 82550 -54520 82750
rect -54480 82550 -54410 82750
rect -54090 82550 -54020 82750
rect -53980 82550 -53910 82750
rect -53590 82550 -53520 82750
rect -53480 82550 -53410 82750
rect -53090 82550 -53020 82750
rect -52980 82550 -52910 82750
rect -52590 82550 -52520 82750
rect -52480 82550 -52410 82750
rect -52090 82550 -52020 82750
rect -51980 82550 -51910 82750
rect -51590 82550 -51520 82750
rect -51480 82550 -51410 82750
rect -51090 82550 -51020 82750
rect -50980 82550 -50910 82750
rect -50590 82550 -50520 82750
rect -50480 82550 -50410 82750
rect -50090 82550 -50020 82750
rect -49980 82550 -49910 82750
rect -49590 82550 -49520 82750
rect -49480 82550 -49410 82750
rect -49090 82550 -49020 82750
rect -48980 82550 -48910 82750
rect -48590 82550 -48520 82750
rect -48480 82550 -48410 82750
rect -48090 82550 -48020 82750
rect -47980 82550 -47910 82750
rect -47590 82550 -47520 82750
rect -47480 82550 -47410 82750
rect -47090 82550 -47020 82750
rect -46980 82550 -46910 82750
rect -46590 82550 -46520 82750
rect -46480 82550 -46410 82750
rect -46090 82550 -46020 82750
rect -45980 82550 -45910 82750
rect -45590 82550 -45520 82750
rect -45480 82550 -45410 82750
rect -45090 82550 -45020 82750
rect -44980 82550 -44910 82750
rect -44590 82550 -44520 82750
rect -44480 82550 -44410 82750
rect -44090 82550 -44020 82750
rect -43980 82550 -43910 82750
rect -43590 82550 -43520 82750
rect -43480 82550 -43410 82750
rect -43090 82550 -43020 82750
rect -42980 82550 -42910 82750
rect -42590 82550 -42520 82750
rect -42480 82550 -42410 82750
rect -42090 82550 -42020 82750
rect -41980 82550 -41910 82750
rect -41590 82550 -41520 82750
rect -41480 82550 -41410 82750
rect -41090 82550 -41020 82750
rect -40980 82550 -40910 82750
rect -40590 82550 -40520 82750
rect -40480 82550 -40410 82750
rect -40090 82550 -40020 82750
rect -39980 82550 -39910 82750
rect -39590 82550 -39520 82750
rect -39480 82550 -39410 82750
rect -39090 82550 -39020 82750
rect -38980 82550 -38910 82750
rect -38590 82550 -38520 82750
rect -38480 82550 -38410 82750
rect -38090 82550 -38020 82750
rect -37980 82550 -37910 82750
rect -37590 82550 -37520 82750
rect -37480 82550 -37410 82750
rect -37090 82550 -37020 82750
rect -36980 82550 -36910 82750
rect -36590 82550 -36520 82750
rect -36480 82550 -36410 82750
rect -36090 82550 -36020 82750
rect -35980 82550 -35910 82750
rect -35590 82550 -35520 82750
rect -35480 82550 -35410 82750
rect -35090 82550 -35020 82750
rect -34980 82550 -34910 82750
rect -34590 82550 -34520 82750
rect -34480 82550 -34410 82750
rect -34090 82550 -34020 82750
rect -33980 82550 -33910 82750
rect -33590 82550 -33520 82750
rect -33480 82550 -33410 82750
rect -33090 82550 -33020 82750
rect -32980 82550 -32910 82750
rect -32590 82550 -32520 82750
rect -32480 82550 -32410 82750
rect -32090 82550 -32020 82750
rect -31980 82550 -31910 82750
rect -31590 82550 -31520 82750
rect -31480 82550 -31410 82750
rect -31090 82550 -31020 82750
rect -30980 82550 -30910 82750
rect -30590 82550 -30520 82750
rect -30480 82550 -30410 82750
rect -30090 82550 -30020 82750
rect -29980 82550 -29910 82750
rect -29590 82550 -29520 82750
rect -29480 82550 -29410 82750
rect -29090 82550 -29020 82750
rect -28980 82550 -28910 82750
rect -28590 82550 -28520 82750
rect -28480 82550 -28410 82750
rect -28090 82550 -28020 82750
rect -27980 82550 -27910 82750
rect -27590 82550 -27520 82750
rect -27480 82550 -27410 82750
rect -27090 82550 -27020 82750
rect -26980 82550 -26910 82750
rect -26590 82550 -26520 82750
rect -26480 82550 -26410 82750
rect -26090 82550 -26020 82750
rect -25980 82550 -25910 82750
rect -25590 82550 -25520 82750
rect -25480 82550 -25410 82750
rect -25090 82550 -25020 82750
rect -24980 82550 -24910 82750
rect -24590 82550 -24520 82750
rect -24480 82550 -24410 82750
rect -24090 82550 -24020 82750
rect -23980 82550 -23910 82750
rect -23590 82550 -23520 82750
rect -23480 82550 -23410 82750
rect -23090 82550 -23020 82750
rect -22980 82550 -22910 82750
rect -22590 82550 -22520 82750
rect -22480 82550 -22410 82750
rect -22090 82550 -22020 82750
rect -21980 82550 -21910 82750
rect -21590 82550 -21520 82750
rect -21480 82550 -21410 82750
rect -21090 82550 -21020 82750
rect -20980 82550 -20910 82750
rect -20590 82550 -20520 82750
rect -20480 82550 -20410 82750
rect -20090 82550 -20020 82750
rect -19980 82550 -19910 82750
rect -19590 82550 -19520 82750
rect -19480 82550 -19410 82750
rect -19090 82550 -19020 82750
rect -18980 82550 -18910 82750
rect -18590 82550 -18520 82750
rect -18480 82550 -18410 82750
rect -18090 82550 -18020 82750
rect -17980 82550 -17910 82750
rect -17590 82550 -17520 82750
rect -17480 82550 -17410 82750
rect -17090 82550 -17020 82750
rect -16980 82550 -16910 82750
rect -16590 82550 -16520 82750
rect -16480 82550 -16410 82750
rect -16090 82550 -16020 82750
rect -15980 82550 -15910 82750
rect -15590 82550 -15520 82750
rect -15480 82550 -15410 82750
rect -15090 82550 -15020 82750
rect -14980 82550 -14910 82750
rect -14590 82550 -14520 82750
rect -14480 82550 -14410 82750
rect -14090 82550 -14020 82750
rect -13980 82550 -13910 82750
rect -13590 82550 -13520 82750
rect -13480 82550 -13410 82750
rect -13090 82550 -13020 82750
rect -12980 82550 -12910 82750
rect -12590 82550 -12520 82750
rect -12480 82550 -12410 82750
rect -12090 82550 -12020 82750
rect -11980 82550 -11910 82750
rect -11590 82550 -11520 82750
rect -11480 82550 -11410 82750
rect -11090 82550 -11020 82750
rect -10980 82550 -10910 82750
rect -10590 82550 -10520 82750
rect -10480 82550 -10410 82750
rect -10090 82550 -10020 82750
rect -9980 82550 -9910 82750
rect -9590 82550 -9520 82750
rect -9480 82550 -9410 82750
rect -9090 82550 -9020 82750
rect -8980 82550 -8910 82750
rect -8590 82550 -8520 82750
rect -8480 82550 -8410 82750
rect -8090 82550 -8020 82750
rect -7980 82550 -7910 82750
rect -7590 82550 -7520 82750
rect -7480 82550 -7410 82750
rect -7090 82550 -7020 82750
rect -6980 82550 -6910 82750
rect -6590 82550 -6520 82750
rect -6480 82550 -6410 82750
rect -6090 82550 -6020 82750
rect -5980 82550 -5910 82750
rect -5590 82550 -5520 82750
rect -5480 82550 -5410 82750
rect -5090 82550 -5020 82750
rect -4980 82550 -4910 82750
rect -4590 82550 -4520 82750
rect -4480 82550 -4410 82750
rect -4090 82550 -4020 82750
rect -3980 82550 -3910 82750
rect -3590 82550 -3520 82750
rect -3480 82550 -3410 82750
rect -3090 82550 -3020 82750
rect -2980 82550 -2910 82750
rect -2590 82550 -2520 82750
rect -2480 82550 -2410 82750
rect -2090 82550 -2020 82750
rect -1980 82550 -1910 82750
rect -1590 82550 -1520 82750
rect -1480 82550 -1410 82750
rect -1090 82550 -1020 82750
rect -980 82550 -910 82750
rect -590 82550 -520 82750
rect -480 82550 -410 82750
rect -90 82550 -20 82750
rect 20 82550 90 82750
rect 410 82550 480 82750
rect 520 82550 590 82750
rect 910 82550 980 82750
rect 1020 82550 1090 82750
rect 1410 82550 1480 82750
rect 1520 82550 1590 82750
rect 1910 82550 1980 82750
rect 2020 82550 2090 82750
rect 2410 82550 2480 82750
rect 2520 82550 2590 82750
rect 2910 82550 2980 82750
rect 3020 82550 3090 82750
rect 3410 82550 3480 82750
rect 3520 82550 3590 82750
rect 3910 82550 3980 82750
rect 4020 82550 4090 82750
rect 4410 82550 4480 82750
rect 4520 82550 4590 82750
rect 4910 82550 4980 82750
rect 5020 82550 5090 82750
rect 5410 82550 5480 82750
rect 5520 82550 5590 82750
rect 5910 82550 5980 82750
rect 6020 82550 6090 82750
rect 6410 82550 6480 82750
rect 6520 82550 6590 82750
rect 6910 82550 6980 82750
rect 7020 82550 7090 82750
rect 7410 82550 7480 82750
rect 7520 82550 7590 82750
rect 7910 82550 7980 82750
rect 8020 82550 8090 82750
rect 8410 82550 8480 82750
rect 8520 82550 8590 82750
rect 8910 82550 8980 82750
rect 9020 82550 9090 82750
rect 9410 82550 9480 82750
rect 9520 82550 9590 82750
rect 9910 82550 9980 82750
rect 10020 82550 10090 82750
rect 10410 82550 10480 82750
rect 10520 82550 10590 82750
rect 10910 82550 10980 82750
rect 11020 82550 11090 82750
rect 11410 82550 11480 82750
rect 11520 82550 11590 82750
rect 11910 82550 11980 82750
rect 12020 82550 12090 82750
rect 12410 82550 12480 82750
rect 12520 82550 12590 82750
rect 12910 82550 12980 82750
rect 13020 82550 13090 82750
rect 13410 82550 13480 82750
rect 13520 82550 13590 82750
rect 13910 82550 13980 82750
rect 14020 82550 14090 82750
rect 14410 82550 14480 82750
rect 14520 82550 14590 82750
rect 14910 82550 14980 82750
rect 15020 82550 15090 82750
rect 15410 82550 15480 82750
rect 15520 82550 15590 82750
rect 15910 82550 15980 82750
rect 16020 82550 16090 82750
rect 16410 82550 16480 82750
rect 16520 82550 16590 82750
rect 16910 82550 16980 82750
rect 17020 82550 17090 82750
rect 17410 82550 17480 82750
rect 17520 82550 17590 82750
rect 17910 82550 17980 82750
rect 18020 82550 18090 82750
rect 18410 82550 18480 82750
rect 18520 82550 18590 82750
rect 18910 82550 18980 82750
rect 19020 82550 19090 82750
rect 19410 82550 19480 82750
rect 19520 82550 19590 82750
rect 19910 82550 19980 82750
rect 20020 82550 20090 82750
rect 20410 82550 20480 82750
rect 20520 82550 20590 82750
rect 20910 82550 20980 82750
rect 21020 82550 21090 82750
rect 21410 82550 21480 82750
rect 21520 82550 21590 82750
rect 21910 82550 21980 82750
rect 22020 82550 22090 82750
rect 22410 82550 22480 82750
rect 22520 82550 22590 82750
rect 22910 82550 22980 82750
rect 23020 82550 23090 82750
rect 23410 82550 23480 82750
rect 23520 82550 23590 82750
rect 23910 82550 23980 82750
rect 24020 82550 24090 82750
rect 24410 82550 24480 82750
rect 24520 82550 24590 82750
rect 24910 82550 24980 82750
rect 25020 82550 25090 82750
rect 25410 82550 25480 82750
rect 25520 82550 25590 82750
rect 25910 82550 25980 82750
rect 26020 82550 26090 82750
rect 26410 82550 26480 82750
rect 26520 82550 26590 82750
rect 26910 82550 26980 82750
rect 27020 82550 27090 82750
rect 27410 82550 27480 82750
rect 27520 82550 27590 82750
rect 27910 82550 27980 82750
rect 28020 82550 28090 82750
rect 28410 82550 28480 82750
rect 28520 82550 28590 82750
rect 28910 82550 28980 82750
rect 29020 82550 29090 82750
rect 29410 82550 29480 82750
rect 29520 82550 29590 82750
rect 29910 82550 29980 82750
rect 30020 82550 30090 82750
rect 30410 82550 30480 82750
rect 30520 82550 30590 82750
rect 30910 82550 30980 82750
rect 31020 82550 31090 82750
rect 31410 82550 31480 82750
rect 31520 82550 31590 82750
rect 31910 82550 31980 82750
rect 32020 82550 32090 82750
rect 32410 82550 32480 82750
rect 32520 82550 32590 82750
rect 32910 82550 32980 82750
rect 33020 82550 33090 82750
rect 33410 82550 33480 82750
rect 33520 82550 33590 82750
rect 33910 82550 33980 82750
rect 34020 82550 34090 82750
rect 34410 82550 34480 82750
rect 34520 82550 34590 82750
rect 34910 82550 34980 82750
rect 35020 82550 35090 82750
rect 35410 82550 35480 82750
rect 35520 82550 35590 82750
rect 35910 82550 35980 82750
rect 36020 82550 36090 82750
rect 36410 82550 36480 82750
rect 36520 82550 36590 82750
rect 36910 82550 36980 82750
rect 37020 82550 37090 82750
rect 37410 82550 37480 82750
rect 37520 82550 37590 82750
rect 37910 82550 37980 82750
rect 38020 82550 38090 82750
rect 38410 82550 38480 82750
rect 38520 82550 38590 82750
rect 38910 82550 38980 82750
rect 39020 82550 39090 82750
rect 39410 82550 39480 82750
rect 39520 82550 39590 82750
rect 39910 82550 39980 82750
rect 40020 82550 40090 82750
rect 40410 82550 40480 82750
rect 40520 82550 40590 82750
rect 40910 82550 40980 82750
rect 41020 82550 41090 82750
rect 41410 82550 41480 82750
rect 41520 82550 41590 82750
rect 41910 82550 41980 82750
rect 42020 82550 42090 82750
rect 42410 82550 42480 82750
rect 42520 82550 42590 82750
rect 42910 82550 42980 82750
rect 43020 82550 43090 82750
rect 43410 82550 43480 82750
rect 43520 82550 43590 82750
rect 43910 82550 43980 82750
rect 44020 82550 44090 82750
rect 44410 82550 44480 82750
rect 44520 82550 44590 82750
rect 44910 82550 44980 82750
rect 45020 82550 45090 82750
rect 45410 82550 45480 82750
rect 45520 82550 45590 82750
rect 45910 82550 45980 82750
rect 46020 82550 46090 82750
rect 46410 82550 46480 82750
rect 46520 82550 46590 82750
rect 46910 82550 46980 82750
rect 47020 82550 47090 82750
rect 47410 82550 47480 82750
rect 47520 82550 47590 82750
rect 47910 82550 47980 82750
rect 48020 82550 48090 82750
rect 48410 82550 48480 82750
rect 48520 82550 48590 82750
rect 48910 82550 48980 82750
rect 49020 82550 49090 82750
rect 49410 82550 49480 82750
rect 49520 82550 49590 82750
rect 49910 82550 49980 82750
rect 50020 82550 50090 82750
rect 50410 82550 50480 82750
rect 50520 82550 50590 82750
rect 50910 82550 50980 82750
rect 51020 82550 51090 82750
rect 51410 82550 51480 82750
rect 51520 82550 51590 82750
rect 51910 82550 51980 82750
rect 52020 82550 52090 82750
rect 52410 82550 52480 82750
rect 52520 82550 52590 82750
rect 52910 82550 52980 82750
rect 53020 82550 53090 82750
rect 53410 82550 53480 82750
rect 53520 82550 53590 82750
rect 53910 82550 53980 82750
rect 54020 82550 54090 82750
rect 54410 82550 54480 82750
rect 54520 82550 54590 82750
rect 54910 82550 54980 82750
rect 55020 82550 55090 82750
rect 55410 82550 55480 82750
rect 55520 82550 55590 82750
rect 55910 82550 55980 82750
rect 56020 82550 56090 82750
rect 56410 82550 56480 82750
rect 56520 82550 56590 82750
rect 56910 82550 56980 82750
rect 57020 82550 57090 82750
rect 57410 82550 57480 82750
rect 57520 82550 57590 82750
rect 57910 82550 57980 82750
rect 58020 82550 58090 82750
rect 58410 82550 58480 82750
rect 58520 82550 58590 82750
rect 58910 82550 58980 82750
rect 59020 82550 59090 82750
rect 59410 82550 59480 82750
rect 59520 82550 59590 82750
rect 59910 82550 59980 82750
rect 60020 82550 60090 82750
rect 60410 82550 60480 82750
rect 60520 82550 60590 82750
rect 60910 82550 60980 82750
rect 61020 82550 61090 82750
rect 61410 82550 61480 82750
rect 61520 82550 61590 82750
rect 61910 82550 61980 82750
rect 62020 82550 62090 82750
rect 62410 82550 62480 82750
rect 62520 82550 62590 82750
rect 62910 82550 62980 82750
rect 63020 82550 63090 82750
rect 63410 82550 63480 82750
rect 63520 82550 63590 82750
rect 63910 82550 63980 82750
rect 64020 82550 64090 82750
rect 64410 82550 64480 82750
rect 64520 82550 64590 82750
rect 64910 82550 64980 82750
rect 65020 82550 65090 82750
rect 65410 82550 65480 82750
rect 65520 82550 65590 82750
rect 65910 82550 65980 82750
rect 66020 82550 66090 82750
rect 66410 82550 66480 82750
rect 66520 82550 66590 82750
rect 66910 82550 66980 82750
rect 67020 82550 67090 82750
rect 67410 82550 67480 82750
rect 67520 82550 67590 82750
rect 67910 82550 67980 82750
rect 68020 82550 68090 82750
rect 68410 82550 68480 82750
rect 68520 82550 68590 82750
rect 68910 82550 68980 82750
rect 69020 82550 69090 82750
rect 69410 82550 69480 82750
rect 69520 82550 69590 82750
rect 69910 82550 69980 82750
rect 70020 82550 70090 82750
rect 70410 82550 70480 82750
rect 70520 82550 70590 82750
rect 70910 82550 70980 82750
rect 71020 82550 71090 82750
rect 71410 82550 71480 82750
rect 71520 82550 71590 82750
rect 71910 82550 71980 82750
rect 72020 82550 72090 82750
rect 72410 82550 72480 82750
rect 72520 82550 72590 82750
rect 72910 82550 72980 82750
rect 73020 82550 73090 82750
rect 73410 82550 73480 82750
rect 73520 82550 73590 82750
rect 73910 82550 73980 82750
rect 74020 82550 74090 82750
rect 74410 82550 74480 82750
rect 74520 82550 74590 82750
rect 74910 82550 74980 82750
rect 75020 82550 75090 82750
rect 75410 82550 75480 82750
rect 75520 82550 75590 82750
rect 75910 82550 75980 82750
rect 76020 82550 76090 82750
rect 76410 82550 76480 82750
rect 76520 82550 76590 82750
rect 76910 82550 76980 82750
rect 77020 82550 77090 82750
rect 77410 82550 77480 82750
rect 77520 82550 77590 82750
rect 77910 82550 77980 82750
rect 78020 82550 78090 82750
rect 78410 82550 78480 82750
rect 78520 82550 78590 82750
rect 78910 82550 78980 82750
rect 79020 82550 79090 82750
rect 79410 82550 79480 82750
rect 79520 82550 79590 82750
rect 79910 82550 79980 82750
rect 80020 82550 80090 82750
rect 80410 82550 80480 82750
rect 80520 82550 80590 82750
rect 80910 82550 80980 82750
rect 81020 82550 81090 82750
rect 81410 82550 81480 82750
rect 81520 82550 81590 82750
rect 81910 82550 81980 82750
rect 82020 82550 82090 82750
rect 82410 82550 82480 82750
rect 82520 82550 82590 82750
rect 82910 82550 82980 82750
rect 83020 82550 83090 82750
rect 83410 82550 83480 82750
rect 83520 82550 83590 82750
rect 83910 82550 83980 82750
rect 84020 82550 84090 82750
rect 84410 82550 84480 82750
rect 84520 82550 84590 82750
rect 84910 82550 84980 82750
rect 85020 82550 85090 82750
rect 85410 82550 85480 82750
rect 85520 82550 85590 82750
rect 85910 82550 85980 82750
rect 86020 82550 86090 82750
rect 86410 82550 86480 82750
rect 86520 82550 86590 82750
rect 86910 82550 86980 82750
rect 87020 82550 87090 82750
rect 87410 82550 87480 82750
rect 87520 82550 87590 82750
rect 87910 82550 87980 82750
rect 88020 82550 88090 82750
rect 88410 82550 88480 82750
rect 88520 82550 88590 82750
rect 88910 82550 88980 82750
rect 89020 82550 89090 82750
rect 89410 82550 89480 82750
rect 89520 82550 89590 82750
rect 89910 82550 89980 82750
rect 90020 82550 90090 82750
rect 90410 82550 90480 82750
rect 90520 82550 90590 82750
rect 90910 82550 90980 82750
rect 91020 82550 91090 82750
rect 91410 82550 91480 82750
rect 91520 82550 91590 82750
rect 91910 82550 91980 82750
rect 92020 82550 92090 82750
rect 92410 82550 92480 82750
rect 92520 82550 92590 82750
rect 92910 82550 92980 82750
rect 93020 82550 93090 82750
rect 93410 82550 93480 82750
rect 93520 82550 93590 82750
rect 93910 82550 93980 82750
rect 94020 82550 94090 82750
rect 94410 82550 94480 82750
rect 94520 82550 94590 82750
rect 94910 82550 94980 82750
rect 95020 82550 95090 82750
rect 95410 82550 95480 82750
rect 95520 82550 95590 82750
rect 95910 82550 95980 82750
rect 96020 82550 96090 82750
rect 96410 82550 96480 82750
rect 96520 82550 96590 82750
rect 96910 82550 96980 82750
rect 97020 82550 97090 82750
rect 97410 82550 97480 82750
rect 97520 82550 97590 82750
rect 97910 82550 97980 82750
rect 98020 82550 98090 82750
rect 98410 82550 98480 82750
rect 98520 82550 98590 82750
rect 98910 82550 98980 82750
rect 99020 82550 99090 82750
rect 99410 82550 99480 82750
rect 99520 82550 99590 82750
rect 99910 82550 99980 82750
rect 100020 82550 100090 82750
rect 100410 82550 100480 82750
rect -83350 82420 -83150 82490
rect -82850 82420 -82650 82490
rect -82350 82420 -82150 82490
rect -81850 82420 -81650 82490
rect -81350 82420 -81150 82490
rect -80850 82420 -80650 82490
rect -80350 82420 -80150 82490
rect -79850 82420 -79650 82490
rect -79350 82420 -79150 82490
rect -78850 82420 -78650 82490
rect -78350 82420 -78150 82490
rect -77850 82420 -77650 82490
rect -77350 82420 -77150 82490
rect -76850 82420 -76650 82490
rect -76350 82420 -76150 82490
rect -75850 82420 -75650 82490
rect -75350 82420 -75150 82490
rect -74850 82420 -74650 82490
rect -74350 82420 -74150 82490
rect -73850 82420 -73650 82490
rect -73350 82420 -73150 82490
rect -72850 82420 -72650 82490
rect -72350 82420 -72150 82490
rect -71850 82420 -71650 82490
rect -71350 82420 -71150 82490
rect -70850 82420 -70650 82490
rect -70350 82420 -70150 82490
rect -69850 82420 -69650 82490
rect -69350 82420 -69150 82490
rect -68850 82420 -68650 82490
rect -68350 82420 -68150 82490
rect -67850 82420 -67650 82490
rect -67350 82420 -67150 82490
rect -66850 82420 -66650 82490
rect -66350 82420 -66150 82490
rect -65850 82420 -65650 82490
rect -65350 82420 -65150 82490
rect -64850 82420 -64650 82490
rect -64350 82420 -64150 82490
rect -63850 82420 -63650 82490
rect -63350 82420 -63150 82490
rect -62850 82420 -62650 82490
rect -62350 82420 -62150 82490
rect -61850 82420 -61650 82490
rect -61350 82420 -61150 82490
rect -60850 82420 -60650 82490
rect -60350 82420 -60150 82490
rect -59850 82420 -59650 82490
rect -59350 82420 -59150 82490
rect -58850 82420 -58650 82490
rect -58350 82420 -58150 82490
rect -57850 82420 -57650 82490
rect -57350 82420 -57150 82490
rect -56850 82420 -56650 82490
rect -56350 82420 -56150 82490
rect -55850 82420 -55650 82490
rect -55350 82420 -55150 82490
rect -54850 82420 -54650 82490
rect -54350 82420 -54150 82490
rect -53850 82420 -53650 82490
rect -53350 82420 -53150 82490
rect -52850 82420 -52650 82490
rect -52350 82420 -52150 82490
rect -51850 82420 -51650 82490
rect -51350 82420 -51150 82490
rect -50850 82420 -50650 82490
rect -50350 82420 -50150 82490
rect -49850 82420 -49650 82490
rect -49350 82420 -49150 82490
rect -48850 82420 -48650 82490
rect -48350 82420 -48150 82490
rect -47850 82420 -47650 82490
rect -47350 82420 -47150 82490
rect -46850 82420 -46650 82490
rect -46350 82420 -46150 82490
rect -45850 82420 -45650 82490
rect -45350 82420 -45150 82490
rect -44850 82420 -44650 82490
rect -44350 82420 -44150 82490
rect -43850 82420 -43650 82490
rect -43350 82420 -43150 82490
rect -42850 82420 -42650 82490
rect -42350 82420 -42150 82490
rect -41850 82420 -41650 82490
rect -41350 82420 -41150 82490
rect -40850 82420 -40650 82490
rect -40350 82420 -40150 82490
rect -39850 82420 -39650 82490
rect -39350 82420 -39150 82490
rect -38850 82420 -38650 82490
rect -38350 82420 -38150 82490
rect -37850 82420 -37650 82490
rect -37350 82420 -37150 82490
rect -36850 82420 -36650 82490
rect -36350 82420 -36150 82490
rect -35850 82420 -35650 82490
rect -35350 82420 -35150 82490
rect -34850 82420 -34650 82490
rect -34350 82420 -34150 82490
rect -33850 82420 -33650 82490
rect -33350 82420 -33150 82490
rect -32850 82420 -32650 82490
rect -32350 82420 -32150 82490
rect -31850 82420 -31650 82490
rect -31350 82420 -31150 82490
rect -30850 82420 -30650 82490
rect -30350 82420 -30150 82490
rect -29850 82420 -29650 82490
rect -29350 82420 -29150 82490
rect -28850 82420 -28650 82490
rect -28350 82420 -28150 82490
rect -27850 82420 -27650 82490
rect -27350 82420 -27150 82490
rect -26850 82420 -26650 82490
rect -26350 82420 -26150 82490
rect -25850 82420 -25650 82490
rect -25350 82420 -25150 82490
rect -24850 82420 -24650 82490
rect -24350 82420 -24150 82490
rect -23850 82420 -23650 82490
rect -23350 82420 -23150 82490
rect -22850 82420 -22650 82490
rect -22350 82420 -22150 82490
rect -21850 82420 -21650 82490
rect -21350 82420 -21150 82490
rect -20850 82420 -20650 82490
rect -20350 82420 -20150 82490
rect -19850 82420 -19650 82490
rect -19350 82420 -19150 82490
rect -18850 82420 -18650 82490
rect -18350 82420 -18150 82490
rect -17850 82420 -17650 82490
rect -17350 82420 -17150 82490
rect -16850 82420 -16650 82490
rect -16350 82420 -16150 82490
rect -15850 82420 -15650 82490
rect -15350 82420 -15150 82490
rect -14850 82420 -14650 82490
rect -14350 82420 -14150 82490
rect -13850 82420 -13650 82490
rect -13350 82420 -13150 82490
rect -12850 82420 -12650 82490
rect -12350 82420 -12150 82490
rect -11850 82420 -11650 82490
rect -11350 82420 -11150 82490
rect -10850 82420 -10650 82490
rect -10350 82420 -10150 82490
rect -9850 82420 -9650 82490
rect -9350 82420 -9150 82490
rect -8850 82420 -8650 82490
rect -8350 82420 -8150 82490
rect -7850 82420 -7650 82490
rect -7350 82420 -7150 82490
rect -6850 82420 -6650 82490
rect -6350 82420 -6150 82490
rect -5850 82420 -5650 82490
rect -5350 82420 -5150 82490
rect -4850 82420 -4650 82490
rect -4350 82420 -4150 82490
rect -3850 82420 -3650 82490
rect -3350 82420 -3150 82490
rect -2850 82420 -2650 82490
rect -2350 82420 -2150 82490
rect -1850 82420 -1650 82490
rect -1350 82420 -1150 82490
rect -850 82420 -650 82490
rect -350 82420 -150 82490
rect 150 82420 350 82490
rect 650 82420 850 82490
rect 1150 82420 1350 82490
rect 1650 82420 1850 82490
rect 2150 82420 2350 82490
rect 2650 82420 2850 82490
rect 3150 82420 3350 82490
rect 3650 82420 3850 82490
rect 4150 82420 4350 82490
rect 4650 82420 4850 82490
rect 5150 82420 5350 82490
rect 5650 82420 5850 82490
rect 6150 82420 6350 82490
rect 6650 82420 6850 82490
rect 7150 82420 7350 82490
rect 7650 82420 7850 82490
rect 8150 82420 8350 82490
rect 8650 82420 8850 82490
rect 9150 82420 9350 82490
rect 9650 82420 9850 82490
rect 10150 82420 10350 82490
rect 10650 82420 10850 82490
rect 11150 82420 11350 82490
rect 11650 82420 11850 82490
rect 12150 82420 12350 82490
rect 12650 82420 12850 82490
rect 13150 82420 13350 82490
rect 13650 82420 13850 82490
rect 14150 82420 14350 82490
rect 14650 82420 14850 82490
rect 15150 82420 15350 82490
rect 15650 82420 15850 82490
rect 16150 82420 16350 82490
rect 16650 82420 16850 82490
rect 17150 82420 17350 82490
rect 17650 82420 17850 82490
rect 18150 82420 18350 82490
rect 18650 82420 18850 82490
rect 19150 82420 19350 82490
rect 19650 82420 19850 82490
rect 20150 82420 20350 82490
rect 20650 82420 20850 82490
rect 21150 82420 21350 82490
rect 21650 82420 21850 82490
rect 22150 82420 22350 82490
rect 22650 82420 22850 82490
rect 23150 82420 23350 82490
rect 23650 82420 23850 82490
rect 24150 82420 24350 82490
rect 24650 82420 24850 82490
rect 25150 82420 25350 82490
rect 25650 82420 25850 82490
rect 26150 82420 26350 82490
rect 26650 82420 26850 82490
rect 27150 82420 27350 82490
rect 27650 82420 27850 82490
rect 28150 82420 28350 82490
rect 28650 82420 28850 82490
rect 29150 82420 29350 82490
rect 29650 82420 29850 82490
rect 30150 82420 30350 82490
rect 30650 82420 30850 82490
rect 31150 82420 31350 82490
rect 31650 82420 31850 82490
rect 32150 82420 32350 82490
rect 32650 82420 32850 82490
rect 33150 82420 33350 82490
rect 33650 82420 33850 82490
rect 34150 82420 34350 82490
rect 34650 82420 34850 82490
rect 35150 82420 35350 82490
rect 35650 82420 35850 82490
rect 36150 82420 36350 82490
rect 36650 82420 36850 82490
rect 37150 82420 37350 82490
rect 37650 82420 37850 82490
rect 38150 82420 38350 82490
rect 38650 82420 38850 82490
rect 39150 82420 39350 82490
rect 39650 82420 39850 82490
rect 40150 82420 40350 82490
rect 40650 82420 40850 82490
rect 41150 82420 41350 82490
rect 41650 82420 41850 82490
rect 42150 82420 42350 82490
rect 42650 82420 42850 82490
rect 43150 82420 43350 82490
rect 43650 82420 43850 82490
rect 44150 82420 44350 82490
rect 44650 82420 44850 82490
rect 45150 82420 45350 82490
rect 45650 82420 45850 82490
rect 46150 82420 46350 82490
rect 46650 82420 46850 82490
rect 47150 82420 47350 82490
rect 47650 82420 47850 82490
rect 48150 82420 48350 82490
rect 48650 82420 48850 82490
rect 49150 82420 49350 82490
rect 49650 82420 49850 82490
rect 50150 82420 50350 82490
rect 50650 82420 50850 82490
rect 51150 82420 51350 82490
rect 51650 82420 51850 82490
rect 52150 82420 52350 82490
rect 52650 82420 52850 82490
rect 53150 82420 53350 82490
rect 53650 82420 53850 82490
rect 54150 82420 54350 82490
rect 54650 82420 54850 82490
rect 55150 82420 55350 82490
rect 55650 82420 55850 82490
rect 56150 82420 56350 82490
rect 56650 82420 56850 82490
rect 57150 82420 57350 82490
rect 57650 82420 57850 82490
rect 58150 82420 58350 82490
rect 58650 82420 58850 82490
rect 59150 82420 59350 82490
rect 59650 82420 59850 82490
rect 60150 82420 60350 82490
rect 60650 82420 60850 82490
rect 61150 82420 61350 82490
rect 61650 82420 61850 82490
rect 62150 82420 62350 82490
rect 62650 82420 62850 82490
rect 63150 82420 63350 82490
rect 63650 82420 63850 82490
rect 64150 82420 64350 82490
rect 64650 82420 64850 82490
rect 65150 82420 65350 82490
rect 65650 82420 65850 82490
rect 66150 82420 66350 82490
rect 66650 82420 66850 82490
rect 67150 82420 67350 82490
rect 67650 82420 67850 82490
rect 68150 82420 68350 82490
rect 68650 82420 68850 82490
rect 69150 82420 69350 82490
rect 69650 82420 69850 82490
rect 70150 82420 70350 82490
rect 70650 82420 70850 82490
rect 71150 82420 71350 82490
rect 71650 82420 71850 82490
rect 72150 82420 72350 82490
rect 72650 82420 72850 82490
rect 73150 82420 73350 82490
rect 73650 82420 73850 82490
rect 74150 82420 74350 82490
rect 74650 82420 74850 82490
rect 75150 82420 75350 82490
rect 75650 82420 75850 82490
rect 76150 82420 76350 82490
rect 76650 82420 76850 82490
rect 77150 82420 77350 82490
rect 77650 82420 77850 82490
rect 78150 82420 78350 82490
rect 78650 82420 78850 82490
rect 79150 82420 79350 82490
rect 79650 82420 79850 82490
rect 80150 82420 80350 82490
rect 80650 82420 80850 82490
rect 81150 82420 81350 82490
rect 81650 82420 81850 82490
rect 82150 82420 82350 82490
rect 82650 82420 82850 82490
rect 83150 82420 83350 82490
rect 83650 82420 83850 82490
rect 84150 82420 84350 82490
rect 84650 82420 84850 82490
rect 85150 82420 85350 82490
rect 85650 82420 85850 82490
rect 86150 82420 86350 82490
rect 86650 82420 86850 82490
rect 87150 82420 87350 82490
rect 87650 82420 87850 82490
rect 88150 82420 88350 82490
rect 88650 82420 88850 82490
rect 89150 82420 89350 82490
rect 89650 82420 89850 82490
rect 90150 82420 90350 82490
rect 90650 82420 90850 82490
rect 91150 82420 91350 82490
rect 91650 82420 91850 82490
rect 92150 82420 92350 82490
rect 92650 82420 92850 82490
rect 93150 82420 93350 82490
rect 93650 82420 93850 82490
rect 94150 82420 94350 82490
rect 94650 82420 94850 82490
rect 95150 82420 95350 82490
rect 95650 82420 95850 82490
rect 96150 82420 96350 82490
rect 96650 82420 96850 82490
rect 97150 82420 97350 82490
rect 97650 82420 97850 82490
rect 98150 82420 98350 82490
rect 98650 82420 98850 82490
rect 99150 82420 99350 82490
rect 99650 82420 99850 82490
rect 100150 82420 100350 82490
rect -83350 82310 -83150 82380
rect -82850 82310 -82650 82380
rect -82350 82310 -82150 82380
rect -81850 82310 -81650 82380
rect -81350 82310 -81150 82380
rect -80850 82310 -80650 82380
rect -80350 82310 -80150 82380
rect -79850 82310 -79650 82380
rect -79350 82310 -79150 82380
rect -78850 82310 -78650 82380
rect -78350 82310 -78150 82380
rect -77850 82310 -77650 82380
rect -77350 82310 -77150 82380
rect -76850 82310 -76650 82380
rect -76350 82310 -76150 82380
rect -75850 82310 -75650 82380
rect -75350 82310 -75150 82380
rect -74850 82310 -74650 82380
rect -74350 82310 -74150 82380
rect -73850 82310 -73650 82380
rect -73350 82310 -73150 82380
rect -72850 82310 -72650 82380
rect -72350 82310 -72150 82380
rect -71850 82310 -71650 82380
rect -71350 82310 -71150 82380
rect -70850 82310 -70650 82380
rect -70350 82310 -70150 82380
rect -69850 82310 -69650 82380
rect -69350 82310 -69150 82380
rect -68850 82310 -68650 82380
rect -68350 82310 -68150 82380
rect -67850 82310 -67650 82380
rect -67350 82310 -67150 82380
rect -66850 82310 -66650 82380
rect -66350 82310 -66150 82380
rect -65850 82310 -65650 82380
rect -65350 82310 -65150 82380
rect -64850 82310 -64650 82380
rect -64350 82310 -64150 82380
rect -63850 82310 -63650 82380
rect -63350 82310 -63150 82380
rect -62850 82310 -62650 82380
rect -62350 82310 -62150 82380
rect -61850 82310 -61650 82380
rect -61350 82310 -61150 82380
rect -60850 82310 -60650 82380
rect -60350 82310 -60150 82380
rect -59850 82310 -59650 82380
rect -59350 82310 -59150 82380
rect -58850 82310 -58650 82380
rect -58350 82310 -58150 82380
rect -57850 82310 -57650 82380
rect -57350 82310 -57150 82380
rect -56850 82310 -56650 82380
rect -56350 82310 -56150 82380
rect -55850 82310 -55650 82380
rect -55350 82310 -55150 82380
rect -54850 82310 -54650 82380
rect -54350 82310 -54150 82380
rect -53850 82310 -53650 82380
rect -53350 82310 -53150 82380
rect -52850 82310 -52650 82380
rect -52350 82310 -52150 82380
rect -51850 82310 -51650 82380
rect -51350 82310 -51150 82380
rect -50850 82310 -50650 82380
rect -50350 82310 -50150 82380
rect -49850 82310 -49650 82380
rect -49350 82310 -49150 82380
rect -48850 82310 -48650 82380
rect -48350 82310 -48150 82380
rect -47850 82310 -47650 82380
rect -47350 82310 -47150 82380
rect -46850 82310 -46650 82380
rect -46350 82310 -46150 82380
rect -45850 82310 -45650 82380
rect -45350 82310 -45150 82380
rect -44850 82310 -44650 82380
rect -44350 82310 -44150 82380
rect -43850 82310 -43650 82380
rect -43350 82310 -43150 82380
rect -42850 82310 -42650 82380
rect -42350 82310 -42150 82380
rect -41850 82310 -41650 82380
rect -41350 82310 -41150 82380
rect -40850 82310 -40650 82380
rect -40350 82310 -40150 82380
rect -39850 82310 -39650 82380
rect -39350 82310 -39150 82380
rect -38850 82310 -38650 82380
rect -38350 82310 -38150 82380
rect -37850 82310 -37650 82380
rect -37350 82310 -37150 82380
rect -36850 82310 -36650 82380
rect -36350 82310 -36150 82380
rect -35850 82310 -35650 82380
rect -35350 82310 -35150 82380
rect -34850 82310 -34650 82380
rect -34350 82310 -34150 82380
rect -33850 82310 -33650 82380
rect -33350 82310 -33150 82380
rect -32850 82310 -32650 82380
rect -32350 82310 -32150 82380
rect -31850 82310 -31650 82380
rect -31350 82310 -31150 82380
rect -30850 82310 -30650 82380
rect -30350 82310 -30150 82380
rect -29850 82310 -29650 82380
rect -29350 82310 -29150 82380
rect -28850 82310 -28650 82380
rect -28350 82310 -28150 82380
rect -27850 82310 -27650 82380
rect -27350 82310 -27150 82380
rect -26850 82310 -26650 82380
rect -26350 82310 -26150 82380
rect -25850 82310 -25650 82380
rect -25350 82310 -25150 82380
rect -24850 82310 -24650 82380
rect -24350 82310 -24150 82380
rect -23850 82310 -23650 82380
rect -23350 82310 -23150 82380
rect -22850 82310 -22650 82380
rect -22350 82310 -22150 82380
rect -21850 82310 -21650 82380
rect -21350 82310 -21150 82380
rect -20850 82310 -20650 82380
rect -20350 82310 -20150 82380
rect -19850 82310 -19650 82380
rect -19350 82310 -19150 82380
rect -18850 82310 -18650 82380
rect -18350 82310 -18150 82380
rect -17850 82310 -17650 82380
rect -17350 82310 -17150 82380
rect -16850 82310 -16650 82380
rect -16350 82310 -16150 82380
rect -15850 82310 -15650 82380
rect -15350 82310 -15150 82380
rect -14850 82310 -14650 82380
rect -14350 82310 -14150 82380
rect -13850 82310 -13650 82380
rect -13350 82310 -13150 82380
rect -12850 82310 -12650 82380
rect -12350 82310 -12150 82380
rect -11850 82310 -11650 82380
rect -11350 82310 -11150 82380
rect -10850 82310 -10650 82380
rect -10350 82310 -10150 82380
rect -9850 82310 -9650 82380
rect -9350 82310 -9150 82380
rect -8850 82310 -8650 82380
rect -8350 82310 -8150 82380
rect -7850 82310 -7650 82380
rect -7350 82310 -7150 82380
rect -6850 82310 -6650 82380
rect -6350 82310 -6150 82380
rect -5850 82310 -5650 82380
rect -5350 82310 -5150 82380
rect -4850 82310 -4650 82380
rect -4350 82310 -4150 82380
rect -3850 82310 -3650 82380
rect -3350 82310 -3150 82380
rect -2850 82310 -2650 82380
rect -2350 82310 -2150 82380
rect -1850 82310 -1650 82380
rect -1350 82310 -1150 82380
rect -850 82310 -650 82380
rect -350 82310 -150 82380
rect 150 82310 350 82380
rect 650 82310 850 82380
rect 1150 82310 1350 82380
rect 1650 82310 1850 82380
rect 2150 82310 2350 82380
rect 2650 82310 2850 82380
rect 3150 82310 3350 82380
rect 3650 82310 3850 82380
rect 4150 82310 4350 82380
rect 4650 82310 4850 82380
rect 5150 82310 5350 82380
rect 5650 82310 5850 82380
rect 6150 82310 6350 82380
rect 6650 82310 6850 82380
rect 7150 82310 7350 82380
rect 7650 82310 7850 82380
rect 8150 82310 8350 82380
rect 8650 82310 8850 82380
rect 9150 82310 9350 82380
rect 9650 82310 9850 82380
rect 10150 82310 10350 82380
rect 10650 82310 10850 82380
rect 11150 82310 11350 82380
rect 11650 82310 11850 82380
rect 12150 82310 12350 82380
rect 12650 82310 12850 82380
rect 13150 82310 13350 82380
rect 13650 82310 13850 82380
rect 14150 82310 14350 82380
rect 14650 82310 14850 82380
rect 15150 82310 15350 82380
rect 15650 82310 15850 82380
rect 16150 82310 16350 82380
rect 16650 82310 16850 82380
rect 17150 82310 17350 82380
rect 17650 82310 17850 82380
rect 18150 82310 18350 82380
rect 18650 82310 18850 82380
rect 19150 82310 19350 82380
rect 19650 82310 19850 82380
rect 20150 82310 20350 82380
rect 20650 82310 20850 82380
rect 21150 82310 21350 82380
rect 21650 82310 21850 82380
rect 22150 82310 22350 82380
rect 22650 82310 22850 82380
rect 23150 82310 23350 82380
rect 23650 82310 23850 82380
rect 24150 82310 24350 82380
rect 24650 82310 24850 82380
rect 25150 82310 25350 82380
rect 25650 82310 25850 82380
rect 26150 82310 26350 82380
rect 26650 82310 26850 82380
rect 27150 82310 27350 82380
rect 27650 82310 27850 82380
rect 28150 82310 28350 82380
rect 28650 82310 28850 82380
rect 29150 82310 29350 82380
rect 29650 82310 29850 82380
rect 30150 82310 30350 82380
rect 30650 82310 30850 82380
rect 31150 82310 31350 82380
rect 31650 82310 31850 82380
rect 32150 82310 32350 82380
rect 32650 82310 32850 82380
rect 33150 82310 33350 82380
rect 33650 82310 33850 82380
rect 34150 82310 34350 82380
rect 34650 82310 34850 82380
rect 35150 82310 35350 82380
rect 35650 82310 35850 82380
rect 36150 82310 36350 82380
rect 36650 82310 36850 82380
rect 37150 82310 37350 82380
rect 37650 82310 37850 82380
rect 38150 82310 38350 82380
rect 38650 82310 38850 82380
rect 39150 82310 39350 82380
rect 39650 82310 39850 82380
rect 40150 82310 40350 82380
rect 40650 82310 40850 82380
rect 41150 82310 41350 82380
rect 41650 82310 41850 82380
rect 42150 82310 42350 82380
rect 42650 82310 42850 82380
rect 43150 82310 43350 82380
rect 43650 82310 43850 82380
rect 44150 82310 44350 82380
rect 44650 82310 44850 82380
rect 45150 82310 45350 82380
rect 45650 82310 45850 82380
rect 46150 82310 46350 82380
rect 46650 82310 46850 82380
rect 47150 82310 47350 82380
rect 47650 82310 47850 82380
rect 48150 82310 48350 82380
rect 48650 82310 48850 82380
rect 49150 82310 49350 82380
rect 49650 82310 49850 82380
rect 50150 82310 50350 82380
rect 50650 82310 50850 82380
rect 51150 82310 51350 82380
rect 51650 82310 51850 82380
rect 52150 82310 52350 82380
rect 52650 82310 52850 82380
rect 53150 82310 53350 82380
rect 53650 82310 53850 82380
rect 54150 82310 54350 82380
rect 54650 82310 54850 82380
rect 55150 82310 55350 82380
rect 55650 82310 55850 82380
rect 56150 82310 56350 82380
rect 56650 82310 56850 82380
rect 57150 82310 57350 82380
rect 57650 82310 57850 82380
rect 58150 82310 58350 82380
rect 58650 82310 58850 82380
rect 59150 82310 59350 82380
rect 59650 82310 59850 82380
rect 60150 82310 60350 82380
rect 60650 82310 60850 82380
rect 61150 82310 61350 82380
rect 61650 82310 61850 82380
rect 62150 82310 62350 82380
rect 62650 82310 62850 82380
rect 63150 82310 63350 82380
rect 63650 82310 63850 82380
rect 64150 82310 64350 82380
rect 64650 82310 64850 82380
rect 65150 82310 65350 82380
rect 65650 82310 65850 82380
rect 66150 82310 66350 82380
rect 66650 82310 66850 82380
rect 67150 82310 67350 82380
rect 67650 82310 67850 82380
rect 68150 82310 68350 82380
rect 68650 82310 68850 82380
rect 69150 82310 69350 82380
rect 69650 82310 69850 82380
rect 70150 82310 70350 82380
rect 70650 82310 70850 82380
rect 71150 82310 71350 82380
rect 71650 82310 71850 82380
rect 72150 82310 72350 82380
rect 72650 82310 72850 82380
rect 73150 82310 73350 82380
rect 73650 82310 73850 82380
rect 74150 82310 74350 82380
rect 74650 82310 74850 82380
rect 75150 82310 75350 82380
rect 75650 82310 75850 82380
rect 76150 82310 76350 82380
rect 76650 82310 76850 82380
rect 77150 82310 77350 82380
rect 77650 82310 77850 82380
rect 78150 82310 78350 82380
rect 78650 82310 78850 82380
rect 79150 82310 79350 82380
rect 79650 82310 79850 82380
rect 80150 82310 80350 82380
rect 80650 82310 80850 82380
rect 81150 82310 81350 82380
rect 81650 82310 81850 82380
rect 82150 82310 82350 82380
rect 82650 82310 82850 82380
rect 83150 82310 83350 82380
rect 83650 82310 83850 82380
rect 84150 82310 84350 82380
rect 84650 82310 84850 82380
rect 85150 82310 85350 82380
rect 85650 82310 85850 82380
rect 86150 82310 86350 82380
rect 86650 82310 86850 82380
rect 87150 82310 87350 82380
rect 87650 82310 87850 82380
rect 88150 82310 88350 82380
rect 88650 82310 88850 82380
rect 89150 82310 89350 82380
rect 89650 82310 89850 82380
rect 90150 82310 90350 82380
rect 90650 82310 90850 82380
rect 91150 82310 91350 82380
rect 91650 82310 91850 82380
rect 92150 82310 92350 82380
rect 92650 82310 92850 82380
rect 93150 82310 93350 82380
rect 93650 82310 93850 82380
rect 94150 82310 94350 82380
rect 94650 82310 94850 82380
rect 95150 82310 95350 82380
rect 95650 82310 95850 82380
rect 96150 82310 96350 82380
rect 96650 82310 96850 82380
rect 97150 82310 97350 82380
rect 97650 82310 97850 82380
rect 98150 82310 98350 82380
rect 98650 82310 98850 82380
rect 99150 82310 99350 82380
rect 99650 82310 99850 82380
rect 100150 82310 100350 82380
rect -83480 82050 -83410 82250
rect -83090 82050 -83020 82250
rect -82980 82050 -82910 82250
rect -82590 82050 -82520 82250
rect -82480 82050 -82410 82250
rect -82090 82050 -82020 82250
rect -81980 82050 -81910 82250
rect -81590 82050 -81520 82250
rect -81480 82050 -81410 82250
rect -81090 82050 -81020 82250
rect -80980 82050 -80910 82250
rect -80590 82050 -80520 82250
rect -80480 82050 -80410 82250
rect -80090 82050 -80020 82250
rect -79980 82050 -79910 82250
rect -79590 82050 -79520 82250
rect -79480 82050 -79410 82250
rect -79090 82050 -79020 82250
rect -78980 82050 -78910 82250
rect -78590 82050 -78520 82250
rect -78480 82050 -78410 82250
rect -78090 82050 -78020 82250
rect -77980 82050 -77910 82250
rect -77590 82050 -77520 82250
rect -77480 82050 -77410 82250
rect -77090 82050 -77020 82250
rect -76980 82050 -76910 82250
rect -76590 82050 -76520 82250
rect -76480 82050 -76410 82250
rect -76090 82050 -76020 82250
rect -75980 82050 -75910 82250
rect -75590 82050 -75520 82250
rect -75480 82050 -75410 82250
rect -75090 82050 -75020 82250
rect -74980 82050 -74910 82250
rect -74590 82050 -74520 82250
rect -74480 82050 -74410 82250
rect -74090 82050 -74020 82250
rect -73980 82050 -73910 82250
rect -73590 82050 -73520 82250
rect -73480 82050 -73410 82250
rect -73090 82050 -73020 82250
rect -72980 82050 -72910 82250
rect -72590 82050 -72520 82250
rect -72480 82050 -72410 82250
rect -72090 82050 -72020 82250
rect -71980 82050 -71910 82250
rect -71590 82050 -71520 82250
rect -71480 82050 -71410 82250
rect -71090 82050 -71020 82250
rect -70980 82050 -70910 82250
rect -70590 82050 -70520 82250
rect -70480 82050 -70410 82250
rect -70090 82050 -70020 82250
rect -69980 82050 -69910 82250
rect -69590 82050 -69520 82250
rect -69480 82050 -69410 82250
rect -69090 82050 -69020 82250
rect -68980 82050 -68910 82250
rect -68590 82050 -68520 82250
rect -68480 82050 -68410 82250
rect -68090 82050 -68020 82250
rect -67980 82050 -67910 82250
rect -67590 82050 -67520 82250
rect -67480 82050 -67410 82250
rect -67090 82050 -67020 82250
rect -66980 82050 -66910 82250
rect -66590 82050 -66520 82250
rect -66480 82050 -66410 82250
rect -66090 82050 -66020 82250
rect -65980 82050 -65910 82250
rect -65590 82050 -65520 82250
rect -65480 82050 -65410 82250
rect -65090 82050 -65020 82250
rect -64980 82050 -64910 82250
rect -64590 82050 -64520 82250
rect -64480 82050 -64410 82250
rect -64090 82050 -64020 82250
rect -63980 82050 -63910 82250
rect -63590 82050 -63520 82250
rect -63480 82050 -63410 82250
rect -63090 82050 -63020 82250
rect -62980 82050 -62910 82250
rect -62590 82050 -62520 82250
rect -62480 82050 -62410 82250
rect -62090 82050 -62020 82250
rect -61980 82050 -61910 82250
rect -61590 82050 -61520 82250
rect -61480 82050 -61410 82250
rect -61090 82050 -61020 82250
rect -60980 82050 -60910 82250
rect -60590 82050 -60520 82250
rect -60480 82050 -60410 82250
rect -60090 82050 -60020 82250
rect -59980 82050 -59910 82250
rect -59590 82050 -59520 82250
rect -59480 82050 -59410 82250
rect -59090 82050 -59020 82250
rect -58980 82050 -58910 82250
rect -58590 82050 -58520 82250
rect -58480 82050 -58410 82250
rect -58090 82050 -58020 82250
rect -57980 82050 -57910 82250
rect -57590 82050 -57520 82250
rect -57480 82050 -57410 82250
rect -57090 82050 -57020 82250
rect -56980 82050 -56910 82250
rect -56590 82050 -56520 82250
rect -56480 82050 -56410 82250
rect -56090 82050 -56020 82250
rect -55980 82050 -55910 82250
rect -55590 82050 -55520 82250
rect -55480 82050 -55410 82250
rect -55090 82050 -55020 82250
rect -54980 82050 -54910 82250
rect -54590 82050 -54520 82250
rect -54480 82050 -54410 82250
rect -54090 82050 -54020 82250
rect -53980 82050 -53910 82250
rect -53590 82050 -53520 82250
rect -53480 82050 -53410 82250
rect -53090 82050 -53020 82250
rect -52980 82050 -52910 82250
rect -52590 82050 -52520 82250
rect -52480 82050 -52410 82250
rect -52090 82050 -52020 82250
rect -51980 82050 -51910 82250
rect -51590 82050 -51520 82250
rect -51480 82050 -51410 82250
rect -51090 82050 -51020 82250
rect -50980 82050 -50910 82250
rect -50590 82050 -50520 82250
rect -50480 82050 -50410 82250
rect -50090 82050 -50020 82250
rect -49980 82050 -49910 82250
rect -49590 82050 -49520 82250
rect -49480 82050 -49410 82250
rect -49090 82050 -49020 82250
rect -48980 82050 -48910 82250
rect -48590 82050 -48520 82250
rect -48480 82050 -48410 82250
rect -48090 82050 -48020 82250
rect -47980 82050 -47910 82250
rect -47590 82050 -47520 82250
rect -47480 82050 -47410 82250
rect -47090 82050 -47020 82250
rect -46980 82050 -46910 82250
rect -46590 82050 -46520 82250
rect -46480 82050 -46410 82250
rect -46090 82050 -46020 82250
rect -45980 82050 -45910 82250
rect -45590 82050 -45520 82250
rect -45480 82050 -45410 82250
rect -45090 82050 -45020 82250
rect -44980 82050 -44910 82250
rect -44590 82050 -44520 82250
rect -44480 82050 -44410 82250
rect -44090 82050 -44020 82250
rect -43980 82050 -43910 82250
rect -43590 82050 -43520 82250
rect -43480 82050 -43410 82250
rect -43090 82050 -43020 82250
rect -42980 82050 -42910 82250
rect -42590 82050 -42520 82250
rect -42480 82050 -42410 82250
rect -42090 82050 -42020 82250
rect -41980 82050 -41910 82250
rect -41590 82050 -41520 82250
rect -41480 82050 -41410 82250
rect -41090 82050 -41020 82250
rect -40980 82050 -40910 82250
rect -40590 82050 -40520 82250
rect -40480 82050 -40410 82250
rect -40090 82050 -40020 82250
rect -39980 82050 -39910 82250
rect -39590 82050 -39520 82250
rect -39480 82050 -39410 82250
rect -39090 82050 -39020 82250
rect -38980 82050 -38910 82250
rect -38590 82050 -38520 82250
rect -38480 82050 -38410 82250
rect -38090 82050 -38020 82250
rect -37980 82050 -37910 82250
rect -37590 82050 -37520 82250
rect -37480 82050 -37410 82250
rect -37090 82050 -37020 82250
rect -36980 82050 -36910 82250
rect -36590 82050 -36520 82250
rect -36480 82050 -36410 82250
rect -36090 82050 -36020 82250
rect -35980 82050 -35910 82250
rect -35590 82050 -35520 82250
rect -35480 82050 -35410 82250
rect -35090 82050 -35020 82250
rect -34980 82050 -34910 82250
rect -34590 82050 -34520 82250
rect -34480 82050 -34410 82250
rect -34090 82050 -34020 82250
rect -33980 82050 -33910 82250
rect -33590 82050 -33520 82250
rect -33480 82050 -33410 82250
rect -33090 82050 -33020 82250
rect -32980 82050 -32910 82250
rect -32590 82050 -32520 82250
rect -32480 82050 -32410 82250
rect -32090 82050 -32020 82250
rect -31980 82050 -31910 82250
rect -31590 82050 -31520 82250
rect -31480 82050 -31410 82250
rect -31090 82050 -31020 82250
rect -30980 82050 -30910 82250
rect -30590 82050 -30520 82250
rect -30480 82050 -30410 82250
rect -30090 82050 -30020 82250
rect -29980 82050 -29910 82250
rect -29590 82050 -29520 82250
rect -29480 82050 -29410 82250
rect -29090 82050 -29020 82250
rect -28980 82050 -28910 82250
rect -28590 82050 -28520 82250
rect -28480 82050 -28410 82250
rect -28090 82050 -28020 82250
rect -27980 82050 -27910 82250
rect -27590 82050 -27520 82250
rect -27480 82050 -27410 82250
rect -27090 82050 -27020 82250
rect -26980 82050 -26910 82250
rect -26590 82050 -26520 82250
rect -26480 82050 -26410 82250
rect -26090 82050 -26020 82250
rect -25980 82050 -25910 82250
rect -25590 82050 -25520 82250
rect -25480 82050 -25410 82250
rect -25090 82050 -25020 82250
rect -24980 82050 -24910 82250
rect -24590 82050 -24520 82250
rect -24480 82050 -24410 82250
rect -24090 82050 -24020 82250
rect -23980 82050 -23910 82250
rect -23590 82050 -23520 82250
rect -23480 82050 -23410 82250
rect -23090 82050 -23020 82250
rect -22980 82050 -22910 82250
rect -22590 82050 -22520 82250
rect -22480 82050 -22410 82250
rect -22090 82050 -22020 82250
rect -21980 82050 -21910 82250
rect -21590 82050 -21520 82250
rect -21480 82050 -21410 82250
rect -21090 82050 -21020 82250
rect -20980 82050 -20910 82250
rect -20590 82050 -20520 82250
rect -20480 82050 -20410 82250
rect -20090 82050 -20020 82250
rect -19980 82050 -19910 82250
rect -19590 82050 -19520 82250
rect -19480 82050 -19410 82250
rect -19090 82050 -19020 82250
rect -18980 82050 -18910 82250
rect -18590 82050 -18520 82250
rect -18480 82050 -18410 82250
rect -18090 82050 -18020 82250
rect -17980 82050 -17910 82250
rect -17590 82050 -17520 82250
rect -17480 82050 -17410 82250
rect -17090 82050 -17020 82250
rect -16980 82050 -16910 82250
rect -16590 82050 -16520 82250
rect -16480 82050 -16410 82250
rect -16090 82050 -16020 82250
rect -15980 82050 -15910 82250
rect -15590 82050 -15520 82250
rect -15480 82050 -15410 82250
rect -15090 82050 -15020 82250
rect -14980 82050 -14910 82250
rect -14590 82050 -14520 82250
rect -14480 82050 -14410 82250
rect -14090 82050 -14020 82250
rect -13980 82050 -13910 82250
rect -13590 82050 -13520 82250
rect -13480 82050 -13410 82250
rect -13090 82050 -13020 82250
rect -12980 82050 -12910 82250
rect -12590 82050 -12520 82250
rect -12480 82050 -12410 82250
rect -12090 82050 -12020 82250
rect -11980 82050 -11910 82250
rect -11590 82050 -11520 82250
rect -11480 82050 -11410 82250
rect -11090 82050 -11020 82250
rect -10980 82050 -10910 82250
rect -10590 82050 -10520 82250
rect -10480 82050 -10410 82250
rect -10090 82050 -10020 82250
rect -9980 82050 -9910 82250
rect -9590 82050 -9520 82250
rect -9480 82050 -9410 82250
rect -9090 82050 -9020 82250
rect -8980 82050 -8910 82250
rect -8590 82050 -8520 82250
rect -8480 82050 -8410 82250
rect -8090 82050 -8020 82250
rect -7980 82050 -7910 82250
rect -7590 82050 -7520 82250
rect -7480 82050 -7410 82250
rect -7090 82050 -7020 82250
rect -6980 82050 -6910 82250
rect -6590 82050 -6520 82250
rect -6480 82050 -6410 82250
rect -6090 82050 -6020 82250
rect -5980 82050 -5910 82250
rect -5590 82050 -5520 82250
rect -5480 82050 -5410 82250
rect -5090 82050 -5020 82250
rect -4980 82050 -4910 82250
rect -4590 82050 -4520 82250
rect -4480 82050 -4410 82250
rect -4090 82050 -4020 82250
rect -3980 82050 -3910 82250
rect -3590 82050 -3520 82250
rect -3480 82050 -3410 82250
rect -3090 82050 -3020 82250
rect -2980 82050 -2910 82250
rect -2590 82050 -2520 82250
rect -2480 82050 -2410 82250
rect -2090 82050 -2020 82250
rect -1980 82050 -1910 82250
rect -1590 82050 -1520 82250
rect -1480 82050 -1410 82250
rect -1090 82050 -1020 82250
rect -980 82050 -910 82250
rect -590 82050 -520 82250
rect -480 82050 -410 82250
rect -90 82050 -20 82250
rect 20 82050 90 82250
rect 410 82050 480 82250
rect 520 82050 590 82250
rect 910 82050 980 82250
rect 1020 82050 1090 82250
rect 1410 82050 1480 82250
rect 1520 82050 1590 82250
rect 1910 82050 1980 82250
rect 2020 82050 2090 82250
rect 2410 82050 2480 82250
rect 2520 82050 2590 82250
rect 2910 82050 2980 82250
rect 3020 82050 3090 82250
rect 3410 82050 3480 82250
rect 3520 82050 3590 82250
rect 3910 82050 3980 82250
rect 4020 82050 4090 82250
rect 4410 82050 4480 82250
rect 4520 82050 4590 82250
rect 4910 82050 4980 82250
rect 5020 82050 5090 82250
rect 5410 82050 5480 82250
rect 5520 82050 5590 82250
rect 5910 82050 5980 82250
rect 6020 82050 6090 82250
rect 6410 82050 6480 82250
rect 6520 82050 6590 82250
rect 6910 82050 6980 82250
rect 7020 82050 7090 82250
rect 7410 82050 7480 82250
rect 7520 82050 7590 82250
rect 7910 82050 7980 82250
rect 8020 82050 8090 82250
rect 8410 82050 8480 82250
rect 8520 82050 8590 82250
rect 8910 82050 8980 82250
rect 9020 82050 9090 82250
rect 9410 82050 9480 82250
rect 9520 82050 9590 82250
rect 9910 82050 9980 82250
rect 10020 82050 10090 82250
rect 10410 82050 10480 82250
rect 10520 82050 10590 82250
rect 10910 82050 10980 82250
rect 11020 82050 11090 82250
rect 11410 82050 11480 82250
rect 11520 82050 11590 82250
rect 11910 82050 11980 82250
rect 12020 82050 12090 82250
rect 12410 82050 12480 82250
rect 12520 82050 12590 82250
rect 12910 82050 12980 82250
rect 13020 82050 13090 82250
rect 13410 82050 13480 82250
rect 13520 82050 13590 82250
rect 13910 82050 13980 82250
rect 14020 82050 14090 82250
rect 14410 82050 14480 82250
rect 14520 82050 14590 82250
rect 14910 82050 14980 82250
rect 15020 82050 15090 82250
rect 15410 82050 15480 82250
rect 15520 82050 15590 82250
rect 15910 82050 15980 82250
rect 16020 82050 16090 82250
rect 16410 82050 16480 82250
rect 16520 82050 16590 82250
rect 16910 82050 16980 82250
rect 17020 82050 17090 82250
rect 17410 82050 17480 82250
rect 17520 82050 17590 82250
rect 17910 82050 17980 82250
rect 18020 82050 18090 82250
rect 18410 82050 18480 82250
rect 18520 82050 18590 82250
rect 18910 82050 18980 82250
rect 19020 82050 19090 82250
rect 19410 82050 19480 82250
rect 19520 82050 19590 82250
rect 19910 82050 19980 82250
rect 20020 82050 20090 82250
rect 20410 82050 20480 82250
rect 20520 82050 20590 82250
rect 20910 82050 20980 82250
rect 21020 82050 21090 82250
rect 21410 82050 21480 82250
rect 21520 82050 21590 82250
rect 21910 82050 21980 82250
rect 22020 82050 22090 82250
rect 22410 82050 22480 82250
rect 22520 82050 22590 82250
rect 22910 82050 22980 82250
rect 23020 82050 23090 82250
rect 23410 82050 23480 82250
rect 23520 82050 23590 82250
rect 23910 82050 23980 82250
rect 24020 82050 24090 82250
rect 24410 82050 24480 82250
rect 24520 82050 24590 82250
rect 24910 82050 24980 82250
rect 25020 82050 25090 82250
rect 25410 82050 25480 82250
rect 25520 82050 25590 82250
rect 25910 82050 25980 82250
rect 26020 82050 26090 82250
rect 26410 82050 26480 82250
rect 26520 82050 26590 82250
rect 26910 82050 26980 82250
rect 27020 82050 27090 82250
rect 27410 82050 27480 82250
rect 27520 82050 27590 82250
rect 27910 82050 27980 82250
rect 28020 82050 28090 82250
rect 28410 82050 28480 82250
rect 28520 82050 28590 82250
rect 28910 82050 28980 82250
rect 29020 82050 29090 82250
rect 29410 82050 29480 82250
rect 29520 82050 29590 82250
rect 29910 82050 29980 82250
rect 30020 82050 30090 82250
rect 30410 82050 30480 82250
rect 30520 82050 30590 82250
rect 30910 82050 30980 82250
rect 31020 82050 31090 82250
rect 31410 82050 31480 82250
rect 31520 82050 31590 82250
rect 31910 82050 31980 82250
rect 32020 82050 32090 82250
rect 32410 82050 32480 82250
rect 32520 82050 32590 82250
rect 32910 82050 32980 82250
rect 33020 82050 33090 82250
rect 33410 82050 33480 82250
rect 33520 82050 33590 82250
rect 33910 82050 33980 82250
rect 34020 82050 34090 82250
rect 34410 82050 34480 82250
rect 34520 82050 34590 82250
rect 34910 82050 34980 82250
rect 35020 82050 35090 82250
rect 35410 82050 35480 82250
rect 35520 82050 35590 82250
rect 35910 82050 35980 82250
rect 36020 82050 36090 82250
rect 36410 82050 36480 82250
rect 36520 82050 36590 82250
rect 36910 82050 36980 82250
rect 37020 82050 37090 82250
rect 37410 82050 37480 82250
rect 37520 82050 37590 82250
rect 37910 82050 37980 82250
rect 38020 82050 38090 82250
rect 38410 82050 38480 82250
rect 38520 82050 38590 82250
rect 38910 82050 38980 82250
rect 39020 82050 39090 82250
rect 39410 82050 39480 82250
rect 39520 82050 39590 82250
rect 39910 82050 39980 82250
rect 40020 82050 40090 82250
rect 40410 82050 40480 82250
rect 40520 82050 40590 82250
rect 40910 82050 40980 82250
rect 41020 82050 41090 82250
rect 41410 82050 41480 82250
rect 41520 82050 41590 82250
rect 41910 82050 41980 82250
rect 42020 82050 42090 82250
rect 42410 82050 42480 82250
rect 42520 82050 42590 82250
rect 42910 82050 42980 82250
rect 43020 82050 43090 82250
rect 43410 82050 43480 82250
rect 43520 82050 43590 82250
rect 43910 82050 43980 82250
rect 44020 82050 44090 82250
rect 44410 82050 44480 82250
rect 44520 82050 44590 82250
rect 44910 82050 44980 82250
rect 45020 82050 45090 82250
rect 45410 82050 45480 82250
rect 45520 82050 45590 82250
rect 45910 82050 45980 82250
rect 46020 82050 46090 82250
rect 46410 82050 46480 82250
rect 46520 82050 46590 82250
rect 46910 82050 46980 82250
rect 47020 82050 47090 82250
rect 47410 82050 47480 82250
rect 47520 82050 47590 82250
rect 47910 82050 47980 82250
rect 48020 82050 48090 82250
rect 48410 82050 48480 82250
rect 48520 82050 48590 82250
rect 48910 82050 48980 82250
rect 49020 82050 49090 82250
rect 49410 82050 49480 82250
rect 49520 82050 49590 82250
rect 49910 82050 49980 82250
rect 50020 82050 50090 82250
rect 50410 82050 50480 82250
rect 50520 82050 50590 82250
rect 50910 82050 50980 82250
rect 51020 82050 51090 82250
rect 51410 82050 51480 82250
rect 51520 82050 51590 82250
rect 51910 82050 51980 82250
rect 52020 82050 52090 82250
rect 52410 82050 52480 82250
rect 52520 82050 52590 82250
rect 52910 82050 52980 82250
rect 53020 82050 53090 82250
rect 53410 82050 53480 82250
rect 53520 82050 53590 82250
rect 53910 82050 53980 82250
rect 54020 82050 54090 82250
rect 54410 82050 54480 82250
rect 54520 82050 54590 82250
rect 54910 82050 54980 82250
rect 55020 82050 55090 82250
rect 55410 82050 55480 82250
rect 55520 82050 55590 82250
rect 55910 82050 55980 82250
rect 56020 82050 56090 82250
rect 56410 82050 56480 82250
rect 56520 82050 56590 82250
rect 56910 82050 56980 82250
rect 57020 82050 57090 82250
rect 57410 82050 57480 82250
rect 57520 82050 57590 82250
rect 57910 82050 57980 82250
rect 58020 82050 58090 82250
rect 58410 82050 58480 82250
rect 58520 82050 58590 82250
rect 58910 82050 58980 82250
rect 59020 82050 59090 82250
rect 59410 82050 59480 82250
rect 59520 82050 59590 82250
rect 59910 82050 59980 82250
rect 60020 82050 60090 82250
rect 60410 82050 60480 82250
rect 60520 82050 60590 82250
rect 60910 82050 60980 82250
rect 61020 82050 61090 82250
rect 61410 82050 61480 82250
rect 61520 82050 61590 82250
rect 61910 82050 61980 82250
rect 62020 82050 62090 82250
rect 62410 82050 62480 82250
rect 62520 82050 62590 82250
rect 62910 82050 62980 82250
rect 63020 82050 63090 82250
rect 63410 82050 63480 82250
rect 63520 82050 63590 82250
rect 63910 82050 63980 82250
rect 64020 82050 64090 82250
rect 64410 82050 64480 82250
rect 64520 82050 64590 82250
rect 64910 82050 64980 82250
rect 65020 82050 65090 82250
rect 65410 82050 65480 82250
rect 65520 82050 65590 82250
rect 65910 82050 65980 82250
rect 66020 82050 66090 82250
rect 66410 82050 66480 82250
rect 66520 82050 66590 82250
rect 66910 82050 66980 82250
rect 67020 82050 67090 82250
rect 67410 82050 67480 82250
rect 67520 82050 67590 82250
rect 67910 82050 67980 82250
rect 68020 82050 68090 82250
rect 68410 82050 68480 82250
rect 68520 82050 68590 82250
rect 68910 82050 68980 82250
rect 69020 82050 69090 82250
rect 69410 82050 69480 82250
rect 69520 82050 69590 82250
rect 69910 82050 69980 82250
rect 70020 82050 70090 82250
rect 70410 82050 70480 82250
rect 70520 82050 70590 82250
rect 70910 82050 70980 82250
rect 71020 82050 71090 82250
rect 71410 82050 71480 82250
rect 71520 82050 71590 82250
rect 71910 82050 71980 82250
rect 72020 82050 72090 82250
rect 72410 82050 72480 82250
rect 72520 82050 72590 82250
rect 72910 82050 72980 82250
rect 73020 82050 73090 82250
rect 73410 82050 73480 82250
rect 73520 82050 73590 82250
rect 73910 82050 73980 82250
rect 74020 82050 74090 82250
rect 74410 82050 74480 82250
rect 74520 82050 74590 82250
rect 74910 82050 74980 82250
rect 75020 82050 75090 82250
rect 75410 82050 75480 82250
rect 75520 82050 75590 82250
rect 75910 82050 75980 82250
rect 76020 82050 76090 82250
rect 76410 82050 76480 82250
rect 76520 82050 76590 82250
rect 76910 82050 76980 82250
rect 77020 82050 77090 82250
rect 77410 82050 77480 82250
rect 77520 82050 77590 82250
rect 77910 82050 77980 82250
rect 78020 82050 78090 82250
rect 78410 82050 78480 82250
rect 78520 82050 78590 82250
rect 78910 82050 78980 82250
rect 79020 82050 79090 82250
rect 79410 82050 79480 82250
rect 79520 82050 79590 82250
rect 79910 82050 79980 82250
rect 80020 82050 80090 82250
rect 80410 82050 80480 82250
rect 80520 82050 80590 82250
rect 80910 82050 80980 82250
rect 81020 82050 81090 82250
rect 81410 82050 81480 82250
rect 81520 82050 81590 82250
rect 81910 82050 81980 82250
rect 82020 82050 82090 82250
rect 82410 82050 82480 82250
rect 82520 82050 82590 82250
rect 82910 82050 82980 82250
rect 83020 82050 83090 82250
rect 83410 82050 83480 82250
rect 83520 82050 83590 82250
rect 83910 82050 83980 82250
rect 84020 82050 84090 82250
rect 84410 82050 84480 82250
rect 84520 82050 84590 82250
rect 84910 82050 84980 82250
rect 85020 82050 85090 82250
rect 85410 82050 85480 82250
rect 85520 82050 85590 82250
rect 85910 82050 85980 82250
rect 86020 82050 86090 82250
rect 86410 82050 86480 82250
rect 86520 82050 86590 82250
rect 86910 82050 86980 82250
rect 87020 82050 87090 82250
rect 87410 82050 87480 82250
rect 87520 82050 87590 82250
rect 87910 82050 87980 82250
rect 88020 82050 88090 82250
rect 88410 82050 88480 82250
rect 88520 82050 88590 82250
rect 88910 82050 88980 82250
rect 89020 82050 89090 82250
rect 89410 82050 89480 82250
rect 89520 82050 89590 82250
rect 89910 82050 89980 82250
rect 90020 82050 90090 82250
rect 90410 82050 90480 82250
rect 90520 82050 90590 82250
rect 90910 82050 90980 82250
rect 91020 82050 91090 82250
rect 91410 82050 91480 82250
rect 91520 82050 91590 82250
rect 91910 82050 91980 82250
rect 92020 82050 92090 82250
rect 92410 82050 92480 82250
rect 92520 82050 92590 82250
rect 92910 82050 92980 82250
rect 93020 82050 93090 82250
rect 93410 82050 93480 82250
rect 93520 82050 93590 82250
rect 93910 82050 93980 82250
rect 94020 82050 94090 82250
rect 94410 82050 94480 82250
rect 94520 82050 94590 82250
rect 94910 82050 94980 82250
rect 95020 82050 95090 82250
rect 95410 82050 95480 82250
rect 95520 82050 95590 82250
rect 95910 82050 95980 82250
rect 96020 82050 96090 82250
rect 96410 82050 96480 82250
rect 96520 82050 96590 82250
rect 96910 82050 96980 82250
rect 97020 82050 97090 82250
rect 97410 82050 97480 82250
rect 97520 82050 97590 82250
rect 97910 82050 97980 82250
rect 98020 82050 98090 82250
rect 98410 82050 98480 82250
rect 98520 82050 98590 82250
rect 98910 82050 98980 82250
rect 99020 82050 99090 82250
rect 99410 82050 99480 82250
rect 99520 82050 99590 82250
rect 99910 82050 99980 82250
rect 100020 82050 100090 82250
rect 100410 82050 100480 82250
rect -83350 81920 -83150 81990
rect -82850 81920 -82650 81990
rect -82350 81920 -82150 81990
rect -81850 81920 -81650 81990
rect -81350 81920 -81150 81990
rect -80850 81920 -80650 81990
rect -80350 81920 -80150 81990
rect -79850 81920 -79650 81990
rect -79350 81920 -79150 81990
rect -78850 81920 -78650 81990
rect -78350 81920 -78150 81990
rect -77850 81920 -77650 81990
rect -77350 81920 -77150 81990
rect -76850 81920 -76650 81990
rect -76350 81920 -76150 81990
rect -75850 81920 -75650 81990
rect -75350 81920 -75150 81990
rect -74850 81920 -74650 81990
rect -74350 81920 -74150 81990
rect -73850 81920 -73650 81990
rect -73350 81920 -73150 81990
rect -72850 81920 -72650 81990
rect -72350 81920 -72150 81990
rect -71850 81920 -71650 81990
rect -71350 81920 -71150 81990
rect -70850 81920 -70650 81990
rect -70350 81920 -70150 81990
rect -69850 81920 -69650 81990
rect -69350 81920 -69150 81990
rect -68850 81920 -68650 81990
rect -68350 81920 -68150 81990
rect -67850 81920 -67650 81990
rect -67350 81920 -67150 81990
rect -66850 81920 -66650 81990
rect -66350 81920 -66150 81990
rect -65850 81920 -65650 81990
rect -65350 81920 -65150 81990
rect -64850 81920 -64650 81990
rect -64350 81920 -64150 81990
rect -63850 81920 -63650 81990
rect -63350 81920 -63150 81990
rect -62850 81920 -62650 81990
rect -62350 81920 -62150 81990
rect -61850 81920 -61650 81990
rect -61350 81920 -61150 81990
rect -60850 81920 -60650 81990
rect -60350 81920 -60150 81990
rect -59850 81920 -59650 81990
rect -59350 81920 -59150 81990
rect -58850 81920 -58650 81990
rect -58350 81920 -58150 81990
rect -57850 81920 -57650 81990
rect -57350 81920 -57150 81990
rect -56850 81920 -56650 81990
rect -56350 81920 -56150 81990
rect -55850 81920 -55650 81990
rect -55350 81920 -55150 81990
rect -54850 81920 -54650 81990
rect -54350 81920 -54150 81990
rect -53850 81920 -53650 81990
rect -53350 81920 -53150 81990
rect -52850 81920 -52650 81990
rect -52350 81920 -52150 81990
rect -51850 81920 -51650 81990
rect -51350 81920 -51150 81990
rect -50850 81920 -50650 81990
rect -50350 81920 -50150 81990
rect -49850 81920 -49650 81990
rect -49350 81920 -49150 81990
rect -48850 81920 -48650 81990
rect -48350 81920 -48150 81990
rect -47850 81920 -47650 81990
rect -47350 81920 -47150 81990
rect -46850 81920 -46650 81990
rect -46350 81920 -46150 81990
rect -45850 81920 -45650 81990
rect -45350 81920 -45150 81990
rect -44850 81920 -44650 81990
rect -44350 81920 -44150 81990
rect -43850 81920 -43650 81990
rect -43350 81920 -43150 81990
rect -42850 81920 -42650 81990
rect -42350 81920 -42150 81990
rect -41850 81920 -41650 81990
rect -41350 81920 -41150 81990
rect -40850 81920 -40650 81990
rect -40350 81920 -40150 81990
rect -39850 81920 -39650 81990
rect -39350 81920 -39150 81990
rect -38850 81920 -38650 81990
rect -38350 81920 -38150 81990
rect -37850 81920 -37650 81990
rect -37350 81920 -37150 81990
rect -36850 81920 -36650 81990
rect -36350 81920 -36150 81990
rect -35850 81920 -35650 81990
rect -35350 81920 -35150 81990
rect -34850 81920 -34650 81990
rect -34350 81920 -34150 81990
rect -33850 81920 -33650 81990
rect -33350 81920 -33150 81990
rect -32850 81920 -32650 81990
rect -32350 81920 -32150 81990
rect -31850 81920 -31650 81990
rect -31350 81920 -31150 81990
rect -30850 81920 -30650 81990
rect -30350 81920 -30150 81990
rect -29850 81920 -29650 81990
rect -29350 81920 -29150 81990
rect -28850 81920 -28650 81990
rect -28350 81920 -28150 81990
rect -27850 81920 -27650 81990
rect -27350 81920 -27150 81990
rect -26850 81920 -26650 81990
rect -26350 81920 -26150 81990
rect -25850 81920 -25650 81990
rect -25350 81920 -25150 81990
rect -24850 81920 -24650 81990
rect -24350 81920 -24150 81990
rect -23850 81920 -23650 81990
rect -23350 81920 -23150 81990
rect -22850 81920 -22650 81990
rect -22350 81920 -22150 81990
rect -21850 81920 -21650 81990
rect -21350 81920 -21150 81990
rect -20850 81920 -20650 81990
rect -20350 81920 -20150 81990
rect -19850 81920 -19650 81990
rect -19350 81920 -19150 81990
rect -18850 81920 -18650 81990
rect -18350 81920 -18150 81990
rect -17850 81920 -17650 81990
rect -17350 81920 -17150 81990
rect -16850 81920 -16650 81990
rect -16350 81920 -16150 81990
rect -15850 81920 -15650 81990
rect -15350 81920 -15150 81990
rect -14850 81920 -14650 81990
rect -14350 81920 -14150 81990
rect -13850 81920 -13650 81990
rect -13350 81920 -13150 81990
rect -12850 81920 -12650 81990
rect -12350 81920 -12150 81990
rect -11850 81920 -11650 81990
rect -11350 81920 -11150 81990
rect -10850 81920 -10650 81990
rect -10350 81920 -10150 81990
rect -9850 81920 -9650 81990
rect -9350 81920 -9150 81990
rect -8850 81920 -8650 81990
rect -8350 81920 -8150 81990
rect -7850 81920 -7650 81990
rect -7350 81920 -7150 81990
rect -6850 81920 -6650 81990
rect -6350 81920 -6150 81990
rect -5850 81920 -5650 81990
rect -5350 81920 -5150 81990
rect -4850 81920 -4650 81990
rect -4350 81920 -4150 81990
rect -3850 81920 -3650 81990
rect -3350 81920 -3150 81990
rect -2850 81920 -2650 81990
rect -2350 81920 -2150 81990
rect -1850 81920 -1650 81990
rect -1350 81920 -1150 81990
rect -850 81920 -650 81990
rect -350 81920 -150 81990
rect 150 81920 350 81990
rect 650 81920 850 81990
rect 1150 81920 1350 81990
rect 1650 81920 1850 81990
rect 2150 81920 2350 81990
rect 2650 81920 2850 81990
rect 3150 81920 3350 81990
rect 3650 81920 3850 81990
rect 4150 81920 4350 81990
rect 4650 81920 4850 81990
rect 5150 81920 5350 81990
rect 5650 81920 5850 81990
rect 6150 81920 6350 81990
rect 6650 81920 6850 81990
rect 7150 81920 7350 81990
rect 7650 81920 7850 81990
rect 8150 81920 8350 81990
rect 8650 81920 8850 81990
rect 9150 81920 9350 81990
rect 9650 81920 9850 81990
rect 10150 81920 10350 81990
rect 10650 81920 10850 81990
rect 11150 81920 11350 81990
rect 11650 81920 11850 81990
rect 12150 81920 12350 81990
rect 12650 81920 12850 81990
rect 13150 81920 13350 81990
rect 13650 81920 13850 81990
rect 14150 81920 14350 81990
rect 14650 81920 14850 81990
rect 15150 81920 15350 81990
rect 15650 81920 15850 81990
rect 16150 81920 16350 81990
rect 16650 81920 16850 81990
rect 17150 81920 17350 81990
rect 17650 81920 17850 81990
rect 18150 81920 18350 81990
rect 18650 81920 18850 81990
rect 19150 81920 19350 81990
rect 19650 81920 19850 81990
rect 20150 81920 20350 81990
rect 20650 81920 20850 81990
rect 21150 81920 21350 81990
rect 21650 81920 21850 81990
rect 22150 81920 22350 81990
rect 22650 81920 22850 81990
rect 23150 81920 23350 81990
rect 23650 81920 23850 81990
rect 24150 81920 24350 81990
rect 24650 81920 24850 81990
rect 25150 81920 25350 81990
rect 25650 81920 25850 81990
rect 26150 81920 26350 81990
rect 26650 81920 26850 81990
rect 27150 81920 27350 81990
rect 27650 81920 27850 81990
rect 28150 81920 28350 81990
rect 28650 81920 28850 81990
rect 29150 81920 29350 81990
rect 29650 81920 29850 81990
rect 30150 81920 30350 81990
rect 30650 81920 30850 81990
rect 31150 81920 31350 81990
rect 31650 81920 31850 81990
rect 32150 81920 32350 81990
rect 32650 81920 32850 81990
rect 33150 81920 33350 81990
rect 33650 81920 33850 81990
rect 34150 81920 34350 81990
rect 34650 81920 34850 81990
rect 35150 81920 35350 81990
rect 35650 81920 35850 81990
rect 36150 81920 36350 81990
rect 36650 81920 36850 81990
rect 37150 81920 37350 81990
rect 37650 81920 37850 81990
rect 38150 81920 38350 81990
rect 38650 81920 38850 81990
rect 39150 81920 39350 81990
rect 39650 81920 39850 81990
rect 40150 81920 40350 81990
rect 40650 81920 40850 81990
rect 41150 81920 41350 81990
rect 41650 81920 41850 81990
rect 42150 81920 42350 81990
rect 42650 81920 42850 81990
rect 43150 81920 43350 81990
rect 43650 81920 43850 81990
rect 44150 81920 44350 81990
rect 44650 81920 44850 81990
rect 45150 81920 45350 81990
rect 45650 81920 45850 81990
rect 46150 81920 46350 81990
rect 46650 81920 46850 81990
rect 47150 81920 47350 81990
rect 47650 81920 47850 81990
rect 48150 81920 48350 81990
rect 48650 81920 48850 81990
rect 49150 81920 49350 81990
rect 49650 81920 49850 81990
rect 50150 81920 50350 81990
rect 50650 81920 50850 81990
rect 51150 81920 51350 81990
rect 51650 81920 51850 81990
rect 52150 81920 52350 81990
rect 52650 81920 52850 81990
rect 53150 81920 53350 81990
rect 53650 81920 53850 81990
rect 54150 81920 54350 81990
rect 54650 81920 54850 81990
rect 55150 81920 55350 81990
rect 55650 81920 55850 81990
rect 56150 81920 56350 81990
rect 56650 81920 56850 81990
rect 57150 81920 57350 81990
rect 57650 81920 57850 81990
rect 58150 81920 58350 81990
rect 58650 81920 58850 81990
rect 59150 81920 59350 81990
rect 59650 81920 59850 81990
rect 60150 81920 60350 81990
rect 60650 81920 60850 81990
rect 61150 81920 61350 81990
rect 61650 81920 61850 81990
rect 62150 81920 62350 81990
rect 62650 81920 62850 81990
rect 63150 81920 63350 81990
rect 63650 81920 63850 81990
rect 64150 81920 64350 81990
rect 64650 81920 64850 81990
rect 65150 81920 65350 81990
rect 65650 81920 65850 81990
rect 66150 81920 66350 81990
rect 66650 81920 66850 81990
rect 67150 81920 67350 81990
rect 67650 81920 67850 81990
rect 68150 81920 68350 81990
rect 68650 81920 68850 81990
rect 69150 81920 69350 81990
rect 69650 81920 69850 81990
rect 70150 81920 70350 81990
rect 70650 81920 70850 81990
rect 71150 81920 71350 81990
rect 71650 81920 71850 81990
rect 72150 81920 72350 81990
rect 72650 81920 72850 81990
rect 73150 81920 73350 81990
rect 73650 81920 73850 81990
rect 74150 81920 74350 81990
rect 74650 81920 74850 81990
rect 75150 81920 75350 81990
rect 75650 81920 75850 81990
rect 76150 81920 76350 81990
rect 76650 81920 76850 81990
rect 77150 81920 77350 81990
rect 77650 81920 77850 81990
rect 78150 81920 78350 81990
rect 78650 81920 78850 81990
rect 79150 81920 79350 81990
rect 79650 81920 79850 81990
rect 80150 81920 80350 81990
rect 80650 81920 80850 81990
rect 81150 81920 81350 81990
rect 81650 81920 81850 81990
rect 82150 81920 82350 81990
rect 82650 81920 82850 81990
rect 83150 81920 83350 81990
rect 83650 81920 83850 81990
rect 84150 81920 84350 81990
rect 84650 81920 84850 81990
rect 85150 81920 85350 81990
rect 85650 81920 85850 81990
rect 86150 81920 86350 81990
rect 86650 81920 86850 81990
rect 87150 81920 87350 81990
rect 87650 81920 87850 81990
rect 88150 81920 88350 81990
rect 88650 81920 88850 81990
rect 89150 81920 89350 81990
rect 89650 81920 89850 81990
rect 90150 81920 90350 81990
rect 90650 81920 90850 81990
rect 91150 81920 91350 81990
rect 91650 81920 91850 81990
rect 92150 81920 92350 81990
rect 92650 81920 92850 81990
rect 93150 81920 93350 81990
rect 93650 81920 93850 81990
rect 94150 81920 94350 81990
rect 94650 81920 94850 81990
rect 95150 81920 95350 81990
rect 95650 81920 95850 81990
rect 96150 81920 96350 81990
rect 96650 81920 96850 81990
rect 97150 81920 97350 81990
rect 97650 81920 97850 81990
rect 98150 81920 98350 81990
rect 98650 81920 98850 81990
rect 99150 81920 99350 81990
rect 99650 81920 99850 81990
rect 100150 81920 100350 81990
rect -83350 81810 -83150 81880
rect -82850 81810 -82650 81880
rect -82350 81810 -82150 81880
rect -81850 81810 -81650 81880
rect -81350 81810 -81150 81880
rect -80850 81810 -80650 81880
rect -80350 81810 -80150 81880
rect -79850 81810 -79650 81880
rect -79350 81810 -79150 81880
rect -78850 81810 -78650 81880
rect -78350 81810 -78150 81880
rect -77850 81810 -77650 81880
rect -77350 81810 -77150 81880
rect -76850 81810 -76650 81880
rect -76350 81810 -76150 81880
rect -75850 81810 -75650 81880
rect -75350 81810 -75150 81880
rect -74850 81810 -74650 81880
rect -74350 81810 -74150 81880
rect -73850 81810 -73650 81880
rect -73350 81810 -73150 81880
rect -72850 81810 -72650 81880
rect -72350 81810 -72150 81880
rect -71850 81810 -71650 81880
rect -71350 81810 -71150 81880
rect -70850 81810 -70650 81880
rect -70350 81810 -70150 81880
rect -69850 81810 -69650 81880
rect -69350 81810 -69150 81880
rect -68850 81810 -68650 81880
rect -68350 81810 -68150 81880
rect -67850 81810 -67650 81880
rect -67350 81810 -67150 81880
rect -66850 81810 -66650 81880
rect -66350 81810 -66150 81880
rect -65850 81810 -65650 81880
rect -65350 81810 -65150 81880
rect -64850 81810 -64650 81880
rect -64350 81810 -64150 81880
rect -63850 81810 -63650 81880
rect -63350 81810 -63150 81880
rect -62850 81810 -62650 81880
rect -62350 81810 -62150 81880
rect -61850 81810 -61650 81880
rect -61350 81810 -61150 81880
rect -60850 81810 -60650 81880
rect -60350 81810 -60150 81880
rect -59850 81810 -59650 81880
rect -59350 81810 -59150 81880
rect -58850 81810 -58650 81880
rect -58350 81810 -58150 81880
rect -57850 81810 -57650 81880
rect -57350 81810 -57150 81880
rect -56850 81810 -56650 81880
rect -56350 81810 -56150 81880
rect -55850 81810 -55650 81880
rect -55350 81810 -55150 81880
rect -54850 81810 -54650 81880
rect -54350 81810 -54150 81880
rect -53850 81810 -53650 81880
rect -53350 81810 -53150 81880
rect -52850 81810 -52650 81880
rect -52350 81810 -52150 81880
rect -51850 81810 -51650 81880
rect -51350 81810 -51150 81880
rect -50850 81810 -50650 81880
rect -50350 81810 -50150 81880
rect -49850 81810 -49650 81880
rect -49350 81810 -49150 81880
rect -48850 81810 -48650 81880
rect -48350 81810 -48150 81880
rect -47850 81810 -47650 81880
rect -47350 81810 -47150 81880
rect -46850 81810 -46650 81880
rect -46350 81810 -46150 81880
rect -45850 81810 -45650 81880
rect -45350 81810 -45150 81880
rect -44850 81810 -44650 81880
rect -44350 81810 -44150 81880
rect -43850 81810 -43650 81880
rect -43350 81810 -43150 81880
rect -42850 81810 -42650 81880
rect -42350 81810 -42150 81880
rect -41850 81810 -41650 81880
rect -41350 81810 -41150 81880
rect -40850 81810 -40650 81880
rect -40350 81810 -40150 81880
rect -39850 81810 -39650 81880
rect -39350 81810 -39150 81880
rect -38850 81810 -38650 81880
rect -38350 81810 -38150 81880
rect -37850 81810 -37650 81880
rect -37350 81810 -37150 81880
rect -36850 81810 -36650 81880
rect -36350 81810 -36150 81880
rect -35850 81810 -35650 81880
rect -35350 81810 -35150 81880
rect -34850 81810 -34650 81880
rect -34350 81810 -34150 81880
rect -33850 81810 -33650 81880
rect -33350 81810 -33150 81880
rect -32850 81810 -32650 81880
rect -32350 81810 -32150 81880
rect -31850 81810 -31650 81880
rect -31350 81810 -31150 81880
rect -30850 81810 -30650 81880
rect -30350 81810 -30150 81880
rect -29850 81810 -29650 81880
rect -29350 81810 -29150 81880
rect -28850 81810 -28650 81880
rect -28350 81810 -28150 81880
rect -27850 81810 -27650 81880
rect -27350 81810 -27150 81880
rect -26850 81810 -26650 81880
rect -26350 81810 -26150 81880
rect -25850 81810 -25650 81880
rect -25350 81810 -25150 81880
rect -24850 81810 -24650 81880
rect -24350 81810 -24150 81880
rect -23850 81810 -23650 81880
rect -23350 81810 -23150 81880
rect -22850 81810 -22650 81880
rect -22350 81810 -22150 81880
rect -21850 81810 -21650 81880
rect -21350 81810 -21150 81880
rect -20850 81810 -20650 81880
rect -20350 81810 -20150 81880
rect -19850 81810 -19650 81880
rect -19350 81810 -19150 81880
rect -18850 81810 -18650 81880
rect -18350 81810 -18150 81880
rect -17850 81810 -17650 81880
rect -17350 81810 -17150 81880
rect -16850 81810 -16650 81880
rect -16350 81810 -16150 81880
rect -15850 81810 -15650 81880
rect -15350 81810 -15150 81880
rect -14850 81810 -14650 81880
rect -14350 81810 -14150 81880
rect -13850 81810 -13650 81880
rect -13350 81810 -13150 81880
rect -12850 81810 -12650 81880
rect -12350 81810 -12150 81880
rect -11850 81810 -11650 81880
rect -11350 81810 -11150 81880
rect -10850 81810 -10650 81880
rect -10350 81810 -10150 81880
rect -9850 81810 -9650 81880
rect -9350 81810 -9150 81880
rect -8850 81810 -8650 81880
rect -8350 81810 -8150 81880
rect -7850 81810 -7650 81880
rect -7350 81810 -7150 81880
rect -6850 81810 -6650 81880
rect -6350 81810 -6150 81880
rect -5850 81810 -5650 81880
rect -5350 81810 -5150 81880
rect -4850 81810 -4650 81880
rect -4350 81810 -4150 81880
rect -3850 81810 -3650 81880
rect -3350 81810 -3150 81880
rect -2850 81810 -2650 81880
rect -2350 81810 -2150 81880
rect -1850 81810 -1650 81880
rect -1350 81810 -1150 81880
rect -850 81810 -650 81880
rect -350 81810 -150 81880
rect 150 81810 350 81880
rect 650 81810 850 81880
rect 1150 81810 1350 81880
rect 1650 81810 1850 81880
rect 2150 81810 2350 81880
rect 2650 81810 2850 81880
rect 3150 81810 3350 81880
rect 3650 81810 3850 81880
rect 4150 81810 4350 81880
rect 4650 81810 4850 81880
rect 5150 81810 5350 81880
rect 5650 81810 5850 81880
rect 6150 81810 6350 81880
rect 6650 81810 6850 81880
rect 7150 81810 7350 81880
rect 7650 81810 7850 81880
rect 8150 81810 8350 81880
rect 8650 81810 8850 81880
rect 9150 81810 9350 81880
rect 9650 81810 9850 81880
rect 10150 81810 10350 81880
rect 10650 81810 10850 81880
rect 11150 81810 11350 81880
rect 11650 81810 11850 81880
rect 12150 81810 12350 81880
rect 12650 81810 12850 81880
rect 13150 81810 13350 81880
rect 13650 81810 13850 81880
rect 14150 81810 14350 81880
rect 14650 81810 14850 81880
rect 15150 81810 15350 81880
rect 15650 81810 15850 81880
rect 16150 81810 16350 81880
rect 16650 81810 16850 81880
rect 17150 81810 17350 81880
rect 17650 81810 17850 81880
rect 18150 81810 18350 81880
rect 18650 81810 18850 81880
rect 19150 81810 19350 81880
rect 19650 81810 19850 81880
rect 20150 81810 20350 81880
rect 20650 81810 20850 81880
rect 21150 81810 21350 81880
rect 21650 81810 21850 81880
rect 22150 81810 22350 81880
rect 22650 81810 22850 81880
rect 23150 81810 23350 81880
rect 23650 81810 23850 81880
rect 24150 81810 24350 81880
rect 24650 81810 24850 81880
rect 25150 81810 25350 81880
rect 25650 81810 25850 81880
rect 26150 81810 26350 81880
rect 26650 81810 26850 81880
rect 27150 81810 27350 81880
rect 27650 81810 27850 81880
rect 28150 81810 28350 81880
rect 28650 81810 28850 81880
rect 29150 81810 29350 81880
rect 29650 81810 29850 81880
rect 30150 81810 30350 81880
rect 30650 81810 30850 81880
rect 31150 81810 31350 81880
rect 31650 81810 31850 81880
rect 32150 81810 32350 81880
rect 32650 81810 32850 81880
rect 33150 81810 33350 81880
rect 33650 81810 33850 81880
rect 34150 81810 34350 81880
rect 34650 81810 34850 81880
rect 35150 81810 35350 81880
rect 35650 81810 35850 81880
rect 36150 81810 36350 81880
rect 36650 81810 36850 81880
rect 37150 81810 37350 81880
rect 37650 81810 37850 81880
rect 38150 81810 38350 81880
rect 38650 81810 38850 81880
rect 39150 81810 39350 81880
rect 39650 81810 39850 81880
rect 40150 81810 40350 81880
rect 40650 81810 40850 81880
rect 41150 81810 41350 81880
rect 41650 81810 41850 81880
rect 42150 81810 42350 81880
rect 42650 81810 42850 81880
rect 43150 81810 43350 81880
rect 43650 81810 43850 81880
rect 44150 81810 44350 81880
rect 44650 81810 44850 81880
rect 45150 81810 45350 81880
rect 45650 81810 45850 81880
rect 46150 81810 46350 81880
rect 46650 81810 46850 81880
rect 47150 81810 47350 81880
rect 47650 81810 47850 81880
rect 48150 81810 48350 81880
rect 48650 81810 48850 81880
rect 49150 81810 49350 81880
rect 49650 81810 49850 81880
rect 50150 81810 50350 81880
rect 50650 81810 50850 81880
rect 51150 81810 51350 81880
rect 51650 81810 51850 81880
rect 52150 81810 52350 81880
rect 52650 81810 52850 81880
rect 53150 81810 53350 81880
rect 53650 81810 53850 81880
rect 54150 81810 54350 81880
rect 54650 81810 54850 81880
rect 55150 81810 55350 81880
rect 55650 81810 55850 81880
rect 56150 81810 56350 81880
rect 56650 81810 56850 81880
rect 57150 81810 57350 81880
rect 57650 81810 57850 81880
rect 58150 81810 58350 81880
rect 58650 81810 58850 81880
rect 59150 81810 59350 81880
rect 59650 81810 59850 81880
rect 60150 81810 60350 81880
rect 60650 81810 60850 81880
rect 61150 81810 61350 81880
rect 61650 81810 61850 81880
rect 62150 81810 62350 81880
rect 62650 81810 62850 81880
rect 63150 81810 63350 81880
rect 63650 81810 63850 81880
rect 64150 81810 64350 81880
rect 64650 81810 64850 81880
rect 65150 81810 65350 81880
rect 65650 81810 65850 81880
rect 66150 81810 66350 81880
rect 66650 81810 66850 81880
rect 67150 81810 67350 81880
rect 67650 81810 67850 81880
rect 68150 81810 68350 81880
rect 68650 81810 68850 81880
rect 69150 81810 69350 81880
rect 69650 81810 69850 81880
rect 70150 81810 70350 81880
rect 70650 81810 70850 81880
rect 71150 81810 71350 81880
rect 71650 81810 71850 81880
rect 72150 81810 72350 81880
rect 72650 81810 72850 81880
rect 73150 81810 73350 81880
rect 73650 81810 73850 81880
rect 74150 81810 74350 81880
rect 74650 81810 74850 81880
rect 75150 81810 75350 81880
rect 75650 81810 75850 81880
rect 76150 81810 76350 81880
rect 76650 81810 76850 81880
rect 77150 81810 77350 81880
rect 77650 81810 77850 81880
rect 78150 81810 78350 81880
rect 78650 81810 78850 81880
rect 79150 81810 79350 81880
rect 79650 81810 79850 81880
rect 80150 81810 80350 81880
rect 80650 81810 80850 81880
rect 81150 81810 81350 81880
rect 81650 81810 81850 81880
rect 82150 81810 82350 81880
rect 82650 81810 82850 81880
rect 83150 81810 83350 81880
rect 83650 81810 83850 81880
rect 84150 81810 84350 81880
rect 84650 81810 84850 81880
rect 85150 81810 85350 81880
rect 85650 81810 85850 81880
rect 86150 81810 86350 81880
rect 86650 81810 86850 81880
rect 87150 81810 87350 81880
rect 87650 81810 87850 81880
rect 88150 81810 88350 81880
rect 88650 81810 88850 81880
rect 89150 81810 89350 81880
rect 89650 81810 89850 81880
rect 90150 81810 90350 81880
rect 90650 81810 90850 81880
rect 91150 81810 91350 81880
rect 91650 81810 91850 81880
rect 92150 81810 92350 81880
rect 92650 81810 92850 81880
rect 93150 81810 93350 81880
rect 93650 81810 93850 81880
rect 94150 81810 94350 81880
rect 94650 81810 94850 81880
rect 95150 81810 95350 81880
rect 95650 81810 95850 81880
rect 96150 81810 96350 81880
rect 96650 81810 96850 81880
rect 97150 81810 97350 81880
rect 97650 81810 97850 81880
rect 98150 81810 98350 81880
rect 98650 81810 98850 81880
rect 99150 81810 99350 81880
rect 99650 81810 99850 81880
rect 100150 81810 100350 81880
rect -83480 81550 -83410 81750
rect -83090 81550 -83020 81750
rect -82980 81550 -82910 81750
rect -82590 81550 -82520 81750
rect -82480 81550 -82410 81750
rect -82090 81550 -82020 81750
rect -81980 81550 -81910 81750
rect -81590 81550 -81520 81750
rect -81480 81550 -81410 81750
rect -81090 81550 -81020 81750
rect -80980 81550 -80910 81750
rect -80590 81550 -80520 81750
rect -80480 81550 -80410 81750
rect -80090 81550 -80020 81750
rect -79980 81550 -79910 81750
rect -79590 81550 -79520 81750
rect -79480 81550 -79410 81750
rect -79090 81550 -79020 81750
rect -78980 81550 -78910 81750
rect -78590 81550 -78520 81750
rect -78480 81550 -78410 81750
rect -78090 81550 -78020 81750
rect -77980 81550 -77910 81750
rect -77590 81550 -77520 81750
rect -77480 81550 -77410 81750
rect -77090 81550 -77020 81750
rect -76980 81550 -76910 81750
rect -76590 81550 -76520 81750
rect -76480 81550 -76410 81750
rect -76090 81550 -76020 81750
rect -75980 81550 -75910 81750
rect -75590 81550 -75520 81750
rect -75480 81550 -75410 81750
rect -75090 81550 -75020 81750
rect -74980 81550 -74910 81750
rect -74590 81550 -74520 81750
rect -74480 81550 -74410 81750
rect -74090 81550 -74020 81750
rect -73980 81550 -73910 81750
rect -73590 81550 -73520 81750
rect -73480 81550 -73410 81750
rect -73090 81550 -73020 81750
rect -72980 81550 -72910 81750
rect -72590 81550 -72520 81750
rect -72480 81550 -72410 81750
rect -72090 81550 -72020 81750
rect -71980 81550 -71910 81750
rect -71590 81550 -71520 81750
rect -71480 81550 -71410 81750
rect -71090 81550 -71020 81750
rect -70980 81550 -70910 81750
rect -70590 81550 -70520 81750
rect -70480 81550 -70410 81750
rect -70090 81550 -70020 81750
rect -69980 81550 -69910 81750
rect -69590 81550 -69520 81750
rect -69480 81550 -69410 81750
rect -69090 81550 -69020 81750
rect -68980 81550 -68910 81750
rect -68590 81550 -68520 81750
rect -68480 81550 -68410 81750
rect -68090 81550 -68020 81750
rect -67980 81550 -67910 81750
rect -67590 81550 -67520 81750
rect -67480 81550 -67410 81750
rect -67090 81550 -67020 81750
rect -66980 81550 -66910 81750
rect -66590 81550 -66520 81750
rect -66480 81550 -66410 81750
rect -66090 81550 -66020 81750
rect -65980 81550 -65910 81750
rect -65590 81550 -65520 81750
rect -65480 81550 -65410 81750
rect -65090 81550 -65020 81750
rect -64980 81550 -64910 81750
rect -64590 81550 -64520 81750
rect -64480 81550 -64410 81750
rect -64090 81550 -64020 81750
rect -63980 81550 -63910 81750
rect -63590 81550 -63520 81750
rect -63480 81550 -63410 81750
rect -63090 81550 -63020 81750
rect -62980 81550 -62910 81750
rect -62590 81550 -62520 81750
rect -62480 81550 -62410 81750
rect -62090 81550 -62020 81750
rect -61980 81550 -61910 81750
rect -61590 81550 -61520 81750
rect -61480 81550 -61410 81750
rect -61090 81550 -61020 81750
rect -60980 81550 -60910 81750
rect -60590 81550 -60520 81750
rect -60480 81550 -60410 81750
rect -60090 81550 -60020 81750
rect -59980 81550 -59910 81750
rect -59590 81550 -59520 81750
rect -59480 81550 -59410 81750
rect -59090 81550 -59020 81750
rect -58980 81550 -58910 81750
rect -58590 81550 -58520 81750
rect -58480 81550 -58410 81750
rect -58090 81550 -58020 81750
rect -57980 81550 -57910 81750
rect -57590 81550 -57520 81750
rect -57480 81550 -57410 81750
rect -57090 81550 -57020 81750
rect -56980 81550 -56910 81750
rect -56590 81550 -56520 81750
rect -56480 81550 -56410 81750
rect -56090 81550 -56020 81750
rect -55980 81550 -55910 81750
rect -55590 81550 -55520 81750
rect -55480 81550 -55410 81750
rect -55090 81550 -55020 81750
rect -54980 81550 -54910 81750
rect -54590 81550 -54520 81750
rect -54480 81550 -54410 81750
rect -54090 81550 -54020 81750
rect -53980 81550 -53910 81750
rect -53590 81550 -53520 81750
rect -53480 81550 -53410 81750
rect -53090 81550 -53020 81750
rect -52980 81550 -52910 81750
rect -52590 81550 -52520 81750
rect -52480 81550 -52410 81750
rect -52090 81550 -52020 81750
rect -51980 81550 -51910 81750
rect -51590 81550 -51520 81750
rect -51480 81550 -51410 81750
rect -51090 81550 -51020 81750
rect -50980 81550 -50910 81750
rect -50590 81550 -50520 81750
rect -50480 81550 -50410 81750
rect -50090 81550 -50020 81750
rect -49980 81550 -49910 81750
rect -49590 81550 -49520 81750
rect -49480 81550 -49410 81750
rect -49090 81550 -49020 81750
rect -48980 81550 -48910 81750
rect -48590 81550 -48520 81750
rect -48480 81550 -48410 81750
rect -48090 81550 -48020 81750
rect -47980 81550 -47910 81750
rect -47590 81550 -47520 81750
rect -47480 81550 -47410 81750
rect -47090 81550 -47020 81750
rect -46980 81550 -46910 81750
rect -46590 81550 -46520 81750
rect -46480 81550 -46410 81750
rect -46090 81550 -46020 81750
rect -45980 81550 -45910 81750
rect -45590 81550 -45520 81750
rect -45480 81550 -45410 81750
rect -45090 81550 -45020 81750
rect -44980 81550 -44910 81750
rect -44590 81550 -44520 81750
rect -44480 81550 -44410 81750
rect -44090 81550 -44020 81750
rect -43980 81550 -43910 81750
rect -43590 81550 -43520 81750
rect -43480 81550 -43410 81750
rect -43090 81550 -43020 81750
rect -42980 81550 -42910 81750
rect -42590 81550 -42520 81750
rect -42480 81550 -42410 81750
rect -42090 81550 -42020 81750
rect -41980 81550 -41910 81750
rect -41590 81550 -41520 81750
rect -41480 81550 -41410 81750
rect -41090 81550 -41020 81750
rect -40980 81550 -40910 81750
rect -40590 81550 -40520 81750
rect -40480 81550 -40410 81750
rect -40090 81550 -40020 81750
rect -39980 81550 -39910 81750
rect -39590 81550 -39520 81750
rect -39480 81550 -39410 81750
rect -39090 81550 -39020 81750
rect -38980 81550 -38910 81750
rect -38590 81550 -38520 81750
rect -38480 81550 -38410 81750
rect -38090 81550 -38020 81750
rect -37980 81550 -37910 81750
rect -37590 81550 -37520 81750
rect -37480 81550 -37410 81750
rect -37090 81550 -37020 81750
rect -36980 81550 -36910 81750
rect -36590 81550 -36520 81750
rect -36480 81550 -36410 81750
rect -36090 81550 -36020 81750
rect -35980 81550 -35910 81750
rect -35590 81550 -35520 81750
rect -35480 81550 -35410 81750
rect -35090 81550 -35020 81750
rect -34980 81550 -34910 81750
rect -34590 81550 -34520 81750
rect -34480 81550 -34410 81750
rect -34090 81550 -34020 81750
rect -33980 81550 -33910 81750
rect -33590 81550 -33520 81750
rect -33480 81550 -33410 81750
rect -33090 81550 -33020 81750
rect -32980 81550 -32910 81750
rect -32590 81550 -32520 81750
rect -32480 81550 -32410 81750
rect -32090 81550 -32020 81750
rect -31980 81550 -31910 81750
rect -31590 81550 -31520 81750
rect -31480 81550 -31410 81750
rect -31090 81550 -31020 81750
rect -30980 81550 -30910 81750
rect -30590 81550 -30520 81750
rect -30480 81550 -30410 81750
rect -30090 81550 -30020 81750
rect -29980 81550 -29910 81750
rect -29590 81550 -29520 81750
rect -29480 81550 -29410 81750
rect -29090 81550 -29020 81750
rect -28980 81550 -28910 81750
rect -28590 81550 -28520 81750
rect -28480 81550 -28410 81750
rect -28090 81550 -28020 81750
rect -27980 81550 -27910 81750
rect -27590 81550 -27520 81750
rect -27480 81550 -27410 81750
rect -27090 81550 -27020 81750
rect -26980 81550 -26910 81750
rect -26590 81550 -26520 81750
rect -26480 81550 -26410 81750
rect -26090 81550 -26020 81750
rect -25980 81550 -25910 81750
rect -25590 81550 -25520 81750
rect -25480 81550 -25410 81750
rect -25090 81550 -25020 81750
rect -24980 81550 -24910 81750
rect -24590 81550 -24520 81750
rect -24480 81550 -24410 81750
rect -24090 81550 -24020 81750
rect -23980 81550 -23910 81750
rect -23590 81550 -23520 81750
rect -23480 81550 -23410 81750
rect -23090 81550 -23020 81750
rect -22980 81550 -22910 81750
rect -22590 81550 -22520 81750
rect -22480 81550 -22410 81750
rect -22090 81550 -22020 81750
rect -21980 81550 -21910 81750
rect -21590 81550 -21520 81750
rect -21480 81550 -21410 81750
rect -21090 81550 -21020 81750
rect -20980 81550 -20910 81750
rect -20590 81550 -20520 81750
rect -20480 81550 -20410 81750
rect -20090 81550 -20020 81750
rect -19980 81550 -19910 81750
rect -19590 81550 -19520 81750
rect -19480 81550 -19410 81750
rect -19090 81550 -19020 81750
rect -18980 81550 -18910 81750
rect -18590 81550 -18520 81750
rect -18480 81550 -18410 81750
rect -18090 81550 -18020 81750
rect -17980 81550 -17910 81750
rect -17590 81550 -17520 81750
rect -17480 81550 -17410 81750
rect -17090 81550 -17020 81750
rect -16980 81550 -16910 81750
rect -16590 81550 -16520 81750
rect -16480 81550 -16410 81750
rect -16090 81550 -16020 81750
rect -15980 81550 -15910 81750
rect -15590 81550 -15520 81750
rect -15480 81550 -15410 81750
rect -15090 81550 -15020 81750
rect -14980 81550 -14910 81750
rect -14590 81550 -14520 81750
rect -14480 81550 -14410 81750
rect -14090 81550 -14020 81750
rect -13980 81550 -13910 81750
rect -13590 81550 -13520 81750
rect -13480 81550 -13410 81750
rect -13090 81550 -13020 81750
rect -12980 81550 -12910 81750
rect -12590 81550 -12520 81750
rect -12480 81550 -12410 81750
rect -12090 81550 -12020 81750
rect -11980 81550 -11910 81750
rect -11590 81550 -11520 81750
rect -11480 81550 -11410 81750
rect -11090 81550 -11020 81750
rect -10980 81550 -10910 81750
rect -10590 81550 -10520 81750
rect -10480 81550 -10410 81750
rect -10090 81550 -10020 81750
rect -9980 81550 -9910 81750
rect -9590 81550 -9520 81750
rect -9480 81550 -9410 81750
rect -9090 81550 -9020 81750
rect -8980 81550 -8910 81750
rect -8590 81550 -8520 81750
rect -8480 81550 -8410 81750
rect -8090 81550 -8020 81750
rect -7980 81550 -7910 81750
rect -7590 81550 -7520 81750
rect -7480 81550 -7410 81750
rect -7090 81550 -7020 81750
rect -6980 81550 -6910 81750
rect -6590 81550 -6520 81750
rect -6480 81550 -6410 81750
rect -6090 81550 -6020 81750
rect -5980 81550 -5910 81750
rect -5590 81550 -5520 81750
rect -5480 81550 -5410 81750
rect -5090 81550 -5020 81750
rect -4980 81550 -4910 81750
rect -4590 81550 -4520 81750
rect -4480 81550 -4410 81750
rect -4090 81550 -4020 81750
rect -3980 81550 -3910 81750
rect -3590 81550 -3520 81750
rect -3480 81550 -3410 81750
rect -3090 81550 -3020 81750
rect -2980 81550 -2910 81750
rect -2590 81550 -2520 81750
rect -2480 81550 -2410 81750
rect -2090 81550 -2020 81750
rect -1980 81550 -1910 81750
rect -1590 81550 -1520 81750
rect -1480 81550 -1410 81750
rect -1090 81550 -1020 81750
rect -980 81550 -910 81750
rect -590 81550 -520 81750
rect -480 81550 -410 81750
rect -90 81550 -20 81750
rect 20 81550 90 81750
rect 410 81550 480 81750
rect 520 81550 590 81750
rect 910 81550 980 81750
rect 1020 81550 1090 81750
rect 1410 81550 1480 81750
rect 1520 81550 1590 81750
rect 1910 81550 1980 81750
rect 2020 81550 2090 81750
rect 2410 81550 2480 81750
rect 2520 81550 2590 81750
rect 2910 81550 2980 81750
rect 3020 81550 3090 81750
rect 3410 81550 3480 81750
rect 3520 81550 3590 81750
rect 3910 81550 3980 81750
rect 4020 81550 4090 81750
rect 4410 81550 4480 81750
rect 4520 81550 4590 81750
rect 4910 81550 4980 81750
rect 5020 81550 5090 81750
rect 5410 81550 5480 81750
rect 5520 81550 5590 81750
rect 5910 81550 5980 81750
rect 6020 81550 6090 81750
rect 6410 81550 6480 81750
rect 6520 81550 6590 81750
rect 6910 81550 6980 81750
rect 7020 81550 7090 81750
rect 7410 81550 7480 81750
rect 7520 81550 7590 81750
rect 7910 81550 7980 81750
rect 8020 81550 8090 81750
rect 8410 81550 8480 81750
rect 8520 81550 8590 81750
rect 8910 81550 8980 81750
rect 9020 81550 9090 81750
rect 9410 81550 9480 81750
rect 9520 81550 9590 81750
rect 9910 81550 9980 81750
rect 10020 81550 10090 81750
rect 10410 81550 10480 81750
rect 10520 81550 10590 81750
rect 10910 81550 10980 81750
rect 11020 81550 11090 81750
rect 11410 81550 11480 81750
rect 11520 81550 11590 81750
rect 11910 81550 11980 81750
rect 12020 81550 12090 81750
rect 12410 81550 12480 81750
rect 12520 81550 12590 81750
rect 12910 81550 12980 81750
rect 13020 81550 13090 81750
rect 13410 81550 13480 81750
rect 13520 81550 13590 81750
rect 13910 81550 13980 81750
rect 14020 81550 14090 81750
rect 14410 81550 14480 81750
rect 14520 81550 14590 81750
rect 14910 81550 14980 81750
rect 15020 81550 15090 81750
rect 15410 81550 15480 81750
rect 15520 81550 15590 81750
rect 15910 81550 15980 81750
rect 16020 81550 16090 81750
rect 16410 81550 16480 81750
rect 16520 81550 16590 81750
rect 16910 81550 16980 81750
rect 17020 81550 17090 81750
rect 17410 81550 17480 81750
rect 17520 81550 17590 81750
rect 17910 81550 17980 81750
rect 18020 81550 18090 81750
rect 18410 81550 18480 81750
rect 18520 81550 18590 81750
rect 18910 81550 18980 81750
rect 19020 81550 19090 81750
rect 19410 81550 19480 81750
rect 19520 81550 19590 81750
rect 19910 81550 19980 81750
rect 20020 81550 20090 81750
rect 20410 81550 20480 81750
rect 20520 81550 20590 81750
rect 20910 81550 20980 81750
rect 21020 81550 21090 81750
rect 21410 81550 21480 81750
rect 21520 81550 21590 81750
rect 21910 81550 21980 81750
rect 22020 81550 22090 81750
rect 22410 81550 22480 81750
rect 22520 81550 22590 81750
rect 22910 81550 22980 81750
rect 23020 81550 23090 81750
rect 23410 81550 23480 81750
rect 23520 81550 23590 81750
rect 23910 81550 23980 81750
rect 24020 81550 24090 81750
rect 24410 81550 24480 81750
rect 24520 81550 24590 81750
rect 24910 81550 24980 81750
rect 25020 81550 25090 81750
rect 25410 81550 25480 81750
rect 25520 81550 25590 81750
rect 25910 81550 25980 81750
rect 26020 81550 26090 81750
rect 26410 81550 26480 81750
rect 26520 81550 26590 81750
rect 26910 81550 26980 81750
rect 27020 81550 27090 81750
rect 27410 81550 27480 81750
rect 27520 81550 27590 81750
rect 27910 81550 27980 81750
rect 28020 81550 28090 81750
rect 28410 81550 28480 81750
rect 28520 81550 28590 81750
rect 28910 81550 28980 81750
rect 29020 81550 29090 81750
rect 29410 81550 29480 81750
rect 29520 81550 29590 81750
rect 29910 81550 29980 81750
rect 30020 81550 30090 81750
rect 30410 81550 30480 81750
rect 30520 81550 30590 81750
rect 30910 81550 30980 81750
rect 31020 81550 31090 81750
rect 31410 81550 31480 81750
rect 31520 81550 31590 81750
rect 31910 81550 31980 81750
rect 32020 81550 32090 81750
rect 32410 81550 32480 81750
rect 32520 81550 32590 81750
rect 32910 81550 32980 81750
rect 33020 81550 33090 81750
rect 33410 81550 33480 81750
rect 33520 81550 33590 81750
rect 33910 81550 33980 81750
rect 34020 81550 34090 81750
rect 34410 81550 34480 81750
rect 34520 81550 34590 81750
rect 34910 81550 34980 81750
rect 35020 81550 35090 81750
rect 35410 81550 35480 81750
rect 35520 81550 35590 81750
rect 35910 81550 35980 81750
rect 36020 81550 36090 81750
rect 36410 81550 36480 81750
rect 36520 81550 36590 81750
rect 36910 81550 36980 81750
rect 37020 81550 37090 81750
rect 37410 81550 37480 81750
rect 37520 81550 37590 81750
rect 37910 81550 37980 81750
rect 38020 81550 38090 81750
rect 38410 81550 38480 81750
rect 38520 81550 38590 81750
rect 38910 81550 38980 81750
rect 39020 81550 39090 81750
rect 39410 81550 39480 81750
rect 39520 81550 39590 81750
rect 39910 81550 39980 81750
rect 40020 81550 40090 81750
rect 40410 81550 40480 81750
rect 40520 81550 40590 81750
rect 40910 81550 40980 81750
rect 41020 81550 41090 81750
rect 41410 81550 41480 81750
rect 41520 81550 41590 81750
rect 41910 81550 41980 81750
rect 42020 81550 42090 81750
rect 42410 81550 42480 81750
rect 42520 81550 42590 81750
rect 42910 81550 42980 81750
rect 43020 81550 43090 81750
rect 43410 81550 43480 81750
rect 43520 81550 43590 81750
rect 43910 81550 43980 81750
rect 44020 81550 44090 81750
rect 44410 81550 44480 81750
rect 44520 81550 44590 81750
rect 44910 81550 44980 81750
rect 45020 81550 45090 81750
rect 45410 81550 45480 81750
rect 45520 81550 45590 81750
rect 45910 81550 45980 81750
rect 46020 81550 46090 81750
rect 46410 81550 46480 81750
rect 46520 81550 46590 81750
rect 46910 81550 46980 81750
rect 47020 81550 47090 81750
rect 47410 81550 47480 81750
rect 47520 81550 47590 81750
rect 47910 81550 47980 81750
rect 48020 81550 48090 81750
rect 48410 81550 48480 81750
rect 48520 81550 48590 81750
rect 48910 81550 48980 81750
rect 49020 81550 49090 81750
rect 49410 81550 49480 81750
rect 49520 81550 49590 81750
rect 49910 81550 49980 81750
rect 50020 81550 50090 81750
rect 50410 81550 50480 81750
rect 50520 81550 50590 81750
rect 50910 81550 50980 81750
rect 51020 81550 51090 81750
rect 51410 81550 51480 81750
rect 51520 81550 51590 81750
rect 51910 81550 51980 81750
rect 52020 81550 52090 81750
rect 52410 81550 52480 81750
rect 52520 81550 52590 81750
rect 52910 81550 52980 81750
rect 53020 81550 53090 81750
rect 53410 81550 53480 81750
rect 53520 81550 53590 81750
rect 53910 81550 53980 81750
rect 54020 81550 54090 81750
rect 54410 81550 54480 81750
rect 54520 81550 54590 81750
rect 54910 81550 54980 81750
rect 55020 81550 55090 81750
rect 55410 81550 55480 81750
rect 55520 81550 55590 81750
rect 55910 81550 55980 81750
rect 56020 81550 56090 81750
rect 56410 81550 56480 81750
rect 56520 81550 56590 81750
rect 56910 81550 56980 81750
rect 57020 81550 57090 81750
rect 57410 81550 57480 81750
rect 57520 81550 57590 81750
rect 57910 81550 57980 81750
rect 58020 81550 58090 81750
rect 58410 81550 58480 81750
rect 58520 81550 58590 81750
rect 58910 81550 58980 81750
rect 59020 81550 59090 81750
rect 59410 81550 59480 81750
rect 59520 81550 59590 81750
rect 59910 81550 59980 81750
rect 60020 81550 60090 81750
rect 60410 81550 60480 81750
rect 60520 81550 60590 81750
rect 60910 81550 60980 81750
rect 61020 81550 61090 81750
rect 61410 81550 61480 81750
rect 61520 81550 61590 81750
rect 61910 81550 61980 81750
rect 62020 81550 62090 81750
rect 62410 81550 62480 81750
rect 62520 81550 62590 81750
rect 62910 81550 62980 81750
rect 63020 81550 63090 81750
rect 63410 81550 63480 81750
rect 63520 81550 63590 81750
rect 63910 81550 63980 81750
rect 64020 81550 64090 81750
rect 64410 81550 64480 81750
rect 64520 81550 64590 81750
rect 64910 81550 64980 81750
rect 65020 81550 65090 81750
rect 65410 81550 65480 81750
rect 65520 81550 65590 81750
rect 65910 81550 65980 81750
rect 66020 81550 66090 81750
rect 66410 81550 66480 81750
rect 66520 81550 66590 81750
rect 66910 81550 66980 81750
rect 67020 81550 67090 81750
rect 67410 81550 67480 81750
rect 67520 81550 67590 81750
rect 67910 81550 67980 81750
rect 68020 81550 68090 81750
rect 68410 81550 68480 81750
rect 68520 81550 68590 81750
rect 68910 81550 68980 81750
rect 69020 81550 69090 81750
rect 69410 81550 69480 81750
rect 69520 81550 69590 81750
rect 69910 81550 69980 81750
rect 70020 81550 70090 81750
rect 70410 81550 70480 81750
rect 70520 81550 70590 81750
rect 70910 81550 70980 81750
rect 71020 81550 71090 81750
rect 71410 81550 71480 81750
rect 71520 81550 71590 81750
rect 71910 81550 71980 81750
rect 72020 81550 72090 81750
rect 72410 81550 72480 81750
rect 72520 81550 72590 81750
rect 72910 81550 72980 81750
rect 73020 81550 73090 81750
rect 73410 81550 73480 81750
rect 73520 81550 73590 81750
rect 73910 81550 73980 81750
rect 74020 81550 74090 81750
rect 74410 81550 74480 81750
rect 74520 81550 74590 81750
rect 74910 81550 74980 81750
rect 75020 81550 75090 81750
rect 75410 81550 75480 81750
rect 75520 81550 75590 81750
rect 75910 81550 75980 81750
rect 76020 81550 76090 81750
rect 76410 81550 76480 81750
rect 76520 81550 76590 81750
rect 76910 81550 76980 81750
rect 77020 81550 77090 81750
rect 77410 81550 77480 81750
rect 77520 81550 77590 81750
rect 77910 81550 77980 81750
rect 78020 81550 78090 81750
rect 78410 81550 78480 81750
rect 78520 81550 78590 81750
rect 78910 81550 78980 81750
rect 79020 81550 79090 81750
rect 79410 81550 79480 81750
rect 79520 81550 79590 81750
rect 79910 81550 79980 81750
rect 80020 81550 80090 81750
rect 80410 81550 80480 81750
rect 80520 81550 80590 81750
rect 80910 81550 80980 81750
rect 81020 81550 81090 81750
rect 81410 81550 81480 81750
rect 81520 81550 81590 81750
rect 81910 81550 81980 81750
rect 82020 81550 82090 81750
rect 82410 81550 82480 81750
rect 82520 81550 82590 81750
rect 82910 81550 82980 81750
rect 83020 81550 83090 81750
rect 83410 81550 83480 81750
rect 83520 81550 83590 81750
rect 83910 81550 83980 81750
rect 84020 81550 84090 81750
rect 84410 81550 84480 81750
rect 84520 81550 84590 81750
rect 84910 81550 84980 81750
rect 85020 81550 85090 81750
rect 85410 81550 85480 81750
rect 85520 81550 85590 81750
rect 85910 81550 85980 81750
rect 86020 81550 86090 81750
rect 86410 81550 86480 81750
rect 86520 81550 86590 81750
rect 86910 81550 86980 81750
rect 87020 81550 87090 81750
rect 87410 81550 87480 81750
rect 87520 81550 87590 81750
rect 87910 81550 87980 81750
rect 88020 81550 88090 81750
rect 88410 81550 88480 81750
rect 88520 81550 88590 81750
rect 88910 81550 88980 81750
rect 89020 81550 89090 81750
rect 89410 81550 89480 81750
rect 89520 81550 89590 81750
rect 89910 81550 89980 81750
rect 90020 81550 90090 81750
rect 90410 81550 90480 81750
rect 90520 81550 90590 81750
rect 90910 81550 90980 81750
rect 91020 81550 91090 81750
rect 91410 81550 91480 81750
rect 91520 81550 91590 81750
rect 91910 81550 91980 81750
rect 92020 81550 92090 81750
rect 92410 81550 92480 81750
rect 92520 81550 92590 81750
rect 92910 81550 92980 81750
rect 93020 81550 93090 81750
rect 93410 81550 93480 81750
rect 93520 81550 93590 81750
rect 93910 81550 93980 81750
rect 94020 81550 94090 81750
rect 94410 81550 94480 81750
rect 94520 81550 94590 81750
rect 94910 81550 94980 81750
rect 95020 81550 95090 81750
rect 95410 81550 95480 81750
rect 95520 81550 95590 81750
rect 95910 81550 95980 81750
rect 96020 81550 96090 81750
rect 96410 81550 96480 81750
rect 96520 81550 96590 81750
rect 96910 81550 96980 81750
rect 97020 81550 97090 81750
rect 97410 81550 97480 81750
rect 97520 81550 97590 81750
rect 97910 81550 97980 81750
rect 98020 81550 98090 81750
rect 98410 81550 98480 81750
rect 98520 81550 98590 81750
rect 98910 81550 98980 81750
rect 99020 81550 99090 81750
rect 99410 81550 99480 81750
rect 99520 81550 99590 81750
rect 99910 81550 99980 81750
rect 100020 81550 100090 81750
rect 100410 81550 100480 81750
rect -83350 81420 -83150 81490
rect -82850 81420 -82650 81490
rect -82350 81420 -82150 81490
rect -81850 81420 -81650 81490
rect -81350 81420 -81150 81490
rect -80850 81420 -80650 81490
rect -80350 81420 -80150 81490
rect -79850 81420 -79650 81490
rect -79350 81420 -79150 81490
rect -78850 81420 -78650 81490
rect -78350 81420 -78150 81490
rect -77850 81420 -77650 81490
rect -77350 81420 -77150 81490
rect -76850 81420 -76650 81490
rect -76350 81420 -76150 81490
rect -75850 81420 -75650 81490
rect -75350 81420 -75150 81490
rect -74850 81420 -74650 81490
rect -74350 81420 -74150 81490
rect -73850 81420 -73650 81490
rect -73350 81420 -73150 81490
rect -72850 81420 -72650 81490
rect -72350 81420 -72150 81490
rect -71850 81420 -71650 81490
rect -71350 81420 -71150 81490
rect -70850 81420 -70650 81490
rect -70350 81420 -70150 81490
rect -69850 81420 -69650 81490
rect -69350 81420 -69150 81490
rect -68850 81420 -68650 81490
rect -68350 81420 -68150 81490
rect -67850 81420 -67650 81490
rect -67350 81420 -67150 81490
rect -66850 81420 -66650 81490
rect -66350 81420 -66150 81490
rect -65850 81420 -65650 81490
rect -65350 81420 -65150 81490
rect -64850 81420 -64650 81490
rect -64350 81420 -64150 81490
rect -63850 81420 -63650 81490
rect -63350 81420 -63150 81490
rect -62850 81420 -62650 81490
rect -62350 81420 -62150 81490
rect -61850 81420 -61650 81490
rect -61350 81420 -61150 81490
rect -60850 81420 -60650 81490
rect -60350 81420 -60150 81490
rect -59850 81420 -59650 81490
rect -59350 81420 -59150 81490
rect -58850 81420 -58650 81490
rect -58350 81420 -58150 81490
rect -57850 81420 -57650 81490
rect -57350 81420 -57150 81490
rect -56850 81420 -56650 81490
rect -56350 81420 -56150 81490
rect -55850 81420 -55650 81490
rect -55350 81420 -55150 81490
rect -54850 81420 -54650 81490
rect -54350 81420 -54150 81490
rect -53850 81420 -53650 81490
rect -53350 81420 -53150 81490
rect -52850 81420 -52650 81490
rect -52350 81420 -52150 81490
rect -51850 81420 -51650 81490
rect -51350 81420 -51150 81490
rect -50850 81420 -50650 81490
rect -50350 81420 -50150 81490
rect -49850 81420 -49650 81490
rect -49350 81420 -49150 81490
rect -48850 81420 -48650 81490
rect -48350 81420 -48150 81490
rect -47850 81420 -47650 81490
rect -47350 81420 -47150 81490
rect -46850 81420 -46650 81490
rect -46350 81420 -46150 81490
rect -45850 81420 -45650 81490
rect -45350 81420 -45150 81490
rect -44850 81420 -44650 81490
rect -44350 81420 -44150 81490
rect -43850 81420 -43650 81490
rect -43350 81420 -43150 81490
rect -42850 81420 -42650 81490
rect -42350 81420 -42150 81490
rect -41850 81420 -41650 81490
rect -41350 81420 -41150 81490
rect -40850 81420 -40650 81490
rect -40350 81420 -40150 81490
rect -39850 81420 -39650 81490
rect -39350 81420 -39150 81490
rect -38850 81420 -38650 81490
rect -38350 81420 -38150 81490
rect -37850 81420 -37650 81490
rect -37350 81420 -37150 81490
rect -36850 81420 -36650 81490
rect -36350 81420 -36150 81490
rect -35850 81420 -35650 81490
rect -35350 81420 -35150 81490
rect -34850 81420 -34650 81490
rect -34350 81420 -34150 81490
rect -33850 81420 -33650 81490
rect -33350 81420 -33150 81490
rect -32850 81420 -32650 81490
rect -32350 81420 -32150 81490
rect -31850 81420 -31650 81490
rect -31350 81420 -31150 81490
rect -30850 81420 -30650 81490
rect -30350 81420 -30150 81490
rect -29850 81420 -29650 81490
rect -29350 81420 -29150 81490
rect -28850 81420 -28650 81490
rect -28350 81420 -28150 81490
rect -27850 81420 -27650 81490
rect -27350 81420 -27150 81490
rect -26850 81420 -26650 81490
rect -26350 81420 -26150 81490
rect -25850 81420 -25650 81490
rect -25350 81420 -25150 81490
rect -24850 81420 -24650 81490
rect -24350 81420 -24150 81490
rect -23850 81420 -23650 81490
rect -23350 81420 -23150 81490
rect -22850 81420 -22650 81490
rect -22350 81420 -22150 81490
rect -21850 81420 -21650 81490
rect -21350 81420 -21150 81490
rect -20850 81420 -20650 81490
rect -20350 81420 -20150 81490
rect -19850 81420 -19650 81490
rect -19350 81420 -19150 81490
rect -18850 81420 -18650 81490
rect -18350 81420 -18150 81490
rect -17850 81420 -17650 81490
rect -17350 81420 -17150 81490
rect -16850 81420 -16650 81490
rect -16350 81420 -16150 81490
rect -15850 81420 -15650 81490
rect -15350 81420 -15150 81490
rect -14850 81420 -14650 81490
rect -14350 81420 -14150 81490
rect -13850 81420 -13650 81490
rect -13350 81420 -13150 81490
rect -12850 81420 -12650 81490
rect -12350 81420 -12150 81490
rect -11850 81420 -11650 81490
rect -11350 81420 -11150 81490
rect -10850 81420 -10650 81490
rect -10350 81420 -10150 81490
rect -9850 81420 -9650 81490
rect -9350 81420 -9150 81490
rect -8850 81420 -8650 81490
rect -8350 81420 -8150 81490
rect -7850 81420 -7650 81490
rect -7350 81420 -7150 81490
rect -6850 81420 -6650 81490
rect -6350 81420 -6150 81490
rect -5850 81420 -5650 81490
rect -5350 81420 -5150 81490
rect -4850 81420 -4650 81490
rect -4350 81420 -4150 81490
rect -3850 81420 -3650 81490
rect -3350 81420 -3150 81490
rect -2850 81420 -2650 81490
rect -2350 81420 -2150 81490
rect -1850 81420 -1650 81490
rect -1350 81420 -1150 81490
rect -850 81420 -650 81490
rect -350 81420 -150 81490
rect 150 81420 350 81490
rect 650 81420 850 81490
rect 1150 81420 1350 81490
rect 1650 81420 1850 81490
rect 2150 81420 2350 81490
rect 2650 81420 2850 81490
rect 3150 81420 3350 81490
rect 3650 81420 3850 81490
rect 4150 81420 4350 81490
rect 4650 81420 4850 81490
rect 5150 81420 5350 81490
rect 5650 81420 5850 81490
rect 6150 81420 6350 81490
rect 6650 81420 6850 81490
rect 7150 81420 7350 81490
rect 7650 81420 7850 81490
rect 8150 81420 8350 81490
rect 8650 81420 8850 81490
rect 9150 81420 9350 81490
rect 9650 81420 9850 81490
rect 10150 81420 10350 81490
rect 10650 81420 10850 81490
rect 11150 81420 11350 81490
rect 11650 81420 11850 81490
rect 12150 81420 12350 81490
rect 12650 81420 12850 81490
rect 13150 81420 13350 81490
rect 13650 81420 13850 81490
rect 14150 81420 14350 81490
rect 14650 81420 14850 81490
rect 15150 81420 15350 81490
rect 15650 81420 15850 81490
rect 16150 81420 16350 81490
rect 16650 81420 16850 81490
rect 17150 81420 17350 81490
rect 17650 81420 17850 81490
rect 18150 81420 18350 81490
rect 18650 81420 18850 81490
rect 19150 81420 19350 81490
rect 19650 81420 19850 81490
rect 20150 81420 20350 81490
rect 20650 81420 20850 81490
rect 21150 81420 21350 81490
rect 21650 81420 21850 81490
rect 22150 81420 22350 81490
rect 22650 81420 22850 81490
rect 23150 81420 23350 81490
rect 23650 81420 23850 81490
rect 24150 81420 24350 81490
rect 24650 81420 24850 81490
rect 25150 81420 25350 81490
rect 25650 81420 25850 81490
rect 26150 81420 26350 81490
rect 26650 81420 26850 81490
rect 27150 81420 27350 81490
rect 27650 81420 27850 81490
rect 28150 81420 28350 81490
rect 28650 81420 28850 81490
rect 29150 81420 29350 81490
rect 29650 81420 29850 81490
rect 30150 81420 30350 81490
rect 30650 81420 30850 81490
rect 31150 81420 31350 81490
rect 31650 81420 31850 81490
rect 32150 81420 32350 81490
rect 32650 81420 32850 81490
rect 33150 81420 33350 81490
rect 33650 81420 33850 81490
rect 34150 81420 34350 81490
rect 34650 81420 34850 81490
rect 35150 81420 35350 81490
rect 35650 81420 35850 81490
rect 36150 81420 36350 81490
rect 36650 81420 36850 81490
rect 37150 81420 37350 81490
rect 37650 81420 37850 81490
rect 38150 81420 38350 81490
rect 38650 81420 38850 81490
rect 39150 81420 39350 81490
rect 39650 81420 39850 81490
rect 40150 81420 40350 81490
rect 40650 81420 40850 81490
rect 41150 81420 41350 81490
rect 41650 81420 41850 81490
rect 42150 81420 42350 81490
rect 42650 81420 42850 81490
rect 43150 81420 43350 81490
rect 43650 81420 43850 81490
rect 44150 81420 44350 81490
rect 44650 81420 44850 81490
rect 45150 81420 45350 81490
rect 45650 81420 45850 81490
rect 46150 81420 46350 81490
rect 46650 81420 46850 81490
rect 47150 81420 47350 81490
rect 47650 81420 47850 81490
rect 48150 81420 48350 81490
rect 48650 81420 48850 81490
rect 49150 81420 49350 81490
rect 49650 81420 49850 81490
rect 50150 81420 50350 81490
rect 50650 81420 50850 81490
rect 51150 81420 51350 81490
rect 51650 81420 51850 81490
rect 52150 81420 52350 81490
rect 52650 81420 52850 81490
rect 53150 81420 53350 81490
rect 53650 81420 53850 81490
rect 54150 81420 54350 81490
rect 54650 81420 54850 81490
rect 55150 81420 55350 81490
rect 55650 81420 55850 81490
rect 56150 81420 56350 81490
rect 56650 81420 56850 81490
rect 57150 81420 57350 81490
rect 57650 81420 57850 81490
rect 58150 81420 58350 81490
rect 58650 81420 58850 81490
rect 59150 81420 59350 81490
rect 59650 81420 59850 81490
rect 60150 81420 60350 81490
rect 60650 81420 60850 81490
rect 61150 81420 61350 81490
rect 61650 81420 61850 81490
rect 62150 81420 62350 81490
rect 62650 81420 62850 81490
rect 63150 81420 63350 81490
rect 63650 81420 63850 81490
rect 64150 81420 64350 81490
rect 64650 81420 64850 81490
rect 65150 81420 65350 81490
rect 65650 81420 65850 81490
rect 66150 81420 66350 81490
rect 66650 81420 66850 81490
rect 67150 81420 67350 81490
rect 67650 81420 67850 81490
rect 68150 81420 68350 81490
rect 68650 81420 68850 81490
rect 69150 81420 69350 81490
rect 69650 81420 69850 81490
rect 70150 81420 70350 81490
rect 70650 81420 70850 81490
rect 71150 81420 71350 81490
rect 71650 81420 71850 81490
rect 72150 81420 72350 81490
rect 72650 81420 72850 81490
rect 73150 81420 73350 81490
rect 73650 81420 73850 81490
rect 74150 81420 74350 81490
rect 74650 81420 74850 81490
rect 75150 81420 75350 81490
rect 75650 81420 75850 81490
rect 76150 81420 76350 81490
rect 76650 81420 76850 81490
rect 77150 81420 77350 81490
rect 77650 81420 77850 81490
rect 78150 81420 78350 81490
rect 78650 81420 78850 81490
rect 79150 81420 79350 81490
rect 79650 81420 79850 81490
rect 80150 81420 80350 81490
rect 80650 81420 80850 81490
rect 81150 81420 81350 81490
rect 81650 81420 81850 81490
rect 82150 81420 82350 81490
rect 82650 81420 82850 81490
rect 83150 81420 83350 81490
rect 83650 81420 83850 81490
rect 84150 81420 84350 81490
rect 84650 81420 84850 81490
rect 85150 81420 85350 81490
rect 85650 81420 85850 81490
rect 86150 81420 86350 81490
rect 86650 81420 86850 81490
rect 87150 81420 87350 81490
rect 87650 81420 87850 81490
rect 88150 81420 88350 81490
rect 88650 81420 88850 81490
rect 89150 81420 89350 81490
rect 89650 81420 89850 81490
rect 90150 81420 90350 81490
rect 90650 81420 90850 81490
rect 91150 81420 91350 81490
rect 91650 81420 91850 81490
rect 92150 81420 92350 81490
rect 92650 81420 92850 81490
rect 93150 81420 93350 81490
rect 93650 81420 93850 81490
rect 94150 81420 94350 81490
rect 94650 81420 94850 81490
rect 95150 81420 95350 81490
rect 95650 81420 95850 81490
rect 96150 81420 96350 81490
rect 96650 81420 96850 81490
rect 97150 81420 97350 81490
rect 97650 81420 97850 81490
rect 98150 81420 98350 81490
rect 98650 81420 98850 81490
rect 99150 81420 99350 81490
rect 99650 81420 99850 81490
rect 100150 81420 100350 81490
rect -83350 81310 -83150 81380
rect -82850 81310 -82650 81380
rect -82350 81310 -82150 81380
rect -81850 81310 -81650 81380
rect -81350 81310 -81150 81380
rect -80850 81310 -80650 81380
rect -80350 81310 -80150 81380
rect -79850 81310 -79650 81380
rect -79350 81310 -79150 81380
rect -78850 81310 -78650 81380
rect -78350 81310 -78150 81380
rect -77850 81310 -77650 81380
rect -77350 81310 -77150 81380
rect -76850 81310 -76650 81380
rect -76350 81310 -76150 81380
rect -75850 81310 -75650 81380
rect -75350 81310 -75150 81380
rect -74850 81310 -74650 81380
rect -74350 81310 -74150 81380
rect -73850 81310 -73650 81380
rect -73350 81310 -73150 81380
rect -72850 81310 -72650 81380
rect -72350 81310 -72150 81380
rect -71850 81310 -71650 81380
rect -71350 81310 -71150 81380
rect -70850 81310 -70650 81380
rect -70350 81310 -70150 81380
rect -69850 81310 -69650 81380
rect -69350 81310 -69150 81380
rect -68850 81310 -68650 81380
rect -68350 81310 -68150 81380
rect -67850 81310 -67650 81380
rect -67350 81310 -67150 81380
rect -66850 81310 -66650 81380
rect -66350 81310 -66150 81380
rect -65850 81310 -65650 81380
rect -65350 81310 -65150 81380
rect -64850 81310 -64650 81380
rect -64350 81310 -64150 81380
rect -63850 81310 -63650 81380
rect -63350 81310 -63150 81380
rect -62850 81310 -62650 81380
rect -62350 81310 -62150 81380
rect -61850 81310 -61650 81380
rect -61350 81310 -61150 81380
rect -60850 81310 -60650 81380
rect -60350 81310 -60150 81380
rect -59850 81310 -59650 81380
rect -59350 81310 -59150 81380
rect -58850 81310 -58650 81380
rect -58350 81310 -58150 81380
rect -57850 81310 -57650 81380
rect -57350 81310 -57150 81380
rect -56850 81310 -56650 81380
rect -56350 81310 -56150 81380
rect -55850 81310 -55650 81380
rect -55350 81310 -55150 81380
rect -54850 81310 -54650 81380
rect -54350 81310 -54150 81380
rect -53850 81310 -53650 81380
rect -53350 81310 -53150 81380
rect -52850 81310 -52650 81380
rect -52350 81310 -52150 81380
rect -51850 81310 -51650 81380
rect -51350 81310 -51150 81380
rect -50850 81310 -50650 81380
rect -50350 81310 -50150 81380
rect -49850 81310 -49650 81380
rect -49350 81310 -49150 81380
rect -48850 81310 -48650 81380
rect -48350 81310 -48150 81380
rect -47850 81310 -47650 81380
rect -47350 81310 -47150 81380
rect -46850 81310 -46650 81380
rect -46350 81310 -46150 81380
rect -45850 81310 -45650 81380
rect -45350 81310 -45150 81380
rect -44850 81310 -44650 81380
rect -44350 81310 -44150 81380
rect -43850 81310 -43650 81380
rect -43350 81310 -43150 81380
rect -42850 81310 -42650 81380
rect -42350 81310 -42150 81380
rect -41850 81310 -41650 81380
rect -41350 81310 -41150 81380
rect -40850 81310 -40650 81380
rect -40350 81310 -40150 81380
rect -39850 81310 -39650 81380
rect -39350 81310 -39150 81380
rect -38850 81310 -38650 81380
rect -38350 81310 -38150 81380
rect -37850 81310 -37650 81380
rect -37350 81310 -37150 81380
rect -36850 81310 -36650 81380
rect -36350 81310 -36150 81380
rect -35850 81310 -35650 81380
rect -35350 81310 -35150 81380
rect -34850 81310 -34650 81380
rect -34350 81310 -34150 81380
rect -33850 81310 -33650 81380
rect -33350 81310 -33150 81380
rect -32850 81310 -32650 81380
rect -32350 81310 -32150 81380
rect -31850 81310 -31650 81380
rect -31350 81310 -31150 81380
rect -30850 81310 -30650 81380
rect -30350 81310 -30150 81380
rect -29850 81310 -29650 81380
rect -29350 81310 -29150 81380
rect -28850 81310 -28650 81380
rect -28350 81310 -28150 81380
rect -27850 81310 -27650 81380
rect -27350 81310 -27150 81380
rect -26850 81310 -26650 81380
rect -26350 81310 -26150 81380
rect -25850 81310 -25650 81380
rect -25350 81310 -25150 81380
rect -24850 81310 -24650 81380
rect -24350 81310 -24150 81380
rect -23850 81310 -23650 81380
rect -23350 81310 -23150 81380
rect -22850 81310 -22650 81380
rect -22350 81310 -22150 81380
rect -21850 81310 -21650 81380
rect -21350 81310 -21150 81380
rect -20850 81310 -20650 81380
rect -20350 81310 -20150 81380
rect -19850 81310 -19650 81380
rect -19350 81310 -19150 81380
rect -18850 81310 -18650 81380
rect -18350 81310 -18150 81380
rect -17850 81310 -17650 81380
rect -17350 81310 -17150 81380
rect -16850 81310 -16650 81380
rect -16350 81310 -16150 81380
rect -15850 81310 -15650 81380
rect -15350 81310 -15150 81380
rect -14850 81310 -14650 81380
rect -14350 81310 -14150 81380
rect -13850 81310 -13650 81380
rect -13350 81310 -13150 81380
rect -12850 81310 -12650 81380
rect -12350 81310 -12150 81380
rect -11850 81310 -11650 81380
rect -11350 81310 -11150 81380
rect -10850 81310 -10650 81380
rect -10350 81310 -10150 81380
rect -9850 81310 -9650 81380
rect -9350 81310 -9150 81380
rect -8850 81310 -8650 81380
rect -8350 81310 -8150 81380
rect -7850 81310 -7650 81380
rect -7350 81310 -7150 81380
rect -6850 81310 -6650 81380
rect -6350 81310 -6150 81380
rect -5850 81310 -5650 81380
rect -5350 81310 -5150 81380
rect -4850 81310 -4650 81380
rect -4350 81310 -4150 81380
rect -3850 81310 -3650 81380
rect -3350 81310 -3150 81380
rect -2850 81310 -2650 81380
rect -2350 81310 -2150 81380
rect -1850 81310 -1650 81380
rect -1350 81310 -1150 81380
rect -850 81310 -650 81380
rect -350 81310 -150 81380
rect 150 81310 350 81380
rect 650 81310 850 81380
rect 1150 81310 1350 81380
rect 1650 81310 1850 81380
rect 2150 81310 2350 81380
rect 2650 81310 2850 81380
rect 3150 81310 3350 81380
rect 3650 81310 3850 81380
rect 4150 81310 4350 81380
rect 4650 81310 4850 81380
rect 5150 81310 5350 81380
rect 5650 81310 5850 81380
rect 6150 81310 6350 81380
rect 6650 81310 6850 81380
rect 7150 81310 7350 81380
rect 7650 81310 7850 81380
rect 8150 81310 8350 81380
rect 8650 81310 8850 81380
rect 9150 81310 9350 81380
rect 9650 81310 9850 81380
rect 10150 81310 10350 81380
rect 10650 81310 10850 81380
rect 11150 81310 11350 81380
rect 11650 81310 11850 81380
rect 12150 81310 12350 81380
rect 12650 81310 12850 81380
rect 13150 81310 13350 81380
rect 13650 81310 13850 81380
rect 14150 81310 14350 81380
rect 14650 81310 14850 81380
rect 15150 81310 15350 81380
rect 15650 81310 15850 81380
rect 16150 81310 16350 81380
rect 16650 81310 16850 81380
rect 17150 81310 17350 81380
rect 17650 81310 17850 81380
rect 18150 81310 18350 81380
rect 18650 81310 18850 81380
rect 19150 81310 19350 81380
rect 19650 81310 19850 81380
rect 20150 81310 20350 81380
rect 20650 81310 20850 81380
rect 21150 81310 21350 81380
rect 21650 81310 21850 81380
rect 22150 81310 22350 81380
rect 22650 81310 22850 81380
rect 23150 81310 23350 81380
rect 23650 81310 23850 81380
rect 24150 81310 24350 81380
rect 24650 81310 24850 81380
rect 25150 81310 25350 81380
rect 25650 81310 25850 81380
rect 26150 81310 26350 81380
rect 26650 81310 26850 81380
rect 27150 81310 27350 81380
rect 27650 81310 27850 81380
rect 28150 81310 28350 81380
rect 28650 81310 28850 81380
rect 29150 81310 29350 81380
rect 29650 81310 29850 81380
rect 30150 81310 30350 81380
rect 30650 81310 30850 81380
rect 31150 81310 31350 81380
rect 31650 81310 31850 81380
rect 32150 81310 32350 81380
rect 32650 81310 32850 81380
rect 33150 81310 33350 81380
rect 33650 81310 33850 81380
rect 34150 81310 34350 81380
rect 34650 81310 34850 81380
rect 35150 81310 35350 81380
rect 35650 81310 35850 81380
rect 36150 81310 36350 81380
rect 36650 81310 36850 81380
rect 37150 81310 37350 81380
rect 37650 81310 37850 81380
rect 38150 81310 38350 81380
rect 38650 81310 38850 81380
rect 39150 81310 39350 81380
rect 39650 81310 39850 81380
rect 40150 81310 40350 81380
rect 40650 81310 40850 81380
rect 41150 81310 41350 81380
rect 41650 81310 41850 81380
rect 42150 81310 42350 81380
rect 42650 81310 42850 81380
rect 43150 81310 43350 81380
rect 43650 81310 43850 81380
rect 44150 81310 44350 81380
rect 44650 81310 44850 81380
rect 45150 81310 45350 81380
rect 45650 81310 45850 81380
rect 46150 81310 46350 81380
rect 46650 81310 46850 81380
rect 47150 81310 47350 81380
rect 47650 81310 47850 81380
rect 48150 81310 48350 81380
rect 48650 81310 48850 81380
rect 49150 81310 49350 81380
rect 49650 81310 49850 81380
rect 50150 81310 50350 81380
rect 50650 81310 50850 81380
rect 51150 81310 51350 81380
rect 51650 81310 51850 81380
rect 52150 81310 52350 81380
rect 52650 81310 52850 81380
rect 53150 81310 53350 81380
rect 53650 81310 53850 81380
rect 54150 81310 54350 81380
rect 54650 81310 54850 81380
rect 55150 81310 55350 81380
rect 55650 81310 55850 81380
rect 56150 81310 56350 81380
rect 56650 81310 56850 81380
rect 57150 81310 57350 81380
rect 57650 81310 57850 81380
rect 58150 81310 58350 81380
rect 58650 81310 58850 81380
rect 59150 81310 59350 81380
rect 59650 81310 59850 81380
rect 60150 81310 60350 81380
rect 60650 81310 60850 81380
rect 61150 81310 61350 81380
rect 61650 81310 61850 81380
rect 62150 81310 62350 81380
rect 62650 81310 62850 81380
rect 63150 81310 63350 81380
rect 63650 81310 63850 81380
rect 64150 81310 64350 81380
rect 64650 81310 64850 81380
rect 65150 81310 65350 81380
rect 65650 81310 65850 81380
rect 66150 81310 66350 81380
rect 66650 81310 66850 81380
rect 67150 81310 67350 81380
rect 67650 81310 67850 81380
rect 68150 81310 68350 81380
rect 68650 81310 68850 81380
rect 69150 81310 69350 81380
rect 69650 81310 69850 81380
rect 70150 81310 70350 81380
rect 70650 81310 70850 81380
rect 71150 81310 71350 81380
rect 71650 81310 71850 81380
rect 72150 81310 72350 81380
rect 72650 81310 72850 81380
rect 73150 81310 73350 81380
rect 73650 81310 73850 81380
rect 74150 81310 74350 81380
rect 74650 81310 74850 81380
rect 75150 81310 75350 81380
rect 75650 81310 75850 81380
rect 76150 81310 76350 81380
rect 76650 81310 76850 81380
rect 77150 81310 77350 81380
rect 77650 81310 77850 81380
rect 78150 81310 78350 81380
rect 78650 81310 78850 81380
rect 79150 81310 79350 81380
rect 79650 81310 79850 81380
rect 80150 81310 80350 81380
rect 80650 81310 80850 81380
rect 81150 81310 81350 81380
rect 81650 81310 81850 81380
rect 82150 81310 82350 81380
rect 82650 81310 82850 81380
rect 83150 81310 83350 81380
rect 83650 81310 83850 81380
rect 84150 81310 84350 81380
rect 84650 81310 84850 81380
rect 85150 81310 85350 81380
rect 85650 81310 85850 81380
rect 86150 81310 86350 81380
rect 86650 81310 86850 81380
rect 87150 81310 87350 81380
rect 87650 81310 87850 81380
rect 88150 81310 88350 81380
rect 88650 81310 88850 81380
rect 89150 81310 89350 81380
rect 89650 81310 89850 81380
rect 90150 81310 90350 81380
rect 90650 81310 90850 81380
rect 91150 81310 91350 81380
rect 91650 81310 91850 81380
rect 92150 81310 92350 81380
rect 92650 81310 92850 81380
rect 93150 81310 93350 81380
rect 93650 81310 93850 81380
rect 94150 81310 94350 81380
rect 94650 81310 94850 81380
rect 95150 81310 95350 81380
rect 95650 81310 95850 81380
rect 96150 81310 96350 81380
rect 96650 81310 96850 81380
rect 97150 81310 97350 81380
rect 97650 81310 97850 81380
rect 98150 81310 98350 81380
rect 98650 81310 98850 81380
rect 99150 81310 99350 81380
rect 99650 81310 99850 81380
rect 100150 81310 100350 81380
rect -83480 81050 -83410 81250
rect -83090 81050 -83020 81250
rect -82980 81050 -82910 81250
rect -82590 81050 -82520 81250
rect -82480 81050 -82410 81250
rect -82090 81050 -82020 81250
rect -81980 81050 -81910 81250
rect -81590 81050 -81520 81250
rect -81480 81050 -81410 81250
rect -81090 81050 -81020 81250
rect -80980 81050 -80910 81250
rect -80590 81050 -80520 81250
rect -80480 81050 -80410 81250
rect -80090 81050 -80020 81250
rect -79980 81050 -79910 81250
rect -79590 81050 -79520 81250
rect -79480 81050 -79410 81250
rect -79090 81050 -79020 81250
rect -78980 81050 -78910 81250
rect -78590 81050 -78520 81250
rect -78480 81050 -78410 81250
rect -78090 81050 -78020 81250
rect -77980 81050 -77910 81250
rect -77590 81050 -77520 81250
rect -77480 81050 -77410 81250
rect -77090 81050 -77020 81250
rect -76980 81050 -76910 81250
rect -76590 81050 -76520 81250
rect -76480 81050 -76410 81250
rect -76090 81050 -76020 81250
rect -75980 81050 -75910 81250
rect -75590 81050 -75520 81250
rect -75480 81050 -75410 81250
rect -75090 81050 -75020 81250
rect -74980 81050 -74910 81250
rect -74590 81050 -74520 81250
rect -74480 81050 -74410 81250
rect -74090 81050 -74020 81250
rect -73980 81050 -73910 81250
rect -73590 81050 -73520 81250
rect -73480 81050 -73410 81250
rect -73090 81050 -73020 81250
rect -72980 81050 -72910 81250
rect -72590 81050 -72520 81250
rect -72480 81050 -72410 81250
rect -72090 81050 -72020 81250
rect -71980 81050 -71910 81250
rect -71590 81050 -71520 81250
rect -71480 81050 -71410 81250
rect -71090 81050 -71020 81250
rect -70980 81050 -70910 81250
rect -70590 81050 -70520 81250
rect -70480 81050 -70410 81250
rect -70090 81050 -70020 81250
rect -69980 81050 -69910 81250
rect -69590 81050 -69520 81250
rect -69480 81050 -69410 81250
rect -69090 81050 -69020 81250
rect -68980 81050 -68910 81250
rect -68590 81050 -68520 81250
rect -68480 81050 -68410 81250
rect -68090 81050 -68020 81250
rect -67980 81050 -67910 81250
rect -67590 81050 -67520 81250
rect -67480 81050 -67410 81250
rect -67090 81050 -67020 81250
rect -66980 81050 -66910 81250
rect -66590 81050 -66520 81250
rect -66480 81050 -66410 81250
rect -66090 81050 -66020 81250
rect -65980 81050 -65910 81250
rect -65590 81050 -65520 81250
rect -65480 81050 -65410 81250
rect -65090 81050 -65020 81250
rect -64980 81050 -64910 81250
rect -64590 81050 -64520 81250
rect -64480 81050 -64410 81250
rect -64090 81050 -64020 81250
rect -63980 81050 -63910 81250
rect -63590 81050 -63520 81250
rect -63480 81050 -63410 81250
rect -63090 81050 -63020 81250
rect -62980 81050 -62910 81250
rect -62590 81050 -62520 81250
rect -62480 81050 -62410 81250
rect -62090 81050 -62020 81250
rect -61980 81050 -61910 81250
rect -61590 81050 -61520 81250
rect -61480 81050 -61410 81250
rect -61090 81050 -61020 81250
rect -60980 81050 -60910 81250
rect -60590 81050 -60520 81250
rect -60480 81050 -60410 81250
rect -60090 81050 -60020 81250
rect -59980 81050 -59910 81250
rect -59590 81050 -59520 81250
rect -59480 81050 -59410 81250
rect -59090 81050 -59020 81250
rect -58980 81050 -58910 81250
rect -58590 81050 -58520 81250
rect -58480 81050 -58410 81250
rect -58090 81050 -58020 81250
rect -57980 81050 -57910 81250
rect -57590 81050 -57520 81250
rect -57480 81050 -57410 81250
rect -57090 81050 -57020 81250
rect -56980 81050 -56910 81250
rect -56590 81050 -56520 81250
rect -56480 81050 -56410 81250
rect -56090 81050 -56020 81250
rect -55980 81050 -55910 81250
rect -55590 81050 -55520 81250
rect -55480 81050 -55410 81250
rect -55090 81050 -55020 81250
rect -54980 81050 -54910 81250
rect -54590 81050 -54520 81250
rect -54480 81050 -54410 81250
rect -54090 81050 -54020 81250
rect -53980 81050 -53910 81250
rect -53590 81050 -53520 81250
rect -53480 81050 -53410 81250
rect -53090 81050 -53020 81250
rect -52980 81050 -52910 81250
rect -52590 81050 -52520 81250
rect -52480 81050 -52410 81250
rect -52090 81050 -52020 81250
rect -51980 81050 -51910 81250
rect -51590 81050 -51520 81250
rect -51480 81050 -51410 81250
rect -51090 81050 -51020 81250
rect -50980 81050 -50910 81250
rect -50590 81050 -50520 81250
rect -50480 81050 -50410 81250
rect -50090 81050 -50020 81250
rect -49980 81050 -49910 81250
rect -49590 81050 -49520 81250
rect -49480 81050 -49410 81250
rect -49090 81050 -49020 81250
rect -48980 81050 -48910 81250
rect -48590 81050 -48520 81250
rect -48480 81050 -48410 81250
rect -48090 81050 -48020 81250
rect -47980 81050 -47910 81250
rect -47590 81050 -47520 81250
rect -47480 81050 -47410 81250
rect -47090 81050 -47020 81250
rect -46980 81050 -46910 81250
rect -46590 81050 -46520 81250
rect -46480 81050 -46410 81250
rect -46090 81050 -46020 81250
rect -45980 81050 -45910 81250
rect -45590 81050 -45520 81250
rect -45480 81050 -45410 81250
rect -45090 81050 -45020 81250
rect -44980 81050 -44910 81250
rect -44590 81050 -44520 81250
rect -44480 81050 -44410 81250
rect -44090 81050 -44020 81250
rect -43980 81050 -43910 81250
rect -43590 81050 -43520 81250
rect -43480 81050 -43410 81250
rect -43090 81050 -43020 81250
rect -42980 81050 -42910 81250
rect -42590 81050 -42520 81250
rect -42480 81050 -42410 81250
rect -42090 81050 -42020 81250
rect -41980 81050 -41910 81250
rect -41590 81050 -41520 81250
rect -41480 81050 -41410 81250
rect -41090 81050 -41020 81250
rect -40980 81050 -40910 81250
rect -40590 81050 -40520 81250
rect -40480 81050 -40410 81250
rect -40090 81050 -40020 81250
rect -39980 81050 -39910 81250
rect -39590 81050 -39520 81250
rect -39480 81050 -39410 81250
rect -39090 81050 -39020 81250
rect -38980 81050 -38910 81250
rect -38590 81050 -38520 81250
rect -38480 81050 -38410 81250
rect -38090 81050 -38020 81250
rect -37980 81050 -37910 81250
rect -37590 81050 -37520 81250
rect -37480 81050 -37410 81250
rect -37090 81050 -37020 81250
rect -36980 81050 -36910 81250
rect -36590 81050 -36520 81250
rect -36480 81050 -36410 81250
rect -36090 81050 -36020 81250
rect -35980 81050 -35910 81250
rect -35590 81050 -35520 81250
rect -35480 81050 -35410 81250
rect -35090 81050 -35020 81250
rect -34980 81050 -34910 81250
rect -34590 81050 -34520 81250
rect -34480 81050 -34410 81250
rect -34090 81050 -34020 81250
rect -33980 81050 -33910 81250
rect -33590 81050 -33520 81250
rect -33480 81050 -33410 81250
rect -33090 81050 -33020 81250
rect -32980 81050 -32910 81250
rect -32590 81050 -32520 81250
rect -32480 81050 -32410 81250
rect -32090 81050 -32020 81250
rect -31980 81050 -31910 81250
rect -31590 81050 -31520 81250
rect -31480 81050 -31410 81250
rect -31090 81050 -31020 81250
rect -30980 81050 -30910 81250
rect -30590 81050 -30520 81250
rect -30480 81050 -30410 81250
rect -30090 81050 -30020 81250
rect -29980 81050 -29910 81250
rect -29590 81050 -29520 81250
rect -29480 81050 -29410 81250
rect -29090 81050 -29020 81250
rect -28980 81050 -28910 81250
rect -28590 81050 -28520 81250
rect -28480 81050 -28410 81250
rect -28090 81050 -28020 81250
rect -27980 81050 -27910 81250
rect -27590 81050 -27520 81250
rect -27480 81050 -27410 81250
rect -27090 81050 -27020 81250
rect -26980 81050 -26910 81250
rect -26590 81050 -26520 81250
rect -26480 81050 -26410 81250
rect -26090 81050 -26020 81250
rect -25980 81050 -25910 81250
rect -25590 81050 -25520 81250
rect -25480 81050 -25410 81250
rect -25090 81050 -25020 81250
rect -24980 81050 -24910 81250
rect -24590 81050 -24520 81250
rect -24480 81050 -24410 81250
rect -24090 81050 -24020 81250
rect -23980 81050 -23910 81250
rect -23590 81050 -23520 81250
rect -23480 81050 -23410 81250
rect -23090 81050 -23020 81250
rect -22980 81050 -22910 81250
rect -22590 81050 -22520 81250
rect -22480 81050 -22410 81250
rect -22090 81050 -22020 81250
rect -21980 81050 -21910 81250
rect -21590 81050 -21520 81250
rect -21480 81050 -21410 81250
rect -21090 81050 -21020 81250
rect -20980 81050 -20910 81250
rect -20590 81050 -20520 81250
rect -20480 81050 -20410 81250
rect -20090 81050 -20020 81250
rect -19980 81050 -19910 81250
rect -19590 81050 -19520 81250
rect -19480 81050 -19410 81250
rect -19090 81050 -19020 81250
rect -18980 81050 -18910 81250
rect -18590 81050 -18520 81250
rect -18480 81050 -18410 81250
rect -18090 81050 -18020 81250
rect -17980 81050 -17910 81250
rect -17590 81050 -17520 81250
rect -17480 81050 -17410 81250
rect -17090 81050 -17020 81250
rect -16980 81050 -16910 81250
rect -16590 81050 -16520 81250
rect -16480 81050 -16410 81250
rect -16090 81050 -16020 81250
rect -15980 81050 -15910 81250
rect -15590 81050 -15520 81250
rect -15480 81050 -15410 81250
rect -15090 81050 -15020 81250
rect -14980 81050 -14910 81250
rect -14590 81050 -14520 81250
rect -14480 81050 -14410 81250
rect -14090 81050 -14020 81250
rect -13980 81050 -13910 81250
rect -13590 81050 -13520 81250
rect -13480 81050 -13410 81250
rect -13090 81050 -13020 81250
rect -12980 81050 -12910 81250
rect -12590 81050 -12520 81250
rect -12480 81050 -12410 81250
rect -12090 81050 -12020 81250
rect -11980 81050 -11910 81250
rect -11590 81050 -11520 81250
rect -11480 81050 -11410 81250
rect -11090 81050 -11020 81250
rect -10980 81050 -10910 81250
rect -10590 81050 -10520 81250
rect -10480 81050 -10410 81250
rect -10090 81050 -10020 81250
rect -9980 81050 -9910 81250
rect -9590 81050 -9520 81250
rect -9480 81050 -9410 81250
rect -9090 81050 -9020 81250
rect -8980 81050 -8910 81250
rect -8590 81050 -8520 81250
rect -8480 81050 -8410 81250
rect -8090 81050 -8020 81250
rect -7980 81050 -7910 81250
rect -7590 81050 -7520 81250
rect -7480 81050 -7410 81250
rect -7090 81050 -7020 81250
rect -6980 81050 -6910 81250
rect -6590 81050 -6520 81250
rect -6480 81050 -6410 81250
rect -6090 81050 -6020 81250
rect -5980 81050 -5910 81250
rect -5590 81050 -5520 81250
rect -5480 81050 -5410 81250
rect -5090 81050 -5020 81250
rect -4980 81050 -4910 81250
rect -4590 81050 -4520 81250
rect -4480 81050 -4410 81250
rect -4090 81050 -4020 81250
rect -3980 81050 -3910 81250
rect -3590 81050 -3520 81250
rect -3480 81050 -3410 81250
rect -3090 81050 -3020 81250
rect -2980 81050 -2910 81250
rect -2590 81050 -2520 81250
rect -2480 81050 -2410 81250
rect -2090 81050 -2020 81250
rect -1980 81050 -1910 81250
rect -1590 81050 -1520 81250
rect -1480 81050 -1410 81250
rect -1090 81050 -1020 81250
rect -980 81050 -910 81250
rect -590 81050 -520 81250
rect -480 81050 -410 81250
rect -90 81050 -20 81250
rect 20 81050 90 81250
rect 410 81050 480 81250
rect 520 81050 590 81250
rect 910 81050 980 81250
rect 1020 81050 1090 81250
rect 1410 81050 1480 81250
rect 1520 81050 1590 81250
rect 1910 81050 1980 81250
rect 2020 81050 2090 81250
rect 2410 81050 2480 81250
rect 2520 81050 2590 81250
rect 2910 81050 2980 81250
rect 3020 81050 3090 81250
rect 3410 81050 3480 81250
rect 3520 81050 3590 81250
rect 3910 81050 3980 81250
rect 4020 81050 4090 81250
rect 4410 81050 4480 81250
rect 4520 81050 4590 81250
rect 4910 81050 4980 81250
rect 5020 81050 5090 81250
rect 5410 81050 5480 81250
rect 5520 81050 5590 81250
rect 5910 81050 5980 81250
rect 6020 81050 6090 81250
rect 6410 81050 6480 81250
rect 6520 81050 6590 81250
rect 6910 81050 6980 81250
rect 7020 81050 7090 81250
rect 7410 81050 7480 81250
rect 7520 81050 7590 81250
rect 7910 81050 7980 81250
rect 8020 81050 8090 81250
rect 8410 81050 8480 81250
rect 8520 81050 8590 81250
rect 8910 81050 8980 81250
rect 9020 81050 9090 81250
rect 9410 81050 9480 81250
rect 9520 81050 9590 81250
rect 9910 81050 9980 81250
rect 10020 81050 10090 81250
rect 10410 81050 10480 81250
rect 10520 81050 10590 81250
rect 10910 81050 10980 81250
rect 11020 81050 11090 81250
rect 11410 81050 11480 81250
rect 11520 81050 11590 81250
rect 11910 81050 11980 81250
rect 12020 81050 12090 81250
rect 12410 81050 12480 81250
rect 12520 81050 12590 81250
rect 12910 81050 12980 81250
rect 13020 81050 13090 81250
rect 13410 81050 13480 81250
rect 13520 81050 13590 81250
rect 13910 81050 13980 81250
rect 14020 81050 14090 81250
rect 14410 81050 14480 81250
rect 14520 81050 14590 81250
rect 14910 81050 14980 81250
rect 15020 81050 15090 81250
rect 15410 81050 15480 81250
rect 15520 81050 15590 81250
rect 15910 81050 15980 81250
rect 16020 81050 16090 81250
rect 16410 81050 16480 81250
rect 16520 81050 16590 81250
rect 16910 81050 16980 81250
rect 17020 81050 17090 81250
rect 17410 81050 17480 81250
rect 17520 81050 17590 81250
rect 17910 81050 17980 81250
rect 18020 81050 18090 81250
rect 18410 81050 18480 81250
rect 18520 81050 18590 81250
rect 18910 81050 18980 81250
rect 19020 81050 19090 81250
rect 19410 81050 19480 81250
rect 19520 81050 19590 81250
rect 19910 81050 19980 81250
rect 20020 81050 20090 81250
rect 20410 81050 20480 81250
rect 20520 81050 20590 81250
rect 20910 81050 20980 81250
rect 21020 81050 21090 81250
rect 21410 81050 21480 81250
rect 21520 81050 21590 81250
rect 21910 81050 21980 81250
rect 22020 81050 22090 81250
rect 22410 81050 22480 81250
rect 22520 81050 22590 81250
rect 22910 81050 22980 81250
rect 23020 81050 23090 81250
rect 23410 81050 23480 81250
rect 23520 81050 23590 81250
rect 23910 81050 23980 81250
rect 24020 81050 24090 81250
rect 24410 81050 24480 81250
rect 24520 81050 24590 81250
rect 24910 81050 24980 81250
rect 25020 81050 25090 81250
rect 25410 81050 25480 81250
rect 25520 81050 25590 81250
rect 25910 81050 25980 81250
rect 26020 81050 26090 81250
rect 26410 81050 26480 81250
rect 26520 81050 26590 81250
rect 26910 81050 26980 81250
rect 27020 81050 27090 81250
rect 27410 81050 27480 81250
rect 27520 81050 27590 81250
rect 27910 81050 27980 81250
rect 28020 81050 28090 81250
rect 28410 81050 28480 81250
rect 28520 81050 28590 81250
rect 28910 81050 28980 81250
rect 29020 81050 29090 81250
rect 29410 81050 29480 81250
rect 29520 81050 29590 81250
rect 29910 81050 29980 81250
rect 30020 81050 30090 81250
rect 30410 81050 30480 81250
rect 30520 81050 30590 81250
rect 30910 81050 30980 81250
rect 31020 81050 31090 81250
rect 31410 81050 31480 81250
rect 31520 81050 31590 81250
rect 31910 81050 31980 81250
rect 32020 81050 32090 81250
rect 32410 81050 32480 81250
rect 32520 81050 32590 81250
rect 32910 81050 32980 81250
rect 33020 81050 33090 81250
rect 33410 81050 33480 81250
rect 33520 81050 33590 81250
rect 33910 81050 33980 81250
rect 34020 81050 34090 81250
rect 34410 81050 34480 81250
rect 34520 81050 34590 81250
rect 34910 81050 34980 81250
rect 35020 81050 35090 81250
rect 35410 81050 35480 81250
rect 35520 81050 35590 81250
rect 35910 81050 35980 81250
rect 36020 81050 36090 81250
rect 36410 81050 36480 81250
rect 36520 81050 36590 81250
rect 36910 81050 36980 81250
rect 37020 81050 37090 81250
rect 37410 81050 37480 81250
rect 37520 81050 37590 81250
rect 37910 81050 37980 81250
rect 38020 81050 38090 81250
rect 38410 81050 38480 81250
rect 38520 81050 38590 81250
rect 38910 81050 38980 81250
rect 39020 81050 39090 81250
rect 39410 81050 39480 81250
rect 39520 81050 39590 81250
rect 39910 81050 39980 81250
rect 40020 81050 40090 81250
rect 40410 81050 40480 81250
rect 40520 81050 40590 81250
rect 40910 81050 40980 81250
rect 41020 81050 41090 81250
rect 41410 81050 41480 81250
rect 41520 81050 41590 81250
rect 41910 81050 41980 81250
rect 42020 81050 42090 81250
rect 42410 81050 42480 81250
rect 42520 81050 42590 81250
rect 42910 81050 42980 81250
rect 43020 81050 43090 81250
rect 43410 81050 43480 81250
rect 43520 81050 43590 81250
rect 43910 81050 43980 81250
rect 44020 81050 44090 81250
rect 44410 81050 44480 81250
rect 44520 81050 44590 81250
rect 44910 81050 44980 81250
rect 45020 81050 45090 81250
rect 45410 81050 45480 81250
rect 45520 81050 45590 81250
rect 45910 81050 45980 81250
rect 46020 81050 46090 81250
rect 46410 81050 46480 81250
rect 46520 81050 46590 81250
rect 46910 81050 46980 81250
rect 47020 81050 47090 81250
rect 47410 81050 47480 81250
rect 47520 81050 47590 81250
rect 47910 81050 47980 81250
rect 48020 81050 48090 81250
rect 48410 81050 48480 81250
rect 48520 81050 48590 81250
rect 48910 81050 48980 81250
rect 49020 81050 49090 81250
rect 49410 81050 49480 81250
rect 49520 81050 49590 81250
rect 49910 81050 49980 81250
rect 50020 81050 50090 81250
rect 50410 81050 50480 81250
rect 50520 81050 50590 81250
rect 50910 81050 50980 81250
rect 51020 81050 51090 81250
rect 51410 81050 51480 81250
rect 51520 81050 51590 81250
rect 51910 81050 51980 81250
rect 52020 81050 52090 81250
rect 52410 81050 52480 81250
rect 52520 81050 52590 81250
rect 52910 81050 52980 81250
rect 53020 81050 53090 81250
rect 53410 81050 53480 81250
rect 53520 81050 53590 81250
rect 53910 81050 53980 81250
rect 54020 81050 54090 81250
rect 54410 81050 54480 81250
rect 54520 81050 54590 81250
rect 54910 81050 54980 81250
rect 55020 81050 55090 81250
rect 55410 81050 55480 81250
rect 55520 81050 55590 81250
rect 55910 81050 55980 81250
rect 56020 81050 56090 81250
rect 56410 81050 56480 81250
rect 56520 81050 56590 81250
rect 56910 81050 56980 81250
rect 57020 81050 57090 81250
rect 57410 81050 57480 81250
rect 57520 81050 57590 81250
rect 57910 81050 57980 81250
rect 58020 81050 58090 81250
rect 58410 81050 58480 81250
rect 58520 81050 58590 81250
rect 58910 81050 58980 81250
rect 59020 81050 59090 81250
rect 59410 81050 59480 81250
rect 59520 81050 59590 81250
rect 59910 81050 59980 81250
rect 60020 81050 60090 81250
rect 60410 81050 60480 81250
rect 60520 81050 60590 81250
rect 60910 81050 60980 81250
rect 61020 81050 61090 81250
rect 61410 81050 61480 81250
rect 61520 81050 61590 81250
rect 61910 81050 61980 81250
rect 62020 81050 62090 81250
rect 62410 81050 62480 81250
rect 62520 81050 62590 81250
rect 62910 81050 62980 81250
rect 63020 81050 63090 81250
rect 63410 81050 63480 81250
rect 63520 81050 63590 81250
rect 63910 81050 63980 81250
rect 64020 81050 64090 81250
rect 64410 81050 64480 81250
rect 64520 81050 64590 81250
rect 64910 81050 64980 81250
rect 65020 81050 65090 81250
rect 65410 81050 65480 81250
rect 65520 81050 65590 81250
rect 65910 81050 65980 81250
rect 66020 81050 66090 81250
rect 66410 81050 66480 81250
rect 66520 81050 66590 81250
rect 66910 81050 66980 81250
rect 67020 81050 67090 81250
rect 67410 81050 67480 81250
rect 67520 81050 67590 81250
rect 67910 81050 67980 81250
rect 68020 81050 68090 81250
rect 68410 81050 68480 81250
rect 68520 81050 68590 81250
rect 68910 81050 68980 81250
rect 69020 81050 69090 81250
rect 69410 81050 69480 81250
rect 69520 81050 69590 81250
rect 69910 81050 69980 81250
rect 70020 81050 70090 81250
rect 70410 81050 70480 81250
rect 70520 81050 70590 81250
rect 70910 81050 70980 81250
rect 71020 81050 71090 81250
rect 71410 81050 71480 81250
rect 71520 81050 71590 81250
rect 71910 81050 71980 81250
rect 72020 81050 72090 81250
rect 72410 81050 72480 81250
rect 72520 81050 72590 81250
rect 72910 81050 72980 81250
rect 73020 81050 73090 81250
rect 73410 81050 73480 81250
rect 73520 81050 73590 81250
rect 73910 81050 73980 81250
rect 74020 81050 74090 81250
rect 74410 81050 74480 81250
rect 74520 81050 74590 81250
rect 74910 81050 74980 81250
rect 75020 81050 75090 81250
rect 75410 81050 75480 81250
rect 75520 81050 75590 81250
rect 75910 81050 75980 81250
rect 76020 81050 76090 81250
rect 76410 81050 76480 81250
rect 76520 81050 76590 81250
rect 76910 81050 76980 81250
rect 77020 81050 77090 81250
rect 77410 81050 77480 81250
rect 77520 81050 77590 81250
rect 77910 81050 77980 81250
rect 78020 81050 78090 81250
rect 78410 81050 78480 81250
rect 78520 81050 78590 81250
rect 78910 81050 78980 81250
rect 79020 81050 79090 81250
rect 79410 81050 79480 81250
rect 79520 81050 79590 81250
rect 79910 81050 79980 81250
rect 80020 81050 80090 81250
rect 80410 81050 80480 81250
rect 80520 81050 80590 81250
rect 80910 81050 80980 81250
rect 81020 81050 81090 81250
rect 81410 81050 81480 81250
rect 81520 81050 81590 81250
rect 81910 81050 81980 81250
rect 82020 81050 82090 81250
rect 82410 81050 82480 81250
rect 82520 81050 82590 81250
rect 82910 81050 82980 81250
rect 83020 81050 83090 81250
rect 83410 81050 83480 81250
rect 83520 81050 83590 81250
rect 83910 81050 83980 81250
rect 84020 81050 84090 81250
rect 84410 81050 84480 81250
rect 84520 81050 84590 81250
rect 84910 81050 84980 81250
rect 85020 81050 85090 81250
rect 85410 81050 85480 81250
rect 85520 81050 85590 81250
rect 85910 81050 85980 81250
rect 86020 81050 86090 81250
rect 86410 81050 86480 81250
rect 86520 81050 86590 81250
rect 86910 81050 86980 81250
rect 87020 81050 87090 81250
rect 87410 81050 87480 81250
rect 87520 81050 87590 81250
rect 87910 81050 87980 81250
rect 88020 81050 88090 81250
rect 88410 81050 88480 81250
rect 88520 81050 88590 81250
rect 88910 81050 88980 81250
rect 89020 81050 89090 81250
rect 89410 81050 89480 81250
rect 89520 81050 89590 81250
rect 89910 81050 89980 81250
rect 90020 81050 90090 81250
rect 90410 81050 90480 81250
rect 90520 81050 90590 81250
rect 90910 81050 90980 81250
rect 91020 81050 91090 81250
rect 91410 81050 91480 81250
rect 91520 81050 91590 81250
rect 91910 81050 91980 81250
rect 92020 81050 92090 81250
rect 92410 81050 92480 81250
rect 92520 81050 92590 81250
rect 92910 81050 92980 81250
rect 93020 81050 93090 81250
rect 93410 81050 93480 81250
rect 93520 81050 93590 81250
rect 93910 81050 93980 81250
rect 94020 81050 94090 81250
rect 94410 81050 94480 81250
rect 94520 81050 94590 81250
rect 94910 81050 94980 81250
rect 95020 81050 95090 81250
rect 95410 81050 95480 81250
rect 95520 81050 95590 81250
rect 95910 81050 95980 81250
rect 96020 81050 96090 81250
rect 96410 81050 96480 81250
rect 96520 81050 96590 81250
rect 96910 81050 96980 81250
rect 97020 81050 97090 81250
rect 97410 81050 97480 81250
rect 97520 81050 97590 81250
rect 97910 81050 97980 81250
rect 98020 81050 98090 81250
rect 98410 81050 98480 81250
rect 98520 81050 98590 81250
rect 98910 81050 98980 81250
rect 99020 81050 99090 81250
rect 99410 81050 99480 81250
rect 99520 81050 99590 81250
rect 99910 81050 99980 81250
rect 100020 81050 100090 81250
rect 100410 81050 100480 81250
rect -83350 80920 -83150 80990
rect -82850 80920 -82650 80990
rect -82350 80920 -82150 80990
rect -81850 80920 -81650 80990
rect -81350 80920 -81150 80990
rect -80850 80920 -80650 80990
rect -80350 80920 -80150 80990
rect -79850 80920 -79650 80990
rect -79350 80920 -79150 80990
rect -78850 80920 -78650 80990
rect -78350 80920 -78150 80990
rect -77850 80920 -77650 80990
rect -77350 80920 -77150 80990
rect -76850 80920 -76650 80990
rect -76350 80920 -76150 80990
rect -75850 80920 -75650 80990
rect -75350 80920 -75150 80990
rect -74850 80920 -74650 80990
rect -74350 80920 -74150 80990
rect -73850 80920 -73650 80990
rect -73350 80920 -73150 80990
rect -72850 80920 -72650 80990
rect -72350 80920 -72150 80990
rect -71850 80920 -71650 80990
rect -71350 80920 -71150 80990
rect -70850 80920 -70650 80990
rect -70350 80920 -70150 80990
rect -69850 80920 -69650 80990
rect -69350 80920 -69150 80990
rect -68850 80920 -68650 80990
rect -68350 80920 -68150 80990
rect -67850 80920 -67650 80990
rect -67350 80920 -67150 80990
rect -66850 80920 -66650 80990
rect -66350 80920 -66150 80990
rect -65850 80920 -65650 80990
rect -65350 80920 -65150 80990
rect -64850 80920 -64650 80990
rect -64350 80920 -64150 80990
rect -63850 80920 -63650 80990
rect -63350 80920 -63150 80990
rect -62850 80920 -62650 80990
rect -62350 80920 -62150 80990
rect -61850 80920 -61650 80990
rect -61350 80920 -61150 80990
rect -60850 80920 -60650 80990
rect -60350 80920 -60150 80990
rect -59850 80920 -59650 80990
rect -59350 80920 -59150 80990
rect -58850 80920 -58650 80990
rect -58350 80920 -58150 80990
rect -57850 80920 -57650 80990
rect -57350 80920 -57150 80990
rect -56850 80920 -56650 80990
rect -56350 80920 -56150 80990
rect -55850 80920 -55650 80990
rect -55350 80920 -55150 80990
rect -54850 80920 -54650 80990
rect -54350 80920 -54150 80990
rect -53850 80920 -53650 80990
rect -53350 80920 -53150 80990
rect -52850 80920 -52650 80990
rect -52350 80920 -52150 80990
rect -51850 80920 -51650 80990
rect -51350 80920 -51150 80990
rect -50850 80920 -50650 80990
rect -50350 80920 -50150 80990
rect -49850 80920 -49650 80990
rect -49350 80920 -49150 80990
rect -48850 80920 -48650 80990
rect -48350 80920 -48150 80990
rect -47850 80920 -47650 80990
rect -47350 80920 -47150 80990
rect -46850 80920 -46650 80990
rect -46350 80920 -46150 80990
rect -45850 80920 -45650 80990
rect -45350 80920 -45150 80990
rect -44850 80920 -44650 80990
rect -44350 80920 -44150 80990
rect -43850 80920 -43650 80990
rect -43350 80920 -43150 80990
rect -42850 80920 -42650 80990
rect -42350 80920 -42150 80990
rect -41850 80920 -41650 80990
rect -41350 80920 -41150 80990
rect -40850 80920 -40650 80990
rect -40350 80920 -40150 80990
rect -39850 80920 -39650 80990
rect -39350 80920 -39150 80990
rect -38850 80920 -38650 80990
rect -38350 80920 -38150 80990
rect -37850 80920 -37650 80990
rect -37350 80920 -37150 80990
rect -36850 80920 -36650 80990
rect -36350 80920 -36150 80990
rect -35850 80920 -35650 80990
rect -35350 80920 -35150 80990
rect -34850 80920 -34650 80990
rect -34350 80920 -34150 80990
rect -33850 80920 -33650 80990
rect -33350 80920 -33150 80990
rect -32850 80920 -32650 80990
rect -32350 80920 -32150 80990
rect -31850 80920 -31650 80990
rect -31350 80920 -31150 80990
rect -30850 80920 -30650 80990
rect -30350 80920 -30150 80990
rect -29850 80920 -29650 80990
rect -29350 80920 -29150 80990
rect -28850 80920 -28650 80990
rect -28350 80920 -28150 80990
rect -27850 80920 -27650 80990
rect -27350 80920 -27150 80990
rect -26850 80920 -26650 80990
rect -26350 80920 -26150 80990
rect -25850 80920 -25650 80990
rect -25350 80920 -25150 80990
rect -24850 80920 -24650 80990
rect -24350 80920 -24150 80990
rect -23850 80920 -23650 80990
rect -23350 80920 -23150 80990
rect -22850 80920 -22650 80990
rect -22350 80920 -22150 80990
rect -21850 80920 -21650 80990
rect -21350 80920 -21150 80990
rect -20850 80920 -20650 80990
rect -20350 80920 -20150 80990
rect -19850 80920 -19650 80990
rect -19350 80920 -19150 80990
rect -18850 80920 -18650 80990
rect -18350 80920 -18150 80990
rect -17850 80920 -17650 80990
rect -17350 80920 -17150 80990
rect -16850 80920 -16650 80990
rect -16350 80920 -16150 80990
rect -15850 80920 -15650 80990
rect -15350 80920 -15150 80990
rect -14850 80920 -14650 80990
rect -14350 80920 -14150 80990
rect -13850 80920 -13650 80990
rect -13350 80920 -13150 80990
rect -12850 80920 -12650 80990
rect -12350 80920 -12150 80990
rect -11850 80920 -11650 80990
rect -11350 80920 -11150 80990
rect -10850 80920 -10650 80990
rect -10350 80920 -10150 80990
rect -9850 80920 -9650 80990
rect -9350 80920 -9150 80990
rect -8850 80920 -8650 80990
rect -8350 80920 -8150 80990
rect -7850 80920 -7650 80990
rect -7350 80920 -7150 80990
rect -6850 80920 -6650 80990
rect -6350 80920 -6150 80990
rect -5850 80920 -5650 80990
rect -5350 80920 -5150 80990
rect -4850 80920 -4650 80990
rect -4350 80920 -4150 80990
rect -3850 80920 -3650 80990
rect -3350 80920 -3150 80990
rect -2850 80920 -2650 80990
rect -2350 80920 -2150 80990
rect -1850 80920 -1650 80990
rect -1350 80920 -1150 80990
rect -850 80920 -650 80990
rect -350 80920 -150 80990
rect 150 80920 350 80990
rect 650 80920 850 80990
rect 1150 80920 1350 80990
rect 1650 80920 1850 80990
rect 2150 80920 2350 80990
rect 2650 80920 2850 80990
rect 3150 80920 3350 80990
rect 3650 80920 3850 80990
rect 4150 80920 4350 80990
rect 4650 80920 4850 80990
rect 5150 80920 5350 80990
rect 5650 80920 5850 80990
rect 6150 80920 6350 80990
rect 6650 80920 6850 80990
rect 7150 80920 7350 80990
rect 7650 80920 7850 80990
rect 8150 80920 8350 80990
rect 8650 80920 8850 80990
rect 9150 80920 9350 80990
rect 9650 80920 9850 80990
rect 10150 80920 10350 80990
rect 10650 80920 10850 80990
rect 11150 80920 11350 80990
rect 11650 80920 11850 80990
rect 12150 80920 12350 80990
rect 12650 80920 12850 80990
rect 13150 80920 13350 80990
rect 13650 80920 13850 80990
rect 14150 80920 14350 80990
rect 14650 80920 14850 80990
rect 15150 80920 15350 80990
rect 15650 80920 15850 80990
rect 16150 80920 16350 80990
rect 16650 80920 16850 80990
rect 17150 80920 17350 80990
rect 17650 80920 17850 80990
rect 18150 80920 18350 80990
rect 18650 80920 18850 80990
rect 19150 80920 19350 80990
rect 19650 80920 19850 80990
rect 20150 80920 20350 80990
rect 20650 80920 20850 80990
rect 21150 80920 21350 80990
rect 21650 80920 21850 80990
rect 22150 80920 22350 80990
rect 22650 80920 22850 80990
rect 23150 80920 23350 80990
rect 23650 80920 23850 80990
rect 24150 80920 24350 80990
rect 24650 80920 24850 80990
rect 25150 80920 25350 80990
rect 25650 80920 25850 80990
rect 26150 80920 26350 80990
rect 26650 80920 26850 80990
rect 27150 80920 27350 80990
rect 27650 80920 27850 80990
rect 28150 80920 28350 80990
rect 28650 80920 28850 80990
rect 29150 80920 29350 80990
rect 29650 80920 29850 80990
rect 30150 80920 30350 80990
rect 30650 80920 30850 80990
rect 31150 80920 31350 80990
rect 31650 80920 31850 80990
rect 32150 80920 32350 80990
rect 32650 80920 32850 80990
rect 33150 80920 33350 80990
rect 33650 80920 33850 80990
rect 34150 80920 34350 80990
rect 34650 80920 34850 80990
rect 35150 80920 35350 80990
rect 35650 80920 35850 80990
rect 36150 80920 36350 80990
rect 36650 80920 36850 80990
rect 37150 80920 37350 80990
rect 37650 80920 37850 80990
rect 38150 80920 38350 80990
rect 38650 80920 38850 80990
rect 39150 80920 39350 80990
rect 39650 80920 39850 80990
rect 40150 80920 40350 80990
rect 40650 80920 40850 80990
rect 41150 80920 41350 80990
rect 41650 80920 41850 80990
rect 42150 80920 42350 80990
rect 42650 80920 42850 80990
rect 43150 80920 43350 80990
rect 43650 80920 43850 80990
rect 44150 80920 44350 80990
rect 44650 80920 44850 80990
rect 45150 80920 45350 80990
rect 45650 80920 45850 80990
rect 46150 80920 46350 80990
rect 46650 80920 46850 80990
rect 47150 80920 47350 80990
rect 47650 80920 47850 80990
rect 48150 80920 48350 80990
rect 48650 80920 48850 80990
rect 49150 80920 49350 80990
rect 49650 80920 49850 80990
rect 50150 80920 50350 80990
rect 50650 80920 50850 80990
rect 51150 80920 51350 80990
rect 51650 80920 51850 80990
rect 52150 80920 52350 80990
rect 52650 80920 52850 80990
rect 53150 80920 53350 80990
rect 53650 80920 53850 80990
rect 54150 80920 54350 80990
rect 54650 80920 54850 80990
rect 55150 80920 55350 80990
rect 55650 80920 55850 80990
rect 56150 80920 56350 80990
rect 56650 80920 56850 80990
rect 57150 80920 57350 80990
rect 57650 80920 57850 80990
rect 58150 80920 58350 80990
rect 58650 80920 58850 80990
rect 59150 80920 59350 80990
rect 59650 80920 59850 80990
rect 60150 80920 60350 80990
rect 60650 80920 60850 80990
rect 61150 80920 61350 80990
rect 61650 80920 61850 80990
rect 62150 80920 62350 80990
rect 62650 80920 62850 80990
rect 63150 80920 63350 80990
rect 63650 80920 63850 80990
rect 64150 80920 64350 80990
rect 64650 80920 64850 80990
rect 65150 80920 65350 80990
rect 65650 80920 65850 80990
rect 66150 80920 66350 80990
rect 66650 80920 66850 80990
rect 67150 80920 67350 80990
rect 67650 80920 67850 80990
rect 68150 80920 68350 80990
rect 68650 80920 68850 80990
rect 69150 80920 69350 80990
rect 69650 80920 69850 80990
rect 70150 80920 70350 80990
rect 70650 80920 70850 80990
rect 71150 80920 71350 80990
rect 71650 80920 71850 80990
rect 72150 80920 72350 80990
rect 72650 80920 72850 80990
rect 73150 80920 73350 80990
rect 73650 80920 73850 80990
rect 74150 80920 74350 80990
rect 74650 80920 74850 80990
rect 75150 80920 75350 80990
rect 75650 80920 75850 80990
rect 76150 80920 76350 80990
rect 76650 80920 76850 80990
rect 77150 80920 77350 80990
rect 77650 80920 77850 80990
rect 78150 80920 78350 80990
rect 78650 80920 78850 80990
rect 79150 80920 79350 80990
rect 79650 80920 79850 80990
rect 80150 80920 80350 80990
rect 80650 80920 80850 80990
rect 81150 80920 81350 80990
rect 81650 80920 81850 80990
rect 82150 80920 82350 80990
rect 82650 80920 82850 80990
rect 83150 80920 83350 80990
rect 83650 80920 83850 80990
rect 84150 80920 84350 80990
rect 84650 80920 84850 80990
rect 85150 80920 85350 80990
rect 85650 80920 85850 80990
rect 86150 80920 86350 80990
rect 86650 80920 86850 80990
rect 87150 80920 87350 80990
rect 87650 80920 87850 80990
rect 88150 80920 88350 80990
rect 88650 80920 88850 80990
rect 89150 80920 89350 80990
rect 89650 80920 89850 80990
rect 90150 80920 90350 80990
rect 90650 80920 90850 80990
rect 91150 80920 91350 80990
rect 91650 80920 91850 80990
rect 92150 80920 92350 80990
rect 92650 80920 92850 80990
rect 93150 80920 93350 80990
rect 93650 80920 93850 80990
rect 94150 80920 94350 80990
rect 94650 80920 94850 80990
rect 95150 80920 95350 80990
rect 95650 80920 95850 80990
rect 96150 80920 96350 80990
rect 96650 80920 96850 80990
rect 97150 80920 97350 80990
rect 97650 80920 97850 80990
rect 98150 80920 98350 80990
rect 98650 80920 98850 80990
rect 99150 80920 99350 80990
rect 99650 80920 99850 80990
rect 100150 80920 100350 80990
rect -83350 80810 -83150 80880
rect -82850 80810 -82650 80880
rect -82350 80810 -82150 80880
rect -81850 80810 -81650 80880
rect -81350 80810 -81150 80880
rect -80850 80810 -80650 80880
rect -80350 80810 -80150 80880
rect -79850 80810 -79650 80880
rect -79350 80810 -79150 80880
rect -78850 80810 -78650 80880
rect -78350 80810 -78150 80880
rect -77850 80810 -77650 80880
rect -77350 80810 -77150 80880
rect -76850 80810 -76650 80880
rect -76350 80810 -76150 80880
rect -75850 80810 -75650 80880
rect -75350 80810 -75150 80880
rect -74850 80810 -74650 80880
rect -74350 80810 -74150 80880
rect -73850 80810 -73650 80880
rect -73350 80810 -73150 80880
rect -72850 80810 -72650 80880
rect -72350 80810 -72150 80880
rect -71850 80810 -71650 80880
rect -71350 80810 -71150 80880
rect -70850 80810 -70650 80880
rect -70350 80810 -70150 80880
rect -69850 80810 -69650 80880
rect -69350 80810 -69150 80880
rect -68850 80810 -68650 80880
rect -68350 80810 -68150 80880
rect -67850 80810 -67650 80880
rect -67350 80810 -67150 80880
rect -66850 80810 -66650 80880
rect -66350 80810 -66150 80880
rect -65850 80810 -65650 80880
rect -65350 80810 -65150 80880
rect -64850 80810 -64650 80880
rect -64350 80810 -64150 80880
rect -63850 80810 -63650 80880
rect -63350 80810 -63150 80880
rect -62850 80810 -62650 80880
rect -62350 80810 -62150 80880
rect -61850 80810 -61650 80880
rect -61350 80810 -61150 80880
rect -60850 80810 -60650 80880
rect -60350 80810 -60150 80880
rect -59850 80810 -59650 80880
rect -59350 80810 -59150 80880
rect -58850 80810 -58650 80880
rect -58350 80810 -58150 80880
rect -57850 80810 -57650 80880
rect -57350 80810 -57150 80880
rect -56850 80810 -56650 80880
rect -56350 80810 -56150 80880
rect -55850 80810 -55650 80880
rect -55350 80810 -55150 80880
rect -54850 80810 -54650 80880
rect -54350 80810 -54150 80880
rect -53850 80810 -53650 80880
rect -53350 80810 -53150 80880
rect -52850 80810 -52650 80880
rect -52350 80810 -52150 80880
rect -51850 80810 -51650 80880
rect -51350 80810 -51150 80880
rect -50850 80810 -50650 80880
rect -50350 80810 -50150 80880
rect -49850 80810 -49650 80880
rect -49350 80810 -49150 80880
rect -48850 80810 -48650 80880
rect -48350 80810 -48150 80880
rect -47850 80810 -47650 80880
rect -47350 80810 -47150 80880
rect -46850 80810 -46650 80880
rect -46350 80810 -46150 80880
rect -45850 80810 -45650 80880
rect -45350 80810 -45150 80880
rect -44850 80810 -44650 80880
rect -44350 80810 -44150 80880
rect -43850 80810 -43650 80880
rect -43350 80810 -43150 80880
rect -42850 80810 -42650 80880
rect -42350 80810 -42150 80880
rect -41850 80810 -41650 80880
rect -41350 80810 -41150 80880
rect -40850 80810 -40650 80880
rect -40350 80810 -40150 80880
rect -39850 80810 -39650 80880
rect -39350 80810 -39150 80880
rect -38850 80810 -38650 80880
rect -38350 80810 -38150 80880
rect -37850 80810 -37650 80880
rect -37350 80810 -37150 80880
rect -36850 80810 -36650 80880
rect -36350 80810 -36150 80880
rect -35850 80810 -35650 80880
rect -35350 80810 -35150 80880
rect -34850 80810 -34650 80880
rect -34350 80810 -34150 80880
rect -33850 80810 -33650 80880
rect -33350 80810 -33150 80880
rect -32850 80810 -32650 80880
rect -32350 80810 -32150 80880
rect -31850 80810 -31650 80880
rect -31350 80810 -31150 80880
rect -30850 80810 -30650 80880
rect -30350 80810 -30150 80880
rect -29850 80810 -29650 80880
rect -29350 80810 -29150 80880
rect -28850 80810 -28650 80880
rect -28350 80810 -28150 80880
rect -27850 80810 -27650 80880
rect -27350 80810 -27150 80880
rect -26850 80810 -26650 80880
rect -26350 80810 -26150 80880
rect -25850 80810 -25650 80880
rect -25350 80810 -25150 80880
rect -24850 80810 -24650 80880
rect -24350 80810 -24150 80880
rect -23850 80810 -23650 80880
rect -23350 80810 -23150 80880
rect -22850 80810 -22650 80880
rect -22350 80810 -22150 80880
rect -21850 80810 -21650 80880
rect -21350 80810 -21150 80880
rect -20850 80810 -20650 80880
rect -20350 80810 -20150 80880
rect -19850 80810 -19650 80880
rect -19350 80810 -19150 80880
rect -18850 80810 -18650 80880
rect -18350 80810 -18150 80880
rect -17850 80810 -17650 80880
rect -17350 80810 -17150 80880
rect -16850 80810 -16650 80880
rect -16350 80810 -16150 80880
rect -15850 80810 -15650 80880
rect -15350 80810 -15150 80880
rect -14850 80810 -14650 80880
rect -14350 80810 -14150 80880
rect -13850 80810 -13650 80880
rect -13350 80810 -13150 80880
rect -12850 80810 -12650 80880
rect -12350 80810 -12150 80880
rect -11850 80810 -11650 80880
rect -11350 80810 -11150 80880
rect -10850 80810 -10650 80880
rect -10350 80810 -10150 80880
rect -9850 80810 -9650 80880
rect -9350 80810 -9150 80880
rect -8850 80810 -8650 80880
rect -8350 80810 -8150 80880
rect -7850 80810 -7650 80880
rect -7350 80810 -7150 80880
rect -6850 80810 -6650 80880
rect -6350 80810 -6150 80880
rect -5850 80810 -5650 80880
rect -5350 80810 -5150 80880
rect -4850 80810 -4650 80880
rect -4350 80810 -4150 80880
rect -3850 80810 -3650 80880
rect -3350 80810 -3150 80880
rect -2850 80810 -2650 80880
rect -2350 80810 -2150 80880
rect -1850 80810 -1650 80880
rect -1350 80810 -1150 80880
rect -850 80810 -650 80880
rect -350 80810 -150 80880
rect 150 80810 350 80880
rect 650 80810 850 80880
rect 1150 80810 1350 80880
rect 1650 80810 1850 80880
rect 2150 80810 2350 80880
rect 2650 80810 2850 80880
rect 3150 80810 3350 80880
rect 3650 80810 3850 80880
rect 4150 80810 4350 80880
rect 4650 80810 4850 80880
rect 5150 80810 5350 80880
rect 5650 80810 5850 80880
rect 6150 80810 6350 80880
rect 6650 80810 6850 80880
rect 7150 80810 7350 80880
rect 7650 80810 7850 80880
rect 8150 80810 8350 80880
rect 8650 80810 8850 80880
rect 9150 80810 9350 80880
rect 9650 80810 9850 80880
rect 10150 80810 10350 80880
rect 10650 80810 10850 80880
rect 11150 80810 11350 80880
rect 11650 80810 11850 80880
rect 12150 80810 12350 80880
rect 12650 80810 12850 80880
rect 13150 80810 13350 80880
rect 13650 80810 13850 80880
rect 14150 80810 14350 80880
rect 14650 80810 14850 80880
rect 15150 80810 15350 80880
rect 15650 80810 15850 80880
rect 16150 80810 16350 80880
rect 16650 80810 16850 80880
rect 17150 80810 17350 80880
rect 17650 80810 17850 80880
rect 18150 80810 18350 80880
rect 18650 80810 18850 80880
rect 19150 80810 19350 80880
rect 19650 80810 19850 80880
rect 20150 80810 20350 80880
rect 20650 80810 20850 80880
rect 21150 80810 21350 80880
rect 21650 80810 21850 80880
rect 22150 80810 22350 80880
rect 22650 80810 22850 80880
rect 23150 80810 23350 80880
rect 23650 80810 23850 80880
rect 24150 80810 24350 80880
rect 24650 80810 24850 80880
rect 25150 80810 25350 80880
rect 25650 80810 25850 80880
rect 26150 80810 26350 80880
rect 26650 80810 26850 80880
rect 27150 80810 27350 80880
rect 27650 80810 27850 80880
rect 28150 80810 28350 80880
rect 28650 80810 28850 80880
rect 29150 80810 29350 80880
rect 29650 80810 29850 80880
rect 30150 80810 30350 80880
rect 30650 80810 30850 80880
rect 31150 80810 31350 80880
rect 31650 80810 31850 80880
rect 32150 80810 32350 80880
rect 32650 80810 32850 80880
rect 33150 80810 33350 80880
rect 33650 80810 33850 80880
rect 34150 80810 34350 80880
rect 34650 80810 34850 80880
rect 35150 80810 35350 80880
rect 35650 80810 35850 80880
rect 36150 80810 36350 80880
rect 36650 80810 36850 80880
rect 37150 80810 37350 80880
rect 37650 80810 37850 80880
rect 38150 80810 38350 80880
rect 38650 80810 38850 80880
rect 39150 80810 39350 80880
rect 39650 80810 39850 80880
rect 40150 80810 40350 80880
rect 40650 80810 40850 80880
rect 41150 80810 41350 80880
rect 41650 80810 41850 80880
rect 42150 80810 42350 80880
rect 42650 80810 42850 80880
rect 43150 80810 43350 80880
rect 43650 80810 43850 80880
rect 44150 80810 44350 80880
rect 44650 80810 44850 80880
rect 45150 80810 45350 80880
rect 45650 80810 45850 80880
rect 46150 80810 46350 80880
rect 46650 80810 46850 80880
rect 47150 80810 47350 80880
rect 47650 80810 47850 80880
rect 48150 80810 48350 80880
rect 48650 80810 48850 80880
rect 49150 80810 49350 80880
rect 49650 80810 49850 80880
rect 50150 80810 50350 80880
rect 50650 80810 50850 80880
rect 51150 80810 51350 80880
rect 51650 80810 51850 80880
rect 52150 80810 52350 80880
rect 52650 80810 52850 80880
rect 53150 80810 53350 80880
rect 53650 80810 53850 80880
rect 54150 80810 54350 80880
rect 54650 80810 54850 80880
rect 55150 80810 55350 80880
rect 55650 80810 55850 80880
rect 56150 80810 56350 80880
rect 56650 80810 56850 80880
rect 57150 80810 57350 80880
rect 57650 80810 57850 80880
rect 58150 80810 58350 80880
rect 58650 80810 58850 80880
rect 59150 80810 59350 80880
rect 59650 80810 59850 80880
rect 60150 80810 60350 80880
rect 60650 80810 60850 80880
rect 61150 80810 61350 80880
rect 61650 80810 61850 80880
rect 62150 80810 62350 80880
rect 62650 80810 62850 80880
rect 63150 80810 63350 80880
rect 63650 80810 63850 80880
rect 64150 80810 64350 80880
rect 64650 80810 64850 80880
rect 65150 80810 65350 80880
rect 65650 80810 65850 80880
rect 66150 80810 66350 80880
rect 66650 80810 66850 80880
rect 67150 80810 67350 80880
rect 67650 80810 67850 80880
rect 68150 80810 68350 80880
rect 68650 80810 68850 80880
rect 69150 80810 69350 80880
rect 69650 80810 69850 80880
rect 70150 80810 70350 80880
rect 70650 80810 70850 80880
rect 71150 80810 71350 80880
rect 71650 80810 71850 80880
rect 72150 80810 72350 80880
rect 72650 80810 72850 80880
rect 73150 80810 73350 80880
rect 73650 80810 73850 80880
rect 74150 80810 74350 80880
rect 74650 80810 74850 80880
rect 75150 80810 75350 80880
rect 75650 80810 75850 80880
rect 76150 80810 76350 80880
rect 76650 80810 76850 80880
rect 77150 80810 77350 80880
rect 77650 80810 77850 80880
rect 78150 80810 78350 80880
rect 78650 80810 78850 80880
rect 79150 80810 79350 80880
rect 79650 80810 79850 80880
rect 80150 80810 80350 80880
rect 80650 80810 80850 80880
rect 81150 80810 81350 80880
rect 81650 80810 81850 80880
rect 82150 80810 82350 80880
rect 82650 80810 82850 80880
rect 83150 80810 83350 80880
rect 83650 80810 83850 80880
rect 84150 80810 84350 80880
rect 84650 80810 84850 80880
rect 85150 80810 85350 80880
rect 85650 80810 85850 80880
rect 86150 80810 86350 80880
rect 86650 80810 86850 80880
rect 87150 80810 87350 80880
rect 87650 80810 87850 80880
rect 88150 80810 88350 80880
rect 88650 80810 88850 80880
rect 89150 80810 89350 80880
rect 89650 80810 89850 80880
rect 90150 80810 90350 80880
rect 90650 80810 90850 80880
rect 91150 80810 91350 80880
rect 91650 80810 91850 80880
rect 92150 80810 92350 80880
rect 92650 80810 92850 80880
rect 93150 80810 93350 80880
rect 93650 80810 93850 80880
rect 94150 80810 94350 80880
rect 94650 80810 94850 80880
rect 95150 80810 95350 80880
rect 95650 80810 95850 80880
rect 96150 80810 96350 80880
rect 96650 80810 96850 80880
rect 97150 80810 97350 80880
rect 97650 80810 97850 80880
rect 98150 80810 98350 80880
rect 98650 80810 98850 80880
rect 99150 80810 99350 80880
rect 99650 80810 99850 80880
rect 100150 80810 100350 80880
rect -83480 80550 -83410 80750
rect -83090 80550 -83020 80750
rect -82980 80550 -82910 80750
rect -82590 80550 -82520 80750
rect -82480 80550 -82410 80750
rect -82090 80550 -82020 80750
rect -81980 80550 -81910 80750
rect -81590 80550 -81520 80750
rect -81480 80550 -81410 80750
rect -81090 80550 -81020 80750
rect -80980 80550 -80910 80750
rect -80590 80550 -80520 80750
rect -80480 80550 -80410 80750
rect -80090 80550 -80020 80750
rect -79980 80550 -79910 80750
rect -79590 80550 -79520 80750
rect -79480 80550 -79410 80750
rect -79090 80550 -79020 80750
rect -78980 80550 -78910 80750
rect -78590 80550 -78520 80750
rect -78480 80550 -78410 80750
rect -78090 80550 -78020 80750
rect -77980 80550 -77910 80750
rect -77590 80550 -77520 80750
rect -77480 80550 -77410 80750
rect -77090 80550 -77020 80750
rect -76980 80550 -76910 80750
rect -76590 80550 -76520 80750
rect -76480 80550 -76410 80750
rect -76090 80550 -76020 80750
rect -75980 80550 -75910 80750
rect -75590 80550 -75520 80750
rect -75480 80550 -75410 80750
rect -75090 80550 -75020 80750
rect -74980 80550 -74910 80750
rect -74590 80550 -74520 80750
rect -74480 80550 -74410 80750
rect -74090 80550 -74020 80750
rect -73980 80550 -73910 80750
rect -73590 80550 -73520 80750
rect -73480 80550 -73410 80750
rect -73090 80550 -73020 80750
rect -72980 80550 -72910 80750
rect -72590 80550 -72520 80750
rect -72480 80550 -72410 80750
rect -72090 80550 -72020 80750
rect -71980 80550 -71910 80750
rect -71590 80550 -71520 80750
rect -71480 80550 -71410 80750
rect -71090 80550 -71020 80750
rect -70980 80550 -70910 80750
rect -70590 80550 -70520 80750
rect -70480 80550 -70410 80750
rect -70090 80550 -70020 80750
rect -69980 80550 -69910 80750
rect -69590 80550 -69520 80750
rect -69480 80550 -69410 80750
rect -69090 80550 -69020 80750
rect -68980 80550 -68910 80750
rect -68590 80550 -68520 80750
rect -68480 80550 -68410 80750
rect -68090 80550 -68020 80750
rect -67980 80550 -67910 80750
rect -67590 80550 -67520 80750
rect -67480 80550 -67410 80750
rect -67090 80550 -67020 80750
rect -66980 80550 -66910 80750
rect -66590 80550 -66520 80750
rect -66480 80550 -66410 80750
rect -66090 80550 -66020 80750
rect -65980 80550 -65910 80750
rect -65590 80550 -65520 80750
rect -65480 80550 -65410 80750
rect -65090 80550 -65020 80750
rect -64980 80550 -64910 80750
rect -64590 80550 -64520 80750
rect -64480 80550 -64410 80750
rect -64090 80550 -64020 80750
rect -63980 80550 -63910 80750
rect -63590 80550 -63520 80750
rect -63480 80550 -63410 80750
rect -63090 80550 -63020 80750
rect -62980 80550 -62910 80750
rect -62590 80550 -62520 80750
rect -62480 80550 -62410 80750
rect -62090 80550 -62020 80750
rect -61980 80550 -61910 80750
rect -61590 80550 -61520 80750
rect -61480 80550 -61410 80750
rect -61090 80550 -61020 80750
rect -60980 80550 -60910 80750
rect -60590 80550 -60520 80750
rect -60480 80550 -60410 80750
rect -60090 80550 -60020 80750
rect -59980 80550 -59910 80750
rect -59590 80550 -59520 80750
rect -59480 80550 -59410 80750
rect -59090 80550 -59020 80750
rect -58980 80550 -58910 80750
rect -58590 80550 -58520 80750
rect -58480 80550 -58410 80750
rect -58090 80550 -58020 80750
rect -57980 80550 -57910 80750
rect -57590 80550 -57520 80750
rect -57480 80550 -57410 80750
rect -57090 80550 -57020 80750
rect -56980 80550 -56910 80750
rect -56590 80550 -56520 80750
rect -56480 80550 -56410 80750
rect -56090 80550 -56020 80750
rect -55980 80550 -55910 80750
rect -55590 80550 -55520 80750
rect -55480 80550 -55410 80750
rect -55090 80550 -55020 80750
rect -54980 80550 -54910 80750
rect -54590 80550 -54520 80750
rect -54480 80550 -54410 80750
rect -54090 80550 -54020 80750
rect -53980 80550 -53910 80750
rect -53590 80550 -53520 80750
rect -53480 80550 -53410 80750
rect -53090 80550 -53020 80750
rect -52980 80550 -52910 80750
rect -52590 80550 -52520 80750
rect -52480 80550 -52410 80750
rect -52090 80550 -52020 80750
rect -51980 80550 -51910 80750
rect -51590 80550 -51520 80750
rect -51480 80550 -51410 80750
rect -51090 80550 -51020 80750
rect -50980 80550 -50910 80750
rect -50590 80550 -50520 80750
rect -50480 80550 -50410 80750
rect -50090 80550 -50020 80750
rect -49980 80550 -49910 80750
rect -49590 80550 -49520 80750
rect -49480 80550 -49410 80750
rect -49090 80550 -49020 80750
rect -48980 80550 -48910 80750
rect -48590 80550 -48520 80750
rect -48480 80550 -48410 80750
rect -48090 80550 -48020 80750
rect -47980 80550 -47910 80750
rect -47590 80550 -47520 80750
rect -47480 80550 -47410 80750
rect -47090 80550 -47020 80750
rect -46980 80550 -46910 80750
rect -46590 80550 -46520 80750
rect -46480 80550 -46410 80750
rect -46090 80550 -46020 80750
rect -45980 80550 -45910 80750
rect -45590 80550 -45520 80750
rect -45480 80550 -45410 80750
rect -45090 80550 -45020 80750
rect -44980 80550 -44910 80750
rect -44590 80550 -44520 80750
rect -44480 80550 -44410 80750
rect -44090 80550 -44020 80750
rect -43980 80550 -43910 80750
rect -43590 80550 -43520 80750
rect -43480 80550 -43410 80750
rect -43090 80550 -43020 80750
rect -42980 80550 -42910 80750
rect -42590 80550 -42520 80750
rect -42480 80550 -42410 80750
rect -42090 80550 -42020 80750
rect -41980 80550 -41910 80750
rect -41590 80550 -41520 80750
rect -41480 80550 -41410 80750
rect -41090 80550 -41020 80750
rect -40980 80550 -40910 80750
rect -40590 80550 -40520 80750
rect -40480 80550 -40410 80750
rect -40090 80550 -40020 80750
rect -39980 80550 -39910 80750
rect -39590 80550 -39520 80750
rect -39480 80550 -39410 80750
rect -39090 80550 -39020 80750
rect -38980 80550 -38910 80750
rect -38590 80550 -38520 80750
rect -38480 80550 -38410 80750
rect -38090 80550 -38020 80750
rect -37980 80550 -37910 80750
rect -37590 80550 -37520 80750
rect -37480 80550 -37410 80750
rect -37090 80550 -37020 80750
rect -36980 80550 -36910 80750
rect -36590 80550 -36520 80750
rect -36480 80550 -36410 80750
rect -36090 80550 -36020 80750
rect -35980 80550 -35910 80750
rect -35590 80550 -35520 80750
rect -35480 80550 -35410 80750
rect -35090 80550 -35020 80750
rect -34980 80550 -34910 80750
rect -34590 80550 -34520 80750
rect -34480 80550 -34410 80750
rect -34090 80550 -34020 80750
rect -33980 80550 -33910 80750
rect -33590 80550 -33520 80750
rect -33480 80550 -33410 80750
rect -33090 80550 -33020 80750
rect -32980 80550 -32910 80750
rect -32590 80550 -32520 80750
rect -32480 80550 -32410 80750
rect -32090 80550 -32020 80750
rect -31980 80550 -31910 80750
rect -31590 80550 -31520 80750
rect -31480 80550 -31410 80750
rect -31090 80550 -31020 80750
rect -30980 80550 -30910 80750
rect -30590 80550 -30520 80750
rect -30480 80550 -30410 80750
rect -30090 80550 -30020 80750
rect -29980 80550 -29910 80750
rect -29590 80550 -29520 80750
rect -29480 80550 -29410 80750
rect -29090 80550 -29020 80750
rect -28980 80550 -28910 80750
rect -28590 80550 -28520 80750
rect -28480 80550 -28410 80750
rect -28090 80550 -28020 80750
rect -27980 80550 -27910 80750
rect -27590 80550 -27520 80750
rect -27480 80550 -27410 80750
rect -27090 80550 -27020 80750
rect -26980 80550 -26910 80750
rect -26590 80550 -26520 80750
rect -26480 80550 -26410 80750
rect -26090 80550 -26020 80750
rect -25980 80550 -25910 80750
rect -25590 80550 -25520 80750
rect -25480 80550 -25410 80750
rect -25090 80550 -25020 80750
rect -24980 80550 -24910 80750
rect -24590 80550 -24520 80750
rect -24480 80550 -24410 80750
rect -24090 80550 -24020 80750
rect -23980 80550 -23910 80750
rect -23590 80550 -23520 80750
rect -23480 80550 -23410 80750
rect -23090 80550 -23020 80750
rect -22980 80550 -22910 80750
rect -22590 80550 -22520 80750
rect -22480 80550 -22410 80750
rect -22090 80550 -22020 80750
rect -21980 80550 -21910 80750
rect -21590 80550 -21520 80750
rect -21480 80550 -21410 80750
rect -21090 80550 -21020 80750
rect -20980 80550 -20910 80750
rect -20590 80550 -20520 80750
rect -20480 80550 -20410 80750
rect -20090 80550 -20020 80750
rect -19980 80550 -19910 80750
rect -19590 80550 -19520 80750
rect -19480 80550 -19410 80750
rect -19090 80550 -19020 80750
rect -18980 80550 -18910 80750
rect -18590 80550 -18520 80750
rect -18480 80550 -18410 80750
rect -18090 80550 -18020 80750
rect -17980 80550 -17910 80750
rect -17590 80550 -17520 80750
rect -17480 80550 -17410 80750
rect -17090 80550 -17020 80750
rect -16980 80550 -16910 80750
rect -16590 80550 -16520 80750
rect -16480 80550 -16410 80750
rect -16090 80550 -16020 80750
rect -15980 80550 -15910 80750
rect -15590 80550 -15520 80750
rect -15480 80550 -15410 80750
rect -15090 80550 -15020 80750
rect -14980 80550 -14910 80750
rect -14590 80550 -14520 80750
rect -14480 80550 -14410 80750
rect -14090 80550 -14020 80750
rect -13980 80550 -13910 80750
rect -13590 80550 -13520 80750
rect -13480 80550 -13410 80750
rect -13090 80550 -13020 80750
rect -12980 80550 -12910 80750
rect -12590 80550 -12520 80750
rect -12480 80550 -12410 80750
rect -12090 80550 -12020 80750
rect -11980 80550 -11910 80750
rect -11590 80550 -11520 80750
rect -11480 80550 -11410 80750
rect -11090 80550 -11020 80750
rect -10980 80550 -10910 80750
rect -10590 80550 -10520 80750
rect -10480 80550 -10410 80750
rect -10090 80550 -10020 80750
rect -9980 80550 -9910 80750
rect -9590 80550 -9520 80750
rect -9480 80550 -9410 80750
rect -9090 80550 -9020 80750
rect -8980 80550 -8910 80750
rect -8590 80550 -8520 80750
rect -8480 80550 -8410 80750
rect -8090 80550 -8020 80750
rect -7980 80550 -7910 80750
rect -7590 80550 -7520 80750
rect -7480 80550 -7410 80750
rect -7090 80550 -7020 80750
rect -6980 80550 -6910 80750
rect -6590 80550 -6520 80750
rect -6480 80550 -6410 80750
rect -6090 80550 -6020 80750
rect -5980 80550 -5910 80750
rect -5590 80550 -5520 80750
rect -5480 80550 -5410 80750
rect -5090 80550 -5020 80750
rect -4980 80550 -4910 80750
rect -4590 80550 -4520 80750
rect -4480 80550 -4410 80750
rect -4090 80550 -4020 80750
rect -3980 80550 -3910 80750
rect -3590 80550 -3520 80750
rect -3480 80550 -3410 80750
rect -3090 80550 -3020 80750
rect -2980 80550 -2910 80750
rect -2590 80550 -2520 80750
rect -2480 80550 -2410 80750
rect -2090 80550 -2020 80750
rect -1980 80550 -1910 80750
rect -1590 80550 -1520 80750
rect -1480 80550 -1410 80750
rect -1090 80550 -1020 80750
rect -980 80550 -910 80750
rect -590 80550 -520 80750
rect -480 80550 -410 80750
rect -90 80550 -20 80750
rect 20 80550 90 80750
rect 410 80550 480 80750
rect 520 80550 590 80750
rect 910 80550 980 80750
rect 1020 80550 1090 80750
rect 1410 80550 1480 80750
rect 1520 80550 1590 80750
rect 1910 80550 1980 80750
rect 2020 80550 2090 80750
rect 2410 80550 2480 80750
rect 2520 80550 2590 80750
rect 2910 80550 2980 80750
rect 3020 80550 3090 80750
rect 3410 80550 3480 80750
rect 3520 80550 3590 80750
rect 3910 80550 3980 80750
rect 4020 80550 4090 80750
rect 4410 80550 4480 80750
rect 4520 80550 4590 80750
rect 4910 80550 4980 80750
rect 5020 80550 5090 80750
rect 5410 80550 5480 80750
rect 5520 80550 5590 80750
rect 5910 80550 5980 80750
rect 6020 80550 6090 80750
rect 6410 80550 6480 80750
rect 6520 80550 6590 80750
rect 6910 80550 6980 80750
rect 7020 80550 7090 80750
rect 7410 80550 7480 80750
rect 7520 80550 7590 80750
rect 7910 80550 7980 80750
rect 8020 80550 8090 80750
rect 8410 80550 8480 80750
rect 8520 80550 8590 80750
rect 8910 80550 8980 80750
rect 9020 80550 9090 80750
rect 9410 80550 9480 80750
rect 9520 80550 9590 80750
rect 9910 80550 9980 80750
rect 10020 80550 10090 80750
rect 10410 80550 10480 80750
rect 10520 80550 10590 80750
rect 10910 80550 10980 80750
rect 11020 80550 11090 80750
rect 11410 80550 11480 80750
rect 11520 80550 11590 80750
rect 11910 80550 11980 80750
rect 12020 80550 12090 80750
rect 12410 80550 12480 80750
rect 12520 80550 12590 80750
rect 12910 80550 12980 80750
rect 13020 80550 13090 80750
rect 13410 80550 13480 80750
rect 13520 80550 13590 80750
rect 13910 80550 13980 80750
rect 14020 80550 14090 80750
rect 14410 80550 14480 80750
rect 14520 80550 14590 80750
rect 14910 80550 14980 80750
rect 15020 80550 15090 80750
rect 15410 80550 15480 80750
rect 15520 80550 15590 80750
rect 15910 80550 15980 80750
rect 16020 80550 16090 80750
rect 16410 80550 16480 80750
rect 16520 80550 16590 80750
rect 16910 80550 16980 80750
rect 17020 80550 17090 80750
rect 17410 80550 17480 80750
rect 17520 80550 17590 80750
rect 17910 80550 17980 80750
rect 18020 80550 18090 80750
rect 18410 80550 18480 80750
rect 18520 80550 18590 80750
rect 18910 80550 18980 80750
rect 19020 80550 19090 80750
rect 19410 80550 19480 80750
rect 19520 80550 19590 80750
rect 19910 80550 19980 80750
rect 20020 80550 20090 80750
rect 20410 80550 20480 80750
rect 20520 80550 20590 80750
rect 20910 80550 20980 80750
rect 21020 80550 21090 80750
rect 21410 80550 21480 80750
rect 21520 80550 21590 80750
rect 21910 80550 21980 80750
rect 22020 80550 22090 80750
rect 22410 80550 22480 80750
rect 22520 80550 22590 80750
rect 22910 80550 22980 80750
rect 23020 80550 23090 80750
rect 23410 80550 23480 80750
rect 23520 80550 23590 80750
rect 23910 80550 23980 80750
rect 24020 80550 24090 80750
rect 24410 80550 24480 80750
rect 24520 80550 24590 80750
rect 24910 80550 24980 80750
rect 25020 80550 25090 80750
rect 25410 80550 25480 80750
rect 25520 80550 25590 80750
rect 25910 80550 25980 80750
rect 26020 80550 26090 80750
rect 26410 80550 26480 80750
rect 26520 80550 26590 80750
rect 26910 80550 26980 80750
rect 27020 80550 27090 80750
rect 27410 80550 27480 80750
rect 27520 80550 27590 80750
rect 27910 80550 27980 80750
rect 28020 80550 28090 80750
rect 28410 80550 28480 80750
rect 28520 80550 28590 80750
rect 28910 80550 28980 80750
rect 29020 80550 29090 80750
rect 29410 80550 29480 80750
rect 29520 80550 29590 80750
rect 29910 80550 29980 80750
rect 30020 80550 30090 80750
rect 30410 80550 30480 80750
rect 30520 80550 30590 80750
rect 30910 80550 30980 80750
rect 31020 80550 31090 80750
rect 31410 80550 31480 80750
rect 31520 80550 31590 80750
rect 31910 80550 31980 80750
rect 32020 80550 32090 80750
rect 32410 80550 32480 80750
rect 32520 80550 32590 80750
rect 32910 80550 32980 80750
rect 33020 80550 33090 80750
rect 33410 80550 33480 80750
rect 33520 80550 33590 80750
rect 33910 80550 33980 80750
rect 34020 80550 34090 80750
rect 34410 80550 34480 80750
rect 34520 80550 34590 80750
rect 34910 80550 34980 80750
rect 35020 80550 35090 80750
rect 35410 80550 35480 80750
rect 35520 80550 35590 80750
rect 35910 80550 35980 80750
rect 36020 80550 36090 80750
rect 36410 80550 36480 80750
rect 36520 80550 36590 80750
rect 36910 80550 36980 80750
rect 37020 80550 37090 80750
rect 37410 80550 37480 80750
rect 37520 80550 37590 80750
rect 37910 80550 37980 80750
rect 38020 80550 38090 80750
rect 38410 80550 38480 80750
rect 38520 80550 38590 80750
rect 38910 80550 38980 80750
rect 39020 80550 39090 80750
rect 39410 80550 39480 80750
rect 39520 80550 39590 80750
rect 39910 80550 39980 80750
rect 40020 80550 40090 80750
rect 40410 80550 40480 80750
rect 40520 80550 40590 80750
rect 40910 80550 40980 80750
rect 41020 80550 41090 80750
rect 41410 80550 41480 80750
rect 41520 80550 41590 80750
rect 41910 80550 41980 80750
rect 42020 80550 42090 80750
rect 42410 80550 42480 80750
rect 42520 80550 42590 80750
rect 42910 80550 42980 80750
rect 43020 80550 43090 80750
rect 43410 80550 43480 80750
rect 43520 80550 43590 80750
rect 43910 80550 43980 80750
rect 44020 80550 44090 80750
rect 44410 80550 44480 80750
rect 44520 80550 44590 80750
rect 44910 80550 44980 80750
rect 45020 80550 45090 80750
rect 45410 80550 45480 80750
rect 45520 80550 45590 80750
rect 45910 80550 45980 80750
rect 46020 80550 46090 80750
rect 46410 80550 46480 80750
rect 46520 80550 46590 80750
rect 46910 80550 46980 80750
rect 47020 80550 47090 80750
rect 47410 80550 47480 80750
rect 47520 80550 47590 80750
rect 47910 80550 47980 80750
rect 48020 80550 48090 80750
rect 48410 80550 48480 80750
rect 48520 80550 48590 80750
rect 48910 80550 48980 80750
rect 49020 80550 49090 80750
rect 49410 80550 49480 80750
rect 49520 80550 49590 80750
rect 49910 80550 49980 80750
rect 50020 80550 50090 80750
rect 50410 80550 50480 80750
rect 50520 80550 50590 80750
rect 50910 80550 50980 80750
rect 51020 80550 51090 80750
rect 51410 80550 51480 80750
rect 51520 80550 51590 80750
rect 51910 80550 51980 80750
rect 52020 80550 52090 80750
rect 52410 80550 52480 80750
rect 52520 80550 52590 80750
rect 52910 80550 52980 80750
rect 53020 80550 53090 80750
rect 53410 80550 53480 80750
rect 53520 80550 53590 80750
rect 53910 80550 53980 80750
rect 54020 80550 54090 80750
rect 54410 80550 54480 80750
rect 54520 80550 54590 80750
rect 54910 80550 54980 80750
rect 55020 80550 55090 80750
rect 55410 80550 55480 80750
rect 55520 80550 55590 80750
rect 55910 80550 55980 80750
rect 56020 80550 56090 80750
rect 56410 80550 56480 80750
rect 56520 80550 56590 80750
rect 56910 80550 56980 80750
rect 57020 80550 57090 80750
rect 57410 80550 57480 80750
rect 57520 80550 57590 80750
rect 57910 80550 57980 80750
rect 58020 80550 58090 80750
rect 58410 80550 58480 80750
rect 58520 80550 58590 80750
rect 58910 80550 58980 80750
rect 59020 80550 59090 80750
rect 59410 80550 59480 80750
rect 59520 80550 59590 80750
rect 59910 80550 59980 80750
rect 60020 80550 60090 80750
rect 60410 80550 60480 80750
rect 60520 80550 60590 80750
rect 60910 80550 60980 80750
rect 61020 80550 61090 80750
rect 61410 80550 61480 80750
rect 61520 80550 61590 80750
rect 61910 80550 61980 80750
rect 62020 80550 62090 80750
rect 62410 80550 62480 80750
rect 62520 80550 62590 80750
rect 62910 80550 62980 80750
rect 63020 80550 63090 80750
rect 63410 80550 63480 80750
rect 63520 80550 63590 80750
rect 63910 80550 63980 80750
rect 64020 80550 64090 80750
rect 64410 80550 64480 80750
rect 64520 80550 64590 80750
rect 64910 80550 64980 80750
rect 65020 80550 65090 80750
rect 65410 80550 65480 80750
rect 65520 80550 65590 80750
rect 65910 80550 65980 80750
rect 66020 80550 66090 80750
rect 66410 80550 66480 80750
rect 66520 80550 66590 80750
rect 66910 80550 66980 80750
rect 67020 80550 67090 80750
rect 67410 80550 67480 80750
rect 67520 80550 67590 80750
rect 67910 80550 67980 80750
rect 68020 80550 68090 80750
rect 68410 80550 68480 80750
rect 68520 80550 68590 80750
rect 68910 80550 68980 80750
rect 69020 80550 69090 80750
rect 69410 80550 69480 80750
rect 69520 80550 69590 80750
rect 69910 80550 69980 80750
rect 70020 80550 70090 80750
rect 70410 80550 70480 80750
rect 70520 80550 70590 80750
rect 70910 80550 70980 80750
rect 71020 80550 71090 80750
rect 71410 80550 71480 80750
rect 71520 80550 71590 80750
rect 71910 80550 71980 80750
rect 72020 80550 72090 80750
rect 72410 80550 72480 80750
rect 72520 80550 72590 80750
rect 72910 80550 72980 80750
rect 73020 80550 73090 80750
rect 73410 80550 73480 80750
rect 73520 80550 73590 80750
rect 73910 80550 73980 80750
rect 74020 80550 74090 80750
rect 74410 80550 74480 80750
rect 74520 80550 74590 80750
rect 74910 80550 74980 80750
rect 75020 80550 75090 80750
rect 75410 80550 75480 80750
rect 75520 80550 75590 80750
rect 75910 80550 75980 80750
rect 76020 80550 76090 80750
rect 76410 80550 76480 80750
rect 76520 80550 76590 80750
rect 76910 80550 76980 80750
rect 77020 80550 77090 80750
rect 77410 80550 77480 80750
rect 77520 80550 77590 80750
rect 77910 80550 77980 80750
rect 78020 80550 78090 80750
rect 78410 80550 78480 80750
rect 78520 80550 78590 80750
rect 78910 80550 78980 80750
rect 79020 80550 79090 80750
rect 79410 80550 79480 80750
rect 79520 80550 79590 80750
rect 79910 80550 79980 80750
rect 80020 80550 80090 80750
rect 80410 80550 80480 80750
rect 80520 80550 80590 80750
rect 80910 80550 80980 80750
rect 81020 80550 81090 80750
rect 81410 80550 81480 80750
rect 81520 80550 81590 80750
rect 81910 80550 81980 80750
rect 82020 80550 82090 80750
rect 82410 80550 82480 80750
rect 82520 80550 82590 80750
rect 82910 80550 82980 80750
rect 83020 80550 83090 80750
rect 83410 80550 83480 80750
rect 83520 80550 83590 80750
rect 83910 80550 83980 80750
rect 84020 80550 84090 80750
rect 84410 80550 84480 80750
rect 84520 80550 84590 80750
rect 84910 80550 84980 80750
rect 85020 80550 85090 80750
rect 85410 80550 85480 80750
rect 85520 80550 85590 80750
rect 85910 80550 85980 80750
rect 86020 80550 86090 80750
rect 86410 80550 86480 80750
rect 86520 80550 86590 80750
rect 86910 80550 86980 80750
rect 87020 80550 87090 80750
rect 87410 80550 87480 80750
rect 87520 80550 87590 80750
rect 87910 80550 87980 80750
rect 88020 80550 88090 80750
rect 88410 80550 88480 80750
rect 88520 80550 88590 80750
rect 88910 80550 88980 80750
rect 89020 80550 89090 80750
rect 89410 80550 89480 80750
rect 89520 80550 89590 80750
rect 89910 80550 89980 80750
rect 90020 80550 90090 80750
rect 90410 80550 90480 80750
rect 90520 80550 90590 80750
rect 90910 80550 90980 80750
rect 91020 80550 91090 80750
rect 91410 80550 91480 80750
rect 91520 80550 91590 80750
rect 91910 80550 91980 80750
rect 92020 80550 92090 80750
rect 92410 80550 92480 80750
rect 92520 80550 92590 80750
rect 92910 80550 92980 80750
rect 93020 80550 93090 80750
rect 93410 80550 93480 80750
rect 93520 80550 93590 80750
rect 93910 80550 93980 80750
rect 94020 80550 94090 80750
rect 94410 80550 94480 80750
rect 94520 80550 94590 80750
rect 94910 80550 94980 80750
rect 95020 80550 95090 80750
rect 95410 80550 95480 80750
rect 95520 80550 95590 80750
rect 95910 80550 95980 80750
rect 96020 80550 96090 80750
rect 96410 80550 96480 80750
rect 96520 80550 96590 80750
rect 96910 80550 96980 80750
rect 97020 80550 97090 80750
rect 97410 80550 97480 80750
rect 97520 80550 97590 80750
rect 97910 80550 97980 80750
rect 98020 80550 98090 80750
rect 98410 80550 98480 80750
rect 98520 80550 98590 80750
rect 98910 80550 98980 80750
rect 99020 80550 99090 80750
rect 99410 80550 99480 80750
rect 99520 80550 99590 80750
rect 99910 80550 99980 80750
rect 100020 80550 100090 80750
rect 100410 80550 100480 80750
rect -83350 80420 -83150 80490
rect -82850 80420 -82650 80490
rect -82350 80420 -82150 80490
rect -81850 80420 -81650 80490
rect -81350 80420 -81150 80490
rect -80850 80420 -80650 80490
rect -80350 80420 -80150 80490
rect -79850 80420 -79650 80490
rect -79350 80420 -79150 80490
rect -78850 80420 -78650 80490
rect -78350 80420 -78150 80490
rect -77850 80420 -77650 80490
rect -77350 80420 -77150 80490
rect -76850 80420 -76650 80490
rect -76350 80420 -76150 80490
rect -75850 80420 -75650 80490
rect -75350 80420 -75150 80490
rect -74850 80420 -74650 80490
rect -74350 80420 -74150 80490
rect -73850 80420 -73650 80490
rect -73350 80420 -73150 80490
rect -72850 80420 -72650 80490
rect -72350 80420 -72150 80490
rect -71850 80420 -71650 80490
rect -71350 80420 -71150 80490
rect -70850 80420 -70650 80490
rect -70350 80420 -70150 80490
rect -69850 80420 -69650 80490
rect -69350 80420 -69150 80490
rect -68850 80420 -68650 80490
rect -68350 80420 -68150 80490
rect -67850 80420 -67650 80490
rect -67350 80420 -67150 80490
rect -66850 80420 -66650 80490
rect -66350 80420 -66150 80490
rect -65850 80420 -65650 80490
rect -65350 80420 -65150 80490
rect -64850 80420 -64650 80490
rect -64350 80420 -64150 80490
rect -63850 80420 -63650 80490
rect -63350 80420 -63150 80490
rect -62850 80420 -62650 80490
rect -62350 80420 -62150 80490
rect -61850 80420 -61650 80490
rect -61350 80420 -61150 80490
rect -60850 80420 -60650 80490
rect -60350 80420 -60150 80490
rect -59850 80420 -59650 80490
rect -59350 80420 -59150 80490
rect -58850 80420 -58650 80490
rect -58350 80420 -58150 80490
rect -57850 80420 -57650 80490
rect -57350 80420 -57150 80490
rect -56850 80420 -56650 80490
rect -56350 80420 -56150 80490
rect -55850 80420 -55650 80490
rect -55350 80420 -55150 80490
rect -54850 80420 -54650 80490
rect -54350 80420 -54150 80490
rect -53850 80420 -53650 80490
rect -53350 80420 -53150 80490
rect -52850 80420 -52650 80490
rect -52350 80420 -52150 80490
rect -51850 80420 -51650 80490
rect -51350 80420 -51150 80490
rect -50850 80420 -50650 80490
rect -50350 80420 -50150 80490
rect -49850 80420 -49650 80490
rect -49350 80420 -49150 80490
rect -48850 80420 -48650 80490
rect -48350 80420 -48150 80490
rect -47850 80420 -47650 80490
rect -47350 80420 -47150 80490
rect -46850 80420 -46650 80490
rect -46350 80420 -46150 80490
rect -45850 80420 -45650 80490
rect -45350 80420 -45150 80490
rect -44850 80420 -44650 80490
rect -44350 80420 -44150 80490
rect -43850 80420 -43650 80490
rect -43350 80420 -43150 80490
rect -42850 80420 -42650 80490
rect -42350 80420 -42150 80490
rect -41850 80420 -41650 80490
rect -41350 80420 -41150 80490
rect -40850 80420 -40650 80490
rect -40350 80420 -40150 80490
rect -39850 80420 -39650 80490
rect -39350 80420 -39150 80490
rect -38850 80420 -38650 80490
rect -38350 80420 -38150 80490
rect -37850 80420 -37650 80490
rect -37350 80420 -37150 80490
rect -36850 80420 -36650 80490
rect -36350 80420 -36150 80490
rect -35850 80420 -35650 80490
rect -35350 80420 -35150 80490
rect -34850 80420 -34650 80490
rect -34350 80420 -34150 80490
rect -33850 80420 -33650 80490
rect -33350 80420 -33150 80490
rect -32850 80420 -32650 80490
rect -32350 80420 -32150 80490
rect -31850 80420 -31650 80490
rect -31350 80420 -31150 80490
rect -30850 80420 -30650 80490
rect -30350 80420 -30150 80490
rect -29850 80420 -29650 80490
rect -29350 80420 -29150 80490
rect -28850 80420 -28650 80490
rect -28350 80420 -28150 80490
rect -27850 80420 -27650 80490
rect -27350 80420 -27150 80490
rect -26850 80420 -26650 80490
rect -26350 80420 -26150 80490
rect -25850 80420 -25650 80490
rect -25350 80420 -25150 80490
rect -24850 80420 -24650 80490
rect -24350 80420 -24150 80490
rect -23850 80420 -23650 80490
rect -23350 80420 -23150 80490
rect -22850 80420 -22650 80490
rect -22350 80420 -22150 80490
rect -21850 80420 -21650 80490
rect -21350 80420 -21150 80490
rect -20850 80420 -20650 80490
rect -20350 80420 -20150 80490
rect -19850 80420 -19650 80490
rect -19350 80420 -19150 80490
rect -18850 80420 -18650 80490
rect -18350 80420 -18150 80490
rect -17850 80420 -17650 80490
rect -17350 80420 -17150 80490
rect -16850 80420 -16650 80490
rect -16350 80420 -16150 80490
rect -15850 80420 -15650 80490
rect -15350 80420 -15150 80490
rect -14850 80420 -14650 80490
rect -14350 80420 -14150 80490
rect -13850 80420 -13650 80490
rect -13350 80420 -13150 80490
rect -12850 80420 -12650 80490
rect -12350 80420 -12150 80490
rect -11850 80420 -11650 80490
rect -11350 80420 -11150 80490
rect -10850 80420 -10650 80490
rect -10350 80420 -10150 80490
rect -9850 80420 -9650 80490
rect -9350 80420 -9150 80490
rect -8850 80420 -8650 80490
rect -8350 80420 -8150 80490
rect -7850 80420 -7650 80490
rect -7350 80420 -7150 80490
rect -6850 80420 -6650 80490
rect -6350 80420 -6150 80490
rect -5850 80420 -5650 80490
rect -5350 80420 -5150 80490
rect -4850 80420 -4650 80490
rect -4350 80420 -4150 80490
rect -3850 80420 -3650 80490
rect -3350 80420 -3150 80490
rect -2850 80420 -2650 80490
rect -2350 80420 -2150 80490
rect -1850 80420 -1650 80490
rect -1350 80420 -1150 80490
rect -850 80420 -650 80490
rect -350 80420 -150 80490
rect 150 80420 350 80490
rect 650 80420 850 80490
rect 1150 80420 1350 80490
rect 1650 80420 1850 80490
rect 2150 80420 2350 80490
rect 2650 80420 2850 80490
rect 3150 80420 3350 80490
rect 3650 80420 3850 80490
rect 4150 80420 4350 80490
rect 4650 80420 4850 80490
rect 5150 80420 5350 80490
rect 5650 80420 5850 80490
rect 6150 80420 6350 80490
rect 6650 80420 6850 80490
rect 7150 80420 7350 80490
rect 7650 80420 7850 80490
rect 8150 80420 8350 80490
rect 8650 80420 8850 80490
rect 9150 80420 9350 80490
rect 9650 80420 9850 80490
rect 10150 80420 10350 80490
rect 10650 80420 10850 80490
rect 11150 80420 11350 80490
rect 11650 80420 11850 80490
rect 12150 80420 12350 80490
rect 12650 80420 12850 80490
rect 13150 80420 13350 80490
rect 13650 80420 13850 80490
rect 14150 80420 14350 80490
rect 14650 80420 14850 80490
rect 15150 80420 15350 80490
rect 15650 80420 15850 80490
rect 16150 80420 16350 80490
rect 16650 80420 16850 80490
rect 17150 80420 17350 80490
rect 17650 80420 17850 80490
rect 18150 80420 18350 80490
rect 18650 80420 18850 80490
rect 19150 80420 19350 80490
rect 19650 80420 19850 80490
rect 20150 80420 20350 80490
rect 20650 80420 20850 80490
rect 21150 80420 21350 80490
rect 21650 80420 21850 80490
rect 22150 80420 22350 80490
rect 22650 80420 22850 80490
rect 23150 80420 23350 80490
rect 23650 80420 23850 80490
rect 24150 80420 24350 80490
rect 24650 80420 24850 80490
rect 25150 80420 25350 80490
rect 25650 80420 25850 80490
rect 26150 80420 26350 80490
rect 26650 80420 26850 80490
rect 27150 80420 27350 80490
rect 27650 80420 27850 80490
rect 28150 80420 28350 80490
rect 28650 80420 28850 80490
rect 29150 80420 29350 80490
rect 29650 80420 29850 80490
rect 30150 80420 30350 80490
rect 30650 80420 30850 80490
rect 31150 80420 31350 80490
rect 31650 80420 31850 80490
rect 32150 80420 32350 80490
rect 32650 80420 32850 80490
rect 33150 80420 33350 80490
rect 33650 80420 33850 80490
rect 34150 80420 34350 80490
rect 34650 80420 34850 80490
rect 35150 80420 35350 80490
rect 35650 80420 35850 80490
rect 36150 80420 36350 80490
rect 36650 80420 36850 80490
rect 37150 80420 37350 80490
rect 37650 80420 37850 80490
rect 38150 80420 38350 80490
rect 38650 80420 38850 80490
rect 39150 80420 39350 80490
rect 39650 80420 39850 80490
rect 40150 80420 40350 80490
rect 40650 80420 40850 80490
rect 41150 80420 41350 80490
rect 41650 80420 41850 80490
rect 42150 80420 42350 80490
rect 42650 80420 42850 80490
rect 43150 80420 43350 80490
rect 43650 80420 43850 80490
rect 44150 80420 44350 80490
rect 44650 80420 44850 80490
rect 45150 80420 45350 80490
rect 45650 80420 45850 80490
rect 46150 80420 46350 80490
rect 46650 80420 46850 80490
rect 47150 80420 47350 80490
rect 47650 80420 47850 80490
rect 48150 80420 48350 80490
rect 48650 80420 48850 80490
rect 49150 80420 49350 80490
rect 49650 80420 49850 80490
rect 50150 80420 50350 80490
rect 50650 80420 50850 80490
rect 51150 80420 51350 80490
rect 51650 80420 51850 80490
rect 52150 80420 52350 80490
rect 52650 80420 52850 80490
rect 53150 80420 53350 80490
rect 53650 80420 53850 80490
rect 54150 80420 54350 80490
rect 54650 80420 54850 80490
rect 55150 80420 55350 80490
rect 55650 80420 55850 80490
rect 56150 80420 56350 80490
rect 56650 80420 56850 80490
rect 57150 80420 57350 80490
rect 57650 80420 57850 80490
rect 58150 80420 58350 80490
rect 58650 80420 58850 80490
rect 59150 80420 59350 80490
rect 59650 80420 59850 80490
rect 60150 80420 60350 80490
rect 60650 80420 60850 80490
rect 61150 80420 61350 80490
rect 61650 80420 61850 80490
rect 62150 80420 62350 80490
rect 62650 80420 62850 80490
rect 63150 80420 63350 80490
rect 63650 80420 63850 80490
rect 64150 80420 64350 80490
rect 64650 80420 64850 80490
rect 65150 80420 65350 80490
rect 65650 80420 65850 80490
rect 66150 80420 66350 80490
rect 66650 80420 66850 80490
rect 67150 80420 67350 80490
rect 67650 80420 67850 80490
rect 68150 80420 68350 80490
rect 68650 80420 68850 80490
rect 69150 80420 69350 80490
rect 69650 80420 69850 80490
rect 70150 80420 70350 80490
rect 70650 80420 70850 80490
rect 71150 80420 71350 80490
rect 71650 80420 71850 80490
rect 72150 80420 72350 80490
rect 72650 80420 72850 80490
rect 73150 80420 73350 80490
rect 73650 80420 73850 80490
rect 74150 80420 74350 80490
rect 74650 80420 74850 80490
rect 75150 80420 75350 80490
rect 75650 80420 75850 80490
rect 76150 80420 76350 80490
rect 76650 80420 76850 80490
rect 77150 80420 77350 80490
rect 77650 80420 77850 80490
rect 78150 80420 78350 80490
rect 78650 80420 78850 80490
rect 79150 80420 79350 80490
rect 79650 80420 79850 80490
rect 80150 80420 80350 80490
rect 80650 80420 80850 80490
rect 81150 80420 81350 80490
rect 81650 80420 81850 80490
rect 82150 80420 82350 80490
rect 82650 80420 82850 80490
rect 83150 80420 83350 80490
rect 83650 80420 83850 80490
rect 84150 80420 84350 80490
rect 84650 80420 84850 80490
rect 85150 80420 85350 80490
rect 85650 80420 85850 80490
rect 86150 80420 86350 80490
rect 86650 80420 86850 80490
rect 87150 80420 87350 80490
rect 87650 80420 87850 80490
rect 88150 80420 88350 80490
rect 88650 80420 88850 80490
rect 89150 80420 89350 80490
rect 89650 80420 89850 80490
rect 90150 80420 90350 80490
rect 90650 80420 90850 80490
rect 91150 80420 91350 80490
rect 91650 80420 91850 80490
rect 92150 80420 92350 80490
rect 92650 80420 92850 80490
rect 93150 80420 93350 80490
rect 93650 80420 93850 80490
rect 94150 80420 94350 80490
rect 94650 80420 94850 80490
rect 95150 80420 95350 80490
rect 95650 80420 95850 80490
rect 96150 80420 96350 80490
rect 96650 80420 96850 80490
rect 97150 80420 97350 80490
rect 97650 80420 97850 80490
rect 98150 80420 98350 80490
rect 98650 80420 98850 80490
rect 99150 80420 99350 80490
rect 99650 80420 99850 80490
rect 100150 80420 100350 80490
rect -83350 80310 -83150 80380
rect -82850 80310 -82650 80380
rect -82350 80310 -82150 80380
rect -81850 80310 -81650 80380
rect -81350 80310 -81150 80380
rect -80850 80310 -80650 80380
rect -80350 80310 -80150 80380
rect -79850 80310 -79650 80380
rect -79350 80310 -79150 80380
rect -78850 80310 -78650 80380
rect -78350 80310 -78150 80380
rect -77850 80310 -77650 80380
rect -77350 80310 -77150 80380
rect -76850 80310 -76650 80380
rect -76350 80310 -76150 80380
rect -75850 80310 -75650 80380
rect -75350 80310 -75150 80380
rect -74850 80310 -74650 80380
rect -74350 80310 -74150 80380
rect -73850 80310 -73650 80380
rect -73350 80310 -73150 80380
rect -72850 80310 -72650 80380
rect -72350 80310 -72150 80380
rect -71850 80310 -71650 80380
rect -71350 80310 -71150 80380
rect -70850 80310 -70650 80380
rect -70350 80310 -70150 80380
rect -69850 80310 -69650 80380
rect -69350 80310 -69150 80380
rect -68850 80310 -68650 80380
rect -68350 80310 -68150 80380
rect -67850 80310 -67650 80380
rect -67350 80310 -67150 80380
rect -66850 80310 -66650 80380
rect -66350 80310 -66150 80380
rect -65850 80310 -65650 80380
rect -65350 80310 -65150 80380
rect -64850 80310 -64650 80380
rect -64350 80310 -64150 80380
rect -63850 80310 -63650 80380
rect -63350 80310 -63150 80380
rect -62850 80310 -62650 80380
rect -62350 80310 -62150 80380
rect -61850 80310 -61650 80380
rect -61350 80310 -61150 80380
rect -60850 80310 -60650 80380
rect -60350 80310 -60150 80380
rect -59850 80310 -59650 80380
rect -59350 80310 -59150 80380
rect -58850 80310 -58650 80380
rect -58350 80310 -58150 80380
rect -57850 80310 -57650 80380
rect -57350 80310 -57150 80380
rect -56850 80310 -56650 80380
rect -56350 80310 -56150 80380
rect -55850 80310 -55650 80380
rect -55350 80310 -55150 80380
rect -54850 80310 -54650 80380
rect -54350 80310 -54150 80380
rect -53850 80310 -53650 80380
rect -53350 80310 -53150 80380
rect -52850 80310 -52650 80380
rect -52350 80310 -52150 80380
rect -51850 80310 -51650 80380
rect -51350 80310 -51150 80380
rect -50850 80310 -50650 80380
rect -50350 80310 -50150 80380
rect -49850 80310 -49650 80380
rect -49350 80310 -49150 80380
rect -48850 80310 -48650 80380
rect -48350 80310 -48150 80380
rect -47850 80310 -47650 80380
rect -47350 80310 -47150 80380
rect -46850 80310 -46650 80380
rect -46350 80310 -46150 80380
rect -45850 80310 -45650 80380
rect -45350 80310 -45150 80380
rect -44850 80310 -44650 80380
rect -44350 80310 -44150 80380
rect -43850 80310 -43650 80380
rect -43350 80310 -43150 80380
rect -42850 80310 -42650 80380
rect -42350 80310 -42150 80380
rect -41850 80310 -41650 80380
rect -41350 80310 -41150 80380
rect -40850 80310 -40650 80380
rect -40350 80310 -40150 80380
rect -39850 80310 -39650 80380
rect -39350 80310 -39150 80380
rect -38850 80310 -38650 80380
rect -38350 80310 -38150 80380
rect -37850 80310 -37650 80380
rect -37350 80310 -37150 80380
rect -36850 80310 -36650 80380
rect -36350 80310 -36150 80380
rect -35850 80310 -35650 80380
rect -35350 80310 -35150 80380
rect -34850 80310 -34650 80380
rect -34350 80310 -34150 80380
rect -33850 80310 -33650 80380
rect -33350 80310 -33150 80380
rect -32850 80310 -32650 80380
rect -32350 80310 -32150 80380
rect -31850 80310 -31650 80380
rect -31350 80310 -31150 80380
rect -30850 80310 -30650 80380
rect -30350 80310 -30150 80380
rect -29850 80310 -29650 80380
rect -29350 80310 -29150 80380
rect -28850 80310 -28650 80380
rect -28350 80310 -28150 80380
rect -27850 80310 -27650 80380
rect -27350 80310 -27150 80380
rect -26850 80310 -26650 80380
rect -26350 80310 -26150 80380
rect -25850 80310 -25650 80380
rect -25350 80310 -25150 80380
rect -24850 80310 -24650 80380
rect -24350 80310 -24150 80380
rect -23850 80310 -23650 80380
rect -23350 80310 -23150 80380
rect -22850 80310 -22650 80380
rect -22350 80310 -22150 80380
rect -21850 80310 -21650 80380
rect -21350 80310 -21150 80380
rect -20850 80310 -20650 80380
rect -20350 80310 -20150 80380
rect -19850 80310 -19650 80380
rect -19350 80310 -19150 80380
rect -18850 80310 -18650 80380
rect -18350 80310 -18150 80380
rect -17850 80310 -17650 80380
rect -17350 80310 -17150 80380
rect -16850 80310 -16650 80380
rect -16350 80310 -16150 80380
rect -15850 80310 -15650 80380
rect -15350 80310 -15150 80380
rect -14850 80310 -14650 80380
rect -14350 80310 -14150 80380
rect -13850 80310 -13650 80380
rect -13350 80310 -13150 80380
rect -12850 80310 -12650 80380
rect -12350 80310 -12150 80380
rect -11850 80310 -11650 80380
rect -11350 80310 -11150 80380
rect -10850 80310 -10650 80380
rect -10350 80310 -10150 80380
rect -9850 80310 -9650 80380
rect -9350 80310 -9150 80380
rect -8850 80310 -8650 80380
rect -8350 80310 -8150 80380
rect -7850 80310 -7650 80380
rect -7350 80310 -7150 80380
rect -6850 80310 -6650 80380
rect -6350 80310 -6150 80380
rect -5850 80310 -5650 80380
rect -5350 80310 -5150 80380
rect -4850 80310 -4650 80380
rect -4350 80310 -4150 80380
rect -3850 80310 -3650 80380
rect -3350 80310 -3150 80380
rect -2850 80310 -2650 80380
rect -2350 80310 -2150 80380
rect -1850 80310 -1650 80380
rect -1350 80310 -1150 80380
rect -850 80310 -650 80380
rect -350 80310 -150 80380
rect 150 80310 350 80380
rect 650 80310 850 80380
rect 1150 80310 1350 80380
rect 1650 80310 1850 80380
rect 2150 80310 2350 80380
rect 2650 80310 2850 80380
rect 3150 80310 3350 80380
rect 3650 80310 3850 80380
rect 4150 80310 4350 80380
rect 4650 80310 4850 80380
rect 5150 80310 5350 80380
rect 5650 80310 5850 80380
rect 6150 80310 6350 80380
rect 6650 80310 6850 80380
rect 7150 80310 7350 80380
rect 7650 80310 7850 80380
rect 8150 80310 8350 80380
rect 8650 80310 8850 80380
rect 9150 80310 9350 80380
rect 9650 80310 9850 80380
rect 10150 80310 10350 80380
rect 10650 80310 10850 80380
rect 11150 80310 11350 80380
rect 11650 80310 11850 80380
rect 12150 80310 12350 80380
rect 12650 80310 12850 80380
rect 13150 80310 13350 80380
rect 13650 80310 13850 80380
rect 14150 80310 14350 80380
rect 14650 80310 14850 80380
rect 15150 80310 15350 80380
rect 15650 80310 15850 80380
rect 16150 80310 16350 80380
rect 16650 80310 16850 80380
rect 17150 80310 17350 80380
rect 17650 80310 17850 80380
rect 18150 80310 18350 80380
rect 18650 80310 18850 80380
rect 19150 80310 19350 80380
rect 19650 80310 19850 80380
rect 20150 80310 20350 80380
rect 20650 80310 20850 80380
rect 21150 80310 21350 80380
rect 21650 80310 21850 80380
rect 22150 80310 22350 80380
rect 22650 80310 22850 80380
rect 23150 80310 23350 80380
rect 23650 80310 23850 80380
rect 24150 80310 24350 80380
rect 24650 80310 24850 80380
rect 25150 80310 25350 80380
rect 25650 80310 25850 80380
rect 26150 80310 26350 80380
rect 26650 80310 26850 80380
rect 27150 80310 27350 80380
rect 27650 80310 27850 80380
rect 28150 80310 28350 80380
rect 28650 80310 28850 80380
rect 29150 80310 29350 80380
rect 29650 80310 29850 80380
rect 30150 80310 30350 80380
rect 30650 80310 30850 80380
rect 31150 80310 31350 80380
rect 31650 80310 31850 80380
rect 32150 80310 32350 80380
rect 32650 80310 32850 80380
rect 33150 80310 33350 80380
rect 33650 80310 33850 80380
rect 34150 80310 34350 80380
rect 34650 80310 34850 80380
rect 35150 80310 35350 80380
rect 35650 80310 35850 80380
rect 36150 80310 36350 80380
rect 36650 80310 36850 80380
rect 37150 80310 37350 80380
rect 37650 80310 37850 80380
rect 38150 80310 38350 80380
rect 38650 80310 38850 80380
rect 39150 80310 39350 80380
rect 39650 80310 39850 80380
rect 40150 80310 40350 80380
rect 40650 80310 40850 80380
rect 41150 80310 41350 80380
rect 41650 80310 41850 80380
rect 42150 80310 42350 80380
rect 42650 80310 42850 80380
rect 43150 80310 43350 80380
rect 43650 80310 43850 80380
rect 44150 80310 44350 80380
rect 44650 80310 44850 80380
rect 45150 80310 45350 80380
rect 45650 80310 45850 80380
rect 46150 80310 46350 80380
rect 46650 80310 46850 80380
rect 47150 80310 47350 80380
rect 47650 80310 47850 80380
rect 48150 80310 48350 80380
rect 48650 80310 48850 80380
rect 49150 80310 49350 80380
rect 49650 80310 49850 80380
rect 50150 80310 50350 80380
rect 50650 80310 50850 80380
rect 51150 80310 51350 80380
rect 51650 80310 51850 80380
rect 52150 80310 52350 80380
rect 52650 80310 52850 80380
rect 53150 80310 53350 80380
rect 53650 80310 53850 80380
rect 54150 80310 54350 80380
rect 54650 80310 54850 80380
rect 55150 80310 55350 80380
rect 55650 80310 55850 80380
rect 56150 80310 56350 80380
rect 56650 80310 56850 80380
rect 57150 80310 57350 80380
rect 57650 80310 57850 80380
rect 58150 80310 58350 80380
rect 58650 80310 58850 80380
rect 59150 80310 59350 80380
rect 59650 80310 59850 80380
rect 60150 80310 60350 80380
rect 60650 80310 60850 80380
rect 61150 80310 61350 80380
rect 61650 80310 61850 80380
rect 62150 80310 62350 80380
rect 62650 80310 62850 80380
rect 63150 80310 63350 80380
rect 63650 80310 63850 80380
rect 64150 80310 64350 80380
rect 64650 80310 64850 80380
rect 65150 80310 65350 80380
rect 65650 80310 65850 80380
rect 66150 80310 66350 80380
rect 66650 80310 66850 80380
rect 67150 80310 67350 80380
rect 67650 80310 67850 80380
rect 68150 80310 68350 80380
rect 68650 80310 68850 80380
rect 69150 80310 69350 80380
rect 69650 80310 69850 80380
rect 70150 80310 70350 80380
rect 70650 80310 70850 80380
rect 71150 80310 71350 80380
rect 71650 80310 71850 80380
rect 72150 80310 72350 80380
rect 72650 80310 72850 80380
rect 73150 80310 73350 80380
rect 73650 80310 73850 80380
rect 74150 80310 74350 80380
rect 74650 80310 74850 80380
rect 75150 80310 75350 80380
rect 75650 80310 75850 80380
rect 76150 80310 76350 80380
rect 76650 80310 76850 80380
rect 77150 80310 77350 80380
rect 77650 80310 77850 80380
rect 78150 80310 78350 80380
rect 78650 80310 78850 80380
rect 79150 80310 79350 80380
rect 79650 80310 79850 80380
rect 80150 80310 80350 80380
rect 80650 80310 80850 80380
rect 81150 80310 81350 80380
rect 81650 80310 81850 80380
rect 82150 80310 82350 80380
rect 82650 80310 82850 80380
rect 83150 80310 83350 80380
rect 83650 80310 83850 80380
rect 84150 80310 84350 80380
rect 84650 80310 84850 80380
rect 85150 80310 85350 80380
rect 85650 80310 85850 80380
rect 86150 80310 86350 80380
rect 86650 80310 86850 80380
rect 87150 80310 87350 80380
rect 87650 80310 87850 80380
rect 88150 80310 88350 80380
rect 88650 80310 88850 80380
rect 89150 80310 89350 80380
rect 89650 80310 89850 80380
rect 90150 80310 90350 80380
rect 90650 80310 90850 80380
rect 91150 80310 91350 80380
rect 91650 80310 91850 80380
rect 92150 80310 92350 80380
rect 92650 80310 92850 80380
rect 93150 80310 93350 80380
rect 93650 80310 93850 80380
rect 94150 80310 94350 80380
rect 94650 80310 94850 80380
rect 95150 80310 95350 80380
rect 95650 80310 95850 80380
rect 96150 80310 96350 80380
rect 96650 80310 96850 80380
rect 97150 80310 97350 80380
rect 97650 80310 97850 80380
rect 98150 80310 98350 80380
rect 98650 80310 98850 80380
rect 99150 80310 99350 80380
rect 99650 80310 99850 80380
rect 100150 80310 100350 80380
rect -83480 80050 -83410 80250
rect -83090 80050 -83020 80250
rect -82980 80050 -82910 80250
rect -82590 80050 -82520 80250
rect -82480 80050 -82410 80250
rect -82090 80050 -82020 80250
rect -81980 80050 -81910 80250
rect -81590 80050 -81520 80250
rect -81480 80050 -81410 80250
rect -81090 80050 -81020 80250
rect -80980 80050 -80910 80250
rect -80590 80050 -80520 80250
rect -80480 80050 -80410 80250
rect -80090 80050 -80020 80250
rect -79980 80050 -79910 80250
rect -79590 80050 -79520 80250
rect -79480 80050 -79410 80250
rect -79090 80050 -79020 80250
rect -78980 80050 -78910 80250
rect -78590 80050 -78520 80250
rect -78480 80050 -78410 80250
rect -78090 80050 -78020 80250
rect -77980 80050 -77910 80250
rect -77590 80050 -77520 80250
rect -77480 80050 -77410 80250
rect -77090 80050 -77020 80250
rect -76980 80050 -76910 80250
rect -76590 80050 -76520 80250
rect -76480 80050 -76410 80250
rect -76090 80050 -76020 80250
rect -75980 80050 -75910 80250
rect -75590 80050 -75520 80250
rect -75480 80050 -75410 80250
rect -75090 80050 -75020 80250
rect -74980 80050 -74910 80250
rect -74590 80050 -74520 80250
rect -74480 80050 -74410 80250
rect -74090 80050 -74020 80250
rect -73980 80050 -73910 80250
rect -73590 80050 -73520 80250
rect -73480 80050 -73410 80250
rect -73090 80050 -73020 80250
rect -72980 80050 -72910 80250
rect -72590 80050 -72520 80250
rect -72480 80050 -72410 80250
rect -72090 80050 -72020 80250
rect -71980 80050 -71910 80250
rect -71590 80050 -71520 80250
rect -71480 80050 -71410 80250
rect -71090 80050 -71020 80250
rect -70980 80050 -70910 80250
rect -70590 80050 -70520 80250
rect -70480 80050 -70410 80250
rect -70090 80050 -70020 80250
rect -69980 80050 -69910 80250
rect -69590 80050 -69520 80250
rect -69480 80050 -69410 80250
rect -69090 80050 -69020 80250
rect -68980 80050 -68910 80250
rect -68590 80050 -68520 80250
rect -68480 80050 -68410 80250
rect -68090 80050 -68020 80250
rect -67980 80050 -67910 80250
rect -67590 80050 -67520 80250
rect -67480 80050 -67410 80250
rect -67090 80050 -67020 80250
rect -66980 80050 -66910 80250
rect -66590 80050 -66520 80250
rect -66480 80050 -66410 80250
rect -66090 80050 -66020 80250
rect -65980 80050 -65910 80250
rect -65590 80050 -65520 80250
rect -65480 80050 -65410 80250
rect -65090 80050 -65020 80250
rect -64980 80050 -64910 80250
rect -64590 80050 -64520 80250
rect -64480 80050 -64410 80250
rect -64090 80050 -64020 80250
rect -63980 80050 -63910 80250
rect -63590 80050 -63520 80250
rect -63480 80050 -63410 80250
rect -63090 80050 -63020 80250
rect -62980 80050 -62910 80250
rect -62590 80050 -62520 80250
rect -62480 80050 -62410 80250
rect -62090 80050 -62020 80250
rect -61980 80050 -61910 80250
rect -61590 80050 -61520 80250
rect -61480 80050 -61410 80250
rect -61090 80050 -61020 80250
rect -60980 80050 -60910 80250
rect -60590 80050 -60520 80250
rect -60480 80050 -60410 80250
rect -60090 80050 -60020 80250
rect -59980 80050 -59910 80250
rect -59590 80050 -59520 80250
rect -59480 80050 -59410 80250
rect -59090 80050 -59020 80250
rect -58980 80050 -58910 80250
rect -58590 80050 -58520 80250
rect -58480 80050 -58410 80250
rect -58090 80050 -58020 80250
rect -57980 80050 -57910 80250
rect -57590 80050 -57520 80250
rect -57480 80050 -57410 80250
rect -57090 80050 -57020 80250
rect -56980 80050 -56910 80250
rect -56590 80050 -56520 80250
rect -56480 80050 -56410 80250
rect -56090 80050 -56020 80250
rect -55980 80050 -55910 80250
rect -55590 80050 -55520 80250
rect -55480 80050 -55410 80250
rect -55090 80050 -55020 80250
rect -54980 80050 -54910 80250
rect -54590 80050 -54520 80250
rect -54480 80050 -54410 80250
rect -54090 80050 -54020 80250
rect -53980 80050 -53910 80250
rect -53590 80050 -53520 80250
rect -53480 80050 -53410 80250
rect -53090 80050 -53020 80250
rect -52980 80050 -52910 80250
rect -52590 80050 -52520 80250
rect -52480 80050 -52410 80250
rect -52090 80050 -52020 80250
rect -51980 80050 -51910 80250
rect -51590 80050 -51520 80250
rect -51480 80050 -51410 80250
rect -51090 80050 -51020 80250
rect -50980 80050 -50910 80250
rect -50590 80050 -50520 80250
rect -50480 80050 -50410 80250
rect -50090 80050 -50020 80250
rect -49980 80050 -49910 80250
rect -49590 80050 -49520 80250
rect -49480 80050 -49410 80250
rect -49090 80050 -49020 80250
rect -48980 80050 -48910 80250
rect -48590 80050 -48520 80250
rect -48480 80050 -48410 80250
rect -48090 80050 -48020 80250
rect -47980 80050 -47910 80250
rect -47590 80050 -47520 80250
rect -47480 80050 -47410 80250
rect -47090 80050 -47020 80250
rect -46980 80050 -46910 80250
rect -46590 80050 -46520 80250
rect -46480 80050 -46410 80250
rect -46090 80050 -46020 80250
rect -45980 80050 -45910 80250
rect -45590 80050 -45520 80250
rect -45480 80050 -45410 80250
rect -45090 80050 -45020 80250
rect -44980 80050 -44910 80250
rect -44590 80050 -44520 80250
rect -44480 80050 -44410 80250
rect -44090 80050 -44020 80250
rect -43980 80050 -43910 80250
rect -43590 80050 -43520 80250
rect -43480 80050 -43410 80250
rect -43090 80050 -43020 80250
rect -42980 80050 -42910 80250
rect -42590 80050 -42520 80250
rect -42480 80050 -42410 80250
rect -42090 80050 -42020 80250
rect -41980 80050 -41910 80250
rect -41590 80050 -41520 80250
rect -41480 80050 -41410 80250
rect -41090 80050 -41020 80250
rect -40980 80050 -40910 80250
rect -40590 80050 -40520 80250
rect -40480 80050 -40410 80250
rect -40090 80050 -40020 80250
rect -39980 80050 -39910 80250
rect -39590 80050 -39520 80250
rect -39480 80050 -39410 80250
rect -39090 80050 -39020 80250
rect -38980 80050 -38910 80250
rect -38590 80050 -38520 80250
rect -38480 80050 -38410 80250
rect -38090 80050 -38020 80250
rect -37980 80050 -37910 80250
rect -37590 80050 -37520 80250
rect -37480 80050 -37410 80250
rect -37090 80050 -37020 80250
rect -36980 80050 -36910 80250
rect -36590 80050 -36520 80250
rect -36480 80050 -36410 80250
rect -36090 80050 -36020 80250
rect -35980 80050 -35910 80250
rect -35590 80050 -35520 80250
rect -35480 80050 -35410 80250
rect -35090 80050 -35020 80250
rect -34980 80050 -34910 80250
rect -34590 80050 -34520 80250
rect -34480 80050 -34410 80250
rect -34090 80050 -34020 80250
rect -33980 80050 -33910 80250
rect -33590 80050 -33520 80250
rect -33480 80050 -33410 80250
rect -33090 80050 -33020 80250
rect -32980 80050 -32910 80250
rect -32590 80050 -32520 80250
rect -32480 80050 -32410 80250
rect -32090 80050 -32020 80250
rect -31980 80050 -31910 80250
rect -31590 80050 -31520 80250
rect -31480 80050 -31410 80250
rect -31090 80050 -31020 80250
rect -30980 80050 -30910 80250
rect -30590 80050 -30520 80250
rect -30480 80050 -30410 80250
rect -30090 80050 -30020 80250
rect -29980 80050 -29910 80250
rect -29590 80050 -29520 80250
rect -29480 80050 -29410 80250
rect -29090 80050 -29020 80250
rect -28980 80050 -28910 80250
rect -28590 80050 -28520 80250
rect -28480 80050 -28410 80250
rect -28090 80050 -28020 80250
rect -27980 80050 -27910 80250
rect -27590 80050 -27520 80250
rect -27480 80050 -27410 80250
rect -27090 80050 -27020 80250
rect -26980 80050 -26910 80250
rect -26590 80050 -26520 80250
rect -26480 80050 -26410 80250
rect -26090 80050 -26020 80250
rect -25980 80050 -25910 80250
rect -25590 80050 -25520 80250
rect -25480 80050 -25410 80250
rect -25090 80050 -25020 80250
rect -24980 80050 -24910 80250
rect -24590 80050 -24520 80250
rect -24480 80050 -24410 80250
rect -24090 80050 -24020 80250
rect -23980 80050 -23910 80250
rect -23590 80050 -23520 80250
rect -23480 80050 -23410 80250
rect -23090 80050 -23020 80250
rect -22980 80050 -22910 80250
rect -22590 80050 -22520 80250
rect -22480 80050 -22410 80250
rect -22090 80050 -22020 80250
rect -21980 80050 -21910 80250
rect -21590 80050 -21520 80250
rect -21480 80050 -21410 80250
rect -21090 80050 -21020 80250
rect -20980 80050 -20910 80250
rect -20590 80050 -20520 80250
rect -20480 80050 -20410 80250
rect -20090 80050 -20020 80250
rect -19980 80050 -19910 80250
rect -19590 80050 -19520 80250
rect -19480 80050 -19410 80250
rect -19090 80050 -19020 80250
rect -18980 80050 -18910 80250
rect -18590 80050 -18520 80250
rect -18480 80050 -18410 80250
rect -18090 80050 -18020 80250
rect -17980 80050 -17910 80250
rect -17590 80050 -17520 80250
rect -17480 80050 -17410 80250
rect -17090 80050 -17020 80250
rect -16980 80050 -16910 80250
rect -16590 80050 -16520 80250
rect -16480 80050 -16410 80250
rect -16090 80050 -16020 80250
rect -15980 80050 -15910 80250
rect -15590 80050 -15520 80250
rect -15480 80050 -15410 80250
rect -15090 80050 -15020 80250
rect -14980 80050 -14910 80250
rect -14590 80050 -14520 80250
rect -14480 80050 -14410 80250
rect -14090 80050 -14020 80250
rect -13980 80050 -13910 80250
rect -13590 80050 -13520 80250
rect -13480 80050 -13410 80250
rect -13090 80050 -13020 80250
rect -12980 80050 -12910 80250
rect -12590 80050 -12520 80250
rect -12480 80050 -12410 80250
rect -12090 80050 -12020 80250
rect -11980 80050 -11910 80250
rect -11590 80050 -11520 80250
rect -11480 80050 -11410 80250
rect -11090 80050 -11020 80250
rect -10980 80050 -10910 80250
rect -10590 80050 -10520 80250
rect -10480 80050 -10410 80250
rect -10090 80050 -10020 80250
rect -9980 80050 -9910 80250
rect -9590 80050 -9520 80250
rect -9480 80050 -9410 80250
rect -9090 80050 -9020 80250
rect -8980 80050 -8910 80250
rect -8590 80050 -8520 80250
rect -8480 80050 -8410 80250
rect -8090 80050 -8020 80250
rect -7980 80050 -7910 80250
rect -7590 80050 -7520 80250
rect -7480 80050 -7410 80250
rect -7090 80050 -7020 80250
rect -6980 80050 -6910 80250
rect -6590 80050 -6520 80250
rect -6480 80050 -6410 80250
rect -6090 80050 -6020 80250
rect -5980 80050 -5910 80250
rect -5590 80050 -5520 80250
rect -5480 80050 -5410 80250
rect -5090 80050 -5020 80250
rect -4980 80050 -4910 80250
rect -4590 80050 -4520 80250
rect -4480 80050 -4410 80250
rect -4090 80050 -4020 80250
rect -3980 80050 -3910 80250
rect -3590 80050 -3520 80250
rect -3480 80050 -3410 80250
rect -3090 80050 -3020 80250
rect -2980 80050 -2910 80250
rect -2590 80050 -2520 80250
rect -2480 80050 -2410 80250
rect -2090 80050 -2020 80250
rect -1980 80050 -1910 80250
rect -1590 80050 -1520 80250
rect -1480 80050 -1410 80250
rect -1090 80050 -1020 80250
rect -980 80050 -910 80250
rect -590 80050 -520 80250
rect -480 80050 -410 80250
rect -90 80050 -20 80250
rect 20 80050 90 80250
rect 410 80050 480 80250
rect 520 80050 590 80250
rect 910 80050 980 80250
rect 1020 80050 1090 80250
rect 1410 80050 1480 80250
rect 1520 80050 1590 80250
rect 1910 80050 1980 80250
rect 2020 80050 2090 80250
rect 2410 80050 2480 80250
rect 2520 80050 2590 80250
rect 2910 80050 2980 80250
rect 3020 80050 3090 80250
rect 3410 80050 3480 80250
rect 3520 80050 3590 80250
rect 3910 80050 3980 80250
rect 4020 80050 4090 80250
rect 4410 80050 4480 80250
rect 4520 80050 4590 80250
rect 4910 80050 4980 80250
rect 5020 80050 5090 80250
rect 5410 80050 5480 80250
rect 5520 80050 5590 80250
rect 5910 80050 5980 80250
rect 6020 80050 6090 80250
rect 6410 80050 6480 80250
rect 6520 80050 6590 80250
rect 6910 80050 6980 80250
rect 7020 80050 7090 80250
rect 7410 80050 7480 80250
rect 7520 80050 7590 80250
rect 7910 80050 7980 80250
rect 8020 80050 8090 80250
rect 8410 80050 8480 80250
rect 8520 80050 8590 80250
rect 8910 80050 8980 80250
rect 9020 80050 9090 80250
rect 9410 80050 9480 80250
rect 9520 80050 9590 80250
rect 9910 80050 9980 80250
rect 10020 80050 10090 80250
rect 10410 80050 10480 80250
rect 10520 80050 10590 80250
rect 10910 80050 10980 80250
rect 11020 80050 11090 80250
rect 11410 80050 11480 80250
rect 11520 80050 11590 80250
rect 11910 80050 11980 80250
rect 12020 80050 12090 80250
rect 12410 80050 12480 80250
rect 12520 80050 12590 80250
rect 12910 80050 12980 80250
rect 13020 80050 13090 80250
rect 13410 80050 13480 80250
rect 13520 80050 13590 80250
rect 13910 80050 13980 80250
rect 14020 80050 14090 80250
rect 14410 80050 14480 80250
rect 14520 80050 14590 80250
rect 14910 80050 14980 80250
rect 15020 80050 15090 80250
rect 15410 80050 15480 80250
rect 15520 80050 15590 80250
rect 15910 80050 15980 80250
rect 16020 80050 16090 80250
rect 16410 80050 16480 80250
rect 16520 80050 16590 80250
rect 16910 80050 16980 80250
rect 17020 80050 17090 80250
rect 17410 80050 17480 80250
rect 17520 80050 17590 80250
rect 17910 80050 17980 80250
rect 18020 80050 18090 80250
rect 18410 80050 18480 80250
rect 18520 80050 18590 80250
rect 18910 80050 18980 80250
rect 19020 80050 19090 80250
rect 19410 80050 19480 80250
rect 19520 80050 19590 80250
rect 19910 80050 19980 80250
rect 20020 80050 20090 80250
rect 20410 80050 20480 80250
rect 20520 80050 20590 80250
rect 20910 80050 20980 80250
rect 21020 80050 21090 80250
rect 21410 80050 21480 80250
rect 21520 80050 21590 80250
rect 21910 80050 21980 80250
rect 22020 80050 22090 80250
rect 22410 80050 22480 80250
rect 22520 80050 22590 80250
rect 22910 80050 22980 80250
rect 23020 80050 23090 80250
rect 23410 80050 23480 80250
rect 23520 80050 23590 80250
rect 23910 80050 23980 80250
rect 24020 80050 24090 80250
rect 24410 80050 24480 80250
rect 24520 80050 24590 80250
rect 24910 80050 24980 80250
rect 25020 80050 25090 80250
rect 25410 80050 25480 80250
rect 25520 80050 25590 80250
rect 25910 80050 25980 80250
rect 26020 80050 26090 80250
rect 26410 80050 26480 80250
rect 26520 80050 26590 80250
rect 26910 80050 26980 80250
rect 27020 80050 27090 80250
rect 27410 80050 27480 80250
rect 27520 80050 27590 80250
rect 27910 80050 27980 80250
rect 28020 80050 28090 80250
rect 28410 80050 28480 80250
rect 28520 80050 28590 80250
rect 28910 80050 28980 80250
rect 29020 80050 29090 80250
rect 29410 80050 29480 80250
rect 29520 80050 29590 80250
rect 29910 80050 29980 80250
rect 30020 80050 30090 80250
rect 30410 80050 30480 80250
rect 30520 80050 30590 80250
rect 30910 80050 30980 80250
rect 31020 80050 31090 80250
rect 31410 80050 31480 80250
rect 31520 80050 31590 80250
rect 31910 80050 31980 80250
rect 32020 80050 32090 80250
rect 32410 80050 32480 80250
rect 32520 80050 32590 80250
rect 32910 80050 32980 80250
rect 33020 80050 33090 80250
rect 33410 80050 33480 80250
rect 33520 80050 33590 80250
rect 33910 80050 33980 80250
rect 34020 80050 34090 80250
rect 34410 80050 34480 80250
rect 34520 80050 34590 80250
rect 34910 80050 34980 80250
rect 35020 80050 35090 80250
rect 35410 80050 35480 80250
rect 35520 80050 35590 80250
rect 35910 80050 35980 80250
rect 36020 80050 36090 80250
rect 36410 80050 36480 80250
rect 36520 80050 36590 80250
rect 36910 80050 36980 80250
rect 37020 80050 37090 80250
rect 37410 80050 37480 80250
rect 37520 80050 37590 80250
rect 37910 80050 37980 80250
rect 38020 80050 38090 80250
rect 38410 80050 38480 80250
rect 38520 80050 38590 80250
rect 38910 80050 38980 80250
rect 39020 80050 39090 80250
rect 39410 80050 39480 80250
rect 39520 80050 39590 80250
rect 39910 80050 39980 80250
rect 40020 80050 40090 80250
rect 40410 80050 40480 80250
rect 40520 80050 40590 80250
rect 40910 80050 40980 80250
rect 41020 80050 41090 80250
rect 41410 80050 41480 80250
rect 41520 80050 41590 80250
rect 41910 80050 41980 80250
rect 42020 80050 42090 80250
rect 42410 80050 42480 80250
rect 42520 80050 42590 80250
rect 42910 80050 42980 80250
rect 43020 80050 43090 80250
rect 43410 80050 43480 80250
rect 43520 80050 43590 80250
rect 43910 80050 43980 80250
rect 44020 80050 44090 80250
rect 44410 80050 44480 80250
rect 44520 80050 44590 80250
rect 44910 80050 44980 80250
rect 45020 80050 45090 80250
rect 45410 80050 45480 80250
rect 45520 80050 45590 80250
rect 45910 80050 45980 80250
rect 46020 80050 46090 80250
rect 46410 80050 46480 80250
rect 46520 80050 46590 80250
rect 46910 80050 46980 80250
rect 47020 80050 47090 80250
rect 47410 80050 47480 80250
rect 47520 80050 47590 80250
rect 47910 80050 47980 80250
rect 48020 80050 48090 80250
rect 48410 80050 48480 80250
rect 48520 80050 48590 80250
rect 48910 80050 48980 80250
rect 49020 80050 49090 80250
rect 49410 80050 49480 80250
rect 49520 80050 49590 80250
rect 49910 80050 49980 80250
rect 50020 80050 50090 80250
rect 50410 80050 50480 80250
rect 50520 80050 50590 80250
rect 50910 80050 50980 80250
rect 51020 80050 51090 80250
rect 51410 80050 51480 80250
rect 51520 80050 51590 80250
rect 51910 80050 51980 80250
rect 52020 80050 52090 80250
rect 52410 80050 52480 80250
rect 52520 80050 52590 80250
rect 52910 80050 52980 80250
rect 53020 80050 53090 80250
rect 53410 80050 53480 80250
rect 53520 80050 53590 80250
rect 53910 80050 53980 80250
rect 54020 80050 54090 80250
rect 54410 80050 54480 80250
rect 54520 80050 54590 80250
rect 54910 80050 54980 80250
rect 55020 80050 55090 80250
rect 55410 80050 55480 80250
rect 55520 80050 55590 80250
rect 55910 80050 55980 80250
rect 56020 80050 56090 80250
rect 56410 80050 56480 80250
rect 56520 80050 56590 80250
rect 56910 80050 56980 80250
rect 57020 80050 57090 80250
rect 57410 80050 57480 80250
rect 57520 80050 57590 80250
rect 57910 80050 57980 80250
rect 58020 80050 58090 80250
rect 58410 80050 58480 80250
rect 58520 80050 58590 80250
rect 58910 80050 58980 80250
rect 59020 80050 59090 80250
rect 59410 80050 59480 80250
rect 59520 80050 59590 80250
rect 59910 80050 59980 80250
rect 60020 80050 60090 80250
rect 60410 80050 60480 80250
rect 60520 80050 60590 80250
rect 60910 80050 60980 80250
rect 61020 80050 61090 80250
rect 61410 80050 61480 80250
rect 61520 80050 61590 80250
rect 61910 80050 61980 80250
rect 62020 80050 62090 80250
rect 62410 80050 62480 80250
rect 62520 80050 62590 80250
rect 62910 80050 62980 80250
rect 63020 80050 63090 80250
rect 63410 80050 63480 80250
rect 63520 80050 63590 80250
rect 63910 80050 63980 80250
rect 64020 80050 64090 80250
rect 64410 80050 64480 80250
rect 64520 80050 64590 80250
rect 64910 80050 64980 80250
rect 65020 80050 65090 80250
rect 65410 80050 65480 80250
rect 65520 80050 65590 80250
rect 65910 80050 65980 80250
rect 66020 80050 66090 80250
rect 66410 80050 66480 80250
rect 66520 80050 66590 80250
rect 66910 80050 66980 80250
rect 67020 80050 67090 80250
rect 67410 80050 67480 80250
rect 67520 80050 67590 80250
rect 67910 80050 67980 80250
rect 68020 80050 68090 80250
rect 68410 80050 68480 80250
rect 68520 80050 68590 80250
rect 68910 80050 68980 80250
rect 69020 80050 69090 80250
rect 69410 80050 69480 80250
rect 69520 80050 69590 80250
rect 69910 80050 69980 80250
rect 70020 80050 70090 80250
rect 70410 80050 70480 80250
rect 70520 80050 70590 80250
rect 70910 80050 70980 80250
rect 71020 80050 71090 80250
rect 71410 80050 71480 80250
rect 71520 80050 71590 80250
rect 71910 80050 71980 80250
rect 72020 80050 72090 80250
rect 72410 80050 72480 80250
rect 72520 80050 72590 80250
rect 72910 80050 72980 80250
rect 73020 80050 73090 80250
rect 73410 80050 73480 80250
rect 73520 80050 73590 80250
rect 73910 80050 73980 80250
rect 74020 80050 74090 80250
rect 74410 80050 74480 80250
rect 74520 80050 74590 80250
rect 74910 80050 74980 80250
rect 75020 80050 75090 80250
rect 75410 80050 75480 80250
rect 75520 80050 75590 80250
rect 75910 80050 75980 80250
rect 76020 80050 76090 80250
rect 76410 80050 76480 80250
rect 76520 80050 76590 80250
rect 76910 80050 76980 80250
rect 77020 80050 77090 80250
rect 77410 80050 77480 80250
rect 77520 80050 77590 80250
rect 77910 80050 77980 80250
rect 78020 80050 78090 80250
rect 78410 80050 78480 80250
rect 78520 80050 78590 80250
rect 78910 80050 78980 80250
rect 79020 80050 79090 80250
rect 79410 80050 79480 80250
rect 79520 80050 79590 80250
rect 79910 80050 79980 80250
rect 80020 80050 80090 80250
rect 80410 80050 80480 80250
rect 80520 80050 80590 80250
rect 80910 80050 80980 80250
rect 81020 80050 81090 80250
rect 81410 80050 81480 80250
rect 81520 80050 81590 80250
rect 81910 80050 81980 80250
rect 82020 80050 82090 80250
rect 82410 80050 82480 80250
rect 82520 80050 82590 80250
rect 82910 80050 82980 80250
rect 83020 80050 83090 80250
rect 83410 80050 83480 80250
rect 83520 80050 83590 80250
rect 83910 80050 83980 80250
rect 84020 80050 84090 80250
rect 84410 80050 84480 80250
rect 84520 80050 84590 80250
rect 84910 80050 84980 80250
rect 85020 80050 85090 80250
rect 85410 80050 85480 80250
rect 85520 80050 85590 80250
rect 85910 80050 85980 80250
rect 86020 80050 86090 80250
rect 86410 80050 86480 80250
rect 86520 80050 86590 80250
rect 86910 80050 86980 80250
rect 87020 80050 87090 80250
rect 87410 80050 87480 80250
rect 87520 80050 87590 80250
rect 87910 80050 87980 80250
rect 88020 80050 88090 80250
rect 88410 80050 88480 80250
rect 88520 80050 88590 80250
rect 88910 80050 88980 80250
rect 89020 80050 89090 80250
rect 89410 80050 89480 80250
rect 89520 80050 89590 80250
rect 89910 80050 89980 80250
rect 90020 80050 90090 80250
rect 90410 80050 90480 80250
rect 90520 80050 90590 80250
rect 90910 80050 90980 80250
rect 91020 80050 91090 80250
rect 91410 80050 91480 80250
rect 91520 80050 91590 80250
rect 91910 80050 91980 80250
rect 92020 80050 92090 80250
rect 92410 80050 92480 80250
rect 92520 80050 92590 80250
rect 92910 80050 92980 80250
rect 93020 80050 93090 80250
rect 93410 80050 93480 80250
rect 93520 80050 93590 80250
rect 93910 80050 93980 80250
rect 94020 80050 94090 80250
rect 94410 80050 94480 80250
rect 94520 80050 94590 80250
rect 94910 80050 94980 80250
rect 95020 80050 95090 80250
rect 95410 80050 95480 80250
rect 95520 80050 95590 80250
rect 95910 80050 95980 80250
rect 96020 80050 96090 80250
rect 96410 80050 96480 80250
rect 96520 80050 96590 80250
rect 96910 80050 96980 80250
rect 97020 80050 97090 80250
rect 97410 80050 97480 80250
rect 97520 80050 97590 80250
rect 97910 80050 97980 80250
rect 98020 80050 98090 80250
rect 98410 80050 98480 80250
rect 98520 80050 98590 80250
rect 98910 80050 98980 80250
rect 99020 80050 99090 80250
rect 99410 80050 99480 80250
rect 99520 80050 99590 80250
rect 99910 80050 99980 80250
rect 100020 80050 100090 80250
rect 100410 80050 100480 80250
rect -83350 79920 -83150 79990
rect -82850 79920 -82650 79990
rect -82350 79920 -82150 79990
rect -81850 79920 -81650 79990
rect -81350 79920 -81150 79990
rect -80850 79920 -80650 79990
rect -80350 79920 -80150 79990
rect -79850 79920 -79650 79990
rect -79350 79920 -79150 79990
rect -78850 79920 -78650 79990
rect -78350 79920 -78150 79990
rect -77850 79920 -77650 79990
rect -77350 79920 -77150 79990
rect -76850 79920 -76650 79990
rect -76350 79920 -76150 79990
rect -75850 79920 -75650 79990
rect -75350 79920 -75150 79990
rect -74850 79920 -74650 79990
rect -74350 79920 -74150 79990
rect -73850 79920 -73650 79990
rect -73350 79920 -73150 79990
rect -72850 79920 -72650 79990
rect -72350 79920 -72150 79990
rect -71850 79920 -71650 79990
rect -71350 79920 -71150 79990
rect -70850 79920 -70650 79990
rect -70350 79920 -70150 79990
rect -69850 79920 -69650 79990
rect -69350 79920 -69150 79990
rect -68850 79920 -68650 79990
rect -68350 79920 -68150 79990
rect -67850 79920 -67650 79990
rect -67350 79920 -67150 79990
rect -66850 79920 -66650 79990
rect -66350 79920 -66150 79990
rect -65850 79920 -65650 79990
rect -65350 79920 -65150 79990
rect -64850 79920 -64650 79990
rect -64350 79920 -64150 79990
rect -63850 79920 -63650 79990
rect -63350 79920 -63150 79990
rect -62850 79920 -62650 79990
rect -62350 79920 -62150 79990
rect -61850 79920 -61650 79990
rect -61350 79920 -61150 79990
rect -60850 79920 -60650 79990
rect -60350 79920 -60150 79990
rect -59850 79920 -59650 79990
rect -59350 79920 -59150 79990
rect -58850 79920 -58650 79990
rect -58350 79920 -58150 79990
rect -57850 79920 -57650 79990
rect -57350 79920 -57150 79990
rect -56850 79920 -56650 79990
rect -56350 79920 -56150 79990
rect -55850 79920 -55650 79990
rect -55350 79920 -55150 79990
rect -54850 79920 -54650 79990
rect -54350 79920 -54150 79990
rect -53850 79920 -53650 79990
rect -53350 79920 -53150 79990
rect -52850 79920 -52650 79990
rect -52350 79920 -52150 79990
rect -51850 79920 -51650 79990
rect -51350 79920 -51150 79990
rect -50850 79920 -50650 79990
rect -50350 79920 -50150 79990
rect -49850 79920 -49650 79990
rect -49350 79920 -49150 79990
rect -48850 79920 -48650 79990
rect -48350 79920 -48150 79990
rect -47850 79920 -47650 79990
rect -47350 79920 -47150 79990
rect -46850 79920 -46650 79990
rect -46350 79920 -46150 79990
rect -45850 79920 -45650 79990
rect -45350 79920 -45150 79990
rect -44850 79920 -44650 79990
rect -44350 79920 -44150 79990
rect -43850 79920 -43650 79990
rect -43350 79920 -43150 79990
rect -42850 79920 -42650 79990
rect -42350 79920 -42150 79990
rect -41850 79920 -41650 79990
rect -41350 79920 -41150 79990
rect -40850 79920 -40650 79990
rect -40350 79920 -40150 79990
rect -39850 79920 -39650 79990
rect -39350 79920 -39150 79990
rect -38850 79920 -38650 79990
rect -38350 79920 -38150 79990
rect -37850 79920 -37650 79990
rect -37350 79920 -37150 79990
rect -36850 79920 -36650 79990
rect -36350 79920 -36150 79990
rect -35850 79920 -35650 79990
rect -35350 79920 -35150 79990
rect -34850 79920 -34650 79990
rect -34350 79920 -34150 79990
rect -33850 79920 -33650 79990
rect -33350 79920 -33150 79990
rect -32850 79920 -32650 79990
rect -32350 79920 -32150 79990
rect -31850 79920 -31650 79990
rect -31350 79920 -31150 79990
rect -30850 79920 -30650 79990
rect -30350 79920 -30150 79990
rect -29850 79920 -29650 79990
rect -29350 79920 -29150 79990
rect -28850 79920 -28650 79990
rect -28350 79920 -28150 79990
rect -27850 79920 -27650 79990
rect -27350 79920 -27150 79990
rect -26850 79920 -26650 79990
rect -26350 79920 -26150 79990
rect -25850 79920 -25650 79990
rect -25350 79920 -25150 79990
rect -24850 79920 -24650 79990
rect -24350 79920 -24150 79990
rect -23850 79920 -23650 79990
rect -23350 79920 -23150 79990
rect -22850 79920 -22650 79990
rect -22350 79920 -22150 79990
rect -21850 79920 -21650 79990
rect -21350 79920 -21150 79990
rect -20850 79920 -20650 79990
rect -20350 79920 -20150 79990
rect -19850 79920 -19650 79990
rect -19350 79920 -19150 79990
rect -18850 79920 -18650 79990
rect -18350 79920 -18150 79990
rect -17850 79920 -17650 79990
rect -17350 79920 -17150 79990
rect -16850 79920 -16650 79990
rect -16350 79920 -16150 79990
rect -15850 79920 -15650 79990
rect -15350 79920 -15150 79990
rect -14850 79920 -14650 79990
rect -14350 79920 -14150 79990
rect -13850 79920 -13650 79990
rect -13350 79920 -13150 79990
rect -12850 79920 -12650 79990
rect -12350 79920 -12150 79990
rect -11850 79920 -11650 79990
rect -11350 79920 -11150 79990
rect -10850 79920 -10650 79990
rect -10350 79920 -10150 79990
rect -9850 79920 -9650 79990
rect -9350 79920 -9150 79990
rect -8850 79920 -8650 79990
rect -8350 79920 -8150 79990
rect -7850 79920 -7650 79990
rect -7350 79920 -7150 79990
rect -6850 79920 -6650 79990
rect -6350 79920 -6150 79990
rect -5850 79920 -5650 79990
rect -5350 79920 -5150 79990
rect -4850 79920 -4650 79990
rect -4350 79920 -4150 79990
rect -3850 79920 -3650 79990
rect -3350 79920 -3150 79990
rect -2850 79920 -2650 79990
rect -2350 79920 -2150 79990
rect -1850 79920 -1650 79990
rect -1350 79920 -1150 79990
rect -850 79920 -650 79990
rect -350 79920 -150 79990
rect 150 79920 350 79990
rect 650 79920 850 79990
rect 1150 79920 1350 79990
rect 1650 79920 1850 79990
rect 2150 79920 2350 79990
rect 2650 79920 2850 79990
rect 3150 79920 3350 79990
rect 3650 79920 3850 79990
rect 4150 79920 4350 79990
rect 4650 79920 4850 79990
rect 5150 79920 5350 79990
rect 5650 79920 5850 79990
rect 6150 79920 6350 79990
rect 6650 79920 6850 79990
rect 7150 79920 7350 79990
rect 7650 79920 7850 79990
rect 8150 79920 8350 79990
rect 8650 79920 8850 79990
rect 9150 79920 9350 79990
rect 9650 79920 9850 79990
rect 10150 79920 10350 79990
rect 10650 79920 10850 79990
rect 11150 79920 11350 79990
rect 11650 79920 11850 79990
rect 12150 79920 12350 79990
rect 12650 79920 12850 79990
rect 13150 79920 13350 79990
rect 13650 79920 13850 79990
rect 14150 79920 14350 79990
rect 14650 79920 14850 79990
rect 15150 79920 15350 79990
rect 15650 79920 15850 79990
rect 16150 79920 16350 79990
rect 16650 79920 16850 79990
rect 17150 79920 17350 79990
rect 17650 79920 17850 79990
rect 18150 79920 18350 79990
rect 18650 79920 18850 79990
rect 19150 79920 19350 79990
rect 19650 79920 19850 79990
rect 20150 79920 20350 79990
rect 20650 79920 20850 79990
rect 21150 79920 21350 79990
rect 21650 79920 21850 79990
rect 22150 79920 22350 79990
rect 22650 79920 22850 79990
rect 23150 79920 23350 79990
rect 23650 79920 23850 79990
rect 24150 79920 24350 79990
rect 24650 79920 24850 79990
rect 25150 79920 25350 79990
rect 25650 79920 25850 79990
rect 26150 79920 26350 79990
rect 26650 79920 26850 79990
rect 27150 79920 27350 79990
rect 27650 79920 27850 79990
rect 28150 79920 28350 79990
rect 28650 79920 28850 79990
rect 29150 79920 29350 79990
rect 29650 79920 29850 79990
rect 30150 79920 30350 79990
rect 30650 79920 30850 79990
rect 31150 79920 31350 79990
rect 31650 79920 31850 79990
rect 32150 79920 32350 79990
rect 32650 79920 32850 79990
rect 33150 79920 33350 79990
rect 33650 79920 33850 79990
rect 34150 79920 34350 79990
rect 34650 79920 34850 79990
rect 35150 79920 35350 79990
rect 35650 79920 35850 79990
rect 36150 79920 36350 79990
rect 36650 79920 36850 79990
rect 37150 79920 37350 79990
rect 37650 79920 37850 79990
rect 38150 79920 38350 79990
rect 38650 79920 38850 79990
rect 39150 79920 39350 79990
rect 39650 79920 39850 79990
rect 40150 79920 40350 79990
rect 40650 79920 40850 79990
rect 41150 79920 41350 79990
rect 41650 79920 41850 79990
rect 42150 79920 42350 79990
rect 42650 79920 42850 79990
rect 43150 79920 43350 79990
rect 43650 79920 43850 79990
rect 44150 79920 44350 79990
rect 44650 79920 44850 79990
rect 45150 79920 45350 79990
rect 45650 79920 45850 79990
rect 46150 79920 46350 79990
rect 46650 79920 46850 79990
rect 47150 79920 47350 79990
rect 47650 79920 47850 79990
rect 48150 79920 48350 79990
rect 48650 79920 48850 79990
rect 49150 79920 49350 79990
rect 49650 79920 49850 79990
rect 50150 79920 50350 79990
rect 50650 79920 50850 79990
rect 51150 79920 51350 79990
rect 51650 79920 51850 79990
rect 52150 79920 52350 79990
rect 52650 79920 52850 79990
rect 53150 79920 53350 79990
rect 53650 79920 53850 79990
rect 54150 79920 54350 79990
rect 54650 79920 54850 79990
rect 55150 79920 55350 79990
rect 55650 79920 55850 79990
rect 56150 79920 56350 79990
rect 56650 79920 56850 79990
rect 57150 79920 57350 79990
rect 57650 79920 57850 79990
rect 58150 79920 58350 79990
rect 58650 79920 58850 79990
rect 59150 79920 59350 79990
rect 59650 79920 59850 79990
rect 60150 79920 60350 79990
rect 60650 79920 60850 79990
rect 61150 79920 61350 79990
rect 61650 79920 61850 79990
rect 62150 79920 62350 79990
rect 62650 79920 62850 79990
rect 63150 79920 63350 79990
rect 63650 79920 63850 79990
rect 64150 79920 64350 79990
rect 64650 79920 64850 79990
rect 65150 79920 65350 79990
rect 65650 79920 65850 79990
rect 66150 79920 66350 79990
rect 66650 79920 66850 79990
rect 67150 79920 67350 79990
rect 67650 79920 67850 79990
rect 68150 79920 68350 79990
rect 68650 79920 68850 79990
rect 69150 79920 69350 79990
rect 69650 79920 69850 79990
rect 70150 79920 70350 79990
rect 70650 79920 70850 79990
rect 71150 79920 71350 79990
rect 71650 79920 71850 79990
rect 72150 79920 72350 79990
rect 72650 79920 72850 79990
rect 73150 79920 73350 79990
rect 73650 79920 73850 79990
rect 74150 79920 74350 79990
rect 74650 79920 74850 79990
rect 75150 79920 75350 79990
rect 75650 79920 75850 79990
rect 76150 79920 76350 79990
rect 76650 79920 76850 79990
rect 77150 79920 77350 79990
rect 77650 79920 77850 79990
rect 78150 79920 78350 79990
rect 78650 79920 78850 79990
rect 79150 79920 79350 79990
rect 79650 79920 79850 79990
rect 80150 79920 80350 79990
rect 80650 79920 80850 79990
rect 81150 79920 81350 79990
rect 81650 79920 81850 79990
rect 82150 79920 82350 79990
rect 82650 79920 82850 79990
rect 83150 79920 83350 79990
rect 83650 79920 83850 79990
rect 84150 79920 84350 79990
rect 84650 79920 84850 79990
rect 85150 79920 85350 79990
rect 85650 79920 85850 79990
rect 86150 79920 86350 79990
rect 86650 79920 86850 79990
rect 87150 79920 87350 79990
rect 87650 79920 87850 79990
rect 88150 79920 88350 79990
rect 88650 79920 88850 79990
rect 89150 79920 89350 79990
rect 89650 79920 89850 79990
rect 90150 79920 90350 79990
rect 90650 79920 90850 79990
rect 91150 79920 91350 79990
rect 91650 79920 91850 79990
rect 92150 79920 92350 79990
rect 92650 79920 92850 79990
rect 93150 79920 93350 79990
rect 93650 79920 93850 79990
rect 94150 79920 94350 79990
rect 94650 79920 94850 79990
rect 95150 79920 95350 79990
rect 95650 79920 95850 79990
rect 96150 79920 96350 79990
rect 96650 79920 96850 79990
rect 97150 79920 97350 79990
rect 97650 79920 97850 79990
rect 98150 79920 98350 79990
rect 98650 79920 98850 79990
rect 99150 79920 99350 79990
rect 99650 79920 99850 79990
rect 100150 79920 100350 79990
rect 22650 -29190 22850 -29120
rect 23150 -29190 23350 -29120
rect 22520 -29450 22590 -29250
rect 22910 -29450 22980 -29250
rect 23020 -29450 23090 -29250
rect 23410 -29450 23480 -29250
rect 22650 -29580 22850 -29510
rect 23150 -29580 23350 -29510
rect 24200 -33200 25800 -30700
rect 31000 -33200 32600 -30700
<< metal2 >>
rect -83360 82880 -83140 82900
rect -83360 82810 -83350 82880
rect -83150 82810 -83140 82880
rect -83360 82760 -83140 82810
rect -82860 82880 -82640 82900
rect -82860 82810 -82850 82880
rect -82650 82810 -82640 82880
rect -82860 82760 -82640 82810
rect -82360 82880 -82140 82900
rect -82360 82810 -82350 82880
rect -82150 82810 -82140 82880
rect -82360 82760 -82140 82810
rect -81860 82880 -81640 82900
rect -81860 82810 -81850 82880
rect -81650 82810 -81640 82880
rect -81860 82760 -81640 82810
rect -81360 82880 -81140 82900
rect -81360 82810 -81350 82880
rect -81150 82810 -81140 82880
rect -81360 82760 -81140 82810
rect -80860 82880 -80640 82900
rect -80860 82810 -80850 82880
rect -80650 82810 -80640 82880
rect -80860 82760 -80640 82810
rect -80360 82880 -80140 82900
rect -80360 82810 -80350 82880
rect -80150 82810 -80140 82880
rect -80360 82760 -80140 82810
rect -79860 82880 -79640 82900
rect -79860 82810 -79850 82880
rect -79650 82810 -79640 82880
rect -79860 82760 -79640 82810
rect -79360 82880 -79140 82900
rect -79360 82810 -79350 82880
rect -79150 82810 -79140 82880
rect -79360 82760 -79140 82810
rect -78860 82880 -78640 82900
rect -78860 82810 -78850 82880
rect -78650 82810 -78640 82880
rect -78860 82760 -78640 82810
rect -78360 82880 -78140 82900
rect -78360 82810 -78350 82880
rect -78150 82810 -78140 82880
rect -78360 82760 -78140 82810
rect -77860 82880 -77640 82900
rect -77860 82810 -77850 82880
rect -77650 82810 -77640 82880
rect -77860 82760 -77640 82810
rect -77360 82880 -77140 82900
rect -77360 82810 -77350 82880
rect -77150 82810 -77140 82880
rect -77360 82760 -77140 82810
rect -76860 82880 -76640 82900
rect -76860 82810 -76850 82880
rect -76650 82810 -76640 82880
rect -76860 82760 -76640 82810
rect -76360 82880 -76140 82900
rect -76360 82810 -76350 82880
rect -76150 82810 -76140 82880
rect -76360 82760 -76140 82810
rect -75860 82880 -75640 82900
rect -75860 82810 -75850 82880
rect -75650 82810 -75640 82880
rect -75860 82760 -75640 82810
rect -75360 82880 -75140 82900
rect -75360 82810 -75350 82880
rect -75150 82810 -75140 82880
rect -75360 82760 -75140 82810
rect -74860 82880 -74640 82900
rect -74860 82810 -74850 82880
rect -74650 82810 -74640 82880
rect -74860 82760 -74640 82810
rect -74360 82880 -74140 82900
rect -74360 82810 -74350 82880
rect -74150 82810 -74140 82880
rect -74360 82760 -74140 82810
rect -73860 82880 -73640 82900
rect -73860 82810 -73850 82880
rect -73650 82810 -73640 82880
rect -73860 82760 -73640 82810
rect -73360 82880 -73140 82900
rect -73360 82810 -73350 82880
rect -73150 82810 -73140 82880
rect -73360 82760 -73140 82810
rect -72860 82880 -72640 82900
rect -72860 82810 -72850 82880
rect -72650 82810 -72640 82880
rect -72860 82760 -72640 82810
rect -72360 82880 -72140 82900
rect -72360 82810 -72350 82880
rect -72150 82810 -72140 82880
rect -72360 82760 -72140 82810
rect -71860 82880 -71640 82900
rect -71860 82810 -71850 82880
rect -71650 82810 -71640 82880
rect -71860 82760 -71640 82810
rect -71360 82880 -71140 82900
rect -71360 82810 -71350 82880
rect -71150 82810 -71140 82880
rect -71360 82760 -71140 82810
rect -70860 82880 -70640 82900
rect -70860 82810 -70850 82880
rect -70650 82810 -70640 82880
rect -70860 82760 -70640 82810
rect -70360 82880 -70140 82900
rect -70360 82810 -70350 82880
rect -70150 82810 -70140 82880
rect -70360 82760 -70140 82810
rect -69860 82880 -69640 82900
rect -69860 82810 -69850 82880
rect -69650 82810 -69640 82880
rect -69860 82760 -69640 82810
rect -69360 82880 -69140 82900
rect -69360 82810 -69350 82880
rect -69150 82810 -69140 82880
rect -69360 82760 -69140 82810
rect -68860 82880 -68640 82900
rect -68860 82810 -68850 82880
rect -68650 82810 -68640 82880
rect -68860 82760 -68640 82810
rect -68360 82880 -68140 82900
rect -68360 82810 -68350 82880
rect -68150 82810 -68140 82880
rect -68360 82760 -68140 82810
rect -67860 82880 -67640 82900
rect -67860 82810 -67850 82880
rect -67650 82810 -67640 82880
rect -67860 82760 -67640 82810
rect -67360 82880 -67140 82900
rect -67360 82810 -67350 82880
rect -67150 82810 -67140 82880
rect -67360 82760 -67140 82810
rect -66860 82880 -66640 82900
rect -66860 82810 -66850 82880
rect -66650 82810 -66640 82880
rect -66860 82760 -66640 82810
rect -66360 82880 -66140 82900
rect -66360 82810 -66350 82880
rect -66150 82810 -66140 82880
rect -66360 82760 -66140 82810
rect -65860 82880 -65640 82900
rect -65860 82810 -65850 82880
rect -65650 82810 -65640 82880
rect -65860 82760 -65640 82810
rect -65360 82880 -65140 82900
rect -65360 82810 -65350 82880
rect -65150 82810 -65140 82880
rect -65360 82760 -65140 82810
rect -64860 82880 -64640 82900
rect -64860 82810 -64850 82880
rect -64650 82810 -64640 82880
rect -64860 82760 -64640 82810
rect -64360 82880 -64140 82900
rect -64360 82810 -64350 82880
rect -64150 82810 -64140 82880
rect -64360 82760 -64140 82810
rect -63860 82880 -63640 82900
rect -63860 82810 -63850 82880
rect -63650 82810 -63640 82880
rect -63860 82760 -63640 82810
rect -63360 82880 -63140 82900
rect -63360 82810 -63350 82880
rect -63150 82810 -63140 82880
rect -63360 82760 -63140 82810
rect -62860 82880 -62640 82900
rect -62860 82810 -62850 82880
rect -62650 82810 -62640 82880
rect -62860 82760 -62640 82810
rect -62360 82880 -62140 82900
rect -62360 82810 -62350 82880
rect -62150 82810 -62140 82880
rect -62360 82760 -62140 82810
rect -61860 82880 -61640 82900
rect -61860 82810 -61850 82880
rect -61650 82810 -61640 82880
rect -61860 82760 -61640 82810
rect -61360 82880 -61140 82900
rect -61360 82810 -61350 82880
rect -61150 82810 -61140 82880
rect -61360 82760 -61140 82810
rect -60860 82880 -60640 82900
rect -60860 82810 -60850 82880
rect -60650 82810 -60640 82880
rect -60860 82760 -60640 82810
rect -60360 82880 -60140 82900
rect -60360 82810 -60350 82880
rect -60150 82810 -60140 82880
rect -60360 82760 -60140 82810
rect -59860 82880 -59640 82900
rect -59860 82810 -59850 82880
rect -59650 82810 -59640 82880
rect -59860 82760 -59640 82810
rect -59360 82880 -59140 82900
rect -59360 82810 -59350 82880
rect -59150 82810 -59140 82880
rect -59360 82760 -59140 82810
rect -58860 82880 -58640 82900
rect -58860 82810 -58850 82880
rect -58650 82810 -58640 82880
rect -58860 82760 -58640 82810
rect -58360 82880 -58140 82900
rect -58360 82810 -58350 82880
rect -58150 82810 -58140 82880
rect -58360 82760 -58140 82810
rect -57860 82880 -57640 82900
rect -57860 82810 -57850 82880
rect -57650 82810 -57640 82880
rect -57860 82760 -57640 82810
rect -57360 82880 -57140 82900
rect -57360 82810 -57350 82880
rect -57150 82810 -57140 82880
rect -57360 82760 -57140 82810
rect -56860 82880 -56640 82900
rect -56860 82810 -56850 82880
rect -56650 82810 -56640 82880
rect -56860 82760 -56640 82810
rect -56360 82880 -56140 82900
rect -56360 82810 -56350 82880
rect -56150 82810 -56140 82880
rect -56360 82760 -56140 82810
rect -55860 82880 -55640 82900
rect -55860 82810 -55850 82880
rect -55650 82810 -55640 82880
rect -55860 82760 -55640 82810
rect -55360 82880 -55140 82900
rect -55360 82810 -55350 82880
rect -55150 82810 -55140 82880
rect -55360 82760 -55140 82810
rect -54860 82880 -54640 82900
rect -54860 82810 -54850 82880
rect -54650 82810 -54640 82880
rect -54860 82760 -54640 82810
rect -54360 82880 -54140 82900
rect -54360 82810 -54350 82880
rect -54150 82810 -54140 82880
rect -54360 82760 -54140 82810
rect -53860 82880 -53640 82900
rect -53860 82810 -53850 82880
rect -53650 82810 -53640 82880
rect -53860 82760 -53640 82810
rect -53360 82880 -53140 82900
rect -53360 82810 -53350 82880
rect -53150 82810 -53140 82880
rect -53360 82760 -53140 82810
rect -52860 82880 -52640 82900
rect -52860 82810 -52850 82880
rect -52650 82810 -52640 82880
rect -52860 82760 -52640 82810
rect -52360 82880 -52140 82900
rect -52360 82810 -52350 82880
rect -52150 82810 -52140 82880
rect -52360 82760 -52140 82810
rect -51860 82880 -51640 82900
rect -51860 82810 -51850 82880
rect -51650 82810 -51640 82880
rect -51860 82760 -51640 82810
rect -51360 82880 -51140 82900
rect -51360 82810 -51350 82880
rect -51150 82810 -51140 82880
rect -51360 82760 -51140 82810
rect -50860 82880 -50640 82900
rect -50860 82810 -50850 82880
rect -50650 82810 -50640 82880
rect -50860 82760 -50640 82810
rect -50360 82880 -50140 82900
rect -50360 82810 -50350 82880
rect -50150 82810 -50140 82880
rect -50360 82760 -50140 82810
rect -49860 82880 -49640 82900
rect -49860 82810 -49850 82880
rect -49650 82810 -49640 82880
rect -49860 82760 -49640 82810
rect -49360 82880 -49140 82900
rect -49360 82810 -49350 82880
rect -49150 82810 -49140 82880
rect -49360 82760 -49140 82810
rect -48860 82880 -48640 82900
rect -48860 82810 -48850 82880
rect -48650 82810 -48640 82880
rect -48860 82760 -48640 82810
rect -48360 82880 -48140 82900
rect -48360 82810 -48350 82880
rect -48150 82810 -48140 82880
rect -48360 82760 -48140 82810
rect -47860 82880 -47640 82900
rect -47860 82810 -47850 82880
rect -47650 82810 -47640 82880
rect -47860 82760 -47640 82810
rect -47360 82880 -47140 82900
rect -47360 82810 -47350 82880
rect -47150 82810 -47140 82880
rect -47360 82760 -47140 82810
rect -46860 82880 -46640 82900
rect -46860 82810 -46850 82880
rect -46650 82810 -46640 82880
rect -46860 82760 -46640 82810
rect -46360 82880 -46140 82900
rect -46360 82810 -46350 82880
rect -46150 82810 -46140 82880
rect -46360 82760 -46140 82810
rect -45860 82880 -45640 82900
rect -45860 82810 -45850 82880
rect -45650 82810 -45640 82880
rect -45860 82760 -45640 82810
rect -45360 82880 -45140 82900
rect -45360 82810 -45350 82880
rect -45150 82810 -45140 82880
rect -45360 82760 -45140 82810
rect -44860 82880 -44640 82900
rect -44860 82810 -44850 82880
rect -44650 82810 -44640 82880
rect -44860 82760 -44640 82810
rect -44360 82880 -44140 82900
rect -44360 82810 -44350 82880
rect -44150 82810 -44140 82880
rect -44360 82760 -44140 82810
rect -43860 82880 -43640 82900
rect -43860 82810 -43850 82880
rect -43650 82810 -43640 82880
rect -43860 82760 -43640 82810
rect -43360 82880 -43140 82900
rect -43360 82810 -43350 82880
rect -43150 82810 -43140 82880
rect -43360 82760 -43140 82810
rect -42860 82880 -42640 82900
rect -42860 82810 -42850 82880
rect -42650 82810 -42640 82880
rect -42860 82760 -42640 82810
rect -42360 82880 -42140 82900
rect -42360 82810 -42350 82880
rect -42150 82810 -42140 82880
rect -42360 82760 -42140 82810
rect -41860 82880 -41640 82900
rect -41860 82810 -41850 82880
rect -41650 82810 -41640 82880
rect -41860 82760 -41640 82810
rect -41360 82880 -41140 82900
rect -41360 82810 -41350 82880
rect -41150 82810 -41140 82880
rect -41360 82760 -41140 82810
rect -40860 82880 -40640 82900
rect -40860 82810 -40850 82880
rect -40650 82810 -40640 82880
rect -40860 82760 -40640 82810
rect -40360 82880 -40140 82900
rect -40360 82810 -40350 82880
rect -40150 82810 -40140 82880
rect -40360 82760 -40140 82810
rect -39860 82880 -39640 82900
rect -39860 82810 -39850 82880
rect -39650 82810 -39640 82880
rect -39860 82760 -39640 82810
rect -39360 82880 -39140 82900
rect -39360 82810 -39350 82880
rect -39150 82810 -39140 82880
rect -39360 82760 -39140 82810
rect -38860 82880 -38640 82900
rect -38860 82810 -38850 82880
rect -38650 82810 -38640 82880
rect -38860 82760 -38640 82810
rect -38360 82880 -38140 82900
rect -38360 82810 -38350 82880
rect -38150 82810 -38140 82880
rect -38360 82760 -38140 82810
rect -37860 82880 -37640 82900
rect -37860 82810 -37850 82880
rect -37650 82810 -37640 82880
rect -37860 82760 -37640 82810
rect -37360 82880 -37140 82900
rect -37360 82810 -37350 82880
rect -37150 82810 -37140 82880
rect -37360 82760 -37140 82810
rect -36860 82880 -36640 82900
rect -36860 82810 -36850 82880
rect -36650 82810 -36640 82880
rect -36860 82760 -36640 82810
rect -36360 82880 -36140 82900
rect -36360 82810 -36350 82880
rect -36150 82810 -36140 82880
rect -36360 82760 -36140 82810
rect -35860 82880 -35640 82900
rect -35860 82810 -35850 82880
rect -35650 82810 -35640 82880
rect -35860 82760 -35640 82810
rect -35360 82880 -35140 82900
rect -35360 82810 -35350 82880
rect -35150 82810 -35140 82880
rect -35360 82760 -35140 82810
rect -34860 82880 -34640 82900
rect -34860 82810 -34850 82880
rect -34650 82810 -34640 82880
rect -34860 82760 -34640 82810
rect -34360 82880 -34140 82900
rect -34360 82810 -34350 82880
rect -34150 82810 -34140 82880
rect -34360 82760 -34140 82810
rect -33860 82880 -33640 82900
rect -33860 82810 -33850 82880
rect -33650 82810 -33640 82880
rect -33860 82760 -33640 82810
rect -33360 82880 -33140 82900
rect -33360 82810 -33350 82880
rect -33150 82810 -33140 82880
rect -33360 82760 -33140 82810
rect -32860 82880 -32640 82900
rect -32860 82810 -32850 82880
rect -32650 82810 -32640 82880
rect -32860 82760 -32640 82810
rect -32360 82880 -32140 82900
rect -32360 82810 -32350 82880
rect -32150 82810 -32140 82880
rect -32360 82760 -32140 82810
rect -31860 82880 -31640 82900
rect -31860 82810 -31850 82880
rect -31650 82810 -31640 82880
rect -31860 82760 -31640 82810
rect -31360 82880 -31140 82900
rect -31360 82810 -31350 82880
rect -31150 82810 -31140 82880
rect -31360 82760 -31140 82810
rect -30860 82880 -30640 82900
rect -30860 82810 -30850 82880
rect -30650 82810 -30640 82880
rect -30860 82760 -30640 82810
rect -30360 82880 -30140 82900
rect -30360 82810 -30350 82880
rect -30150 82810 -30140 82880
rect -30360 82760 -30140 82810
rect -29860 82880 -29640 82900
rect -29860 82810 -29850 82880
rect -29650 82810 -29640 82880
rect -29860 82760 -29640 82810
rect -29360 82880 -29140 82900
rect -29360 82810 -29350 82880
rect -29150 82810 -29140 82880
rect -29360 82760 -29140 82810
rect -28860 82880 -28640 82900
rect -28860 82810 -28850 82880
rect -28650 82810 -28640 82880
rect -28860 82760 -28640 82810
rect -28360 82880 -28140 82900
rect -28360 82810 -28350 82880
rect -28150 82810 -28140 82880
rect -28360 82760 -28140 82810
rect -27860 82880 -27640 82900
rect -27860 82810 -27850 82880
rect -27650 82810 -27640 82880
rect -27860 82760 -27640 82810
rect -27360 82880 -27140 82900
rect -27360 82810 -27350 82880
rect -27150 82810 -27140 82880
rect -27360 82760 -27140 82810
rect -26860 82880 -26640 82900
rect -26860 82810 -26850 82880
rect -26650 82810 -26640 82880
rect -26860 82760 -26640 82810
rect -26360 82880 -26140 82900
rect -26360 82810 -26350 82880
rect -26150 82810 -26140 82880
rect -26360 82760 -26140 82810
rect -25860 82880 -25640 82900
rect -25860 82810 -25850 82880
rect -25650 82810 -25640 82880
rect -25860 82760 -25640 82810
rect -25360 82880 -25140 82900
rect -25360 82810 -25350 82880
rect -25150 82810 -25140 82880
rect -25360 82760 -25140 82810
rect -24860 82880 -24640 82900
rect -24860 82810 -24850 82880
rect -24650 82810 -24640 82880
rect -24860 82760 -24640 82810
rect -24360 82880 -24140 82900
rect -24360 82810 -24350 82880
rect -24150 82810 -24140 82880
rect -24360 82760 -24140 82810
rect -23860 82880 -23640 82900
rect -23860 82810 -23850 82880
rect -23650 82810 -23640 82880
rect -23860 82760 -23640 82810
rect -23360 82880 -23140 82900
rect -23360 82810 -23350 82880
rect -23150 82810 -23140 82880
rect -23360 82760 -23140 82810
rect -22860 82880 -22640 82900
rect -22860 82810 -22850 82880
rect -22650 82810 -22640 82880
rect -22860 82760 -22640 82810
rect -22360 82880 -22140 82900
rect -22360 82810 -22350 82880
rect -22150 82810 -22140 82880
rect -22360 82760 -22140 82810
rect -21860 82880 -21640 82900
rect -21860 82810 -21850 82880
rect -21650 82810 -21640 82880
rect -21860 82760 -21640 82810
rect -21360 82880 -21140 82900
rect -21360 82810 -21350 82880
rect -21150 82810 -21140 82880
rect -21360 82760 -21140 82810
rect -20860 82880 -20640 82900
rect -20860 82810 -20850 82880
rect -20650 82810 -20640 82880
rect -20860 82760 -20640 82810
rect -20360 82880 -20140 82900
rect -20360 82810 -20350 82880
rect -20150 82810 -20140 82880
rect -20360 82760 -20140 82810
rect -19860 82880 -19640 82900
rect -19860 82810 -19850 82880
rect -19650 82810 -19640 82880
rect -19860 82760 -19640 82810
rect -19360 82880 -19140 82900
rect -19360 82810 -19350 82880
rect -19150 82810 -19140 82880
rect -19360 82760 -19140 82810
rect -18860 82880 -18640 82900
rect -18860 82810 -18850 82880
rect -18650 82810 -18640 82880
rect -18860 82760 -18640 82810
rect -18360 82880 -18140 82900
rect -18360 82810 -18350 82880
rect -18150 82810 -18140 82880
rect -18360 82760 -18140 82810
rect -17860 82880 -17640 82900
rect -17860 82810 -17850 82880
rect -17650 82810 -17640 82880
rect -17860 82760 -17640 82810
rect -17360 82880 -17140 82900
rect -17360 82810 -17350 82880
rect -17150 82810 -17140 82880
rect -17360 82760 -17140 82810
rect -16860 82880 -16640 82900
rect -16860 82810 -16850 82880
rect -16650 82810 -16640 82880
rect -16860 82760 -16640 82810
rect -16360 82880 -16140 82900
rect -16360 82810 -16350 82880
rect -16150 82810 -16140 82880
rect -16360 82760 -16140 82810
rect -15860 82880 -15640 82900
rect -15860 82810 -15850 82880
rect -15650 82810 -15640 82880
rect -15860 82760 -15640 82810
rect -15360 82880 -15140 82900
rect -15360 82810 -15350 82880
rect -15150 82810 -15140 82880
rect -15360 82760 -15140 82810
rect -14860 82880 -14640 82900
rect -14860 82810 -14850 82880
rect -14650 82810 -14640 82880
rect -14860 82760 -14640 82810
rect -14360 82880 -14140 82900
rect -14360 82810 -14350 82880
rect -14150 82810 -14140 82880
rect -14360 82760 -14140 82810
rect -13860 82880 -13640 82900
rect -13860 82810 -13850 82880
rect -13650 82810 -13640 82880
rect -13860 82760 -13640 82810
rect -13360 82880 -13140 82900
rect -13360 82810 -13350 82880
rect -13150 82810 -13140 82880
rect -13360 82760 -13140 82810
rect -12860 82880 -12640 82900
rect -12860 82810 -12850 82880
rect -12650 82810 -12640 82880
rect -12860 82760 -12640 82810
rect -12360 82880 -12140 82900
rect -12360 82810 -12350 82880
rect -12150 82810 -12140 82880
rect -12360 82760 -12140 82810
rect -11860 82880 -11640 82900
rect -11860 82810 -11850 82880
rect -11650 82810 -11640 82880
rect -11860 82760 -11640 82810
rect -11360 82880 -11140 82900
rect -11360 82810 -11350 82880
rect -11150 82810 -11140 82880
rect -11360 82760 -11140 82810
rect -10860 82880 -10640 82900
rect -10860 82810 -10850 82880
rect -10650 82810 -10640 82880
rect -10860 82760 -10640 82810
rect -10360 82880 -10140 82900
rect -10360 82810 -10350 82880
rect -10150 82810 -10140 82880
rect -10360 82760 -10140 82810
rect -9860 82880 -9640 82900
rect -9860 82810 -9850 82880
rect -9650 82810 -9640 82880
rect -9860 82760 -9640 82810
rect -9360 82880 -9140 82900
rect -9360 82810 -9350 82880
rect -9150 82810 -9140 82880
rect -9360 82760 -9140 82810
rect -8860 82880 -8640 82900
rect -8860 82810 -8850 82880
rect -8650 82810 -8640 82880
rect -8860 82760 -8640 82810
rect -8360 82880 -8140 82900
rect -8360 82810 -8350 82880
rect -8150 82810 -8140 82880
rect -8360 82760 -8140 82810
rect -7860 82880 -7640 82900
rect -7860 82810 -7850 82880
rect -7650 82810 -7640 82880
rect -7860 82760 -7640 82810
rect -7360 82880 -7140 82900
rect -7360 82810 -7350 82880
rect -7150 82810 -7140 82880
rect -7360 82760 -7140 82810
rect -6860 82880 -6640 82900
rect -6860 82810 -6850 82880
rect -6650 82810 -6640 82880
rect -6860 82760 -6640 82810
rect -6360 82880 -6140 82900
rect -6360 82810 -6350 82880
rect -6150 82810 -6140 82880
rect -6360 82760 -6140 82810
rect -5860 82880 -5640 82900
rect -5860 82810 -5850 82880
rect -5650 82810 -5640 82880
rect -5860 82760 -5640 82810
rect -5360 82880 -5140 82900
rect -5360 82810 -5350 82880
rect -5150 82810 -5140 82880
rect -5360 82760 -5140 82810
rect -4860 82880 -4640 82900
rect -4860 82810 -4850 82880
rect -4650 82810 -4640 82880
rect -4860 82760 -4640 82810
rect -4360 82880 -4140 82900
rect -4360 82810 -4350 82880
rect -4150 82810 -4140 82880
rect -4360 82760 -4140 82810
rect -3860 82880 -3640 82900
rect -3860 82810 -3850 82880
rect -3650 82810 -3640 82880
rect -3860 82760 -3640 82810
rect -3360 82880 -3140 82900
rect -3360 82810 -3350 82880
rect -3150 82810 -3140 82880
rect -3360 82760 -3140 82810
rect -2860 82880 -2640 82900
rect -2860 82810 -2850 82880
rect -2650 82810 -2640 82880
rect -2860 82760 -2640 82810
rect -2360 82880 -2140 82900
rect -2360 82810 -2350 82880
rect -2150 82810 -2140 82880
rect -2360 82760 -2140 82810
rect -1860 82880 -1640 82900
rect -1860 82810 -1850 82880
rect -1650 82810 -1640 82880
rect -1860 82760 -1640 82810
rect -1360 82880 -1140 82900
rect -1360 82810 -1350 82880
rect -1150 82810 -1140 82880
rect -1360 82760 -1140 82810
rect -860 82880 -640 82900
rect -860 82810 -850 82880
rect -650 82810 -640 82880
rect -860 82760 -640 82810
rect -360 82880 -140 82900
rect -360 82810 -350 82880
rect -150 82810 -140 82880
rect -360 82760 -140 82810
rect 140 82880 360 82900
rect 140 82810 150 82880
rect 350 82810 360 82880
rect 140 82760 360 82810
rect 640 82880 860 82900
rect 640 82810 650 82880
rect 850 82810 860 82880
rect 640 82760 860 82810
rect 1140 82880 1360 82900
rect 1140 82810 1150 82880
rect 1350 82810 1360 82880
rect 1140 82760 1360 82810
rect 1640 82880 1860 82900
rect 1640 82810 1650 82880
rect 1850 82810 1860 82880
rect 1640 82760 1860 82810
rect 2140 82880 2360 82900
rect 2140 82810 2150 82880
rect 2350 82810 2360 82880
rect 2140 82760 2360 82810
rect 2640 82880 2860 82900
rect 2640 82810 2650 82880
rect 2850 82810 2860 82880
rect 2640 82760 2860 82810
rect 3140 82880 3360 82900
rect 3140 82810 3150 82880
rect 3350 82810 3360 82880
rect 3140 82760 3360 82810
rect 3640 82880 3860 82900
rect 3640 82810 3650 82880
rect 3850 82810 3860 82880
rect 3640 82760 3860 82810
rect 4140 82880 4360 82900
rect 4140 82810 4150 82880
rect 4350 82810 4360 82880
rect 4140 82760 4360 82810
rect 4640 82880 4860 82900
rect 4640 82810 4650 82880
rect 4850 82810 4860 82880
rect 4640 82760 4860 82810
rect 5140 82880 5360 82900
rect 5140 82810 5150 82880
rect 5350 82810 5360 82880
rect 5140 82760 5360 82810
rect 5640 82880 5860 82900
rect 5640 82810 5650 82880
rect 5850 82810 5860 82880
rect 5640 82760 5860 82810
rect 6140 82880 6360 82900
rect 6140 82810 6150 82880
rect 6350 82810 6360 82880
rect 6140 82760 6360 82810
rect 6640 82880 6860 82900
rect 6640 82810 6650 82880
rect 6850 82810 6860 82880
rect 6640 82760 6860 82810
rect 7140 82880 7360 82900
rect 7140 82810 7150 82880
rect 7350 82810 7360 82880
rect 7140 82760 7360 82810
rect 7640 82880 7860 82900
rect 7640 82810 7650 82880
rect 7850 82810 7860 82880
rect 7640 82760 7860 82810
rect 8140 82880 8360 82900
rect 8140 82810 8150 82880
rect 8350 82810 8360 82880
rect 8140 82760 8360 82810
rect 8640 82880 8860 82900
rect 8640 82810 8650 82880
rect 8850 82810 8860 82880
rect 8640 82760 8860 82810
rect 9140 82880 9360 82900
rect 9140 82810 9150 82880
rect 9350 82810 9360 82880
rect 9140 82760 9360 82810
rect 9640 82880 9860 82900
rect 9640 82810 9650 82880
rect 9850 82810 9860 82880
rect 9640 82760 9860 82810
rect 10140 82880 10360 82900
rect 10140 82810 10150 82880
rect 10350 82810 10360 82880
rect 10140 82760 10360 82810
rect 10640 82880 10860 82900
rect 10640 82810 10650 82880
rect 10850 82810 10860 82880
rect 10640 82760 10860 82810
rect 11140 82880 11360 82900
rect 11140 82810 11150 82880
rect 11350 82810 11360 82880
rect 11140 82760 11360 82810
rect 11640 82880 11860 82900
rect 11640 82810 11650 82880
rect 11850 82810 11860 82880
rect 11640 82760 11860 82810
rect 12140 82880 12360 82900
rect 12140 82810 12150 82880
rect 12350 82810 12360 82880
rect 12140 82760 12360 82810
rect 12640 82880 12860 82900
rect 12640 82810 12650 82880
rect 12850 82810 12860 82880
rect 12640 82760 12860 82810
rect 13140 82880 13360 82900
rect 13140 82810 13150 82880
rect 13350 82810 13360 82880
rect 13140 82760 13360 82810
rect 13640 82880 13860 82900
rect 13640 82810 13650 82880
rect 13850 82810 13860 82880
rect 13640 82760 13860 82810
rect 14140 82880 14360 82900
rect 14140 82810 14150 82880
rect 14350 82810 14360 82880
rect 14140 82760 14360 82810
rect 14640 82880 14860 82900
rect 14640 82810 14650 82880
rect 14850 82810 14860 82880
rect 14640 82760 14860 82810
rect 15140 82880 15360 82900
rect 15140 82810 15150 82880
rect 15350 82810 15360 82880
rect 15140 82760 15360 82810
rect 15640 82880 15860 82900
rect 15640 82810 15650 82880
rect 15850 82810 15860 82880
rect 15640 82760 15860 82810
rect 16140 82880 16360 82900
rect 16140 82810 16150 82880
rect 16350 82810 16360 82880
rect 16140 82760 16360 82810
rect 16640 82880 16860 82900
rect 16640 82810 16650 82880
rect 16850 82810 16860 82880
rect 16640 82760 16860 82810
rect 17140 82880 17360 82900
rect 17140 82810 17150 82880
rect 17350 82810 17360 82880
rect 17140 82760 17360 82810
rect 17640 82880 17860 82900
rect 17640 82810 17650 82880
rect 17850 82810 17860 82880
rect 17640 82760 17860 82810
rect 18140 82880 18360 82900
rect 18140 82810 18150 82880
rect 18350 82810 18360 82880
rect 18140 82760 18360 82810
rect 18640 82880 18860 82900
rect 18640 82810 18650 82880
rect 18850 82810 18860 82880
rect 18640 82760 18860 82810
rect 19140 82880 19360 82900
rect 19140 82810 19150 82880
rect 19350 82810 19360 82880
rect 19140 82760 19360 82810
rect 19640 82880 19860 82900
rect 19640 82810 19650 82880
rect 19850 82810 19860 82880
rect 19640 82760 19860 82810
rect 20140 82880 20360 82900
rect 20140 82810 20150 82880
rect 20350 82810 20360 82880
rect 20140 82760 20360 82810
rect 20640 82880 20860 82900
rect 20640 82810 20650 82880
rect 20850 82810 20860 82880
rect 20640 82760 20860 82810
rect 21140 82880 21360 82900
rect 21140 82810 21150 82880
rect 21350 82810 21360 82880
rect 21140 82760 21360 82810
rect 21640 82880 21860 82900
rect 21640 82810 21650 82880
rect 21850 82810 21860 82880
rect 21640 82760 21860 82810
rect 22140 82880 22360 82900
rect 22140 82810 22150 82880
rect 22350 82810 22360 82880
rect 22140 82760 22360 82810
rect 22640 82880 22860 82900
rect 22640 82810 22650 82880
rect 22850 82810 22860 82880
rect 22640 82760 22860 82810
rect 23140 82880 23360 82900
rect 23140 82810 23150 82880
rect 23350 82810 23360 82880
rect 23140 82760 23360 82810
rect 23640 82880 23860 82900
rect 23640 82810 23650 82880
rect 23850 82810 23860 82880
rect 23640 82760 23860 82810
rect 24140 82880 24360 82900
rect 24140 82810 24150 82880
rect 24350 82810 24360 82880
rect 24140 82760 24360 82810
rect 24640 82880 24860 82900
rect 24640 82810 24650 82880
rect 24850 82810 24860 82880
rect 24640 82760 24860 82810
rect 25140 82880 25360 82900
rect 25140 82810 25150 82880
rect 25350 82810 25360 82880
rect 25140 82760 25360 82810
rect 25640 82880 25860 82900
rect 25640 82810 25650 82880
rect 25850 82810 25860 82880
rect 25640 82760 25860 82810
rect 26140 82880 26360 82900
rect 26140 82810 26150 82880
rect 26350 82810 26360 82880
rect 26140 82760 26360 82810
rect 26640 82880 26860 82900
rect 26640 82810 26650 82880
rect 26850 82810 26860 82880
rect 26640 82760 26860 82810
rect 27140 82880 27360 82900
rect 27140 82810 27150 82880
rect 27350 82810 27360 82880
rect 27140 82760 27360 82810
rect 27640 82880 27860 82900
rect 27640 82810 27650 82880
rect 27850 82810 27860 82880
rect 27640 82760 27860 82810
rect 28140 82880 28360 82900
rect 28140 82810 28150 82880
rect 28350 82810 28360 82880
rect 28140 82760 28360 82810
rect 28640 82880 28860 82900
rect 28640 82810 28650 82880
rect 28850 82810 28860 82880
rect 28640 82760 28860 82810
rect 29140 82880 29360 82900
rect 29140 82810 29150 82880
rect 29350 82810 29360 82880
rect 29140 82760 29360 82810
rect 29640 82880 29860 82900
rect 29640 82810 29650 82880
rect 29850 82810 29860 82880
rect 29640 82760 29860 82810
rect 30140 82880 30360 82900
rect 30140 82810 30150 82880
rect 30350 82810 30360 82880
rect 30140 82760 30360 82810
rect 30640 82880 30860 82900
rect 30640 82810 30650 82880
rect 30850 82810 30860 82880
rect 30640 82760 30860 82810
rect 31140 82880 31360 82900
rect 31140 82810 31150 82880
rect 31350 82810 31360 82880
rect 31140 82760 31360 82810
rect 31640 82880 31860 82900
rect 31640 82810 31650 82880
rect 31850 82810 31860 82880
rect 31640 82760 31860 82810
rect 32140 82880 32360 82900
rect 32140 82810 32150 82880
rect 32350 82810 32360 82880
rect 32140 82760 32360 82810
rect 32640 82880 32860 82900
rect 32640 82810 32650 82880
rect 32850 82810 32860 82880
rect 32640 82760 32860 82810
rect 33140 82880 33360 82900
rect 33140 82810 33150 82880
rect 33350 82810 33360 82880
rect 33140 82760 33360 82810
rect 33640 82880 33860 82900
rect 33640 82810 33650 82880
rect 33850 82810 33860 82880
rect 33640 82760 33860 82810
rect 34140 82880 34360 82900
rect 34140 82810 34150 82880
rect 34350 82810 34360 82880
rect 34140 82760 34360 82810
rect 34640 82880 34860 82900
rect 34640 82810 34650 82880
rect 34850 82810 34860 82880
rect 34640 82760 34860 82810
rect 35140 82880 35360 82900
rect 35140 82810 35150 82880
rect 35350 82810 35360 82880
rect 35140 82760 35360 82810
rect 35640 82880 35860 82900
rect 35640 82810 35650 82880
rect 35850 82810 35860 82880
rect 35640 82760 35860 82810
rect 36140 82880 36360 82900
rect 36140 82810 36150 82880
rect 36350 82810 36360 82880
rect 36140 82760 36360 82810
rect 36640 82880 36860 82900
rect 36640 82810 36650 82880
rect 36850 82810 36860 82880
rect 36640 82760 36860 82810
rect 37140 82880 37360 82900
rect 37140 82810 37150 82880
rect 37350 82810 37360 82880
rect 37140 82760 37360 82810
rect 37640 82880 37860 82900
rect 37640 82810 37650 82880
rect 37850 82810 37860 82880
rect 37640 82760 37860 82810
rect 38140 82880 38360 82900
rect 38140 82810 38150 82880
rect 38350 82810 38360 82880
rect 38140 82760 38360 82810
rect 38640 82880 38860 82900
rect 38640 82810 38650 82880
rect 38850 82810 38860 82880
rect 38640 82760 38860 82810
rect 39140 82880 39360 82900
rect 39140 82810 39150 82880
rect 39350 82810 39360 82880
rect 39140 82760 39360 82810
rect 39640 82880 39860 82900
rect 39640 82810 39650 82880
rect 39850 82810 39860 82880
rect 39640 82760 39860 82810
rect 40140 82880 40360 82900
rect 40140 82810 40150 82880
rect 40350 82810 40360 82880
rect 40140 82760 40360 82810
rect 40640 82880 40860 82900
rect 40640 82810 40650 82880
rect 40850 82810 40860 82880
rect 40640 82760 40860 82810
rect 41140 82880 41360 82900
rect 41140 82810 41150 82880
rect 41350 82810 41360 82880
rect 41140 82760 41360 82810
rect 41640 82880 41860 82900
rect 41640 82810 41650 82880
rect 41850 82810 41860 82880
rect 41640 82760 41860 82810
rect 42140 82880 42360 82900
rect 42140 82810 42150 82880
rect 42350 82810 42360 82880
rect 42140 82760 42360 82810
rect 42640 82880 42860 82900
rect 42640 82810 42650 82880
rect 42850 82810 42860 82880
rect 42640 82760 42860 82810
rect 43140 82880 43360 82900
rect 43140 82810 43150 82880
rect 43350 82810 43360 82880
rect 43140 82760 43360 82810
rect 43640 82880 43860 82900
rect 43640 82810 43650 82880
rect 43850 82810 43860 82880
rect 43640 82760 43860 82810
rect 44140 82880 44360 82900
rect 44140 82810 44150 82880
rect 44350 82810 44360 82880
rect 44140 82760 44360 82810
rect 44640 82880 44860 82900
rect 44640 82810 44650 82880
rect 44850 82810 44860 82880
rect 44640 82760 44860 82810
rect 45140 82880 45360 82900
rect 45140 82810 45150 82880
rect 45350 82810 45360 82880
rect 45140 82760 45360 82810
rect 45640 82880 45860 82900
rect 45640 82810 45650 82880
rect 45850 82810 45860 82880
rect 45640 82760 45860 82810
rect 46140 82880 46360 82900
rect 46140 82810 46150 82880
rect 46350 82810 46360 82880
rect 46140 82760 46360 82810
rect 46640 82880 46860 82900
rect 46640 82810 46650 82880
rect 46850 82810 46860 82880
rect 46640 82760 46860 82810
rect 47140 82880 47360 82900
rect 47140 82810 47150 82880
rect 47350 82810 47360 82880
rect 47140 82760 47360 82810
rect 47640 82880 47860 82900
rect 47640 82810 47650 82880
rect 47850 82810 47860 82880
rect 47640 82760 47860 82810
rect 48140 82880 48360 82900
rect 48140 82810 48150 82880
rect 48350 82810 48360 82880
rect 48140 82760 48360 82810
rect 48640 82880 48860 82900
rect 48640 82810 48650 82880
rect 48850 82810 48860 82880
rect 48640 82760 48860 82810
rect 49140 82880 49360 82900
rect 49140 82810 49150 82880
rect 49350 82810 49360 82880
rect 49140 82760 49360 82810
rect 49640 82880 49860 82900
rect 49640 82810 49650 82880
rect 49850 82810 49860 82880
rect 49640 82760 49860 82810
rect 50140 82880 50360 82900
rect 50140 82810 50150 82880
rect 50350 82810 50360 82880
rect 50140 82760 50360 82810
rect 50640 82880 50860 82900
rect 50640 82810 50650 82880
rect 50850 82810 50860 82880
rect 50640 82760 50860 82810
rect 51140 82880 51360 82900
rect 51140 82810 51150 82880
rect 51350 82810 51360 82880
rect 51140 82760 51360 82810
rect 51640 82880 51860 82900
rect 51640 82810 51650 82880
rect 51850 82810 51860 82880
rect 51640 82760 51860 82810
rect 52140 82880 52360 82900
rect 52140 82810 52150 82880
rect 52350 82810 52360 82880
rect 52140 82760 52360 82810
rect 52640 82880 52860 82900
rect 52640 82810 52650 82880
rect 52850 82810 52860 82880
rect 52640 82760 52860 82810
rect 53140 82880 53360 82900
rect 53140 82810 53150 82880
rect 53350 82810 53360 82880
rect 53140 82760 53360 82810
rect 53640 82880 53860 82900
rect 53640 82810 53650 82880
rect 53850 82810 53860 82880
rect 53640 82760 53860 82810
rect 54140 82880 54360 82900
rect 54140 82810 54150 82880
rect 54350 82810 54360 82880
rect 54140 82760 54360 82810
rect 54640 82880 54860 82900
rect 54640 82810 54650 82880
rect 54850 82810 54860 82880
rect 54640 82760 54860 82810
rect 55140 82880 55360 82900
rect 55140 82810 55150 82880
rect 55350 82810 55360 82880
rect 55140 82760 55360 82810
rect 55640 82880 55860 82900
rect 55640 82810 55650 82880
rect 55850 82810 55860 82880
rect 55640 82760 55860 82810
rect 56140 82880 56360 82900
rect 56140 82810 56150 82880
rect 56350 82810 56360 82880
rect 56140 82760 56360 82810
rect 56640 82880 56860 82900
rect 56640 82810 56650 82880
rect 56850 82810 56860 82880
rect 56640 82760 56860 82810
rect 57140 82880 57360 82900
rect 57140 82810 57150 82880
rect 57350 82810 57360 82880
rect 57140 82760 57360 82810
rect 57640 82880 57860 82900
rect 57640 82810 57650 82880
rect 57850 82810 57860 82880
rect 57640 82760 57860 82810
rect 58140 82880 58360 82900
rect 58140 82810 58150 82880
rect 58350 82810 58360 82880
rect 58140 82760 58360 82810
rect 58640 82880 58860 82900
rect 58640 82810 58650 82880
rect 58850 82810 58860 82880
rect 58640 82760 58860 82810
rect 59140 82880 59360 82900
rect 59140 82810 59150 82880
rect 59350 82810 59360 82880
rect 59140 82760 59360 82810
rect 59640 82880 59860 82900
rect 59640 82810 59650 82880
rect 59850 82810 59860 82880
rect 59640 82760 59860 82810
rect 60140 82880 60360 82900
rect 60140 82810 60150 82880
rect 60350 82810 60360 82880
rect 60140 82760 60360 82810
rect 60640 82880 60860 82900
rect 60640 82810 60650 82880
rect 60850 82810 60860 82880
rect 60640 82760 60860 82810
rect 61140 82880 61360 82900
rect 61140 82810 61150 82880
rect 61350 82810 61360 82880
rect 61140 82760 61360 82810
rect 61640 82880 61860 82900
rect 61640 82810 61650 82880
rect 61850 82810 61860 82880
rect 61640 82760 61860 82810
rect 62140 82880 62360 82900
rect 62140 82810 62150 82880
rect 62350 82810 62360 82880
rect 62140 82760 62360 82810
rect 62640 82880 62860 82900
rect 62640 82810 62650 82880
rect 62850 82810 62860 82880
rect 62640 82760 62860 82810
rect 63140 82880 63360 82900
rect 63140 82810 63150 82880
rect 63350 82810 63360 82880
rect 63140 82760 63360 82810
rect 63640 82880 63860 82900
rect 63640 82810 63650 82880
rect 63850 82810 63860 82880
rect 63640 82760 63860 82810
rect 64140 82880 64360 82900
rect 64140 82810 64150 82880
rect 64350 82810 64360 82880
rect 64140 82760 64360 82810
rect 64640 82880 64860 82900
rect 64640 82810 64650 82880
rect 64850 82810 64860 82880
rect 64640 82760 64860 82810
rect 65140 82880 65360 82900
rect 65140 82810 65150 82880
rect 65350 82810 65360 82880
rect 65140 82760 65360 82810
rect 65640 82880 65860 82900
rect 65640 82810 65650 82880
rect 65850 82810 65860 82880
rect 65640 82760 65860 82810
rect 66140 82880 66360 82900
rect 66140 82810 66150 82880
rect 66350 82810 66360 82880
rect 66140 82760 66360 82810
rect 66640 82880 66860 82900
rect 66640 82810 66650 82880
rect 66850 82810 66860 82880
rect 66640 82760 66860 82810
rect 67140 82880 67360 82900
rect 67140 82810 67150 82880
rect 67350 82810 67360 82880
rect 67140 82760 67360 82810
rect 67640 82880 67860 82900
rect 67640 82810 67650 82880
rect 67850 82810 67860 82880
rect 67640 82760 67860 82810
rect 68140 82880 68360 82900
rect 68140 82810 68150 82880
rect 68350 82810 68360 82880
rect 68140 82760 68360 82810
rect 68640 82880 68860 82900
rect 68640 82810 68650 82880
rect 68850 82810 68860 82880
rect 68640 82760 68860 82810
rect 69140 82880 69360 82900
rect 69140 82810 69150 82880
rect 69350 82810 69360 82880
rect 69140 82760 69360 82810
rect 69640 82880 69860 82900
rect 69640 82810 69650 82880
rect 69850 82810 69860 82880
rect 69640 82760 69860 82810
rect 70140 82880 70360 82900
rect 70140 82810 70150 82880
rect 70350 82810 70360 82880
rect 70140 82760 70360 82810
rect 70640 82880 70860 82900
rect 70640 82810 70650 82880
rect 70850 82810 70860 82880
rect 70640 82760 70860 82810
rect 71140 82880 71360 82900
rect 71140 82810 71150 82880
rect 71350 82810 71360 82880
rect 71140 82760 71360 82810
rect 71640 82880 71860 82900
rect 71640 82810 71650 82880
rect 71850 82810 71860 82880
rect 71640 82760 71860 82810
rect 72140 82880 72360 82900
rect 72140 82810 72150 82880
rect 72350 82810 72360 82880
rect 72140 82760 72360 82810
rect 72640 82880 72860 82900
rect 72640 82810 72650 82880
rect 72850 82810 72860 82880
rect 72640 82760 72860 82810
rect 73140 82880 73360 82900
rect 73140 82810 73150 82880
rect 73350 82810 73360 82880
rect 73140 82760 73360 82810
rect 73640 82880 73860 82900
rect 73640 82810 73650 82880
rect 73850 82810 73860 82880
rect 73640 82760 73860 82810
rect 74140 82880 74360 82900
rect 74140 82810 74150 82880
rect 74350 82810 74360 82880
rect 74140 82760 74360 82810
rect 74640 82880 74860 82900
rect 74640 82810 74650 82880
rect 74850 82810 74860 82880
rect 74640 82760 74860 82810
rect 75140 82880 75360 82900
rect 75140 82810 75150 82880
rect 75350 82810 75360 82880
rect 75140 82760 75360 82810
rect 75640 82880 75860 82900
rect 75640 82810 75650 82880
rect 75850 82810 75860 82880
rect 75640 82760 75860 82810
rect 76140 82880 76360 82900
rect 76140 82810 76150 82880
rect 76350 82810 76360 82880
rect 76140 82760 76360 82810
rect 76640 82880 76860 82900
rect 76640 82810 76650 82880
rect 76850 82810 76860 82880
rect 76640 82760 76860 82810
rect 77140 82880 77360 82900
rect 77140 82810 77150 82880
rect 77350 82810 77360 82880
rect 77140 82760 77360 82810
rect 77640 82880 77860 82900
rect 77640 82810 77650 82880
rect 77850 82810 77860 82880
rect 77640 82760 77860 82810
rect 78140 82880 78360 82900
rect 78140 82810 78150 82880
rect 78350 82810 78360 82880
rect 78140 82760 78360 82810
rect 78640 82880 78860 82900
rect 78640 82810 78650 82880
rect 78850 82810 78860 82880
rect 78640 82760 78860 82810
rect 79140 82880 79360 82900
rect 79140 82810 79150 82880
rect 79350 82810 79360 82880
rect 79140 82760 79360 82810
rect 79640 82880 79860 82900
rect 79640 82810 79650 82880
rect 79850 82810 79860 82880
rect 79640 82760 79860 82810
rect 80140 82880 80360 82900
rect 80140 82810 80150 82880
rect 80350 82810 80360 82880
rect 80140 82760 80360 82810
rect 80640 82880 80860 82900
rect 80640 82810 80650 82880
rect 80850 82810 80860 82880
rect 80640 82760 80860 82810
rect 81140 82880 81360 82900
rect 81140 82810 81150 82880
rect 81350 82810 81360 82880
rect 81140 82760 81360 82810
rect 81640 82880 81860 82900
rect 81640 82810 81650 82880
rect 81850 82810 81860 82880
rect 81640 82760 81860 82810
rect 82140 82880 82360 82900
rect 82140 82810 82150 82880
rect 82350 82810 82360 82880
rect 82140 82760 82360 82810
rect 82640 82880 82860 82900
rect 82640 82810 82650 82880
rect 82850 82810 82860 82880
rect 82640 82760 82860 82810
rect 83140 82880 83360 82900
rect 83140 82810 83150 82880
rect 83350 82810 83360 82880
rect 83140 82760 83360 82810
rect 83640 82880 83860 82900
rect 83640 82810 83650 82880
rect 83850 82810 83860 82880
rect 83640 82760 83860 82810
rect 84140 82880 84360 82900
rect 84140 82810 84150 82880
rect 84350 82810 84360 82880
rect 84140 82760 84360 82810
rect 84640 82880 84860 82900
rect 84640 82810 84650 82880
rect 84850 82810 84860 82880
rect 84640 82760 84860 82810
rect 85140 82880 85360 82900
rect 85140 82810 85150 82880
rect 85350 82810 85360 82880
rect 85140 82760 85360 82810
rect 85640 82880 85860 82900
rect 85640 82810 85650 82880
rect 85850 82810 85860 82880
rect 85640 82760 85860 82810
rect 86140 82880 86360 82900
rect 86140 82810 86150 82880
rect 86350 82810 86360 82880
rect 86140 82760 86360 82810
rect 86640 82880 86860 82900
rect 86640 82810 86650 82880
rect 86850 82810 86860 82880
rect 86640 82760 86860 82810
rect 87140 82880 87360 82900
rect 87140 82810 87150 82880
rect 87350 82810 87360 82880
rect 87140 82760 87360 82810
rect 87640 82880 87860 82900
rect 87640 82810 87650 82880
rect 87850 82810 87860 82880
rect 87640 82760 87860 82810
rect 88140 82880 88360 82900
rect 88140 82810 88150 82880
rect 88350 82810 88360 82880
rect 88140 82760 88360 82810
rect 88640 82880 88860 82900
rect 88640 82810 88650 82880
rect 88850 82810 88860 82880
rect 88640 82760 88860 82810
rect 89140 82880 89360 82900
rect 89140 82810 89150 82880
rect 89350 82810 89360 82880
rect 89140 82760 89360 82810
rect 89640 82880 89860 82900
rect 89640 82810 89650 82880
rect 89850 82810 89860 82880
rect 89640 82760 89860 82810
rect 90140 82880 90360 82900
rect 90140 82810 90150 82880
rect 90350 82810 90360 82880
rect 90140 82760 90360 82810
rect 90640 82880 90860 82900
rect 90640 82810 90650 82880
rect 90850 82810 90860 82880
rect 90640 82760 90860 82810
rect 91140 82880 91360 82900
rect 91140 82810 91150 82880
rect 91350 82810 91360 82880
rect 91140 82760 91360 82810
rect 91640 82880 91860 82900
rect 91640 82810 91650 82880
rect 91850 82810 91860 82880
rect 91640 82760 91860 82810
rect 92140 82880 92360 82900
rect 92140 82810 92150 82880
rect 92350 82810 92360 82880
rect 92140 82760 92360 82810
rect 92640 82880 92860 82900
rect 92640 82810 92650 82880
rect 92850 82810 92860 82880
rect 92640 82760 92860 82810
rect 93140 82880 93360 82900
rect 93140 82810 93150 82880
rect 93350 82810 93360 82880
rect 93140 82760 93360 82810
rect 93640 82880 93860 82900
rect 93640 82810 93650 82880
rect 93850 82810 93860 82880
rect 93640 82760 93860 82810
rect 94140 82880 94360 82900
rect 94140 82810 94150 82880
rect 94350 82810 94360 82880
rect 94140 82760 94360 82810
rect 94640 82880 94860 82900
rect 94640 82810 94650 82880
rect 94850 82810 94860 82880
rect 94640 82760 94860 82810
rect 95140 82880 95360 82900
rect 95140 82810 95150 82880
rect 95350 82810 95360 82880
rect 95140 82760 95360 82810
rect 95640 82880 95860 82900
rect 95640 82810 95650 82880
rect 95850 82810 95860 82880
rect 95640 82760 95860 82810
rect 96140 82880 96360 82900
rect 96140 82810 96150 82880
rect 96350 82810 96360 82880
rect 96140 82760 96360 82810
rect 96640 82880 96860 82900
rect 96640 82810 96650 82880
rect 96850 82810 96860 82880
rect 96640 82760 96860 82810
rect 97140 82880 97360 82900
rect 97140 82810 97150 82880
rect 97350 82810 97360 82880
rect 97140 82760 97360 82810
rect 97640 82880 97860 82900
rect 97640 82810 97650 82880
rect 97850 82810 97860 82880
rect 97640 82760 97860 82810
rect 98140 82880 98360 82900
rect 98140 82810 98150 82880
rect 98350 82810 98360 82880
rect 98140 82760 98360 82810
rect 98640 82880 98860 82900
rect 98640 82810 98650 82880
rect 98850 82810 98860 82880
rect 98640 82760 98860 82810
rect 99140 82880 99360 82900
rect 99140 82810 99150 82880
rect 99350 82810 99360 82880
rect 99140 82760 99360 82810
rect 99640 82880 99860 82900
rect 99640 82810 99650 82880
rect 99850 82810 99860 82880
rect 99640 82760 99860 82810
rect 100140 82880 100360 82900
rect 100140 82810 100150 82880
rect 100350 82810 100360 82880
rect 100140 82760 100360 82810
rect -83500 82750 100500 82760
rect -83500 82550 -83480 82750
rect -83410 82550 -83090 82750
rect -83020 82550 -82980 82750
rect -82910 82550 -82590 82750
rect -82520 82550 -82480 82750
rect -82410 82550 -82090 82750
rect -82020 82550 -81980 82750
rect -81910 82550 -81590 82750
rect -81520 82550 -81480 82750
rect -81410 82550 -81090 82750
rect -81020 82550 -80980 82750
rect -80910 82550 -80590 82750
rect -80520 82550 -80480 82750
rect -80410 82550 -80090 82750
rect -80020 82550 -79980 82750
rect -79910 82550 -79590 82750
rect -79520 82550 -79480 82750
rect -79410 82550 -79090 82750
rect -79020 82550 -78980 82750
rect -78910 82550 -78590 82750
rect -78520 82550 -78480 82750
rect -78410 82550 -78090 82750
rect -78020 82550 -77980 82750
rect -77910 82550 -77590 82750
rect -77520 82550 -77480 82750
rect -77410 82550 -77090 82750
rect -77020 82550 -76980 82750
rect -76910 82550 -76590 82750
rect -76520 82550 -76480 82750
rect -76410 82550 -76090 82750
rect -76020 82550 -75980 82750
rect -75910 82550 -75590 82750
rect -75520 82550 -75480 82750
rect -75410 82550 -75090 82750
rect -75020 82550 -74980 82750
rect -74910 82550 -74590 82750
rect -74520 82550 -74480 82750
rect -74410 82550 -74090 82750
rect -74020 82550 -73980 82750
rect -73910 82550 -73590 82750
rect -73520 82550 -73480 82750
rect -73410 82550 -73090 82750
rect -73020 82550 -72980 82750
rect -72910 82550 -72590 82750
rect -72520 82550 -72480 82750
rect -72410 82550 -72090 82750
rect -72020 82550 -71980 82750
rect -71910 82550 -71590 82750
rect -71520 82550 -71480 82750
rect -71410 82550 -71090 82750
rect -71020 82550 -70980 82750
rect -70910 82550 -70590 82750
rect -70520 82550 -70480 82750
rect -70410 82550 -70090 82750
rect -70020 82550 -69980 82750
rect -69910 82550 -69590 82750
rect -69520 82550 -69480 82750
rect -69410 82550 -69090 82750
rect -69020 82550 -68980 82750
rect -68910 82550 -68590 82750
rect -68520 82550 -68480 82750
rect -68410 82550 -68090 82750
rect -68020 82550 -67980 82750
rect -67910 82550 -67590 82750
rect -67520 82550 -67480 82750
rect -67410 82550 -67090 82750
rect -67020 82550 -66980 82750
rect -66910 82550 -66590 82750
rect -66520 82550 -66480 82750
rect -66410 82550 -66090 82750
rect -66020 82550 -65980 82750
rect -65910 82550 -65590 82750
rect -65520 82550 -65480 82750
rect -65410 82550 -65090 82750
rect -65020 82550 -64980 82750
rect -64910 82550 -64590 82750
rect -64520 82550 -64480 82750
rect -64410 82550 -64090 82750
rect -64020 82550 -63980 82750
rect -63910 82550 -63590 82750
rect -63520 82550 -63480 82750
rect -63410 82550 -63090 82750
rect -63020 82550 -62980 82750
rect -62910 82550 -62590 82750
rect -62520 82550 -62480 82750
rect -62410 82550 -62090 82750
rect -62020 82550 -61980 82750
rect -61910 82550 -61590 82750
rect -61520 82550 -61480 82750
rect -61410 82550 -61090 82750
rect -61020 82550 -60980 82750
rect -60910 82550 -60590 82750
rect -60520 82550 -60480 82750
rect -60410 82550 -60090 82750
rect -60020 82550 -59980 82750
rect -59910 82550 -59590 82750
rect -59520 82550 -59480 82750
rect -59410 82550 -59090 82750
rect -59020 82550 -58980 82750
rect -58910 82550 -58590 82750
rect -58520 82550 -58480 82750
rect -58410 82550 -58090 82750
rect -58020 82550 -57980 82750
rect -57910 82550 -57590 82750
rect -57520 82550 -57480 82750
rect -57410 82550 -57090 82750
rect -57020 82550 -56980 82750
rect -56910 82550 -56590 82750
rect -56520 82550 -56480 82750
rect -56410 82550 -56090 82750
rect -56020 82550 -55980 82750
rect -55910 82550 -55590 82750
rect -55520 82550 -55480 82750
rect -55410 82550 -55090 82750
rect -55020 82550 -54980 82750
rect -54910 82550 -54590 82750
rect -54520 82550 -54480 82750
rect -54410 82550 -54090 82750
rect -54020 82550 -53980 82750
rect -53910 82550 -53590 82750
rect -53520 82550 -53480 82750
rect -53410 82550 -53090 82750
rect -53020 82550 -52980 82750
rect -52910 82550 -52590 82750
rect -52520 82550 -52480 82750
rect -52410 82550 -52090 82750
rect -52020 82550 -51980 82750
rect -51910 82550 -51590 82750
rect -51520 82550 -51480 82750
rect -51410 82550 -51090 82750
rect -51020 82550 -50980 82750
rect -50910 82550 -50590 82750
rect -50520 82550 -50480 82750
rect -50410 82550 -50090 82750
rect -50020 82550 -49980 82750
rect -49910 82550 -49590 82750
rect -49520 82550 -49480 82750
rect -49410 82550 -49090 82750
rect -49020 82550 -48980 82750
rect -48910 82550 -48590 82750
rect -48520 82550 -48480 82750
rect -48410 82550 -48090 82750
rect -48020 82550 -47980 82750
rect -47910 82550 -47590 82750
rect -47520 82550 -47480 82750
rect -47410 82550 -47090 82750
rect -47020 82550 -46980 82750
rect -46910 82550 -46590 82750
rect -46520 82550 -46480 82750
rect -46410 82550 -46090 82750
rect -46020 82550 -45980 82750
rect -45910 82550 -45590 82750
rect -45520 82550 -45480 82750
rect -45410 82550 -45090 82750
rect -45020 82550 -44980 82750
rect -44910 82550 -44590 82750
rect -44520 82550 -44480 82750
rect -44410 82550 -44090 82750
rect -44020 82550 -43980 82750
rect -43910 82550 -43590 82750
rect -43520 82550 -43480 82750
rect -43410 82550 -43090 82750
rect -43020 82550 -42980 82750
rect -42910 82550 -42590 82750
rect -42520 82550 -42480 82750
rect -42410 82550 -42090 82750
rect -42020 82550 -41980 82750
rect -41910 82550 -41590 82750
rect -41520 82550 -41480 82750
rect -41410 82550 -41090 82750
rect -41020 82550 -40980 82750
rect -40910 82550 -40590 82750
rect -40520 82550 -40480 82750
rect -40410 82550 -40090 82750
rect -40020 82550 -39980 82750
rect -39910 82550 -39590 82750
rect -39520 82550 -39480 82750
rect -39410 82550 -39090 82750
rect -39020 82550 -38980 82750
rect -38910 82550 -38590 82750
rect -38520 82550 -38480 82750
rect -38410 82550 -38090 82750
rect -38020 82550 -37980 82750
rect -37910 82550 -37590 82750
rect -37520 82550 -37480 82750
rect -37410 82550 -37090 82750
rect -37020 82550 -36980 82750
rect -36910 82550 -36590 82750
rect -36520 82550 -36480 82750
rect -36410 82550 -36090 82750
rect -36020 82550 -35980 82750
rect -35910 82550 -35590 82750
rect -35520 82550 -35480 82750
rect -35410 82550 -35090 82750
rect -35020 82550 -34980 82750
rect -34910 82550 -34590 82750
rect -34520 82550 -34480 82750
rect -34410 82550 -34090 82750
rect -34020 82550 -33980 82750
rect -33910 82550 -33590 82750
rect -33520 82550 -33480 82750
rect -33410 82550 -33090 82750
rect -33020 82550 -32980 82750
rect -32910 82550 -32590 82750
rect -32520 82550 -32480 82750
rect -32410 82550 -32090 82750
rect -32020 82550 -31980 82750
rect -31910 82550 -31590 82750
rect -31520 82550 -31480 82750
rect -31410 82550 -31090 82750
rect -31020 82550 -30980 82750
rect -30910 82550 -30590 82750
rect -30520 82550 -30480 82750
rect -30410 82550 -30090 82750
rect -30020 82550 -29980 82750
rect -29910 82550 -29590 82750
rect -29520 82550 -29480 82750
rect -29410 82550 -29090 82750
rect -29020 82550 -28980 82750
rect -28910 82550 -28590 82750
rect -28520 82550 -28480 82750
rect -28410 82550 -28090 82750
rect -28020 82550 -27980 82750
rect -27910 82550 -27590 82750
rect -27520 82550 -27480 82750
rect -27410 82550 -27090 82750
rect -27020 82550 -26980 82750
rect -26910 82550 -26590 82750
rect -26520 82550 -26480 82750
rect -26410 82550 -26090 82750
rect -26020 82550 -25980 82750
rect -25910 82550 -25590 82750
rect -25520 82550 -25480 82750
rect -25410 82550 -25090 82750
rect -25020 82550 -24980 82750
rect -24910 82550 -24590 82750
rect -24520 82550 -24480 82750
rect -24410 82550 -24090 82750
rect -24020 82550 -23980 82750
rect -23910 82550 -23590 82750
rect -23520 82550 -23480 82750
rect -23410 82550 -23090 82750
rect -23020 82550 -22980 82750
rect -22910 82550 -22590 82750
rect -22520 82550 -22480 82750
rect -22410 82550 -22090 82750
rect -22020 82550 -21980 82750
rect -21910 82550 -21590 82750
rect -21520 82550 -21480 82750
rect -21410 82550 -21090 82750
rect -21020 82550 -20980 82750
rect -20910 82550 -20590 82750
rect -20520 82550 -20480 82750
rect -20410 82550 -20090 82750
rect -20020 82550 -19980 82750
rect -19910 82550 -19590 82750
rect -19520 82550 -19480 82750
rect -19410 82550 -19090 82750
rect -19020 82550 -18980 82750
rect -18910 82550 -18590 82750
rect -18520 82550 -18480 82750
rect -18410 82550 -18090 82750
rect -18020 82550 -17980 82750
rect -17910 82550 -17590 82750
rect -17520 82550 -17480 82750
rect -17410 82550 -17090 82750
rect -17020 82550 -16980 82750
rect -16910 82550 -16590 82750
rect -16520 82550 -16480 82750
rect -16410 82550 -16090 82750
rect -16020 82550 -15980 82750
rect -15910 82550 -15590 82750
rect -15520 82550 -15480 82750
rect -15410 82550 -15090 82750
rect -15020 82550 -14980 82750
rect -14910 82550 -14590 82750
rect -14520 82550 -14480 82750
rect -14410 82550 -14090 82750
rect -14020 82550 -13980 82750
rect -13910 82550 -13590 82750
rect -13520 82550 -13480 82750
rect -13410 82550 -13090 82750
rect -13020 82550 -12980 82750
rect -12910 82550 -12590 82750
rect -12520 82550 -12480 82750
rect -12410 82550 -12090 82750
rect -12020 82550 -11980 82750
rect -11910 82550 -11590 82750
rect -11520 82550 -11480 82750
rect -11410 82550 -11090 82750
rect -11020 82550 -10980 82750
rect -10910 82550 -10590 82750
rect -10520 82550 -10480 82750
rect -10410 82550 -10090 82750
rect -10020 82550 -9980 82750
rect -9910 82550 -9590 82750
rect -9520 82550 -9480 82750
rect -9410 82550 -9090 82750
rect -9020 82550 -8980 82750
rect -8910 82550 -8590 82750
rect -8520 82550 -8480 82750
rect -8410 82550 -8090 82750
rect -8020 82550 -7980 82750
rect -7910 82550 -7590 82750
rect -7520 82550 -7480 82750
rect -7410 82550 -7090 82750
rect -7020 82550 -6980 82750
rect -6910 82550 -6590 82750
rect -6520 82550 -6480 82750
rect -6410 82550 -6090 82750
rect -6020 82550 -5980 82750
rect -5910 82550 -5590 82750
rect -5520 82550 -5480 82750
rect -5410 82550 -5090 82750
rect -5020 82550 -4980 82750
rect -4910 82550 -4590 82750
rect -4520 82550 -4480 82750
rect -4410 82550 -4090 82750
rect -4020 82550 -3980 82750
rect -3910 82550 -3590 82750
rect -3520 82550 -3480 82750
rect -3410 82550 -3090 82750
rect -3020 82550 -2980 82750
rect -2910 82550 -2590 82750
rect -2520 82550 -2480 82750
rect -2410 82550 -2090 82750
rect -2020 82550 -1980 82750
rect -1910 82550 -1590 82750
rect -1520 82550 -1480 82750
rect -1410 82550 -1090 82750
rect -1020 82550 -980 82750
rect -910 82550 -590 82750
rect -520 82550 -480 82750
rect -410 82550 -90 82750
rect -20 82550 20 82750
rect 90 82550 410 82750
rect 480 82550 520 82750
rect 590 82550 910 82750
rect 980 82550 1020 82750
rect 1090 82550 1410 82750
rect 1480 82550 1520 82750
rect 1590 82550 1910 82750
rect 1980 82550 2020 82750
rect 2090 82550 2410 82750
rect 2480 82550 2520 82750
rect 2590 82550 2910 82750
rect 2980 82550 3020 82750
rect 3090 82550 3410 82750
rect 3480 82550 3520 82750
rect 3590 82550 3910 82750
rect 3980 82550 4020 82750
rect 4090 82550 4410 82750
rect 4480 82550 4520 82750
rect 4590 82550 4910 82750
rect 4980 82550 5020 82750
rect 5090 82550 5410 82750
rect 5480 82550 5520 82750
rect 5590 82550 5910 82750
rect 5980 82550 6020 82750
rect 6090 82550 6410 82750
rect 6480 82550 6520 82750
rect 6590 82550 6910 82750
rect 6980 82550 7020 82750
rect 7090 82550 7410 82750
rect 7480 82550 7520 82750
rect 7590 82550 7910 82750
rect 7980 82550 8020 82750
rect 8090 82550 8410 82750
rect 8480 82550 8520 82750
rect 8590 82550 8910 82750
rect 8980 82550 9020 82750
rect 9090 82550 9410 82750
rect 9480 82550 9520 82750
rect 9590 82550 9910 82750
rect 9980 82550 10020 82750
rect 10090 82550 10410 82750
rect 10480 82550 10520 82750
rect 10590 82550 10910 82750
rect 10980 82550 11020 82750
rect 11090 82550 11410 82750
rect 11480 82550 11520 82750
rect 11590 82550 11910 82750
rect 11980 82550 12020 82750
rect 12090 82550 12410 82750
rect 12480 82550 12520 82750
rect 12590 82550 12910 82750
rect 12980 82550 13020 82750
rect 13090 82550 13410 82750
rect 13480 82550 13520 82750
rect 13590 82550 13910 82750
rect 13980 82550 14020 82750
rect 14090 82550 14410 82750
rect 14480 82550 14520 82750
rect 14590 82550 14910 82750
rect 14980 82550 15020 82750
rect 15090 82550 15410 82750
rect 15480 82550 15520 82750
rect 15590 82550 15910 82750
rect 15980 82550 16020 82750
rect 16090 82550 16410 82750
rect 16480 82550 16520 82750
rect 16590 82550 16910 82750
rect 16980 82550 17020 82750
rect 17090 82550 17410 82750
rect 17480 82550 17520 82750
rect 17590 82550 17910 82750
rect 17980 82550 18020 82750
rect 18090 82550 18410 82750
rect 18480 82550 18520 82750
rect 18590 82550 18910 82750
rect 18980 82550 19020 82750
rect 19090 82550 19410 82750
rect 19480 82550 19520 82750
rect 19590 82550 19910 82750
rect 19980 82550 20020 82750
rect 20090 82550 20410 82750
rect 20480 82550 20520 82750
rect 20590 82550 20910 82750
rect 20980 82550 21020 82750
rect 21090 82550 21410 82750
rect 21480 82550 21520 82750
rect 21590 82550 21910 82750
rect 21980 82550 22020 82750
rect 22090 82550 22410 82750
rect 22480 82550 22520 82750
rect 22590 82550 22910 82750
rect 22980 82550 23020 82750
rect 23090 82550 23410 82750
rect 23480 82550 23520 82750
rect 23590 82550 23910 82750
rect 23980 82550 24020 82750
rect 24090 82550 24410 82750
rect 24480 82550 24520 82750
rect 24590 82550 24910 82750
rect 24980 82550 25020 82750
rect 25090 82550 25410 82750
rect 25480 82550 25520 82750
rect 25590 82550 25910 82750
rect 25980 82550 26020 82750
rect 26090 82550 26410 82750
rect 26480 82550 26520 82750
rect 26590 82550 26910 82750
rect 26980 82550 27020 82750
rect 27090 82550 27410 82750
rect 27480 82550 27520 82750
rect 27590 82550 27910 82750
rect 27980 82550 28020 82750
rect 28090 82550 28410 82750
rect 28480 82550 28520 82750
rect 28590 82550 28910 82750
rect 28980 82550 29020 82750
rect 29090 82550 29410 82750
rect 29480 82550 29520 82750
rect 29590 82550 29910 82750
rect 29980 82550 30020 82750
rect 30090 82550 30410 82750
rect 30480 82550 30520 82750
rect 30590 82550 30910 82750
rect 30980 82550 31020 82750
rect 31090 82550 31410 82750
rect 31480 82550 31520 82750
rect 31590 82550 31910 82750
rect 31980 82550 32020 82750
rect 32090 82550 32410 82750
rect 32480 82550 32520 82750
rect 32590 82550 32910 82750
rect 32980 82550 33020 82750
rect 33090 82550 33410 82750
rect 33480 82550 33520 82750
rect 33590 82550 33910 82750
rect 33980 82550 34020 82750
rect 34090 82550 34410 82750
rect 34480 82550 34520 82750
rect 34590 82550 34910 82750
rect 34980 82550 35020 82750
rect 35090 82550 35410 82750
rect 35480 82550 35520 82750
rect 35590 82550 35910 82750
rect 35980 82550 36020 82750
rect 36090 82550 36410 82750
rect 36480 82550 36520 82750
rect 36590 82550 36910 82750
rect 36980 82550 37020 82750
rect 37090 82550 37410 82750
rect 37480 82550 37520 82750
rect 37590 82550 37910 82750
rect 37980 82550 38020 82750
rect 38090 82550 38410 82750
rect 38480 82550 38520 82750
rect 38590 82550 38910 82750
rect 38980 82550 39020 82750
rect 39090 82550 39410 82750
rect 39480 82550 39520 82750
rect 39590 82550 39910 82750
rect 39980 82550 40020 82750
rect 40090 82550 40410 82750
rect 40480 82550 40520 82750
rect 40590 82550 40910 82750
rect 40980 82550 41020 82750
rect 41090 82550 41410 82750
rect 41480 82550 41520 82750
rect 41590 82550 41910 82750
rect 41980 82550 42020 82750
rect 42090 82550 42410 82750
rect 42480 82550 42520 82750
rect 42590 82550 42910 82750
rect 42980 82550 43020 82750
rect 43090 82550 43410 82750
rect 43480 82550 43520 82750
rect 43590 82550 43910 82750
rect 43980 82550 44020 82750
rect 44090 82550 44410 82750
rect 44480 82550 44520 82750
rect 44590 82550 44910 82750
rect 44980 82550 45020 82750
rect 45090 82550 45410 82750
rect 45480 82550 45520 82750
rect 45590 82550 45910 82750
rect 45980 82550 46020 82750
rect 46090 82550 46410 82750
rect 46480 82550 46520 82750
rect 46590 82550 46910 82750
rect 46980 82550 47020 82750
rect 47090 82550 47410 82750
rect 47480 82550 47520 82750
rect 47590 82550 47910 82750
rect 47980 82550 48020 82750
rect 48090 82550 48410 82750
rect 48480 82550 48520 82750
rect 48590 82550 48910 82750
rect 48980 82550 49020 82750
rect 49090 82550 49410 82750
rect 49480 82550 49520 82750
rect 49590 82550 49910 82750
rect 49980 82550 50020 82750
rect 50090 82550 50410 82750
rect 50480 82550 50520 82750
rect 50590 82550 50910 82750
rect 50980 82550 51020 82750
rect 51090 82550 51410 82750
rect 51480 82550 51520 82750
rect 51590 82550 51910 82750
rect 51980 82550 52020 82750
rect 52090 82550 52410 82750
rect 52480 82550 52520 82750
rect 52590 82550 52910 82750
rect 52980 82550 53020 82750
rect 53090 82550 53410 82750
rect 53480 82550 53520 82750
rect 53590 82550 53910 82750
rect 53980 82550 54020 82750
rect 54090 82550 54410 82750
rect 54480 82550 54520 82750
rect 54590 82550 54910 82750
rect 54980 82550 55020 82750
rect 55090 82550 55410 82750
rect 55480 82550 55520 82750
rect 55590 82550 55910 82750
rect 55980 82550 56020 82750
rect 56090 82550 56410 82750
rect 56480 82550 56520 82750
rect 56590 82550 56910 82750
rect 56980 82550 57020 82750
rect 57090 82550 57410 82750
rect 57480 82550 57520 82750
rect 57590 82550 57910 82750
rect 57980 82550 58020 82750
rect 58090 82550 58410 82750
rect 58480 82550 58520 82750
rect 58590 82550 58910 82750
rect 58980 82550 59020 82750
rect 59090 82550 59410 82750
rect 59480 82550 59520 82750
rect 59590 82550 59910 82750
rect 59980 82550 60020 82750
rect 60090 82550 60410 82750
rect 60480 82550 60520 82750
rect 60590 82550 60910 82750
rect 60980 82550 61020 82750
rect 61090 82550 61410 82750
rect 61480 82550 61520 82750
rect 61590 82550 61910 82750
rect 61980 82550 62020 82750
rect 62090 82550 62410 82750
rect 62480 82550 62520 82750
rect 62590 82550 62910 82750
rect 62980 82550 63020 82750
rect 63090 82550 63410 82750
rect 63480 82550 63520 82750
rect 63590 82550 63910 82750
rect 63980 82550 64020 82750
rect 64090 82550 64410 82750
rect 64480 82550 64520 82750
rect 64590 82550 64910 82750
rect 64980 82550 65020 82750
rect 65090 82550 65410 82750
rect 65480 82550 65520 82750
rect 65590 82550 65910 82750
rect 65980 82550 66020 82750
rect 66090 82550 66410 82750
rect 66480 82550 66520 82750
rect 66590 82550 66910 82750
rect 66980 82550 67020 82750
rect 67090 82550 67410 82750
rect 67480 82550 67520 82750
rect 67590 82550 67910 82750
rect 67980 82550 68020 82750
rect 68090 82550 68410 82750
rect 68480 82550 68520 82750
rect 68590 82550 68910 82750
rect 68980 82550 69020 82750
rect 69090 82550 69410 82750
rect 69480 82550 69520 82750
rect 69590 82550 69910 82750
rect 69980 82550 70020 82750
rect 70090 82550 70410 82750
rect 70480 82550 70520 82750
rect 70590 82550 70910 82750
rect 70980 82550 71020 82750
rect 71090 82550 71410 82750
rect 71480 82550 71520 82750
rect 71590 82550 71910 82750
rect 71980 82550 72020 82750
rect 72090 82550 72410 82750
rect 72480 82550 72520 82750
rect 72590 82550 72910 82750
rect 72980 82550 73020 82750
rect 73090 82550 73410 82750
rect 73480 82550 73520 82750
rect 73590 82550 73910 82750
rect 73980 82550 74020 82750
rect 74090 82550 74410 82750
rect 74480 82550 74520 82750
rect 74590 82550 74910 82750
rect 74980 82550 75020 82750
rect 75090 82550 75410 82750
rect 75480 82550 75520 82750
rect 75590 82550 75910 82750
rect 75980 82550 76020 82750
rect 76090 82550 76410 82750
rect 76480 82550 76520 82750
rect 76590 82550 76910 82750
rect 76980 82550 77020 82750
rect 77090 82550 77410 82750
rect 77480 82550 77520 82750
rect 77590 82550 77910 82750
rect 77980 82550 78020 82750
rect 78090 82550 78410 82750
rect 78480 82550 78520 82750
rect 78590 82550 78910 82750
rect 78980 82550 79020 82750
rect 79090 82550 79410 82750
rect 79480 82550 79520 82750
rect 79590 82550 79910 82750
rect 79980 82550 80020 82750
rect 80090 82550 80410 82750
rect 80480 82550 80520 82750
rect 80590 82550 80910 82750
rect 80980 82550 81020 82750
rect 81090 82550 81410 82750
rect 81480 82550 81520 82750
rect 81590 82550 81910 82750
rect 81980 82550 82020 82750
rect 82090 82550 82410 82750
rect 82480 82550 82520 82750
rect 82590 82550 82910 82750
rect 82980 82550 83020 82750
rect 83090 82550 83410 82750
rect 83480 82550 83520 82750
rect 83590 82550 83910 82750
rect 83980 82550 84020 82750
rect 84090 82550 84410 82750
rect 84480 82550 84520 82750
rect 84590 82550 84910 82750
rect 84980 82550 85020 82750
rect 85090 82550 85410 82750
rect 85480 82550 85520 82750
rect 85590 82550 85910 82750
rect 85980 82550 86020 82750
rect 86090 82550 86410 82750
rect 86480 82550 86520 82750
rect 86590 82550 86910 82750
rect 86980 82550 87020 82750
rect 87090 82550 87410 82750
rect 87480 82550 87520 82750
rect 87590 82550 87910 82750
rect 87980 82550 88020 82750
rect 88090 82550 88410 82750
rect 88480 82550 88520 82750
rect 88590 82550 88910 82750
rect 88980 82550 89020 82750
rect 89090 82550 89410 82750
rect 89480 82550 89520 82750
rect 89590 82550 89910 82750
rect 89980 82550 90020 82750
rect 90090 82550 90410 82750
rect 90480 82550 90520 82750
rect 90590 82550 90910 82750
rect 90980 82550 91020 82750
rect 91090 82550 91410 82750
rect 91480 82550 91520 82750
rect 91590 82550 91910 82750
rect 91980 82550 92020 82750
rect 92090 82550 92410 82750
rect 92480 82550 92520 82750
rect 92590 82550 92910 82750
rect 92980 82550 93020 82750
rect 93090 82550 93410 82750
rect 93480 82550 93520 82750
rect 93590 82550 93910 82750
rect 93980 82550 94020 82750
rect 94090 82550 94410 82750
rect 94480 82550 94520 82750
rect 94590 82550 94910 82750
rect 94980 82550 95020 82750
rect 95090 82550 95410 82750
rect 95480 82550 95520 82750
rect 95590 82550 95910 82750
rect 95980 82550 96020 82750
rect 96090 82550 96410 82750
rect 96480 82550 96520 82750
rect 96590 82550 96910 82750
rect 96980 82550 97020 82750
rect 97090 82550 97410 82750
rect 97480 82550 97520 82750
rect 97590 82550 97910 82750
rect 97980 82550 98020 82750
rect 98090 82550 98410 82750
rect 98480 82550 98520 82750
rect 98590 82550 98910 82750
rect 98980 82550 99020 82750
rect 99090 82550 99410 82750
rect 99480 82550 99520 82750
rect 99590 82550 99910 82750
rect 99980 82550 100020 82750
rect 100090 82550 100410 82750
rect 100480 82550 100500 82750
rect -83500 82540 100500 82550
rect -83360 82490 -83140 82540
rect -83360 82420 -83350 82490
rect -83150 82420 -83140 82490
rect -83360 82380 -83140 82420
rect -83360 82310 -83350 82380
rect -83150 82310 -83140 82380
rect -83360 82260 -83140 82310
rect -82860 82490 -82640 82540
rect -82860 82420 -82850 82490
rect -82650 82420 -82640 82490
rect -82860 82380 -82640 82420
rect -82860 82310 -82850 82380
rect -82650 82310 -82640 82380
rect -82860 82260 -82640 82310
rect -82360 82490 -82140 82540
rect -82360 82420 -82350 82490
rect -82150 82420 -82140 82490
rect -82360 82380 -82140 82420
rect -82360 82310 -82350 82380
rect -82150 82310 -82140 82380
rect -82360 82260 -82140 82310
rect -81860 82490 -81640 82540
rect -81860 82420 -81850 82490
rect -81650 82420 -81640 82490
rect -81860 82380 -81640 82420
rect -81860 82310 -81850 82380
rect -81650 82310 -81640 82380
rect -81860 82260 -81640 82310
rect -81360 82490 -81140 82540
rect -81360 82420 -81350 82490
rect -81150 82420 -81140 82490
rect -81360 82380 -81140 82420
rect -81360 82310 -81350 82380
rect -81150 82310 -81140 82380
rect -81360 82260 -81140 82310
rect -80860 82490 -80640 82540
rect -80860 82420 -80850 82490
rect -80650 82420 -80640 82490
rect -80860 82380 -80640 82420
rect -80860 82310 -80850 82380
rect -80650 82310 -80640 82380
rect -80860 82260 -80640 82310
rect -80360 82490 -80140 82540
rect -80360 82420 -80350 82490
rect -80150 82420 -80140 82490
rect -80360 82380 -80140 82420
rect -80360 82310 -80350 82380
rect -80150 82310 -80140 82380
rect -80360 82260 -80140 82310
rect -79860 82490 -79640 82540
rect -79860 82420 -79850 82490
rect -79650 82420 -79640 82490
rect -79860 82380 -79640 82420
rect -79860 82310 -79850 82380
rect -79650 82310 -79640 82380
rect -79860 82260 -79640 82310
rect -79360 82490 -79140 82540
rect -79360 82420 -79350 82490
rect -79150 82420 -79140 82490
rect -79360 82380 -79140 82420
rect -79360 82310 -79350 82380
rect -79150 82310 -79140 82380
rect -79360 82260 -79140 82310
rect -78860 82490 -78640 82540
rect -78860 82420 -78850 82490
rect -78650 82420 -78640 82490
rect -78860 82380 -78640 82420
rect -78860 82310 -78850 82380
rect -78650 82310 -78640 82380
rect -78860 82260 -78640 82310
rect -78360 82490 -78140 82540
rect -78360 82420 -78350 82490
rect -78150 82420 -78140 82490
rect -78360 82380 -78140 82420
rect -78360 82310 -78350 82380
rect -78150 82310 -78140 82380
rect -78360 82260 -78140 82310
rect -77860 82490 -77640 82540
rect -77860 82420 -77850 82490
rect -77650 82420 -77640 82490
rect -77860 82380 -77640 82420
rect -77860 82310 -77850 82380
rect -77650 82310 -77640 82380
rect -77860 82260 -77640 82310
rect -77360 82490 -77140 82540
rect -77360 82420 -77350 82490
rect -77150 82420 -77140 82490
rect -77360 82380 -77140 82420
rect -77360 82310 -77350 82380
rect -77150 82310 -77140 82380
rect -77360 82260 -77140 82310
rect -76860 82490 -76640 82540
rect -76860 82420 -76850 82490
rect -76650 82420 -76640 82490
rect -76860 82380 -76640 82420
rect -76860 82310 -76850 82380
rect -76650 82310 -76640 82380
rect -76860 82260 -76640 82310
rect -76360 82490 -76140 82540
rect -76360 82420 -76350 82490
rect -76150 82420 -76140 82490
rect -76360 82380 -76140 82420
rect -76360 82310 -76350 82380
rect -76150 82310 -76140 82380
rect -76360 82260 -76140 82310
rect -75860 82490 -75640 82540
rect -75860 82420 -75850 82490
rect -75650 82420 -75640 82490
rect -75860 82380 -75640 82420
rect -75860 82310 -75850 82380
rect -75650 82310 -75640 82380
rect -75860 82260 -75640 82310
rect -75360 82490 -75140 82540
rect -75360 82420 -75350 82490
rect -75150 82420 -75140 82490
rect -75360 82380 -75140 82420
rect -75360 82310 -75350 82380
rect -75150 82310 -75140 82380
rect -75360 82260 -75140 82310
rect -74860 82490 -74640 82540
rect -74860 82420 -74850 82490
rect -74650 82420 -74640 82490
rect -74860 82380 -74640 82420
rect -74860 82310 -74850 82380
rect -74650 82310 -74640 82380
rect -74860 82260 -74640 82310
rect -74360 82490 -74140 82540
rect -74360 82420 -74350 82490
rect -74150 82420 -74140 82490
rect -74360 82380 -74140 82420
rect -74360 82310 -74350 82380
rect -74150 82310 -74140 82380
rect -74360 82260 -74140 82310
rect -73860 82490 -73640 82540
rect -73860 82420 -73850 82490
rect -73650 82420 -73640 82490
rect -73860 82380 -73640 82420
rect -73860 82310 -73850 82380
rect -73650 82310 -73640 82380
rect -73860 82260 -73640 82310
rect -73360 82490 -73140 82540
rect -73360 82420 -73350 82490
rect -73150 82420 -73140 82490
rect -73360 82380 -73140 82420
rect -73360 82310 -73350 82380
rect -73150 82310 -73140 82380
rect -73360 82260 -73140 82310
rect -72860 82490 -72640 82540
rect -72860 82420 -72850 82490
rect -72650 82420 -72640 82490
rect -72860 82380 -72640 82420
rect -72860 82310 -72850 82380
rect -72650 82310 -72640 82380
rect -72860 82260 -72640 82310
rect -72360 82490 -72140 82540
rect -72360 82420 -72350 82490
rect -72150 82420 -72140 82490
rect -72360 82380 -72140 82420
rect -72360 82310 -72350 82380
rect -72150 82310 -72140 82380
rect -72360 82260 -72140 82310
rect -71860 82490 -71640 82540
rect -71860 82420 -71850 82490
rect -71650 82420 -71640 82490
rect -71860 82380 -71640 82420
rect -71860 82310 -71850 82380
rect -71650 82310 -71640 82380
rect -71860 82260 -71640 82310
rect -71360 82490 -71140 82540
rect -71360 82420 -71350 82490
rect -71150 82420 -71140 82490
rect -71360 82380 -71140 82420
rect -71360 82310 -71350 82380
rect -71150 82310 -71140 82380
rect -71360 82260 -71140 82310
rect -70860 82490 -70640 82540
rect -70860 82420 -70850 82490
rect -70650 82420 -70640 82490
rect -70860 82380 -70640 82420
rect -70860 82310 -70850 82380
rect -70650 82310 -70640 82380
rect -70860 82260 -70640 82310
rect -70360 82490 -70140 82540
rect -70360 82420 -70350 82490
rect -70150 82420 -70140 82490
rect -70360 82380 -70140 82420
rect -70360 82310 -70350 82380
rect -70150 82310 -70140 82380
rect -70360 82260 -70140 82310
rect -69860 82490 -69640 82540
rect -69860 82420 -69850 82490
rect -69650 82420 -69640 82490
rect -69860 82380 -69640 82420
rect -69860 82310 -69850 82380
rect -69650 82310 -69640 82380
rect -69860 82260 -69640 82310
rect -69360 82490 -69140 82540
rect -69360 82420 -69350 82490
rect -69150 82420 -69140 82490
rect -69360 82380 -69140 82420
rect -69360 82310 -69350 82380
rect -69150 82310 -69140 82380
rect -69360 82260 -69140 82310
rect -68860 82490 -68640 82540
rect -68860 82420 -68850 82490
rect -68650 82420 -68640 82490
rect -68860 82380 -68640 82420
rect -68860 82310 -68850 82380
rect -68650 82310 -68640 82380
rect -68860 82260 -68640 82310
rect -68360 82490 -68140 82540
rect -68360 82420 -68350 82490
rect -68150 82420 -68140 82490
rect -68360 82380 -68140 82420
rect -68360 82310 -68350 82380
rect -68150 82310 -68140 82380
rect -68360 82260 -68140 82310
rect -67860 82490 -67640 82540
rect -67860 82420 -67850 82490
rect -67650 82420 -67640 82490
rect -67860 82380 -67640 82420
rect -67860 82310 -67850 82380
rect -67650 82310 -67640 82380
rect -67860 82260 -67640 82310
rect -67360 82490 -67140 82540
rect -67360 82420 -67350 82490
rect -67150 82420 -67140 82490
rect -67360 82380 -67140 82420
rect -67360 82310 -67350 82380
rect -67150 82310 -67140 82380
rect -67360 82260 -67140 82310
rect -66860 82490 -66640 82540
rect -66860 82420 -66850 82490
rect -66650 82420 -66640 82490
rect -66860 82380 -66640 82420
rect -66860 82310 -66850 82380
rect -66650 82310 -66640 82380
rect -66860 82260 -66640 82310
rect -66360 82490 -66140 82540
rect -66360 82420 -66350 82490
rect -66150 82420 -66140 82490
rect -66360 82380 -66140 82420
rect -66360 82310 -66350 82380
rect -66150 82310 -66140 82380
rect -66360 82260 -66140 82310
rect -65860 82490 -65640 82540
rect -65860 82420 -65850 82490
rect -65650 82420 -65640 82490
rect -65860 82380 -65640 82420
rect -65860 82310 -65850 82380
rect -65650 82310 -65640 82380
rect -65860 82260 -65640 82310
rect -65360 82490 -65140 82540
rect -65360 82420 -65350 82490
rect -65150 82420 -65140 82490
rect -65360 82380 -65140 82420
rect -65360 82310 -65350 82380
rect -65150 82310 -65140 82380
rect -65360 82260 -65140 82310
rect -64860 82490 -64640 82540
rect -64860 82420 -64850 82490
rect -64650 82420 -64640 82490
rect -64860 82380 -64640 82420
rect -64860 82310 -64850 82380
rect -64650 82310 -64640 82380
rect -64860 82260 -64640 82310
rect -64360 82490 -64140 82540
rect -64360 82420 -64350 82490
rect -64150 82420 -64140 82490
rect -64360 82380 -64140 82420
rect -64360 82310 -64350 82380
rect -64150 82310 -64140 82380
rect -64360 82260 -64140 82310
rect -63860 82490 -63640 82540
rect -63860 82420 -63850 82490
rect -63650 82420 -63640 82490
rect -63860 82380 -63640 82420
rect -63860 82310 -63850 82380
rect -63650 82310 -63640 82380
rect -63860 82260 -63640 82310
rect -63360 82490 -63140 82540
rect -63360 82420 -63350 82490
rect -63150 82420 -63140 82490
rect -63360 82380 -63140 82420
rect -63360 82310 -63350 82380
rect -63150 82310 -63140 82380
rect -63360 82260 -63140 82310
rect -62860 82490 -62640 82540
rect -62860 82420 -62850 82490
rect -62650 82420 -62640 82490
rect -62860 82380 -62640 82420
rect -62860 82310 -62850 82380
rect -62650 82310 -62640 82380
rect -62860 82260 -62640 82310
rect -62360 82490 -62140 82540
rect -62360 82420 -62350 82490
rect -62150 82420 -62140 82490
rect -62360 82380 -62140 82420
rect -62360 82310 -62350 82380
rect -62150 82310 -62140 82380
rect -62360 82260 -62140 82310
rect -61860 82490 -61640 82540
rect -61860 82420 -61850 82490
rect -61650 82420 -61640 82490
rect -61860 82380 -61640 82420
rect -61860 82310 -61850 82380
rect -61650 82310 -61640 82380
rect -61860 82260 -61640 82310
rect -61360 82490 -61140 82540
rect -61360 82420 -61350 82490
rect -61150 82420 -61140 82490
rect -61360 82380 -61140 82420
rect -61360 82310 -61350 82380
rect -61150 82310 -61140 82380
rect -61360 82260 -61140 82310
rect -60860 82490 -60640 82540
rect -60860 82420 -60850 82490
rect -60650 82420 -60640 82490
rect -60860 82380 -60640 82420
rect -60860 82310 -60850 82380
rect -60650 82310 -60640 82380
rect -60860 82260 -60640 82310
rect -60360 82490 -60140 82540
rect -60360 82420 -60350 82490
rect -60150 82420 -60140 82490
rect -60360 82380 -60140 82420
rect -60360 82310 -60350 82380
rect -60150 82310 -60140 82380
rect -60360 82260 -60140 82310
rect -59860 82490 -59640 82540
rect -59860 82420 -59850 82490
rect -59650 82420 -59640 82490
rect -59860 82380 -59640 82420
rect -59860 82310 -59850 82380
rect -59650 82310 -59640 82380
rect -59860 82260 -59640 82310
rect -59360 82490 -59140 82540
rect -59360 82420 -59350 82490
rect -59150 82420 -59140 82490
rect -59360 82380 -59140 82420
rect -59360 82310 -59350 82380
rect -59150 82310 -59140 82380
rect -59360 82260 -59140 82310
rect -58860 82490 -58640 82540
rect -58860 82420 -58850 82490
rect -58650 82420 -58640 82490
rect -58860 82380 -58640 82420
rect -58860 82310 -58850 82380
rect -58650 82310 -58640 82380
rect -58860 82260 -58640 82310
rect -58360 82490 -58140 82540
rect -58360 82420 -58350 82490
rect -58150 82420 -58140 82490
rect -58360 82380 -58140 82420
rect -58360 82310 -58350 82380
rect -58150 82310 -58140 82380
rect -58360 82260 -58140 82310
rect -57860 82490 -57640 82540
rect -57860 82420 -57850 82490
rect -57650 82420 -57640 82490
rect -57860 82380 -57640 82420
rect -57860 82310 -57850 82380
rect -57650 82310 -57640 82380
rect -57860 82260 -57640 82310
rect -57360 82490 -57140 82540
rect -57360 82420 -57350 82490
rect -57150 82420 -57140 82490
rect -57360 82380 -57140 82420
rect -57360 82310 -57350 82380
rect -57150 82310 -57140 82380
rect -57360 82260 -57140 82310
rect -56860 82490 -56640 82540
rect -56860 82420 -56850 82490
rect -56650 82420 -56640 82490
rect -56860 82380 -56640 82420
rect -56860 82310 -56850 82380
rect -56650 82310 -56640 82380
rect -56860 82260 -56640 82310
rect -56360 82490 -56140 82540
rect -56360 82420 -56350 82490
rect -56150 82420 -56140 82490
rect -56360 82380 -56140 82420
rect -56360 82310 -56350 82380
rect -56150 82310 -56140 82380
rect -56360 82260 -56140 82310
rect -55860 82490 -55640 82540
rect -55860 82420 -55850 82490
rect -55650 82420 -55640 82490
rect -55860 82380 -55640 82420
rect -55860 82310 -55850 82380
rect -55650 82310 -55640 82380
rect -55860 82260 -55640 82310
rect -55360 82490 -55140 82540
rect -55360 82420 -55350 82490
rect -55150 82420 -55140 82490
rect -55360 82380 -55140 82420
rect -55360 82310 -55350 82380
rect -55150 82310 -55140 82380
rect -55360 82260 -55140 82310
rect -54860 82490 -54640 82540
rect -54860 82420 -54850 82490
rect -54650 82420 -54640 82490
rect -54860 82380 -54640 82420
rect -54860 82310 -54850 82380
rect -54650 82310 -54640 82380
rect -54860 82260 -54640 82310
rect -54360 82490 -54140 82540
rect -54360 82420 -54350 82490
rect -54150 82420 -54140 82490
rect -54360 82380 -54140 82420
rect -54360 82310 -54350 82380
rect -54150 82310 -54140 82380
rect -54360 82260 -54140 82310
rect -53860 82490 -53640 82540
rect -53860 82420 -53850 82490
rect -53650 82420 -53640 82490
rect -53860 82380 -53640 82420
rect -53860 82310 -53850 82380
rect -53650 82310 -53640 82380
rect -53860 82260 -53640 82310
rect -53360 82490 -53140 82540
rect -53360 82420 -53350 82490
rect -53150 82420 -53140 82490
rect -53360 82380 -53140 82420
rect -53360 82310 -53350 82380
rect -53150 82310 -53140 82380
rect -53360 82260 -53140 82310
rect -52860 82490 -52640 82540
rect -52860 82420 -52850 82490
rect -52650 82420 -52640 82490
rect -52860 82380 -52640 82420
rect -52860 82310 -52850 82380
rect -52650 82310 -52640 82380
rect -52860 82260 -52640 82310
rect -52360 82490 -52140 82540
rect -52360 82420 -52350 82490
rect -52150 82420 -52140 82490
rect -52360 82380 -52140 82420
rect -52360 82310 -52350 82380
rect -52150 82310 -52140 82380
rect -52360 82260 -52140 82310
rect -51860 82490 -51640 82540
rect -51860 82420 -51850 82490
rect -51650 82420 -51640 82490
rect -51860 82380 -51640 82420
rect -51860 82310 -51850 82380
rect -51650 82310 -51640 82380
rect -51860 82260 -51640 82310
rect -51360 82490 -51140 82540
rect -51360 82420 -51350 82490
rect -51150 82420 -51140 82490
rect -51360 82380 -51140 82420
rect -51360 82310 -51350 82380
rect -51150 82310 -51140 82380
rect -51360 82260 -51140 82310
rect -50860 82490 -50640 82540
rect -50860 82420 -50850 82490
rect -50650 82420 -50640 82490
rect -50860 82380 -50640 82420
rect -50860 82310 -50850 82380
rect -50650 82310 -50640 82380
rect -50860 82260 -50640 82310
rect -50360 82490 -50140 82540
rect -50360 82420 -50350 82490
rect -50150 82420 -50140 82490
rect -50360 82380 -50140 82420
rect -50360 82310 -50350 82380
rect -50150 82310 -50140 82380
rect -50360 82260 -50140 82310
rect -49860 82490 -49640 82540
rect -49860 82420 -49850 82490
rect -49650 82420 -49640 82490
rect -49860 82380 -49640 82420
rect -49860 82310 -49850 82380
rect -49650 82310 -49640 82380
rect -49860 82260 -49640 82310
rect -49360 82490 -49140 82540
rect -49360 82420 -49350 82490
rect -49150 82420 -49140 82490
rect -49360 82380 -49140 82420
rect -49360 82310 -49350 82380
rect -49150 82310 -49140 82380
rect -49360 82260 -49140 82310
rect -48860 82490 -48640 82540
rect -48860 82420 -48850 82490
rect -48650 82420 -48640 82490
rect -48860 82380 -48640 82420
rect -48860 82310 -48850 82380
rect -48650 82310 -48640 82380
rect -48860 82260 -48640 82310
rect -48360 82490 -48140 82540
rect -48360 82420 -48350 82490
rect -48150 82420 -48140 82490
rect -48360 82380 -48140 82420
rect -48360 82310 -48350 82380
rect -48150 82310 -48140 82380
rect -48360 82260 -48140 82310
rect -47860 82490 -47640 82540
rect -47860 82420 -47850 82490
rect -47650 82420 -47640 82490
rect -47860 82380 -47640 82420
rect -47860 82310 -47850 82380
rect -47650 82310 -47640 82380
rect -47860 82260 -47640 82310
rect -47360 82490 -47140 82540
rect -47360 82420 -47350 82490
rect -47150 82420 -47140 82490
rect -47360 82380 -47140 82420
rect -47360 82310 -47350 82380
rect -47150 82310 -47140 82380
rect -47360 82260 -47140 82310
rect -46860 82490 -46640 82540
rect -46860 82420 -46850 82490
rect -46650 82420 -46640 82490
rect -46860 82380 -46640 82420
rect -46860 82310 -46850 82380
rect -46650 82310 -46640 82380
rect -46860 82260 -46640 82310
rect -46360 82490 -46140 82540
rect -46360 82420 -46350 82490
rect -46150 82420 -46140 82490
rect -46360 82380 -46140 82420
rect -46360 82310 -46350 82380
rect -46150 82310 -46140 82380
rect -46360 82260 -46140 82310
rect -45860 82490 -45640 82540
rect -45860 82420 -45850 82490
rect -45650 82420 -45640 82490
rect -45860 82380 -45640 82420
rect -45860 82310 -45850 82380
rect -45650 82310 -45640 82380
rect -45860 82260 -45640 82310
rect -45360 82490 -45140 82540
rect -45360 82420 -45350 82490
rect -45150 82420 -45140 82490
rect -45360 82380 -45140 82420
rect -45360 82310 -45350 82380
rect -45150 82310 -45140 82380
rect -45360 82260 -45140 82310
rect -44860 82490 -44640 82540
rect -44860 82420 -44850 82490
rect -44650 82420 -44640 82490
rect -44860 82380 -44640 82420
rect -44860 82310 -44850 82380
rect -44650 82310 -44640 82380
rect -44860 82260 -44640 82310
rect -44360 82490 -44140 82540
rect -44360 82420 -44350 82490
rect -44150 82420 -44140 82490
rect -44360 82380 -44140 82420
rect -44360 82310 -44350 82380
rect -44150 82310 -44140 82380
rect -44360 82260 -44140 82310
rect -43860 82490 -43640 82540
rect -43860 82420 -43850 82490
rect -43650 82420 -43640 82490
rect -43860 82380 -43640 82420
rect -43860 82310 -43850 82380
rect -43650 82310 -43640 82380
rect -43860 82260 -43640 82310
rect -43360 82490 -43140 82540
rect -43360 82420 -43350 82490
rect -43150 82420 -43140 82490
rect -43360 82380 -43140 82420
rect -43360 82310 -43350 82380
rect -43150 82310 -43140 82380
rect -43360 82260 -43140 82310
rect -42860 82490 -42640 82540
rect -42860 82420 -42850 82490
rect -42650 82420 -42640 82490
rect -42860 82380 -42640 82420
rect -42860 82310 -42850 82380
rect -42650 82310 -42640 82380
rect -42860 82260 -42640 82310
rect -42360 82490 -42140 82540
rect -42360 82420 -42350 82490
rect -42150 82420 -42140 82490
rect -42360 82380 -42140 82420
rect -42360 82310 -42350 82380
rect -42150 82310 -42140 82380
rect -42360 82260 -42140 82310
rect -41860 82490 -41640 82540
rect -41860 82420 -41850 82490
rect -41650 82420 -41640 82490
rect -41860 82380 -41640 82420
rect -41860 82310 -41850 82380
rect -41650 82310 -41640 82380
rect -41860 82260 -41640 82310
rect -41360 82490 -41140 82540
rect -41360 82420 -41350 82490
rect -41150 82420 -41140 82490
rect -41360 82380 -41140 82420
rect -41360 82310 -41350 82380
rect -41150 82310 -41140 82380
rect -41360 82260 -41140 82310
rect -40860 82490 -40640 82540
rect -40860 82420 -40850 82490
rect -40650 82420 -40640 82490
rect -40860 82380 -40640 82420
rect -40860 82310 -40850 82380
rect -40650 82310 -40640 82380
rect -40860 82260 -40640 82310
rect -40360 82490 -40140 82540
rect -40360 82420 -40350 82490
rect -40150 82420 -40140 82490
rect -40360 82380 -40140 82420
rect -40360 82310 -40350 82380
rect -40150 82310 -40140 82380
rect -40360 82260 -40140 82310
rect -39860 82490 -39640 82540
rect -39860 82420 -39850 82490
rect -39650 82420 -39640 82490
rect -39860 82380 -39640 82420
rect -39860 82310 -39850 82380
rect -39650 82310 -39640 82380
rect -39860 82260 -39640 82310
rect -39360 82490 -39140 82540
rect -39360 82420 -39350 82490
rect -39150 82420 -39140 82490
rect -39360 82380 -39140 82420
rect -39360 82310 -39350 82380
rect -39150 82310 -39140 82380
rect -39360 82260 -39140 82310
rect -38860 82490 -38640 82540
rect -38860 82420 -38850 82490
rect -38650 82420 -38640 82490
rect -38860 82380 -38640 82420
rect -38860 82310 -38850 82380
rect -38650 82310 -38640 82380
rect -38860 82260 -38640 82310
rect -38360 82490 -38140 82540
rect -38360 82420 -38350 82490
rect -38150 82420 -38140 82490
rect -38360 82380 -38140 82420
rect -38360 82310 -38350 82380
rect -38150 82310 -38140 82380
rect -38360 82260 -38140 82310
rect -37860 82490 -37640 82540
rect -37860 82420 -37850 82490
rect -37650 82420 -37640 82490
rect -37860 82380 -37640 82420
rect -37860 82310 -37850 82380
rect -37650 82310 -37640 82380
rect -37860 82260 -37640 82310
rect -37360 82490 -37140 82540
rect -37360 82420 -37350 82490
rect -37150 82420 -37140 82490
rect -37360 82380 -37140 82420
rect -37360 82310 -37350 82380
rect -37150 82310 -37140 82380
rect -37360 82260 -37140 82310
rect -36860 82490 -36640 82540
rect -36860 82420 -36850 82490
rect -36650 82420 -36640 82490
rect -36860 82380 -36640 82420
rect -36860 82310 -36850 82380
rect -36650 82310 -36640 82380
rect -36860 82260 -36640 82310
rect -36360 82490 -36140 82540
rect -36360 82420 -36350 82490
rect -36150 82420 -36140 82490
rect -36360 82380 -36140 82420
rect -36360 82310 -36350 82380
rect -36150 82310 -36140 82380
rect -36360 82260 -36140 82310
rect -35860 82490 -35640 82540
rect -35860 82420 -35850 82490
rect -35650 82420 -35640 82490
rect -35860 82380 -35640 82420
rect -35860 82310 -35850 82380
rect -35650 82310 -35640 82380
rect -35860 82260 -35640 82310
rect -35360 82490 -35140 82540
rect -35360 82420 -35350 82490
rect -35150 82420 -35140 82490
rect -35360 82380 -35140 82420
rect -35360 82310 -35350 82380
rect -35150 82310 -35140 82380
rect -35360 82260 -35140 82310
rect -34860 82490 -34640 82540
rect -34860 82420 -34850 82490
rect -34650 82420 -34640 82490
rect -34860 82380 -34640 82420
rect -34860 82310 -34850 82380
rect -34650 82310 -34640 82380
rect -34860 82260 -34640 82310
rect -34360 82490 -34140 82540
rect -34360 82420 -34350 82490
rect -34150 82420 -34140 82490
rect -34360 82380 -34140 82420
rect -34360 82310 -34350 82380
rect -34150 82310 -34140 82380
rect -34360 82260 -34140 82310
rect -33860 82490 -33640 82540
rect -33860 82420 -33850 82490
rect -33650 82420 -33640 82490
rect -33860 82380 -33640 82420
rect -33860 82310 -33850 82380
rect -33650 82310 -33640 82380
rect -33860 82260 -33640 82310
rect -33360 82490 -33140 82540
rect -33360 82420 -33350 82490
rect -33150 82420 -33140 82490
rect -33360 82380 -33140 82420
rect -33360 82310 -33350 82380
rect -33150 82310 -33140 82380
rect -33360 82260 -33140 82310
rect -32860 82490 -32640 82540
rect -32860 82420 -32850 82490
rect -32650 82420 -32640 82490
rect -32860 82380 -32640 82420
rect -32860 82310 -32850 82380
rect -32650 82310 -32640 82380
rect -32860 82260 -32640 82310
rect -32360 82490 -32140 82540
rect -32360 82420 -32350 82490
rect -32150 82420 -32140 82490
rect -32360 82380 -32140 82420
rect -32360 82310 -32350 82380
rect -32150 82310 -32140 82380
rect -32360 82260 -32140 82310
rect -31860 82490 -31640 82540
rect -31860 82420 -31850 82490
rect -31650 82420 -31640 82490
rect -31860 82380 -31640 82420
rect -31860 82310 -31850 82380
rect -31650 82310 -31640 82380
rect -31860 82260 -31640 82310
rect -31360 82490 -31140 82540
rect -31360 82420 -31350 82490
rect -31150 82420 -31140 82490
rect -31360 82380 -31140 82420
rect -31360 82310 -31350 82380
rect -31150 82310 -31140 82380
rect -31360 82260 -31140 82310
rect -30860 82490 -30640 82540
rect -30860 82420 -30850 82490
rect -30650 82420 -30640 82490
rect -30860 82380 -30640 82420
rect -30860 82310 -30850 82380
rect -30650 82310 -30640 82380
rect -30860 82260 -30640 82310
rect -30360 82490 -30140 82540
rect -30360 82420 -30350 82490
rect -30150 82420 -30140 82490
rect -30360 82380 -30140 82420
rect -30360 82310 -30350 82380
rect -30150 82310 -30140 82380
rect -30360 82260 -30140 82310
rect -29860 82490 -29640 82540
rect -29860 82420 -29850 82490
rect -29650 82420 -29640 82490
rect -29860 82380 -29640 82420
rect -29860 82310 -29850 82380
rect -29650 82310 -29640 82380
rect -29860 82260 -29640 82310
rect -29360 82490 -29140 82540
rect -29360 82420 -29350 82490
rect -29150 82420 -29140 82490
rect -29360 82380 -29140 82420
rect -29360 82310 -29350 82380
rect -29150 82310 -29140 82380
rect -29360 82260 -29140 82310
rect -28860 82490 -28640 82540
rect -28860 82420 -28850 82490
rect -28650 82420 -28640 82490
rect -28860 82380 -28640 82420
rect -28860 82310 -28850 82380
rect -28650 82310 -28640 82380
rect -28860 82260 -28640 82310
rect -28360 82490 -28140 82540
rect -28360 82420 -28350 82490
rect -28150 82420 -28140 82490
rect -28360 82380 -28140 82420
rect -28360 82310 -28350 82380
rect -28150 82310 -28140 82380
rect -28360 82260 -28140 82310
rect -27860 82490 -27640 82540
rect -27860 82420 -27850 82490
rect -27650 82420 -27640 82490
rect -27860 82380 -27640 82420
rect -27860 82310 -27850 82380
rect -27650 82310 -27640 82380
rect -27860 82260 -27640 82310
rect -27360 82490 -27140 82540
rect -27360 82420 -27350 82490
rect -27150 82420 -27140 82490
rect -27360 82380 -27140 82420
rect -27360 82310 -27350 82380
rect -27150 82310 -27140 82380
rect -27360 82260 -27140 82310
rect -26860 82490 -26640 82540
rect -26860 82420 -26850 82490
rect -26650 82420 -26640 82490
rect -26860 82380 -26640 82420
rect -26860 82310 -26850 82380
rect -26650 82310 -26640 82380
rect -26860 82260 -26640 82310
rect -26360 82490 -26140 82540
rect -26360 82420 -26350 82490
rect -26150 82420 -26140 82490
rect -26360 82380 -26140 82420
rect -26360 82310 -26350 82380
rect -26150 82310 -26140 82380
rect -26360 82260 -26140 82310
rect -25860 82490 -25640 82540
rect -25860 82420 -25850 82490
rect -25650 82420 -25640 82490
rect -25860 82380 -25640 82420
rect -25860 82310 -25850 82380
rect -25650 82310 -25640 82380
rect -25860 82260 -25640 82310
rect -25360 82490 -25140 82540
rect -25360 82420 -25350 82490
rect -25150 82420 -25140 82490
rect -25360 82380 -25140 82420
rect -25360 82310 -25350 82380
rect -25150 82310 -25140 82380
rect -25360 82260 -25140 82310
rect -24860 82490 -24640 82540
rect -24860 82420 -24850 82490
rect -24650 82420 -24640 82490
rect -24860 82380 -24640 82420
rect -24860 82310 -24850 82380
rect -24650 82310 -24640 82380
rect -24860 82260 -24640 82310
rect -24360 82490 -24140 82540
rect -24360 82420 -24350 82490
rect -24150 82420 -24140 82490
rect -24360 82380 -24140 82420
rect -24360 82310 -24350 82380
rect -24150 82310 -24140 82380
rect -24360 82260 -24140 82310
rect -23860 82490 -23640 82540
rect -23860 82420 -23850 82490
rect -23650 82420 -23640 82490
rect -23860 82380 -23640 82420
rect -23860 82310 -23850 82380
rect -23650 82310 -23640 82380
rect -23860 82260 -23640 82310
rect -23360 82490 -23140 82540
rect -23360 82420 -23350 82490
rect -23150 82420 -23140 82490
rect -23360 82380 -23140 82420
rect -23360 82310 -23350 82380
rect -23150 82310 -23140 82380
rect -23360 82260 -23140 82310
rect -22860 82490 -22640 82540
rect -22860 82420 -22850 82490
rect -22650 82420 -22640 82490
rect -22860 82380 -22640 82420
rect -22860 82310 -22850 82380
rect -22650 82310 -22640 82380
rect -22860 82260 -22640 82310
rect -22360 82490 -22140 82540
rect -22360 82420 -22350 82490
rect -22150 82420 -22140 82490
rect -22360 82380 -22140 82420
rect -22360 82310 -22350 82380
rect -22150 82310 -22140 82380
rect -22360 82260 -22140 82310
rect -21860 82490 -21640 82540
rect -21860 82420 -21850 82490
rect -21650 82420 -21640 82490
rect -21860 82380 -21640 82420
rect -21860 82310 -21850 82380
rect -21650 82310 -21640 82380
rect -21860 82260 -21640 82310
rect -21360 82490 -21140 82540
rect -21360 82420 -21350 82490
rect -21150 82420 -21140 82490
rect -21360 82380 -21140 82420
rect -21360 82310 -21350 82380
rect -21150 82310 -21140 82380
rect -21360 82260 -21140 82310
rect -20860 82490 -20640 82540
rect -20860 82420 -20850 82490
rect -20650 82420 -20640 82490
rect -20860 82380 -20640 82420
rect -20860 82310 -20850 82380
rect -20650 82310 -20640 82380
rect -20860 82260 -20640 82310
rect -20360 82490 -20140 82540
rect -20360 82420 -20350 82490
rect -20150 82420 -20140 82490
rect -20360 82380 -20140 82420
rect -20360 82310 -20350 82380
rect -20150 82310 -20140 82380
rect -20360 82260 -20140 82310
rect -19860 82490 -19640 82540
rect -19860 82420 -19850 82490
rect -19650 82420 -19640 82490
rect -19860 82380 -19640 82420
rect -19860 82310 -19850 82380
rect -19650 82310 -19640 82380
rect -19860 82260 -19640 82310
rect -19360 82490 -19140 82540
rect -19360 82420 -19350 82490
rect -19150 82420 -19140 82490
rect -19360 82380 -19140 82420
rect -19360 82310 -19350 82380
rect -19150 82310 -19140 82380
rect -19360 82260 -19140 82310
rect -18860 82490 -18640 82540
rect -18860 82420 -18850 82490
rect -18650 82420 -18640 82490
rect -18860 82380 -18640 82420
rect -18860 82310 -18850 82380
rect -18650 82310 -18640 82380
rect -18860 82260 -18640 82310
rect -18360 82490 -18140 82540
rect -18360 82420 -18350 82490
rect -18150 82420 -18140 82490
rect -18360 82380 -18140 82420
rect -18360 82310 -18350 82380
rect -18150 82310 -18140 82380
rect -18360 82260 -18140 82310
rect -17860 82490 -17640 82540
rect -17860 82420 -17850 82490
rect -17650 82420 -17640 82490
rect -17860 82380 -17640 82420
rect -17860 82310 -17850 82380
rect -17650 82310 -17640 82380
rect -17860 82260 -17640 82310
rect -17360 82490 -17140 82540
rect -17360 82420 -17350 82490
rect -17150 82420 -17140 82490
rect -17360 82380 -17140 82420
rect -17360 82310 -17350 82380
rect -17150 82310 -17140 82380
rect -17360 82260 -17140 82310
rect -16860 82490 -16640 82540
rect -16860 82420 -16850 82490
rect -16650 82420 -16640 82490
rect -16860 82380 -16640 82420
rect -16860 82310 -16850 82380
rect -16650 82310 -16640 82380
rect -16860 82260 -16640 82310
rect -16360 82490 -16140 82540
rect -16360 82420 -16350 82490
rect -16150 82420 -16140 82490
rect -16360 82380 -16140 82420
rect -16360 82310 -16350 82380
rect -16150 82310 -16140 82380
rect -16360 82260 -16140 82310
rect -15860 82490 -15640 82540
rect -15860 82420 -15850 82490
rect -15650 82420 -15640 82490
rect -15860 82380 -15640 82420
rect -15860 82310 -15850 82380
rect -15650 82310 -15640 82380
rect -15860 82260 -15640 82310
rect -15360 82490 -15140 82540
rect -15360 82420 -15350 82490
rect -15150 82420 -15140 82490
rect -15360 82380 -15140 82420
rect -15360 82310 -15350 82380
rect -15150 82310 -15140 82380
rect -15360 82260 -15140 82310
rect -14860 82490 -14640 82540
rect -14860 82420 -14850 82490
rect -14650 82420 -14640 82490
rect -14860 82380 -14640 82420
rect -14860 82310 -14850 82380
rect -14650 82310 -14640 82380
rect -14860 82260 -14640 82310
rect -14360 82490 -14140 82540
rect -14360 82420 -14350 82490
rect -14150 82420 -14140 82490
rect -14360 82380 -14140 82420
rect -14360 82310 -14350 82380
rect -14150 82310 -14140 82380
rect -14360 82260 -14140 82310
rect -13860 82490 -13640 82540
rect -13860 82420 -13850 82490
rect -13650 82420 -13640 82490
rect -13860 82380 -13640 82420
rect -13860 82310 -13850 82380
rect -13650 82310 -13640 82380
rect -13860 82260 -13640 82310
rect -13360 82490 -13140 82540
rect -13360 82420 -13350 82490
rect -13150 82420 -13140 82490
rect -13360 82380 -13140 82420
rect -13360 82310 -13350 82380
rect -13150 82310 -13140 82380
rect -13360 82260 -13140 82310
rect -12860 82490 -12640 82540
rect -12860 82420 -12850 82490
rect -12650 82420 -12640 82490
rect -12860 82380 -12640 82420
rect -12860 82310 -12850 82380
rect -12650 82310 -12640 82380
rect -12860 82260 -12640 82310
rect -12360 82490 -12140 82540
rect -12360 82420 -12350 82490
rect -12150 82420 -12140 82490
rect -12360 82380 -12140 82420
rect -12360 82310 -12350 82380
rect -12150 82310 -12140 82380
rect -12360 82260 -12140 82310
rect -11860 82490 -11640 82540
rect -11860 82420 -11850 82490
rect -11650 82420 -11640 82490
rect -11860 82380 -11640 82420
rect -11860 82310 -11850 82380
rect -11650 82310 -11640 82380
rect -11860 82260 -11640 82310
rect -11360 82490 -11140 82540
rect -11360 82420 -11350 82490
rect -11150 82420 -11140 82490
rect -11360 82380 -11140 82420
rect -11360 82310 -11350 82380
rect -11150 82310 -11140 82380
rect -11360 82260 -11140 82310
rect -10860 82490 -10640 82540
rect -10860 82420 -10850 82490
rect -10650 82420 -10640 82490
rect -10860 82380 -10640 82420
rect -10860 82310 -10850 82380
rect -10650 82310 -10640 82380
rect -10860 82260 -10640 82310
rect -10360 82490 -10140 82540
rect -10360 82420 -10350 82490
rect -10150 82420 -10140 82490
rect -10360 82380 -10140 82420
rect -10360 82310 -10350 82380
rect -10150 82310 -10140 82380
rect -10360 82260 -10140 82310
rect -9860 82490 -9640 82540
rect -9860 82420 -9850 82490
rect -9650 82420 -9640 82490
rect -9860 82380 -9640 82420
rect -9860 82310 -9850 82380
rect -9650 82310 -9640 82380
rect -9860 82260 -9640 82310
rect -9360 82490 -9140 82540
rect -9360 82420 -9350 82490
rect -9150 82420 -9140 82490
rect -9360 82380 -9140 82420
rect -9360 82310 -9350 82380
rect -9150 82310 -9140 82380
rect -9360 82260 -9140 82310
rect -8860 82490 -8640 82540
rect -8860 82420 -8850 82490
rect -8650 82420 -8640 82490
rect -8860 82380 -8640 82420
rect -8860 82310 -8850 82380
rect -8650 82310 -8640 82380
rect -8860 82260 -8640 82310
rect -8360 82490 -8140 82540
rect -8360 82420 -8350 82490
rect -8150 82420 -8140 82490
rect -8360 82380 -8140 82420
rect -8360 82310 -8350 82380
rect -8150 82310 -8140 82380
rect -8360 82260 -8140 82310
rect -7860 82490 -7640 82540
rect -7860 82420 -7850 82490
rect -7650 82420 -7640 82490
rect -7860 82380 -7640 82420
rect -7860 82310 -7850 82380
rect -7650 82310 -7640 82380
rect -7860 82260 -7640 82310
rect -7360 82490 -7140 82540
rect -7360 82420 -7350 82490
rect -7150 82420 -7140 82490
rect -7360 82380 -7140 82420
rect -7360 82310 -7350 82380
rect -7150 82310 -7140 82380
rect -7360 82260 -7140 82310
rect -6860 82490 -6640 82540
rect -6860 82420 -6850 82490
rect -6650 82420 -6640 82490
rect -6860 82380 -6640 82420
rect -6860 82310 -6850 82380
rect -6650 82310 -6640 82380
rect -6860 82260 -6640 82310
rect -6360 82490 -6140 82540
rect -6360 82420 -6350 82490
rect -6150 82420 -6140 82490
rect -6360 82380 -6140 82420
rect -6360 82310 -6350 82380
rect -6150 82310 -6140 82380
rect -6360 82260 -6140 82310
rect -5860 82490 -5640 82540
rect -5860 82420 -5850 82490
rect -5650 82420 -5640 82490
rect -5860 82380 -5640 82420
rect -5860 82310 -5850 82380
rect -5650 82310 -5640 82380
rect -5860 82260 -5640 82310
rect -5360 82490 -5140 82540
rect -5360 82420 -5350 82490
rect -5150 82420 -5140 82490
rect -5360 82380 -5140 82420
rect -5360 82310 -5350 82380
rect -5150 82310 -5140 82380
rect -5360 82260 -5140 82310
rect -4860 82490 -4640 82540
rect -4860 82420 -4850 82490
rect -4650 82420 -4640 82490
rect -4860 82380 -4640 82420
rect -4860 82310 -4850 82380
rect -4650 82310 -4640 82380
rect -4860 82260 -4640 82310
rect -4360 82490 -4140 82540
rect -4360 82420 -4350 82490
rect -4150 82420 -4140 82490
rect -4360 82380 -4140 82420
rect -4360 82310 -4350 82380
rect -4150 82310 -4140 82380
rect -4360 82260 -4140 82310
rect -3860 82490 -3640 82540
rect -3860 82420 -3850 82490
rect -3650 82420 -3640 82490
rect -3860 82380 -3640 82420
rect -3860 82310 -3850 82380
rect -3650 82310 -3640 82380
rect -3860 82260 -3640 82310
rect -3360 82490 -3140 82540
rect -3360 82420 -3350 82490
rect -3150 82420 -3140 82490
rect -3360 82380 -3140 82420
rect -3360 82310 -3350 82380
rect -3150 82310 -3140 82380
rect -3360 82260 -3140 82310
rect -2860 82490 -2640 82540
rect -2860 82420 -2850 82490
rect -2650 82420 -2640 82490
rect -2860 82380 -2640 82420
rect -2860 82310 -2850 82380
rect -2650 82310 -2640 82380
rect -2860 82260 -2640 82310
rect -2360 82490 -2140 82540
rect -2360 82420 -2350 82490
rect -2150 82420 -2140 82490
rect -2360 82380 -2140 82420
rect -2360 82310 -2350 82380
rect -2150 82310 -2140 82380
rect -2360 82260 -2140 82310
rect -1860 82490 -1640 82540
rect -1860 82420 -1850 82490
rect -1650 82420 -1640 82490
rect -1860 82380 -1640 82420
rect -1860 82310 -1850 82380
rect -1650 82310 -1640 82380
rect -1860 82260 -1640 82310
rect -1360 82490 -1140 82540
rect -1360 82420 -1350 82490
rect -1150 82420 -1140 82490
rect -1360 82380 -1140 82420
rect -1360 82310 -1350 82380
rect -1150 82310 -1140 82380
rect -1360 82260 -1140 82310
rect -860 82490 -640 82540
rect -860 82420 -850 82490
rect -650 82420 -640 82490
rect -860 82380 -640 82420
rect -860 82310 -850 82380
rect -650 82310 -640 82380
rect -860 82260 -640 82310
rect -360 82490 -140 82540
rect -360 82420 -350 82490
rect -150 82420 -140 82490
rect -360 82380 -140 82420
rect -360 82310 -350 82380
rect -150 82310 -140 82380
rect -360 82260 -140 82310
rect 140 82490 360 82540
rect 140 82420 150 82490
rect 350 82420 360 82490
rect 140 82380 360 82420
rect 140 82310 150 82380
rect 350 82310 360 82380
rect 140 82260 360 82310
rect 640 82490 860 82540
rect 640 82420 650 82490
rect 850 82420 860 82490
rect 640 82380 860 82420
rect 640 82310 650 82380
rect 850 82310 860 82380
rect 640 82260 860 82310
rect 1140 82490 1360 82540
rect 1140 82420 1150 82490
rect 1350 82420 1360 82490
rect 1140 82380 1360 82420
rect 1140 82310 1150 82380
rect 1350 82310 1360 82380
rect 1140 82260 1360 82310
rect 1640 82490 1860 82540
rect 1640 82420 1650 82490
rect 1850 82420 1860 82490
rect 1640 82380 1860 82420
rect 1640 82310 1650 82380
rect 1850 82310 1860 82380
rect 1640 82260 1860 82310
rect 2140 82490 2360 82540
rect 2140 82420 2150 82490
rect 2350 82420 2360 82490
rect 2140 82380 2360 82420
rect 2140 82310 2150 82380
rect 2350 82310 2360 82380
rect 2140 82260 2360 82310
rect 2640 82490 2860 82540
rect 2640 82420 2650 82490
rect 2850 82420 2860 82490
rect 2640 82380 2860 82420
rect 2640 82310 2650 82380
rect 2850 82310 2860 82380
rect 2640 82260 2860 82310
rect 3140 82490 3360 82540
rect 3140 82420 3150 82490
rect 3350 82420 3360 82490
rect 3140 82380 3360 82420
rect 3140 82310 3150 82380
rect 3350 82310 3360 82380
rect 3140 82260 3360 82310
rect 3640 82490 3860 82540
rect 3640 82420 3650 82490
rect 3850 82420 3860 82490
rect 3640 82380 3860 82420
rect 3640 82310 3650 82380
rect 3850 82310 3860 82380
rect 3640 82260 3860 82310
rect 4140 82490 4360 82540
rect 4140 82420 4150 82490
rect 4350 82420 4360 82490
rect 4140 82380 4360 82420
rect 4140 82310 4150 82380
rect 4350 82310 4360 82380
rect 4140 82260 4360 82310
rect 4640 82490 4860 82540
rect 4640 82420 4650 82490
rect 4850 82420 4860 82490
rect 4640 82380 4860 82420
rect 4640 82310 4650 82380
rect 4850 82310 4860 82380
rect 4640 82260 4860 82310
rect 5140 82490 5360 82540
rect 5140 82420 5150 82490
rect 5350 82420 5360 82490
rect 5140 82380 5360 82420
rect 5140 82310 5150 82380
rect 5350 82310 5360 82380
rect 5140 82260 5360 82310
rect 5640 82490 5860 82540
rect 5640 82420 5650 82490
rect 5850 82420 5860 82490
rect 5640 82380 5860 82420
rect 5640 82310 5650 82380
rect 5850 82310 5860 82380
rect 5640 82260 5860 82310
rect 6140 82490 6360 82540
rect 6140 82420 6150 82490
rect 6350 82420 6360 82490
rect 6140 82380 6360 82420
rect 6140 82310 6150 82380
rect 6350 82310 6360 82380
rect 6140 82260 6360 82310
rect 6640 82490 6860 82540
rect 6640 82420 6650 82490
rect 6850 82420 6860 82490
rect 6640 82380 6860 82420
rect 6640 82310 6650 82380
rect 6850 82310 6860 82380
rect 6640 82260 6860 82310
rect 7140 82490 7360 82540
rect 7140 82420 7150 82490
rect 7350 82420 7360 82490
rect 7140 82380 7360 82420
rect 7140 82310 7150 82380
rect 7350 82310 7360 82380
rect 7140 82260 7360 82310
rect 7640 82490 7860 82540
rect 7640 82420 7650 82490
rect 7850 82420 7860 82490
rect 7640 82380 7860 82420
rect 7640 82310 7650 82380
rect 7850 82310 7860 82380
rect 7640 82260 7860 82310
rect 8140 82490 8360 82540
rect 8140 82420 8150 82490
rect 8350 82420 8360 82490
rect 8140 82380 8360 82420
rect 8140 82310 8150 82380
rect 8350 82310 8360 82380
rect 8140 82260 8360 82310
rect 8640 82490 8860 82540
rect 8640 82420 8650 82490
rect 8850 82420 8860 82490
rect 8640 82380 8860 82420
rect 8640 82310 8650 82380
rect 8850 82310 8860 82380
rect 8640 82260 8860 82310
rect 9140 82490 9360 82540
rect 9140 82420 9150 82490
rect 9350 82420 9360 82490
rect 9140 82380 9360 82420
rect 9140 82310 9150 82380
rect 9350 82310 9360 82380
rect 9140 82260 9360 82310
rect 9640 82490 9860 82540
rect 9640 82420 9650 82490
rect 9850 82420 9860 82490
rect 9640 82380 9860 82420
rect 9640 82310 9650 82380
rect 9850 82310 9860 82380
rect 9640 82260 9860 82310
rect 10140 82490 10360 82540
rect 10140 82420 10150 82490
rect 10350 82420 10360 82490
rect 10140 82380 10360 82420
rect 10140 82310 10150 82380
rect 10350 82310 10360 82380
rect 10140 82260 10360 82310
rect 10640 82490 10860 82540
rect 10640 82420 10650 82490
rect 10850 82420 10860 82490
rect 10640 82380 10860 82420
rect 10640 82310 10650 82380
rect 10850 82310 10860 82380
rect 10640 82260 10860 82310
rect 11140 82490 11360 82540
rect 11140 82420 11150 82490
rect 11350 82420 11360 82490
rect 11140 82380 11360 82420
rect 11140 82310 11150 82380
rect 11350 82310 11360 82380
rect 11140 82260 11360 82310
rect 11640 82490 11860 82540
rect 11640 82420 11650 82490
rect 11850 82420 11860 82490
rect 11640 82380 11860 82420
rect 11640 82310 11650 82380
rect 11850 82310 11860 82380
rect 11640 82260 11860 82310
rect 12140 82490 12360 82540
rect 12140 82420 12150 82490
rect 12350 82420 12360 82490
rect 12140 82380 12360 82420
rect 12140 82310 12150 82380
rect 12350 82310 12360 82380
rect 12140 82260 12360 82310
rect 12640 82490 12860 82540
rect 12640 82420 12650 82490
rect 12850 82420 12860 82490
rect 12640 82380 12860 82420
rect 12640 82310 12650 82380
rect 12850 82310 12860 82380
rect 12640 82260 12860 82310
rect 13140 82490 13360 82540
rect 13140 82420 13150 82490
rect 13350 82420 13360 82490
rect 13140 82380 13360 82420
rect 13140 82310 13150 82380
rect 13350 82310 13360 82380
rect 13140 82260 13360 82310
rect 13640 82490 13860 82540
rect 13640 82420 13650 82490
rect 13850 82420 13860 82490
rect 13640 82380 13860 82420
rect 13640 82310 13650 82380
rect 13850 82310 13860 82380
rect 13640 82260 13860 82310
rect 14140 82490 14360 82540
rect 14140 82420 14150 82490
rect 14350 82420 14360 82490
rect 14140 82380 14360 82420
rect 14140 82310 14150 82380
rect 14350 82310 14360 82380
rect 14140 82260 14360 82310
rect 14640 82490 14860 82540
rect 14640 82420 14650 82490
rect 14850 82420 14860 82490
rect 14640 82380 14860 82420
rect 14640 82310 14650 82380
rect 14850 82310 14860 82380
rect 14640 82260 14860 82310
rect 15140 82490 15360 82540
rect 15140 82420 15150 82490
rect 15350 82420 15360 82490
rect 15140 82380 15360 82420
rect 15140 82310 15150 82380
rect 15350 82310 15360 82380
rect 15140 82260 15360 82310
rect 15640 82490 15860 82540
rect 15640 82420 15650 82490
rect 15850 82420 15860 82490
rect 15640 82380 15860 82420
rect 15640 82310 15650 82380
rect 15850 82310 15860 82380
rect 15640 82260 15860 82310
rect 16140 82490 16360 82540
rect 16140 82420 16150 82490
rect 16350 82420 16360 82490
rect 16140 82380 16360 82420
rect 16140 82310 16150 82380
rect 16350 82310 16360 82380
rect 16140 82260 16360 82310
rect 16640 82490 16860 82540
rect 16640 82420 16650 82490
rect 16850 82420 16860 82490
rect 16640 82380 16860 82420
rect 16640 82310 16650 82380
rect 16850 82310 16860 82380
rect 16640 82260 16860 82310
rect 17140 82490 17360 82540
rect 17140 82420 17150 82490
rect 17350 82420 17360 82490
rect 17140 82380 17360 82420
rect 17140 82310 17150 82380
rect 17350 82310 17360 82380
rect 17140 82260 17360 82310
rect 17640 82490 17860 82540
rect 17640 82420 17650 82490
rect 17850 82420 17860 82490
rect 17640 82380 17860 82420
rect 17640 82310 17650 82380
rect 17850 82310 17860 82380
rect 17640 82260 17860 82310
rect 18140 82490 18360 82540
rect 18140 82420 18150 82490
rect 18350 82420 18360 82490
rect 18140 82380 18360 82420
rect 18140 82310 18150 82380
rect 18350 82310 18360 82380
rect 18140 82260 18360 82310
rect 18640 82490 18860 82540
rect 18640 82420 18650 82490
rect 18850 82420 18860 82490
rect 18640 82380 18860 82420
rect 18640 82310 18650 82380
rect 18850 82310 18860 82380
rect 18640 82260 18860 82310
rect 19140 82490 19360 82540
rect 19140 82420 19150 82490
rect 19350 82420 19360 82490
rect 19140 82380 19360 82420
rect 19140 82310 19150 82380
rect 19350 82310 19360 82380
rect 19140 82260 19360 82310
rect 19640 82490 19860 82540
rect 19640 82420 19650 82490
rect 19850 82420 19860 82490
rect 19640 82380 19860 82420
rect 19640 82310 19650 82380
rect 19850 82310 19860 82380
rect 19640 82260 19860 82310
rect 20140 82490 20360 82540
rect 20140 82420 20150 82490
rect 20350 82420 20360 82490
rect 20140 82380 20360 82420
rect 20140 82310 20150 82380
rect 20350 82310 20360 82380
rect 20140 82260 20360 82310
rect 20640 82490 20860 82540
rect 20640 82420 20650 82490
rect 20850 82420 20860 82490
rect 20640 82380 20860 82420
rect 20640 82310 20650 82380
rect 20850 82310 20860 82380
rect 20640 82260 20860 82310
rect 21140 82490 21360 82540
rect 21140 82420 21150 82490
rect 21350 82420 21360 82490
rect 21140 82380 21360 82420
rect 21140 82310 21150 82380
rect 21350 82310 21360 82380
rect 21140 82260 21360 82310
rect 21640 82490 21860 82540
rect 21640 82420 21650 82490
rect 21850 82420 21860 82490
rect 21640 82380 21860 82420
rect 21640 82310 21650 82380
rect 21850 82310 21860 82380
rect 21640 82260 21860 82310
rect 22140 82490 22360 82540
rect 22140 82420 22150 82490
rect 22350 82420 22360 82490
rect 22140 82380 22360 82420
rect 22140 82310 22150 82380
rect 22350 82310 22360 82380
rect 22140 82260 22360 82310
rect 22640 82490 22860 82540
rect 22640 82420 22650 82490
rect 22850 82420 22860 82490
rect 22640 82380 22860 82420
rect 22640 82310 22650 82380
rect 22850 82310 22860 82380
rect 22640 82260 22860 82310
rect 23140 82490 23360 82540
rect 23140 82420 23150 82490
rect 23350 82420 23360 82490
rect 23140 82380 23360 82420
rect 23140 82310 23150 82380
rect 23350 82310 23360 82380
rect 23140 82260 23360 82310
rect 23640 82490 23860 82540
rect 23640 82420 23650 82490
rect 23850 82420 23860 82490
rect 23640 82380 23860 82420
rect 23640 82310 23650 82380
rect 23850 82310 23860 82380
rect 23640 82260 23860 82310
rect 24140 82490 24360 82540
rect 24140 82420 24150 82490
rect 24350 82420 24360 82490
rect 24140 82380 24360 82420
rect 24140 82310 24150 82380
rect 24350 82310 24360 82380
rect 24140 82260 24360 82310
rect 24640 82490 24860 82540
rect 24640 82420 24650 82490
rect 24850 82420 24860 82490
rect 24640 82380 24860 82420
rect 24640 82310 24650 82380
rect 24850 82310 24860 82380
rect 24640 82260 24860 82310
rect 25140 82490 25360 82540
rect 25140 82420 25150 82490
rect 25350 82420 25360 82490
rect 25140 82380 25360 82420
rect 25140 82310 25150 82380
rect 25350 82310 25360 82380
rect 25140 82260 25360 82310
rect 25640 82490 25860 82540
rect 25640 82420 25650 82490
rect 25850 82420 25860 82490
rect 25640 82380 25860 82420
rect 25640 82310 25650 82380
rect 25850 82310 25860 82380
rect 25640 82260 25860 82310
rect 26140 82490 26360 82540
rect 26140 82420 26150 82490
rect 26350 82420 26360 82490
rect 26140 82380 26360 82420
rect 26140 82310 26150 82380
rect 26350 82310 26360 82380
rect 26140 82260 26360 82310
rect 26640 82490 26860 82540
rect 26640 82420 26650 82490
rect 26850 82420 26860 82490
rect 26640 82380 26860 82420
rect 26640 82310 26650 82380
rect 26850 82310 26860 82380
rect 26640 82260 26860 82310
rect 27140 82490 27360 82540
rect 27140 82420 27150 82490
rect 27350 82420 27360 82490
rect 27140 82380 27360 82420
rect 27140 82310 27150 82380
rect 27350 82310 27360 82380
rect 27140 82260 27360 82310
rect 27640 82490 27860 82540
rect 27640 82420 27650 82490
rect 27850 82420 27860 82490
rect 27640 82380 27860 82420
rect 27640 82310 27650 82380
rect 27850 82310 27860 82380
rect 27640 82260 27860 82310
rect 28140 82490 28360 82540
rect 28140 82420 28150 82490
rect 28350 82420 28360 82490
rect 28140 82380 28360 82420
rect 28140 82310 28150 82380
rect 28350 82310 28360 82380
rect 28140 82260 28360 82310
rect 28640 82490 28860 82540
rect 28640 82420 28650 82490
rect 28850 82420 28860 82490
rect 28640 82380 28860 82420
rect 28640 82310 28650 82380
rect 28850 82310 28860 82380
rect 28640 82260 28860 82310
rect 29140 82490 29360 82540
rect 29140 82420 29150 82490
rect 29350 82420 29360 82490
rect 29140 82380 29360 82420
rect 29140 82310 29150 82380
rect 29350 82310 29360 82380
rect 29140 82260 29360 82310
rect 29640 82490 29860 82540
rect 29640 82420 29650 82490
rect 29850 82420 29860 82490
rect 29640 82380 29860 82420
rect 29640 82310 29650 82380
rect 29850 82310 29860 82380
rect 29640 82260 29860 82310
rect 30140 82490 30360 82540
rect 30140 82420 30150 82490
rect 30350 82420 30360 82490
rect 30140 82380 30360 82420
rect 30140 82310 30150 82380
rect 30350 82310 30360 82380
rect 30140 82260 30360 82310
rect 30640 82490 30860 82540
rect 30640 82420 30650 82490
rect 30850 82420 30860 82490
rect 30640 82380 30860 82420
rect 30640 82310 30650 82380
rect 30850 82310 30860 82380
rect 30640 82260 30860 82310
rect 31140 82490 31360 82540
rect 31140 82420 31150 82490
rect 31350 82420 31360 82490
rect 31140 82380 31360 82420
rect 31140 82310 31150 82380
rect 31350 82310 31360 82380
rect 31140 82260 31360 82310
rect 31640 82490 31860 82540
rect 31640 82420 31650 82490
rect 31850 82420 31860 82490
rect 31640 82380 31860 82420
rect 31640 82310 31650 82380
rect 31850 82310 31860 82380
rect 31640 82260 31860 82310
rect 32140 82490 32360 82540
rect 32140 82420 32150 82490
rect 32350 82420 32360 82490
rect 32140 82380 32360 82420
rect 32140 82310 32150 82380
rect 32350 82310 32360 82380
rect 32140 82260 32360 82310
rect 32640 82490 32860 82540
rect 32640 82420 32650 82490
rect 32850 82420 32860 82490
rect 32640 82380 32860 82420
rect 32640 82310 32650 82380
rect 32850 82310 32860 82380
rect 32640 82260 32860 82310
rect 33140 82490 33360 82540
rect 33140 82420 33150 82490
rect 33350 82420 33360 82490
rect 33140 82380 33360 82420
rect 33140 82310 33150 82380
rect 33350 82310 33360 82380
rect 33140 82260 33360 82310
rect 33640 82490 33860 82540
rect 33640 82420 33650 82490
rect 33850 82420 33860 82490
rect 33640 82380 33860 82420
rect 33640 82310 33650 82380
rect 33850 82310 33860 82380
rect 33640 82260 33860 82310
rect 34140 82490 34360 82540
rect 34140 82420 34150 82490
rect 34350 82420 34360 82490
rect 34140 82380 34360 82420
rect 34140 82310 34150 82380
rect 34350 82310 34360 82380
rect 34140 82260 34360 82310
rect 34640 82490 34860 82540
rect 34640 82420 34650 82490
rect 34850 82420 34860 82490
rect 34640 82380 34860 82420
rect 34640 82310 34650 82380
rect 34850 82310 34860 82380
rect 34640 82260 34860 82310
rect 35140 82490 35360 82540
rect 35140 82420 35150 82490
rect 35350 82420 35360 82490
rect 35140 82380 35360 82420
rect 35140 82310 35150 82380
rect 35350 82310 35360 82380
rect 35140 82260 35360 82310
rect 35640 82490 35860 82540
rect 35640 82420 35650 82490
rect 35850 82420 35860 82490
rect 35640 82380 35860 82420
rect 35640 82310 35650 82380
rect 35850 82310 35860 82380
rect 35640 82260 35860 82310
rect 36140 82490 36360 82540
rect 36140 82420 36150 82490
rect 36350 82420 36360 82490
rect 36140 82380 36360 82420
rect 36140 82310 36150 82380
rect 36350 82310 36360 82380
rect 36140 82260 36360 82310
rect 36640 82490 36860 82540
rect 36640 82420 36650 82490
rect 36850 82420 36860 82490
rect 36640 82380 36860 82420
rect 36640 82310 36650 82380
rect 36850 82310 36860 82380
rect 36640 82260 36860 82310
rect 37140 82490 37360 82540
rect 37140 82420 37150 82490
rect 37350 82420 37360 82490
rect 37140 82380 37360 82420
rect 37140 82310 37150 82380
rect 37350 82310 37360 82380
rect 37140 82260 37360 82310
rect 37640 82490 37860 82540
rect 37640 82420 37650 82490
rect 37850 82420 37860 82490
rect 37640 82380 37860 82420
rect 37640 82310 37650 82380
rect 37850 82310 37860 82380
rect 37640 82260 37860 82310
rect 38140 82490 38360 82540
rect 38140 82420 38150 82490
rect 38350 82420 38360 82490
rect 38140 82380 38360 82420
rect 38140 82310 38150 82380
rect 38350 82310 38360 82380
rect 38140 82260 38360 82310
rect 38640 82490 38860 82540
rect 38640 82420 38650 82490
rect 38850 82420 38860 82490
rect 38640 82380 38860 82420
rect 38640 82310 38650 82380
rect 38850 82310 38860 82380
rect 38640 82260 38860 82310
rect 39140 82490 39360 82540
rect 39140 82420 39150 82490
rect 39350 82420 39360 82490
rect 39140 82380 39360 82420
rect 39140 82310 39150 82380
rect 39350 82310 39360 82380
rect 39140 82260 39360 82310
rect 39640 82490 39860 82540
rect 39640 82420 39650 82490
rect 39850 82420 39860 82490
rect 39640 82380 39860 82420
rect 39640 82310 39650 82380
rect 39850 82310 39860 82380
rect 39640 82260 39860 82310
rect 40140 82490 40360 82540
rect 40140 82420 40150 82490
rect 40350 82420 40360 82490
rect 40140 82380 40360 82420
rect 40140 82310 40150 82380
rect 40350 82310 40360 82380
rect 40140 82260 40360 82310
rect 40640 82490 40860 82540
rect 40640 82420 40650 82490
rect 40850 82420 40860 82490
rect 40640 82380 40860 82420
rect 40640 82310 40650 82380
rect 40850 82310 40860 82380
rect 40640 82260 40860 82310
rect 41140 82490 41360 82540
rect 41140 82420 41150 82490
rect 41350 82420 41360 82490
rect 41140 82380 41360 82420
rect 41140 82310 41150 82380
rect 41350 82310 41360 82380
rect 41140 82260 41360 82310
rect 41640 82490 41860 82540
rect 41640 82420 41650 82490
rect 41850 82420 41860 82490
rect 41640 82380 41860 82420
rect 41640 82310 41650 82380
rect 41850 82310 41860 82380
rect 41640 82260 41860 82310
rect 42140 82490 42360 82540
rect 42140 82420 42150 82490
rect 42350 82420 42360 82490
rect 42140 82380 42360 82420
rect 42140 82310 42150 82380
rect 42350 82310 42360 82380
rect 42140 82260 42360 82310
rect 42640 82490 42860 82540
rect 42640 82420 42650 82490
rect 42850 82420 42860 82490
rect 42640 82380 42860 82420
rect 42640 82310 42650 82380
rect 42850 82310 42860 82380
rect 42640 82260 42860 82310
rect 43140 82490 43360 82540
rect 43140 82420 43150 82490
rect 43350 82420 43360 82490
rect 43140 82380 43360 82420
rect 43140 82310 43150 82380
rect 43350 82310 43360 82380
rect 43140 82260 43360 82310
rect 43640 82490 43860 82540
rect 43640 82420 43650 82490
rect 43850 82420 43860 82490
rect 43640 82380 43860 82420
rect 43640 82310 43650 82380
rect 43850 82310 43860 82380
rect 43640 82260 43860 82310
rect 44140 82490 44360 82540
rect 44140 82420 44150 82490
rect 44350 82420 44360 82490
rect 44140 82380 44360 82420
rect 44140 82310 44150 82380
rect 44350 82310 44360 82380
rect 44140 82260 44360 82310
rect 44640 82490 44860 82540
rect 44640 82420 44650 82490
rect 44850 82420 44860 82490
rect 44640 82380 44860 82420
rect 44640 82310 44650 82380
rect 44850 82310 44860 82380
rect 44640 82260 44860 82310
rect 45140 82490 45360 82540
rect 45140 82420 45150 82490
rect 45350 82420 45360 82490
rect 45140 82380 45360 82420
rect 45140 82310 45150 82380
rect 45350 82310 45360 82380
rect 45140 82260 45360 82310
rect 45640 82490 45860 82540
rect 45640 82420 45650 82490
rect 45850 82420 45860 82490
rect 45640 82380 45860 82420
rect 45640 82310 45650 82380
rect 45850 82310 45860 82380
rect 45640 82260 45860 82310
rect 46140 82490 46360 82540
rect 46140 82420 46150 82490
rect 46350 82420 46360 82490
rect 46140 82380 46360 82420
rect 46140 82310 46150 82380
rect 46350 82310 46360 82380
rect 46140 82260 46360 82310
rect 46640 82490 46860 82540
rect 46640 82420 46650 82490
rect 46850 82420 46860 82490
rect 46640 82380 46860 82420
rect 46640 82310 46650 82380
rect 46850 82310 46860 82380
rect 46640 82260 46860 82310
rect 47140 82490 47360 82540
rect 47140 82420 47150 82490
rect 47350 82420 47360 82490
rect 47140 82380 47360 82420
rect 47140 82310 47150 82380
rect 47350 82310 47360 82380
rect 47140 82260 47360 82310
rect 47640 82490 47860 82540
rect 47640 82420 47650 82490
rect 47850 82420 47860 82490
rect 47640 82380 47860 82420
rect 47640 82310 47650 82380
rect 47850 82310 47860 82380
rect 47640 82260 47860 82310
rect 48140 82490 48360 82540
rect 48140 82420 48150 82490
rect 48350 82420 48360 82490
rect 48140 82380 48360 82420
rect 48140 82310 48150 82380
rect 48350 82310 48360 82380
rect 48140 82260 48360 82310
rect 48640 82490 48860 82540
rect 48640 82420 48650 82490
rect 48850 82420 48860 82490
rect 48640 82380 48860 82420
rect 48640 82310 48650 82380
rect 48850 82310 48860 82380
rect 48640 82260 48860 82310
rect 49140 82490 49360 82540
rect 49140 82420 49150 82490
rect 49350 82420 49360 82490
rect 49140 82380 49360 82420
rect 49140 82310 49150 82380
rect 49350 82310 49360 82380
rect 49140 82260 49360 82310
rect 49640 82490 49860 82540
rect 49640 82420 49650 82490
rect 49850 82420 49860 82490
rect 49640 82380 49860 82420
rect 49640 82310 49650 82380
rect 49850 82310 49860 82380
rect 49640 82260 49860 82310
rect 50140 82490 50360 82540
rect 50140 82420 50150 82490
rect 50350 82420 50360 82490
rect 50140 82380 50360 82420
rect 50140 82310 50150 82380
rect 50350 82310 50360 82380
rect 50140 82260 50360 82310
rect 50640 82490 50860 82540
rect 50640 82420 50650 82490
rect 50850 82420 50860 82490
rect 50640 82380 50860 82420
rect 50640 82310 50650 82380
rect 50850 82310 50860 82380
rect 50640 82260 50860 82310
rect 51140 82490 51360 82540
rect 51140 82420 51150 82490
rect 51350 82420 51360 82490
rect 51140 82380 51360 82420
rect 51140 82310 51150 82380
rect 51350 82310 51360 82380
rect 51140 82260 51360 82310
rect 51640 82490 51860 82540
rect 51640 82420 51650 82490
rect 51850 82420 51860 82490
rect 51640 82380 51860 82420
rect 51640 82310 51650 82380
rect 51850 82310 51860 82380
rect 51640 82260 51860 82310
rect 52140 82490 52360 82540
rect 52140 82420 52150 82490
rect 52350 82420 52360 82490
rect 52140 82380 52360 82420
rect 52140 82310 52150 82380
rect 52350 82310 52360 82380
rect 52140 82260 52360 82310
rect 52640 82490 52860 82540
rect 52640 82420 52650 82490
rect 52850 82420 52860 82490
rect 52640 82380 52860 82420
rect 52640 82310 52650 82380
rect 52850 82310 52860 82380
rect 52640 82260 52860 82310
rect 53140 82490 53360 82540
rect 53140 82420 53150 82490
rect 53350 82420 53360 82490
rect 53140 82380 53360 82420
rect 53140 82310 53150 82380
rect 53350 82310 53360 82380
rect 53140 82260 53360 82310
rect 53640 82490 53860 82540
rect 53640 82420 53650 82490
rect 53850 82420 53860 82490
rect 53640 82380 53860 82420
rect 53640 82310 53650 82380
rect 53850 82310 53860 82380
rect 53640 82260 53860 82310
rect 54140 82490 54360 82540
rect 54140 82420 54150 82490
rect 54350 82420 54360 82490
rect 54140 82380 54360 82420
rect 54140 82310 54150 82380
rect 54350 82310 54360 82380
rect 54140 82260 54360 82310
rect 54640 82490 54860 82540
rect 54640 82420 54650 82490
rect 54850 82420 54860 82490
rect 54640 82380 54860 82420
rect 54640 82310 54650 82380
rect 54850 82310 54860 82380
rect 54640 82260 54860 82310
rect 55140 82490 55360 82540
rect 55140 82420 55150 82490
rect 55350 82420 55360 82490
rect 55140 82380 55360 82420
rect 55140 82310 55150 82380
rect 55350 82310 55360 82380
rect 55140 82260 55360 82310
rect 55640 82490 55860 82540
rect 55640 82420 55650 82490
rect 55850 82420 55860 82490
rect 55640 82380 55860 82420
rect 55640 82310 55650 82380
rect 55850 82310 55860 82380
rect 55640 82260 55860 82310
rect 56140 82490 56360 82540
rect 56140 82420 56150 82490
rect 56350 82420 56360 82490
rect 56140 82380 56360 82420
rect 56140 82310 56150 82380
rect 56350 82310 56360 82380
rect 56140 82260 56360 82310
rect 56640 82490 56860 82540
rect 56640 82420 56650 82490
rect 56850 82420 56860 82490
rect 56640 82380 56860 82420
rect 56640 82310 56650 82380
rect 56850 82310 56860 82380
rect 56640 82260 56860 82310
rect 57140 82490 57360 82540
rect 57140 82420 57150 82490
rect 57350 82420 57360 82490
rect 57140 82380 57360 82420
rect 57140 82310 57150 82380
rect 57350 82310 57360 82380
rect 57140 82260 57360 82310
rect 57640 82490 57860 82540
rect 57640 82420 57650 82490
rect 57850 82420 57860 82490
rect 57640 82380 57860 82420
rect 57640 82310 57650 82380
rect 57850 82310 57860 82380
rect 57640 82260 57860 82310
rect 58140 82490 58360 82540
rect 58140 82420 58150 82490
rect 58350 82420 58360 82490
rect 58140 82380 58360 82420
rect 58140 82310 58150 82380
rect 58350 82310 58360 82380
rect 58140 82260 58360 82310
rect 58640 82490 58860 82540
rect 58640 82420 58650 82490
rect 58850 82420 58860 82490
rect 58640 82380 58860 82420
rect 58640 82310 58650 82380
rect 58850 82310 58860 82380
rect 58640 82260 58860 82310
rect 59140 82490 59360 82540
rect 59140 82420 59150 82490
rect 59350 82420 59360 82490
rect 59140 82380 59360 82420
rect 59140 82310 59150 82380
rect 59350 82310 59360 82380
rect 59140 82260 59360 82310
rect 59640 82490 59860 82540
rect 59640 82420 59650 82490
rect 59850 82420 59860 82490
rect 59640 82380 59860 82420
rect 59640 82310 59650 82380
rect 59850 82310 59860 82380
rect 59640 82260 59860 82310
rect 60140 82490 60360 82540
rect 60140 82420 60150 82490
rect 60350 82420 60360 82490
rect 60140 82380 60360 82420
rect 60140 82310 60150 82380
rect 60350 82310 60360 82380
rect 60140 82260 60360 82310
rect 60640 82490 60860 82540
rect 60640 82420 60650 82490
rect 60850 82420 60860 82490
rect 60640 82380 60860 82420
rect 60640 82310 60650 82380
rect 60850 82310 60860 82380
rect 60640 82260 60860 82310
rect 61140 82490 61360 82540
rect 61140 82420 61150 82490
rect 61350 82420 61360 82490
rect 61140 82380 61360 82420
rect 61140 82310 61150 82380
rect 61350 82310 61360 82380
rect 61140 82260 61360 82310
rect 61640 82490 61860 82540
rect 61640 82420 61650 82490
rect 61850 82420 61860 82490
rect 61640 82380 61860 82420
rect 61640 82310 61650 82380
rect 61850 82310 61860 82380
rect 61640 82260 61860 82310
rect 62140 82490 62360 82540
rect 62140 82420 62150 82490
rect 62350 82420 62360 82490
rect 62140 82380 62360 82420
rect 62140 82310 62150 82380
rect 62350 82310 62360 82380
rect 62140 82260 62360 82310
rect 62640 82490 62860 82540
rect 62640 82420 62650 82490
rect 62850 82420 62860 82490
rect 62640 82380 62860 82420
rect 62640 82310 62650 82380
rect 62850 82310 62860 82380
rect 62640 82260 62860 82310
rect 63140 82490 63360 82540
rect 63140 82420 63150 82490
rect 63350 82420 63360 82490
rect 63140 82380 63360 82420
rect 63140 82310 63150 82380
rect 63350 82310 63360 82380
rect 63140 82260 63360 82310
rect 63640 82490 63860 82540
rect 63640 82420 63650 82490
rect 63850 82420 63860 82490
rect 63640 82380 63860 82420
rect 63640 82310 63650 82380
rect 63850 82310 63860 82380
rect 63640 82260 63860 82310
rect 64140 82490 64360 82540
rect 64140 82420 64150 82490
rect 64350 82420 64360 82490
rect 64140 82380 64360 82420
rect 64140 82310 64150 82380
rect 64350 82310 64360 82380
rect 64140 82260 64360 82310
rect 64640 82490 64860 82540
rect 64640 82420 64650 82490
rect 64850 82420 64860 82490
rect 64640 82380 64860 82420
rect 64640 82310 64650 82380
rect 64850 82310 64860 82380
rect 64640 82260 64860 82310
rect 65140 82490 65360 82540
rect 65140 82420 65150 82490
rect 65350 82420 65360 82490
rect 65140 82380 65360 82420
rect 65140 82310 65150 82380
rect 65350 82310 65360 82380
rect 65140 82260 65360 82310
rect 65640 82490 65860 82540
rect 65640 82420 65650 82490
rect 65850 82420 65860 82490
rect 65640 82380 65860 82420
rect 65640 82310 65650 82380
rect 65850 82310 65860 82380
rect 65640 82260 65860 82310
rect 66140 82490 66360 82540
rect 66140 82420 66150 82490
rect 66350 82420 66360 82490
rect 66140 82380 66360 82420
rect 66140 82310 66150 82380
rect 66350 82310 66360 82380
rect 66140 82260 66360 82310
rect 66640 82490 66860 82540
rect 66640 82420 66650 82490
rect 66850 82420 66860 82490
rect 66640 82380 66860 82420
rect 66640 82310 66650 82380
rect 66850 82310 66860 82380
rect 66640 82260 66860 82310
rect 67140 82490 67360 82540
rect 67140 82420 67150 82490
rect 67350 82420 67360 82490
rect 67140 82380 67360 82420
rect 67140 82310 67150 82380
rect 67350 82310 67360 82380
rect 67140 82260 67360 82310
rect 67640 82490 67860 82540
rect 67640 82420 67650 82490
rect 67850 82420 67860 82490
rect 67640 82380 67860 82420
rect 67640 82310 67650 82380
rect 67850 82310 67860 82380
rect 67640 82260 67860 82310
rect 68140 82490 68360 82540
rect 68140 82420 68150 82490
rect 68350 82420 68360 82490
rect 68140 82380 68360 82420
rect 68140 82310 68150 82380
rect 68350 82310 68360 82380
rect 68140 82260 68360 82310
rect 68640 82490 68860 82540
rect 68640 82420 68650 82490
rect 68850 82420 68860 82490
rect 68640 82380 68860 82420
rect 68640 82310 68650 82380
rect 68850 82310 68860 82380
rect 68640 82260 68860 82310
rect 69140 82490 69360 82540
rect 69140 82420 69150 82490
rect 69350 82420 69360 82490
rect 69140 82380 69360 82420
rect 69140 82310 69150 82380
rect 69350 82310 69360 82380
rect 69140 82260 69360 82310
rect 69640 82490 69860 82540
rect 69640 82420 69650 82490
rect 69850 82420 69860 82490
rect 69640 82380 69860 82420
rect 69640 82310 69650 82380
rect 69850 82310 69860 82380
rect 69640 82260 69860 82310
rect 70140 82490 70360 82540
rect 70140 82420 70150 82490
rect 70350 82420 70360 82490
rect 70140 82380 70360 82420
rect 70140 82310 70150 82380
rect 70350 82310 70360 82380
rect 70140 82260 70360 82310
rect 70640 82490 70860 82540
rect 70640 82420 70650 82490
rect 70850 82420 70860 82490
rect 70640 82380 70860 82420
rect 70640 82310 70650 82380
rect 70850 82310 70860 82380
rect 70640 82260 70860 82310
rect 71140 82490 71360 82540
rect 71140 82420 71150 82490
rect 71350 82420 71360 82490
rect 71140 82380 71360 82420
rect 71140 82310 71150 82380
rect 71350 82310 71360 82380
rect 71140 82260 71360 82310
rect 71640 82490 71860 82540
rect 71640 82420 71650 82490
rect 71850 82420 71860 82490
rect 71640 82380 71860 82420
rect 71640 82310 71650 82380
rect 71850 82310 71860 82380
rect 71640 82260 71860 82310
rect 72140 82490 72360 82540
rect 72140 82420 72150 82490
rect 72350 82420 72360 82490
rect 72140 82380 72360 82420
rect 72140 82310 72150 82380
rect 72350 82310 72360 82380
rect 72140 82260 72360 82310
rect 72640 82490 72860 82540
rect 72640 82420 72650 82490
rect 72850 82420 72860 82490
rect 72640 82380 72860 82420
rect 72640 82310 72650 82380
rect 72850 82310 72860 82380
rect 72640 82260 72860 82310
rect 73140 82490 73360 82540
rect 73140 82420 73150 82490
rect 73350 82420 73360 82490
rect 73140 82380 73360 82420
rect 73140 82310 73150 82380
rect 73350 82310 73360 82380
rect 73140 82260 73360 82310
rect 73640 82490 73860 82540
rect 73640 82420 73650 82490
rect 73850 82420 73860 82490
rect 73640 82380 73860 82420
rect 73640 82310 73650 82380
rect 73850 82310 73860 82380
rect 73640 82260 73860 82310
rect 74140 82490 74360 82540
rect 74140 82420 74150 82490
rect 74350 82420 74360 82490
rect 74140 82380 74360 82420
rect 74140 82310 74150 82380
rect 74350 82310 74360 82380
rect 74140 82260 74360 82310
rect 74640 82490 74860 82540
rect 74640 82420 74650 82490
rect 74850 82420 74860 82490
rect 74640 82380 74860 82420
rect 74640 82310 74650 82380
rect 74850 82310 74860 82380
rect 74640 82260 74860 82310
rect 75140 82490 75360 82540
rect 75140 82420 75150 82490
rect 75350 82420 75360 82490
rect 75140 82380 75360 82420
rect 75140 82310 75150 82380
rect 75350 82310 75360 82380
rect 75140 82260 75360 82310
rect 75640 82490 75860 82540
rect 75640 82420 75650 82490
rect 75850 82420 75860 82490
rect 75640 82380 75860 82420
rect 75640 82310 75650 82380
rect 75850 82310 75860 82380
rect 75640 82260 75860 82310
rect 76140 82490 76360 82540
rect 76140 82420 76150 82490
rect 76350 82420 76360 82490
rect 76140 82380 76360 82420
rect 76140 82310 76150 82380
rect 76350 82310 76360 82380
rect 76140 82260 76360 82310
rect 76640 82490 76860 82540
rect 76640 82420 76650 82490
rect 76850 82420 76860 82490
rect 76640 82380 76860 82420
rect 76640 82310 76650 82380
rect 76850 82310 76860 82380
rect 76640 82260 76860 82310
rect 77140 82490 77360 82540
rect 77140 82420 77150 82490
rect 77350 82420 77360 82490
rect 77140 82380 77360 82420
rect 77140 82310 77150 82380
rect 77350 82310 77360 82380
rect 77140 82260 77360 82310
rect 77640 82490 77860 82540
rect 77640 82420 77650 82490
rect 77850 82420 77860 82490
rect 77640 82380 77860 82420
rect 77640 82310 77650 82380
rect 77850 82310 77860 82380
rect 77640 82260 77860 82310
rect 78140 82490 78360 82540
rect 78140 82420 78150 82490
rect 78350 82420 78360 82490
rect 78140 82380 78360 82420
rect 78140 82310 78150 82380
rect 78350 82310 78360 82380
rect 78140 82260 78360 82310
rect 78640 82490 78860 82540
rect 78640 82420 78650 82490
rect 78850 82420 78860 82490
rect 78640 82380 78860 82420
rect 78640 82310 78650 82380
rect 78850 82310 78860 82380
rect 78640 82260 78860 82310
rect 79140 82490 79360 82540
rect 79140 82420 79150 82490
rect 79350 82420 79360 82490
rect 79140 82380 79360 82420
rect 79140 82310 79150 82380
rect 79350 82310 79360 82380
rect 79140 82260 79360 82310
rect 79640 82490 79860 82540
rect 79640 82420 79650 82490
rect 79850 82420 79860 82490
rect 79640 82380 79860 82420
rect 79640 82310 79650 82380
rect 79850 82310 79860 82380
rect 79640 82260 79860 82310
rect 80140 82490 80360 82540
rect 80140 82420 80150 82490
rect 80350 82420 80360 82490
rect 80140 82380 80360 82420
rect 80140 82310 80150 82380
rect 80350 82310 80360 82380
rect 80140 82260 80360 82310
rect 80640 82490 80860 82540
rect 80640 82420 80650 82490
rect 80850 82420 80860 82490
rect 80640 82380 80860 82420
rect 80640 82310 80650 82380
rect 80850 82310 80860 82380
rect 80640 82260 80860 82310
rect 81140 82490 81360 82540
rect 81140 82420 81150 82490
rect 81350 82420 81360 82490
rect 81140 82380 81360 82420
rect 81140 82310 81150 82380
rect 81350 82310 81360 82380
rect 81140 82260 81360 82310
rect 81640 82490 81860 82540
rect 81640 82420 81650 82490
rect 81850 82420 81860 82490
rect 81640 82380 81860 82420
rect 81640 82310 81650 82380
rect 81850 82310 81860 82380
rect 81640 82260 81860 82310
rect 82140 82490 82360 82540
rect 82140 82420 82150 82490
rect 82350 82420 82360 82490
rect 82140 82380 82360 82420
rect 82140 82310 82150 82380
rect 82350 82310 82360 82380
rect 82140 82260 82360 82310
rect 82640 82490 82860 82540
rect 82640 82420 82650 82490
rect 82850 82420 82860 82490
rect 82640 82380 82860 82420
rect 82640 82310 82650 82380
rect 82850 82310 82860 82380
rect 82640 82260 82860 82310
rect 83140 82490 83360 82540
rect 83140 82420 83150 82490
rect 83350 82420 83360 82490
rect 83140 82380 83360 82420
rect 83140 82310 83150 82380
rect 83350 82310 83360 82380
rect 83140 82260 83360 82310
rect 83640 82490 83860 82540
rect 83640 82420 83650 82490
rect 83850 82420 83860 82490
rect 83640 82380 83860 82420
rect 83640 82310 83650 82380
rect 83850 82310 83860 82380
rect 83640 82260 83860 82310
rect 84140 82490 84360 82540
rect 84140 82420 84150 82490
rect 84350 82420 84360 82490
rect 84140 82380 84360 82420
rect 84140 82310 84150 82380
rect 84350 82310 84360 82380
rect 84140 82260 84360 82310
rect 84640 82490 84860 82540
rect 84640 82420 84650 82490
rect 84850 82420 84860 82490
rect 84640 82380 84860 82420
rect 84640 82310 84650 82380
rect 84850 82310 84860 82380
rect 84640 82260 84860 82310
rect 85140 82490 85360 82540
rect 85140 82420 85150 82490
rect 85350 82420 85360 82490
rect 85140 82380 85360 82420
rect 85140 82310 85150 82380
rect 85350 82310 85360 82380
rect 85140 82260 85360 82310
rect 85640 82490 85860 82540
rect 85640 82420 85650 82490
rect 85850 82420 85860 82490
rect 85640 82380 85860 82420
rect 85640 82310 85650 82380
rect 85850 82310 85860 82380
rect 85640 82260 85860 82310
rect 86140 82490 86360 82540
rect 86140 82420 86150 82490
rect 86350 82420 86360 82490
rect 86140 82380 86360 82420
rect 86140 82310 86150 82380
rect 86350 82310 86360 82380
rect 86140 82260 86360 82310
rect 86640 82490 86860 82540
rect 86640 82420 86650 82490
rect 86850 82420 86860 82490
rect 86640 82380 86860 82420
rect 86640 82310 86650 82380
rect 86850 82310 86860 82380
rect 86640 82260 86860 82310
rect 87140 82490 87360 82540
rect 87140 82420 87150 82490
rect 87350 82420 87360 82490
rect 87140 82380 87360 82420
rect 87140 82310 87150 82380
rect 87350 82310 87360 82380
rect 87140 82260 87360 82310
rect 87640 82490 87860 82540
rect 87640 82420 87650 82490
rect 87850 82420 87860 82490
rect 87640 82380 87860 82420
rect 87640 82310 87650 82380
rect 87850 82310 87860 82380
rect 87640 82260 87860 82310
rect 88140 82490 88360 82540
rect 88140 82420 88150 82490
rect 88350 82420 88360 82490
rect 88140 82380 88360 82420
rect 88140 82310 88150 82380
rect 88350 82310 88360 82380
rect 88140 82260 88360 82310
rect 88640 82490 88860 82540
rect 88640 82420 88650 82490
rect 88850 82420 88860 82490
rect 88640 82380 88860 82420
rect 88640 82310 88650 82380
rect 88850 82310 88860 82380
rect 88640 82260 88860 82310
rect 89140 82490 89360 82540
rect 89140 82420 89150 82490
rect 89350 82420 89360 82490
rect 89140 82380 89360 82420
rect 89140 82310 89150 82380
rect 89350 82310 89360 82380
rect 89140 82260 89360 82310
rect 89640 82490 89860 82540
rect 89640 82420 89650 82490
rect 89850 82420 89860 82490
rect 89640 82380 89860 82420
rect 89640 82310 89650 82380
rect 89850 82310 89860 82380
rect 89640 82260 89860 82310
rect 90140 82490 90360 82540
rect 90140 82420 90150 82490
rect 90350 82420 90360 82490
rect 90140 82380 90360 82420
rect 90140 82310 90150 82380
rect 90350 82310 90360 82380
rect 90140 82260 90360 82310
rect 90640 82490 90860 82540
rect 90640 82420 90650 82490
rect 90850 82420 90860 82490
rect 90640 82380 90860 82420
rect 90640 82310 90650 82380
rect 90850 82310 90860 82380
rect 90640 82260 90860 82310
rect 91140 82490 91360 82540
rect 91140 82420 91150 82490
rect 91350 82420 91360 82490
rect 91140 82380 91360 82420
rect 91140 82310 91150 82380
rect 91350 82310 91360 82380
rect 91140 82260 91360 82310
rect 91640 82490 91860 82540
rect 91640 82420 91650 82490
rect 91850 82420 91860 82490
rect 91640 82380 91860 82420
rect 91640 82310 91650 82380
rect 91850 82310 91860 82380
rect 91640 82260 91860 82310
rect 92140 82490 92360 82540
rect 92140 82420 92150 82490
rect 92350 82420 92360 82490
rect 92140 82380 92360 82420
rect 92140 82310 92150 82380
rect 92350 82310 92360 82380
rect 92140 82260 92360 82310
rect 92640 82490 92860 82540
rect 92640 82420 92650 82490
rect 92850 82420 92860 82490
rect 92640 82380 92860 82420
rect 92640 82310 92650 82380
rect 92850 82310 92860 82380
rect 92640 82260 92860 82310
rect 93140 82490 93360 82540
rect 93140 82420 93150 82490
rect 93350 82420 93360 82490
rect 93140 82380 93360 82420
rect 93140 82310 93150 82380
rect 93350 82310 93360 82380
rect 93140 82260 93360 82310
rect 93640 82490 93860 82540
rect 93640 82420 93650 82490
rect 93850 82420 93860 82490
rect 93640 82380 93860 82420
rect 93640 82310 93650 82380
rect 93850 82310 93860 82380
rect 93640 82260 93860 82310
rect 94140 82490 94360 82540
rect 94140 82420 94150 82490
rect 94350 82420 94360 82490
rect 94140 82380 94360 82420
rect 94140 82310 94150 82380
rect 94350 82310 94360 82380
rect 94140 82260 94360 82310
rect 94640 82490 94860 82540
rect 94640 82420 94650 82490
rect 94850 82420 94860 82490
rect 94640 82380 94860 82420
rect 94640 82310 94650 82380
rect 94850 82310 94860 82380
rect 94640 82260 94860 82310
rect 95140 82490 95360 82540
rect 95140 82420 95150 82490
rect 95350 82420 95360 82490
rect 95140 82380 95360 82420
rect 95140 82310 95150 82380
rect 95350 82310 95360 82380
rect 95140 82260 95360 82310
rect 95640 82490 95860 82540
rect 95640 82420 95650 82490
rect 95850 82420 95860 82490
rect 95640 82380 95860 82420
rect 95640 82310 95650 82380
rect 95850 82310 95860 82380
rect 95640 82260 95860 82310
rect 96140 82490 96360 82540
rect 96140 82420 96150 82490
rect 96350 82420 96360 82490
rect 96140 82380 96360 82420
rect 96140 82310 96150 82380
rect 96350 82310 96360 82380
rect 96140 82260 96360 82310
rect 96640 82490 96860 82540
rect 96640 82420 96650 82490
rect 96850 82420 96860 82490
rect 96640 82380 96860 82420
rect 96640 82310 96650 82380
rect 96850 82310 96860 82380
rect 96640 82260 96860 82310
rect 97140 82490 97360 82540
rect 97140 82420 97150 82490
rect 97350 82420 97360 82490
rect 97140 82380 97360 82420
rect 97140 82310 97150 82380
rect 97350 82310 97360 82380
rect 97140 82260 97360 82310
rect 97640 82490 97860 82540
rect 97640 82420 97650 82490
rect 97850 82420 97860 82490
rect 97640 82380 97860 82420
rect 97640 82310 97650 82380
rect 97850 82310 97860 82380
rect 97640 82260 97860 82310
rect 98140 82490 98360 82540
rect 98140 82420 98150 82490
rect 98350 82420 98360 82490
rect 98140 82380 98360 82420
rect 98140 82310 98150 82380
rect 98350 82310 98360 82380
rect 98140 82260 98360 82310
rect 98640 82490 98860 82540
rect 98640 82420 98650 82490
rect 98850 82420 98860 82490
rect 98640 82380 98860 82420
rect 98640 82310 98650 82380
rect 98850 82310 98860 82380
rect 98640 82260 98860 82310
rect 99140 82490 99360 82540
rect 99140 82420 99150 82490
rect 99350 82420 99360 82490
rect 99140 82380 99360 82420
rect 99140 82310 99150 82380
rect 99350 82310 99360 82380
rect 99140 82260 99360 82310
rect 99640 82490 99860 82540
rect 99640 82420 99650 82490
rect 99850 82420 99860 82490
rect 99640 82380 99860 82420
rect 99640 82310 99650 82380
rect 99850 82310 99860 82380
rect 99640 82260 99860 82310
rect 100140 82490 100360 82540
rect 100140 82420 100150 82490
rect 100350 82420 100360 82490
rect 100140 82380 100360 82420
rect 100140 82310 100150 82380
rect 100350 82310 100360 82380
rect 100140 82260 100360 82310
rect -83500 82250 100500 82260
rect -83500 82050 -83480 82250
rect -83410 82050 -83090 82250
rect -83020 82050 -82980 82250
rect -82910 82050 -82590 82250
rect -82520 82050 -82480 82250
rect -82410 82050 -82090 82250
rect -82020 82050 -81980 82250
rect -81910 82050 -81590 82250
rect -81520 82050 -81480 82250
rect -81410 82050 -81090 82250
rect -81020 82050 -80980 82250
rect -80910 82050 -80590 82250
rect -80520 82050 -80480 82250
rect -80410 82050 -80090 82250
rect -80020 82050 -79980 82250
rect -79910 82050 -79590 82250
rect -79520 82050 -79480 82250
rect -79410 82050 -79090 82250
rect -79020 82050 -78980 82250
rect -78910 82050 -78590 82250
rect -78520 82050 -78480 82250
rect -78410 82050 -78090 82250
rect -78020 82050 -77980 82250
rect -77910 82050 -77590 82250
rect -77520 82050 -77480 82250
rect -77410 82050 -77090 82250
rect -77020 82050 -76980 82250
rect -76910 82050 -76590 82250
rect -76520 82050 -76480 82250
rect -76410 82050 -76090 82250
rect -76020 82050 -75980 82250
rect -75910 82050 -75590 82250
rect -75520 82050 -75480 82250
rect -75410 82050 -75090 82250
rect -75020 82050 -74980 82250
rect -74910 82050 -74590 82250
rect -74520 82050 -74480 82250
rect -74410 82050 -74090 82250
rect -74020 82050 -73980 82250
rect -73910 82050 -73590 82250
rect -73520 82050 -73480 82250
rect -73410 82050 -73090 82250
rect -73020 82050 -72980 82250
rect -72910 82050 -72590 82250
rect -72520 82050 -72480 82250
rect -72410 82050 -72090 82250
rect -72020 82050 -71980 82250
rect -71910 82050 -71590 82250
rect -71520 82050 -71480 82250
rect -71410 82050 -71090 82250
rect -71020 82050 -70980 82250
rect -70910 82050 -70590 82250
rect -70520 82050 -70480 82250
rect -70410 82050 -70090 82250
rect -70020 82050 -69980 82250
rect -69910 82050 -69590 82250
rect -69520 82050 -69480 82250
rect -69410 82050 -69090 82250
rect -69020 82050 -68980 82250
rect -68910 82050 -68590 82250
rect -68520 82050 -68480 82250
rect -68410 82050 -68090 82250
rect -68020 82050 -67980 82250
rect -67910 82050 -67590 82250
rect -67520 82050 -67480 82250
rect -67410 82050 -67090 82250
rect -67020 82050 -66980 82250
rect -66910 82050 -66590 82250
rect -66520 82050 -66480 82250
rect -66410 82050 -66090 82250
rect -66020 82050 -65980 82250
rect -65910 82050 -65590 82250
rect -65520 82050 -65480 82250
rect -65410 82050 -65090 82250
rect -65020 82050 -64980 82250
rect -64910 82050 -64590 82250
rect -64520 82050 -64480 82250
rect -64410 82050 -64090 82250
rect -64020 82050 -63980 82250
rect -63910 82050 -63590 82250
rect -63520 82050 -63480 82250
rect -63410 82050 -63090 82250
rect -63020 82050 -62980 82250
rect -62910 82050 -62590 82250
rect -62520 82050 -62480 82250
rect -62410 82050 -62090 82250
rect -62020 82050 -61980 82250
rect -61910 82050 -61590 82250
rect -61520 82050 -61480 82250
rect -61410 82050 -61090 82250
rect -61020 82050 -60980 82250
rect -60910 82050 -60590 82250
rect -60520 82050 -60480 82250
rect -60410 82050 -60090 82250
rect -60020 82050 -59980 82250
rect -59910 82050 -59590 82250
rect -59520 82050 -59480 82250
rect -59410 82050 -59090 82250
rect -59020 82050 -58980 82250
rect -58910 82050 -58590 82250
rect -58520 82050 -58480 82250
rect -58410 82050 -58090 82250
rect -58020 82050 -57980 82250
rect -57910 82050 -57590 82250
rect -57520 82050 -57480 82250
rect -57410 82050 -57090 82250
rect -57020 82050 -56980 82250
rect -56910 82050 -56590 82250
rect -56520 82050 -56480 82250
rect -56410 82050 -56090 82250
rect -56020 82050 -55980 82250
rect -55910 82050 -55590 82250
rect -55520 82050 -55480 82250
rect -55410 82050 -55090 82250
rect -55020 82050 -54980 82250
rect -54910 82050 -54590 82250
rect -54520 82050 -54480 82250
rect -54410 82050 -54090 82250
rect -54020 82050 -53980 82250
rect -53910 82050 -53590 82250
rect -53520 82050 -53480 82250
rect -53410 82050 -53090 82250
rect -53020 82050 -52980 82250
rect -52910 82050 -52590 82250
rect -52520 82050 -52480 82250
rect -52410 82050 -52090 82250
rect -52020 82050 -51980 82250
rect -51910 82050 -51590 82250
rect -51520 82050 -51480 82250
rect -51410 82050 -51090 82250
rect -51020 82050 -50980 82250
rect -50910 82050 -50590 82250
rect -50520 82050 -50480 82250
rect -50410 82050 -50090 82250
rect -50020 82050 -49980 82250
rect -49910 82050 -49590 82250
rect -49520 82050 -49480 82250
rect -49410 82050 -49090 82250
rect -49020 82050 -48980 82250
rect -48910 82050 -48590 82250
rect -48520 82050 -48480 82250
rect -48410 82050 -48090 82250
rect -48020 82050 -47980 82250
rect -47910 82050 -47590 82250
rect -47520 82050 -47480 82250
rect -47410 82050 -47090 82250
rect -47020 82050 -46980 82250
rect -46910 82050 -46590 82250
rect -46520 82050 -46480 82250
rect -46410 82050 -46090 82250
rect -46020 82050 -45980 82250
rect -45910 82050 -45590 82250
rect -45520 82050 -45480 82250
rect -45410 82050 -45090 82250
rect -45020 82050 -44980 82250
rect -44910 82050 -44590 82250
rect -44520 82050 -44480 82250
rect -44410 82050 -44090 82250
rect -44020 82050 -43980 82250
rect -43910 82050 -43590 82250
rect -43520 82050 -43480 82250
rect -43410 82050 -43090 82250
rect -43020 82050 -42980 82250
rect -42910 82050 -42590 82250
rect -42520 82050 -42480 82250
rect -42410 82050 -42090 82250
rect -42020 82050 -41980 82250
rect -41910 82050 -41590 82250
rect -41520 82050 -41480 82250
rect -41410 82050 -41090 82250
rect -41020 82050 -40980 82250
rect -40910 82050 -40590 82250
rect -40520 82050 -40480 82250
rect -40410 82050 -40090 82250
rect -40020 82050 -39980 82250
rect -39910 82050 -39590 82250
rect -39520 82050 -39480 82250
rect -39410 82050 -39090 82250
rect -39020 82050 -38980 82250
rect -38910 82050 -38590 82250
rect -38520 82050 -38480 82250
rect -38410 82050 -38090 82250
rect -38020 82050 -37980 82250
rect -37910 82050 -37590 82250
rect -37520 82050 -37480 82250
rect -37410 82050 -37090 82250
rect -37020 82050 -36980 82250
rect -36910 82050 -36590 82250
rect -36520 82050 -36480 82250
rect -36410 82050 -36090 82250
rect -36020 82050 -35980 82250
rect -35910 82050 -35590 82250
rect -35520 82050 -35480 82250
rect -35410 82050 -35090 82250
rect -35020 82050 -34980 82250
rect -34910 82050 -34590 82250
rect -34520 82050 -34480 82250
rect -34410 82050 -34090 82250
rect -34020 82050 -33980 82250
rect -33910 82050 -33590 82250
rect -33520 82050 -33480 82250
rect -33410 82050 -33090 82250
rect -33020 82050 -32980 82250
rect -32910 82050 -32590 82250
rect -32520 82050 -32480 82250
rect -32410 82050 -32090 82250
rect -32020 82050 -31980 82250
rect -31910 82050 -31590 82250
rect -31520 82050 -31480 82250
rect -31410 82050 -31090 82250
rect -31020 82050 -30980 82250
rect -30910 82050 -30590 82250
rect -30520 82050 -30480 82250
rect -30410 82050 -30090 82250
rect -30020 82050 -29980 82250
rect -29910 82050 -29590 82250
rect -29520 82050 -29480 82250
rect -29410 82050 -29090 82250
rect -29020 82050 -28980 82250
rect -28910 82050 -28590 82250
rect -28520 82050 -28480 82250
rect -28410 82050 -28090 82250
rect -28020 82050 -27980 82250
rect -27910 82050 -27590 82250
rect -27520 82050 -27480 82250
rect -27410 82050 -27090 82250
rect -27020 82050 -26980 82250
rect -26910 82050 -26590 82250
rect -26520 82050 -26480 82250
rect -26410 82050 -26090 82250
rect -26020 82050 -25980 82250
rect -25910 82050 -25590 82250
rect -25520 82050 -25480 82250
rect -25410 82050 -25090 82250
rect -25020 82050 -24980 82250
rect -24910 82050 -24590 82250
rect -24520 82050 -24480 82250
rect -24410 82050 -24090 82250
rect -24020 82050 -23980 82250
rect -23910 82050 -23590 82250
rect -23520 82050 -23480 82250
rect -23410 82050 -23090 82250
rect -23020 82050 -22980 82250
rect -22910 82050 -22590 82250
rect -22520 82050 -22480 82250
rect -22410 82050 -22090 82250
rect -22020 82050 -21980 82250
rect -21910 82050 -21590 82250
rect -21520 82050 -21480 82250
rect -21410 82050 -21090 82250
rect -21020 82050 -20980 82250
rect -20910 82050 -20590 82250
rect -20520 82050 -20480 82250
rect -20410 82050 -20090 82250
rect -20020 82050 -19980 82250
rect -19910 82050 -19590 82250
rect -19520 82050 -19480 82250
rect -19410 82050 -19090 82250
rect -19020 82050 -18980 82250
rect -18910 82050 -18590 82250
rect -18520 82050 -18480 82250
rect -18410 82050 -18090 82250
rect -18020 82050 -17980 82250
rect -17910 82050 -17590 82250
rect -17520 82050 -17480 82250
rect -17410 82050 -17090 82250
rect -17020 82050 -16980 82250
rect -16910 82050 -16590 82250
rect -16520 82050 -16480 82250
rect -16410 82050 -16090 82250
rect -16020 82050 -15980 82250
rect -15910 82050 -15590 82250
rect -15520 82050 -15480 82250
rect -15410 82050 -15090 82250
rect -15020 82050 -14980 82250
rect -14910 82050 -14590 82250
rect -14520 82050 -14480 82250
rect -14410 82050 -14090 82250
rect -14020 82050 -13980 82250
rect -13910 82050 -13590 82250
rect -13520 82050 -13480 82250
rect -13410 82050 -13090 82250
rect -13020 82050 -12980 82250
rect -12910 82050 -12590 82250
rect -12520 82050 -12480 82250
rect -12410 82050 -12090 82250
rect -12020 82050 -11980 82250
rect -11910 82050 -11590 82250
rect -11520 82050 -11480 82250
rect -11410 82050 -11090 82250
rect -11020 82050 -10980 82250
rect -10910 82050 -10590 82250
rect -10520 82050 -10480 82250
rect -10410 82050 -10090 82250
rect -10020 82050 -9980 82250
rect -9910 82050 -9590 82250
rect -9520 82050 -9480 82250
rect -9410 82050 -9090 82250
rect -9020 82050 -8980 82250
rect -8910 82050 -8590 82250
rect -8520 82050 -8480 82250
rect -8410 82050 -8090 82250
rect -8020 82050 -7980 82250
rect -7910 82050 -7590 82250
rect -7520 82050 -7480 82250
rect -7410 82050 -7090 82250
rect -7020 82050 -6980 82250
rect -6910 82050 -6590 82250
rect -6520 82050 -6480 82250
rect -6410 82050 -6090 82250
rect -6020 82050 -5980 82250
rect -5910 82050 -5590 82250
rect -5520 82050 -5480 82250
rect -5410 82050 -5090 82250
rect -5020 82050 -4980 82250
rect -4910 82050 -4590 82250
rect -4520 82050 -4480 82250
rect -4410 82050 -4090 82250
rect -4020 82050 -3980 82250
rect -3910 82050 -3590 82250
rect -3520 82050 -3480 82250
rect -3410 82050 -3090 82250
rect -3020 82050 -2980 82250
rect -2910 82050 -2590 82250
rect -2520 82050 -2480 82250
rect -2410 82050 -2090 82250
rect -2020 82050 -1980 82250
rect -1910 82050 -1590 82250
rect -1520 82050 -1480 82250
rect -1410 82050 -1090 82250
rect -1020 82050 -980 82250
rect -910 82050 -590 82250
rect -520 82050 -480 82250
rect -410 82050 -90 82250
rect -20 82050 20 82250
rect 90 82050 410 82250
rect 480 82050 520 82250
rect 590 82050 910 82250
rect 980 82050 1020 82250
rect 1090 82050 1410 82250
rect 1480 82050 1520 82250
rect 1590 82050 1910 82250
rect 1980 82050 2020 82250
rect 2090 82050 2410 82250
rect 2480 82050 2520 82250
rect 2590 82050 2910 82250
rect 2980 82050 3020 82250
rect 3090 82050 3410 82250
rect 3480 82050 3520 82250
rect 3590 82050 3910 82250
rect 3980 82050 4020 82250
rect 4090 82050 4410 82250
rect 4480 82050 4520 82250
rect 4590 82050 4910 82250
rect 4980 82050 5020 82250
rect 5090 82050 5410 82250
rect 5480 82050 5520 82250
rect 5590 82050 5910 82250
rect 5980 82050 6020 82250
rect 6090 82050 6410 82250
rect 6480 82050 6520 82250
rect 6590 82050 6910 82250
rect 6980 82050 7020 82250
rect 7090 82050 7410 82250
rect 7480 82050 7520 82250
rect 7590 82050 7910 82250
rect 7980 82050 8020 82250
rect 8090 82050 8410 82250
rect 8480 82050 8520 82250
rect 8590 82050 8910 82250
rect 8980 82050 9020 82250
rect 9090 82050 9410 82250
rect 9480 82050 9520 82250
rect 9590 82050 9910 82250
rect 9980 82050 10020 82250
rect 10090 82050 10410 82250
rect 10480 82050 10520 82250
rect 10590 82050 10910 82250
rect 10980 82050 11020 82250
rect 11090 82050 11410 82250
rect 11480 82050 11520 82250
rect 11590 82050 11910 82250
rect 11980 82050 12020 82250
rect 12090 82050 12410 82250
rect 12480 82050 12520 82250
rect 12590 82050 12910 82250
rect 12980 82050 13020 82250
rect 13090 82050 13410 82250
rect 13480 82050 13520 82250
rect 13590 82050 13910 82250
rect 13980 82050 14020 82250
rect 14090 82050 14410 82250
rect 14480 82050 14520 82250
rect 14590 82050 14910 82250
rect 14980 82050 15020 82250
rect 15090 82050 15410 82250
rect 15480 82050 15520 82250
rect 15590 82050 15910 82250
rect 15980 82050 16020 82250
rect 16090 82050 16410 82250
rect 16480 82050 16520 82250
rect 16590 82050 16910 82250
rect 16980 82050 17020 82250
rect 17090 82050 17410 82250
rect 17480 82050 17520 82250
rect 17590 82050 17910 82250
rect 17980 82050 18020 82250
rect 18090 82050 18410 82250
rect 18480 82050 18520 82250
rect 18590 82050 18910 82250
rect 18980 82050 19020 82250
rect 19090 82050 19410 82250
rect 19480 82050 19520 82250
rect 19590 82050 19910 82250
rect 19980 82050 20020 82250
rect 20090 82050 20410 82250
rect 20480 82050 20520 82250
rect 20590 82050 20910 82250
rect 20980 82050 21020 82250
rect 21090 82050 21410 82250
rect 21480 82050 21520 82250
rect 21590 82050 21910 82250
rect 21980 82050 22020 82250
rect 22090 82050 22410 82250
rect 22480 82050 22520 82250
rect 22590 82050 22910 82250
rect 22980 82050 23020 82250
rect 23090 82050 23410 82250
rect 23480 82050 23520 82250
rect 23590 82050 23910 82250
rect 23980 82050 24020 82250
rect 24090 82050 24410 82250
rect 24480 82050 24520 82250
rect 24590 82050 24910 82250
rect 24980 82050 25020 82250
rect 25090 82050 25410 82250
rect 25480 82050 25520 82250
rect 25590 82050 25910 82250
rect 25980 82050 26020 82250
rect 26090 82050 26410 82250
rect 26480 82050 26520 82250
rect 26590 82050 26910 82250
rect 26980 82050 27020 82250
rect 27090 82050 27410 82250
rect 27480 82050 27520 82250
rect 27590 82050 27910 82250
rect 27980 82050 28020 82250
rect 28090 82050 28410 82250
rect 28480 82050 28520 82250
rect 28590 82050 28910 82250
rect 28980 82050 29020 82250
rect 29090 82050 29410 82250
rect 29480 82050 29520 82250
rect 29590 82050 29910 82250
rect 29980 82050 30020 82250
rect 30090 82050 30410 82250
rect 30480 82050 30520 82250
rect 30590 82050 30910 82250
rect 30980 82050 31020 82250
rect 31090 82050 31410 82250
rect 31480 82050 31520 82250
rect 31590 82050 31910 82250
rect 31980 82050 32020 82250
rect 32090 82050 32410 82250
rect 32480 82050 32520 82250
rect 32590 82050 32910 82250
rect 32980 82050 33020 82250
rect 33090 82050 33410 82250
rect 33480 82050 33520 82250
rect 33590 82050 33910 82250
rect 33980 82050 34020 82250
rect 34090 82050 34410 82250
rect 34480 82050 34520 82250
rect 34590 82050 34910 82250
rect 34980 82050 35020 82250
rect 35090 82050 35410 82250
rect 35480 82050 35520 82250
rect 35590 82050 35910 82250
rect 35980 82050 36020 82250
rect 36090 82050 36410 82250
rect 36480 82050 36520 82250
rect 36590 82050 36910 82250
rect 36980 82050 37020 82250
rect 37090 82050 37410 82250
rect 37480 82050 37520 82250
rect 37590 82050 37910 82250
rect 37980 82050 38020 82250
rect 38090 82050 38410 82250
rect 38480 82050 38520 82250
rect 38590 82050 38910 82250
rect 38980 82050 39020 82250
rect 39090 82050 39410 82250
rect 39480 82050 39520 82250
rect 39590 82050 39910 82250
rect 39980 82050 40020 82250
rect 40090 82050 40410 82250
rect 40480 82050 40520 82250
rect 40590 82050 40910 82250
rect 40980 82050 41020 82250
rect 41090 82050 41410 82250
rect 41480 82050 41520 82250
rect 41590 82050 41910 82250
rect 41980 82050 42020 82250
rect 42090 82050 42410 82250
rect 42480 82050 42520 82250
rect 42590 82050 42910 82250
rect 42980 82050 43020 82250
rect 43090 82050 43410 82250
rect 43480 82050 43520 82250
rect 43590 82050 43910 82250
rect 43980 82050 44020 82250
rect 44090 82050 44410 82250
rect 44480 82050 44520 82250
rect 44590 82050 44910 82250
rect 44980 82050 45020 82250
rect 45090 82050 45410 82250
rect 45480 82050 45520 82250
rect 45590 82050 45910 82250
rect 45980 82050 46020 82250
rect 46090 82050 46410 82250
rect 46480 82050 46520 82250
rect 46590 82050 46910 82250
rect 46980 82050 47020 82250
rect 47090 82050 47410 82250
rect 47480 82050 47520 82250
rect 47590 82050 47910 82250
rect 47980 82050 48020 82250
rect 48090 82050 48410 82250
rect 48480 82050 48520 82250
rect 48590 82050 48910 82250
rect 48980 82050 49020 82250
rect 49090 82050 49410 82250
rect 49480 82050 49520 82250
rect 49590 82050 49910 82250
rect 49980 82050 50020 82250
rect 50090 82050 50410 82250
rect 50480 82050 50520 82250
rect 50590 82050 50910 82250
rect 50980 82050 51020 82250
rect 51090 82050 51410 82250
rect 51480 82050 51520 82250
rect 51590 82050 51910 82250
rect 51980 82050 52020 82250
rect 52090 82050 52410 82250
rect 52480 82050 52520 82250
rect 52590 82050 52910 82250
rect 52980 82050 53020 82250
rect 53090 82050 53410 82250
rect 53480 82050 53520 82250
rect 53590 82050 53910 82250
rect 53980 82050 54020 82250
rect 54090 82050 54410 82250
rect 54480 82050 54520 82250
rect 54590 82050 54910 82250
rect 54980 82050 55020 82250
rect 55090 82050 55410 82250
rect 55480 82050 55520 82250
rect 55590 82050 55910 82250
rect 55980 82050 56020 82250
rect 56090 82050 56410 82250
rect 56480 82050 56520 82250
rect 56590 82050 56910 82250
rect 56980 82050 57020 82250
rect 57090 82050 57410 82250
rect 57480 82050 57520 82250
rect 57590 82050 57910 82250
rect 57980 82050 58020 82250
rect 58090 82050 58410 82250
rect 58480 82050 58520 82250
rect 58590 82050 58910 82250
rect 58980 82050 59020 82250
rect 59090 82050 59410 82250
rect 59480 82050 59520 82250
rect 59590 82050 59910 82250
rect 59980 82050 60020 82250
rect 60090 82050 60410 82250
rect 60480 82050 60520 82250
rect 60590 82050 60910 82250
rect 60980 82050 61020 82250
rect 61090 82050 61410 82250
rect 61480 82050 61520 82250
rect 61590 82050 61910 82250
rect 61980 82050 62020 82250
rect 62090 82050 62410 82250
rect 62480 82050 62520 82250
rect 62590 82050 62910 82250
rect 62980 82050 63020 82250
rect 63090 82050 63410 82250
rect 63480 82050 63520 82250
rect 63590 82050 63910 82250
rect 63980 82050 64020 82250
rect 64090 82050 64410 82250
rect 64480 82050 64520 82250
rect 64590 82050 64910 82250
rect 64980 82050 65020 82250
rect 65090 82050 65410 82250
rect 65480 82050 65520 82250
rect 65590 82050 65910 82250
rect 65980 82050 66020 82250
rect 66090 82050 66410 82250
rect 66480 82050 66520 82250
rect 66590 82050 66910 82250
rect 66980 82050 67020 82250
rect 67090 82050 67410 82250
rect 67480 82050 67520 82250
rect 67590 82050 67910 82250
rect 67980 82050 68020 82250
rect 68090 82050 68410 82250
rect 68480 82050 68520 82250
rect 68590 82050 68910 82250
rect 68980 82050 69020 82250
rect 69090 82050 69410 82250
rect 69480 82050 69520 82250
rect 69590 82050 69910 82250
rect 69980 82050 70020 82250
rect 70090 82050 70410 82250
rect 70480 82050 70520 82250
rect 70590 82050 70910 82250
rect 70980 82050 71020 82250
rect 71090 82050 71410 82250
rect 71480 82050 71520 82250
rect 71590 82050 71910 82250
rect 71980 82050 72020 82250
rect 72090 82050 72410 82250
rect 72480 82050 72520 82250
rect 72590 82050 72910 82250
rect 72980 82050 73020 82250
rect 73090 82050 73410 82250
rect 73480 82050 73520 82250
rect 73590 82050 73910 82250
rect 73980 82050 74020 82250
rect 74090 82050 74410 82250
rect 74480 82050 74520 82250
rect 74590 82050 74910 82250
rect 74980 82050 75020 82250
rect 75090 82050 75410 82250
rect 75480 82050 75520 82250
rect 75590 82050 75910 82250
rect 75980 82050 76020 82250
rect 76090 82050 76410 82250
rect 76480 82050 76520 82250
rect 76590 82050 76910 82250
rect 76980 82050 77020 82250
rect 77090 82050 77410 82250
rect 77480 82050 77520 82250
rect 77590 82050 77910 82250
rect 77980 82050 78020 82250
rect 78090 82050 78410 82250
rect 78480 82050 78520 82250
rect 78590 82050 78910 82250
rect 78980 82050 79020 82250
rect 79090 82050 79410 82250
rect 79480 82050 79520 82250
rect 79590 82050 79910 82250
rect 79980 82050 80020 82250
rect 80090 82050 80410 82250
rect 80480 82050 80520 82250
rect 80590 82050 80910 82250
rect 80980 82050 81020 82250
rect 81090 82050 81410 82250
rect 81480 82050 81520 82250
rect 81590 82050 81910 82250
rect 81980 82050 82020 82250
rect 82090 82050 82410 82250
rect 82480 82050 82520 82250
rect 82590 82050 82910 82250
rect 82980 82050 83020 82250
rect 83090 82050 83410 82250
rect 83480 82050 83520 82250
rect 83590 82050 83910 82250
rect 83980 82050 84020 82250
rect 84090 82050 84410 82250
rect 84480 82050 84520 82250
rect 84590 82050 84910 82250
rect 84980 82050 85020 82250
rect 85090 82050 85410 82250
rect 85480 82050 85520 82250
rect 85590 82050 85910 82250
rect 85980 82050 86020 82250
rect 86090 82050 86410 82250
rect 86480 82050 86520 82250
rect 86590 82050 86910 82250
rect 86980 82050 87020 82250
rect 87090 82050 87410 82250
rect 87480 82050 87520 82250
rect 87590 82050 87910 82250
rect 87980 82050 88020 82250
rect 88090 82050 88410 82250
rect 88480 82050 88520 82250
rect 88590 82050 88910 82250
rect 88980 82050 89020 82250
rect 89090 82050 89410 82250
rect 89480 82050 89520 82250
rect 89590 82050 89910 82250
rect 89980 82050 90020 82250
rect 90090 82050 90410 82250
rect 90480 82050 90520 82250
rect 90590 82050 90910 82250
rect 90980 82050 91020 82250
rect 91090 82050 91410 82250
rect 91480 82050 91520 82250
rect 91590 82050 91910 82250
rect 91980 82050 92020 82250
rect 92090 82050 92410 82250
rect 92480 82050 92520 82250
rect 92590 82050 92910 82250
rect 92980 82050 93020 82250
rect 93090 82050 93410 82250
rect 93480 82050 93520 82250
rect 93590 82050 93910 82250
rect 93980 82050 94020 82250
rect 94090 82050 94410 82250
rect 94480 82050 94520 82250
rect 94590 82050 94910 82250
rect 94980 82050 95020 82250
rect 95090 82050 95410 82250
rect 95480 82050 95520 82250
rect 95590 82050 95910 82250
rect 95980 82050 96020 82250
rect 96090 82050 96410 82250
rect 96480 82050 96520 82250
rect 96590 82050 96910 82250
rect 96980 82050 97020 82250
rect 97090 82050 97410 82250
rect 97480 82050 97520 82250
rect 97590 82050 97910 82250
rect 97980 82050 98020 82250
rect 98090 82050 98410 82250
rect 98480 82050 98520 82250
rect 98590 82050 98910 82250
rect 98980 82050 99020 82250
rect 99090 82050 99410 82250
rect 99480 82050 99520 82250
rect 99590 82050 99910 82250
rect 99980 82050 100020 82250
rect 100090 82050 100410 82250
rect 100480 82050 100500 82250
rect -83500 82040 100500 82050
rect -83360 81990 -83140 82040
rect -83360 81920 -83350 81990
rect -83150 81920 -83140 81990
rect -83360 81880 -83140 81920
rect -83360 81810 -83350 81880
rect -83150 81810 -83140 81880
rect -83360 81760 -83140 81810
rect -82860 81990 -82640 82040
rect -82860 81920 -82850 81990
rect -82650 81920 -82640 81990
rect -82860 81880 -82640 81920
rect -82860 81810 -82850 81880
rect -82650 81810 -82640 81880
rect -82860 81760 -82640 81810
rect -82360 81990 -82140 82040
rect -82360 81920 -82350 81990
rect -82150 81920 -82140 81990
rect -82360 81880 -82140 81920
rect -82360 81810 -82350 81880
rect -82150 81810 -82140 81880
rect -82360 81760 -82140 81810
rect -81860 81990 -81640 82040
rect -81860 81920 -81850 81990
rect -81650 81920 -81640 81990
rect -81860 81880 -81640 81920
rect -81860 81810 -81850 81880
rect -81650 81810 -81640 81880
rect -81860 81760 -81640 81810
rect -81360 81990 -81140 82040
rect -81360 81920 -81350 81990
rect -81150 81920 -81140 81990
rect -81360 81880 -81140 81920
rect -81360 81810 -81350 81880
rect -81150 81810 -81140 81880
rect -81360 81760 -81140 81810
rect -80860 81990 -80640 82040
rect -80860 81920 -80850 81990
rect -80650 81920 -80640 81990
rect -80860 81880 -80640 81920
rect -80860 81810 -80850 81880
rect -80650 81810 -80640 81880
rect -80860 81760 -80640 81810
rect -80360 81990 -80140 82040
rect -80360 81920 -80350 81990
rect -80150 81920 -80140 81990
rect -80360 81880 -80140 81920
rect -80360 81810 -80350 81880
rect -80150 81810 -80140 81880
rect -80360 81760 -80140 81810
rect -79860 81990 -79640 82040
rect -79860 81920 -79850 81990
rect -79650 81920 -79640 81990
rect -79860 81880 -79640 81920
rect -79860 81810 -79850 81880
rect -79650 81810 -79640 81880
rect -79860 81760 -79640 81810
rect -79360 81990 -79140 82040
rect -79360 81920 -79350 81990
rect -79150 81920 -79140 81990
rect -79360 81880 -79140 81920
rect -79360 81810 -79350 81880
rect -79150 81810 -79140 81880
rect -79360 81760 -79140 81810
rect -78860 81990 -78640 82040
rect -78860 81920 -78850 81990
rect -78650 81920 -78640 81990
rect -78860 81880 -78640 81920
rect -78860 81810 -78850 81880
rect -78650 81810 -78640 81880
rect -78860 81760 -78640 81810
rect -78360 81990 -78140 82040
rect -78360 81920 -78350 81990
rect -78150 81920 -78140 81990
rect -78360 81880 -78140 81920
rect -78360 81810 -78350 81880
rect -78150 81810 -78140 81880
rect -78360 81760 -78140 81810
rect -77860 81990 -77640 82040
rect -77860 81920 -77850 81990
rect -77650 81920 -77640 81990
rect -77860 81880 -77640 81920
rect -77860 81810 -77850 81880
rect -77650 81810 -77640 81880
rect -77860 81760 -77640 81810
rect -77360 81990 -77140 82040
rect -77360 81920 -77350 81990
rect -77150 81920 -77140 81990
rect -77360 81880 -77140 81920
rect -77360 81810 -77350 81880
rect -77150 81810 -77140 81880
rect -77360 81760 -77140 81810
rect -76860 81990 -76640 82040
rect -76860 81920 -76850 81990
rect -76650 81920 -76640 81990
rect -76860 81880 -76640 81920
rect -76860 81810 -76850 81880
rect -76650 81810 -76640 81880
rect -76860 81760 -76640 81810
rect -76360 81990 -76140 82040
rect -76360 81920 -76350 81990
rect -76150 81920 -76140 81990
rect -76360 81880 -76140 81920
rect -76360 81810 -76350 81880
rect -76150 81810 -76140 81880
rect -76360 81760 -76140 81810
rect -75860 81990 -75640 82040
rect -75860 81920 -75850 81990
rect -75650 81920 -75640 81990
rect -75860 81880 -75640 81920
rect -75860 81810 -75850 81880
rect -75650 81810 -75640 81880
rect -75860 81760 -75640 81810
rect -75360 81990 -75140 82040
rect -75360 81920 -75350 81990
rect -75150 81920 -75140 81990
rect -75360 81880 -75140 81920
rect -75360 81810 -75350 81880
rect -75150 81810 -75140 81880
rect -75360 81760 -75140 81810
rect -74860 81990 -74640 82040
rect -74860 81920 -74850 81990
rect -74650 81920 -74640 81990
rect -74860 81880 -74640 81920
rect -74860 81810 -74850 81880
rect -74650 81810 -74640 81880
rect -74860 81760 -74640 81810
rect -74360 81990 -74140 82040
rect -74360 81920 -74350 81990
rect -74150 81920 -74140 81990
rect -74360 81880 -74140 81920
rect -74360 81810 -74350 81880
rect -74150 81810 -74140 81880
rect -74360 81760 -74140 81810
rect -73860 81990 -73640 82040
rect -73860 81920 -73850 81990
rect -73650 81920 -73640 81990
rect -73860 81880 -73640 81920
rect -73860 81810 -73850 81880
rect -73650 81810 -73640 81880
rect -73860 81760 -73640 81810
rect -73360 81990 -73140 82040
rect -73360 81920 -73350 81990
rect -73150 81920 -73140 81990
rect -73360 81880 -73140 81920
rect -73360 81810 -73350 81880
rect -73150 81810 -73140 81880
rect -73360 81760 -73140 81810
rect -72860 81990 -72640 82040
rect -72860 81920 -72850 81990
rect -72650 81920 -72640 81990
rect -72860 81880 -72640 81920
rect -72860 81810 -72850 81880
rect -72650 81810 -72640 81880
rect -72860 81760 -72640 81810
rect -72360 81990 -72140 82040
rect -72360 81920 -72350 81990
rect -72150 81920 -72140 81990
rect -72360 81880 -72140 81920
rect -72360 81810 -72350 81880
rect -72150 81810 -72140 81880
rect -72360 81760 -72140 81810
rect -71860 81990 -71640 82040
rect -71860 81920 -71850 81990
rect -71650 81920 -71640 81990
rect -71860 81880 -71640 81920
rect -71860 81810 -71850 81880
rect -71650 81810 -71640 81880
rect -71860 81760 -71640 81810
rect -71360 81990 -71140 82040
rect -71360 81920 -71350 81990
rect -71150 81920 -71140 81990
rect -71360 81880 -71140 81920
rect -71360 81810 -71350 81880
rect -71150 81810 -71140 81880
rect -71360 81760 -71140 81810
rect -70860 81990 -70640 82040
rect -70860 81920 -70850 81990
rect -70650 81920 -70640 81990
rect -70860 81880 -70640 81920
rect -70860 81810 -70850 81880
rect -70650 81810 -70640 81880
rect -70860 81760 -70640 81810
rect -70360 81990 -70140 82040
rect -70360 81920 -70350 81990
rect -70150 81920 -70140 81990
rect -70360 81880 -70140 81920
rect -70360 81810 -70350 81880
rect -70150 81810 -70140 81880
rect -70360 81760 -70140 81810
rect -69860 81990 -69640 82040
rect -69860 81920 -69850 81990
rect -69650 81920 -69640 81990
rect -69860 81880 -69640 81920
rect -69860 81810 -69850 81880
rect -69650 81810 -69640 81880
rect -69860 81760 -69640 81810
rect -69360 81990 -69140 82040
rect -69360 81920 -69350 81990
rect -69150 81920 -69140 81990
rect -69360 81880 -69140 81920
rect -69360 81810 -69350 81880
rect -69150 81810 -69140 81880
rect -69360 81760 -69140 81810
rect -68860 81990 -68640 82040
rect -68860 81920 -68850 81990
rect -68650 81920 -68640 81990
rect -68860 81880 -68640 81920
rect -68860 81810 -68850 81880
rect -68650 81810 -68640 81880
rect -68860 81760 -68640 81810
rect -68360 81990 -68140 82040
rect -68360 81920 -68350 81990
rect -68150 81920 -68140 81990
rect -68360 81880 -68140 81920
rect -68360 81810 -68350 81880
rect -68150 81810 -68140 81880
rect -68360 81760 -68140 81810
rect -67860 81990 -67640 82040
rect -67860 81920 -67850 81990
rect -67650 81920 -67640 81990
rect -67860 81880 -67640 81920
rect -67860 81810 -67850 81880
rect -67650 81810 -67640 81880
rect -67860 81760 -67640 81810
rect -67360 81990 -67140 82040
rect -67360 81920 -67350 81990
rect -67150 81920 -67140 81990
rect -67360 81880 -67140 81920
rect -67360 81810 -67350 81880
rect -67150 81810 -67140 81880
rect -67360 81760 -67140 81810
rect -66860 81990 -66640 82040
rect -66860 81920 -66850 81990
rect -66650 81920 -66640 81990
rect -66860 81880 -66640 81920
rect -66860 81810 -66850 81880
rect -66650 81810 -66640 81880
rect -66860 81760 -66640 81810
rect -66360 81990 -66140 82040
rect -66360 81920 -66350 81990
rect -66150 81920 -66140 81990
rect -66360 81880 -66140 81920
rect -66360 81810 -66350 81880
rect -66150 81810 -66140 81880
rect -66360 81760 -66140 81810
rect -65860 81990 -65640 82040
rect -65860 81920 -65850 81990
rect -65650 81920 -65640 81990
rect -65860 81880 -65640 81920
rect -65860 81810 -65850 81880
rect -65650 81810 -65640 81880
rect -65860 81760 -65640 81810
rect -65360 81990 -65140 82040
rect -65360 81920 -65350 81990
rect -65150 81920 -65140 81990
rect -65360 81880 -65140 81920
rect -65360 81810 -65350 81880
rect -65150 81810 -65140 81880
rect -65360 81760 -65140 81810
rect -64860 81990 -64640 82040
rect -64860 81920 -64850 81990
rect -64650 81920 -64640 81990
rect -64860 81880 -64640 81920
rect -64860 81810 -64850 81880
rect -64650 81810 -64640 81880
rect -64860 81760 -64640 81810
rect -64360 81990 -64140 82040
rect -64360 81920 -64350 81990
rect -64150 81920 -64140 81990
rect -64360 81880 -64140 81920
rect -64360 81810 -64350 81880
rect -64150 81810 -64140 81880
rect -64360 81760 -64140 81810
rect -63860 81990 -63640 82040
rect -63860 81920 -63850 81990
rect -63650 81920 -63640 81990
rect -63860 81880 -63640 81920
rect -63860 81810 -63850 81880
rect -63650 81810 -63640 81880
rect -63860 81760 -63640 81810
rect -63360 81990 -63140 82040
rect -63360 81920 -63350 81990
rect -63150 81920 -63140 81990
rect -63360 81880 -63140 81920
rect -63360 81810 -63350 81880
rect -63150 81810 -63140 81880
rect -63360 81760 -63140 81810
rect -62860 81990 -62640 82040
rect -62860 81920 -62850 81990
rect -62650 81920 -62640 81990
rect -62860 81880 -62640 81920
rect -62860 81810 -62850 81880
rect -62650 81810 -62640 81880
rect -62860 81760 -62640 81810
rect -62360 81990 -62140 82040
rect -62360 81920 -62350 81990
rect -62150 81920 -62140 81990
rect -62360 81880 -62140 81920
rect -62360 81810 -62350 81880
rect -62150 81810 -62140 81880
rect -62360 81760 -62140 81810
rect -61860 81990 -61640 82040
rect -61860 81920 -61850 81990
rect -61650 81920 -61640 81990
rect -61860 81880 -61640 81920
rect -61860 81810 -61850 81880
rect -61650 81810 -61640 81880
rect -61860 81760 -61640 81810
rect -61360 81990 -61140 82040
rect -61360 81920 -61350 81990
rect -61150 81920 -61140 81990
rect -61360 81880 -61140 81920
rect -61360 81810 -61350 81880
rect -61150 81810 -61140 81880
rect -61360 81760 -61140 81810
rect -60860 81990 -60640 82040
rect -60860 81920 -60850 81990
rect -60650 81920 -60640 81990
rect -60860 81880 -60640 81920
rect -60860 81810 -60850 81880
rect -60650 81810 -60640 81880
rect -60860 81760 -60640 81810
rect -60360 81990 -60140 82040
rect -60360 81920 -60350 81990
rect -60150 81920 -60140 81990
rect -60360 81880 -60140 81920
rect -60360 81810 -60350 81880
rect -60150 81810 -60140 81880
rect -60360 81760 -60140 81810
rect -59860 81990 -59640 82040
rect -59860 81920 -59850 81990
rect -59650 81920 -59640 81990
rect -59860 81880 -59640 81920
rect -59860 81810 -59850 81880
rect -59650 81810 -59640 81880
rect -59860 81760 -59640 81810
rect -59360 81990 -59140 82040
rect -59360 81920 -59350 81990
rect -59150 81920 -59140 81990
rect -59360 81880 -59140 81920
rect -59360 81810 -59350 81880
rect -59150 81810 -59140 81880
rect -59360 81760 -59140 81810
rect -58860 81990 -58640 82040
rect -58860 81920 -58850 81990
rect -58650 81920 -58640 81990
rect -58860 81880 -58640 81920
rect -58860 81810 -58850 81880
rect -58650 81810 -58640 81880
rect -58860 81760 -58640 81810
rect -58360 81990 -58140 82040
rect -58360 81920 -58350 81990
rect -58150 81920 -58140 81990
rect -58360 81880 -58140 81920
rect -58360 81810 -58350 81880
rect -58150 81810 -58140 81880
rect -58360 81760 -58140 81810
rect -57860 81990 -57640 82040
rect -57860 81920 -57850 81990
rect -57650 81920 -57640 81990
rect -57860 81880 -57640 81920
rect -57860 81810 -57850 81880
rect -57650 81810 -57640 81880
rect -57860 81760 -57640 81810
rect -57360 81990 -57140 82040
rect -57360 81920 -57350 81990
rect -57150 81920 -57140 81990
rect -57360 81880 -57140 81920
rect -57360 81810 -57350 81880
rect -57150 81810 -57140 81880
rect -57360 81760 -57140 81810
rect -56860 81990 -56640 82040
rect -56860 81920 -56850 81990
rect -56650 81920 -56640 81990
rect -56860 81880 -56640 81920
rect -56860 81810 -56850 81880
rect -56650 81810 -56640 81880
rect -56860 81760 -56640 81810
rect -56360 81990 -56140 82040
rect -56360 81920 -56350 81990
rect -56150 81920 -56140 81990
rect -56360 81880 -56140 81920
rect -56360 81810 -56350 81880
rect -56150 81810 -56140 81880
rect -56360 81760 -56140 81810
rect -55860 81990 -55640 82040
rect -55860 81920 -55850 81990
rect -55650 81920 -55640 81990
rect -55860 81880 -55640 81920
rect -55860 81810 -55850 81880
rect -55650 81810 -55640 81880
rect -55860 81760 -55640 81810
rect -55360 81990 -55140 82040
rect -55360 81920 -55350 81990
rect -55150 81920 -55140 81990
rect -55360 81880 -55140 81920
rect -55360 81810 -55350 81880
rect -55150 81810 -55140 81880
rect -55360 81760 -55140 81810
rect -54860 81990 -54640 82040
rect -54860 81920 -54850 81990
rect -54650 81920 -54640 81990
rect -54860 81880 -54640 81920
rect -54860 81810 -54850 81880
rect -54650 81810 -54640 81880
rect -54860 81760 -54640 81810
rect -54360 81990 -54140 82040
rect -54360 81920 -54350 81990
rect -54150 81920 -54140 81990
rect -54360 81880 -54140 81920
rect -54360 81810 -54350 81880
rect -54150 81810 -54140 81880
rect -54360 81760 -54140 81810
rect -53860 81990 -53640 82040
rect -53860 81920 -53850 81990
rect -53650 81920 -53640 81990
rect -53860 81880 -53640 81920
rect -53860 81810 -53850 81880
rect -53650 81810 -53640 81880
rect -53860 81760 -53640 81810
rect -53360 81990 -53140 82040
rect -53360 81920 -53350 81990
rect -53150 81920 -53140 81990
rect -53360 81880 -53140 81920
rect -53360 81810 -53350 81880
rect -53150 81810 -53140 81880
rect -53360 81760 -53140 81810
rect -52860 81990 -52640 82040
rect -52860 81920 -52850 81990
rect -52650 81920 -52640 81990
rect -52860 81880 -52640 81920
rect -52860 81810 -52850 81880
rect -52650 81810 -52640 81880
rect -52860 81760 -52640 81810
rect -52360 81990 -52140 82040
rect -52360 81920 -52350 81990
rect -52150 81920 -52140 81990
rect -52360 81880 -52140 81920
rect -52360 81810 -52350 81880
rect -52150 81810 -52140 81880
rect -52360 81760 -52140 81810
rect -51860 81990 -51640 82040
rect -51860 81920 -51850 81990
rect -51650 81920 -51640 81990
rect -51860 81880 -51640 81920
rect -51860 81810 -51850 81880
rect -51650 81810 -51640 81880
rect -51860 81760 -51640 81810
rect -51360 81990 -51140 82040
rect -51360 81920 -51350 81990
rect -51150 81920 -51140 81990
rect -51360 81880 -51140 81920
rect -51360 81810 -51350 81880
rect -51150 81810 -51140 81880
rect -51360 81760 -51140 81810
rect -50860 81990 -50640 82040
rect -50860 81920 -50850 81990
rect -50650 81920 -50640 81990
rect -50860 81880 -50640 81920
rect -50860 81810 -50850 81880
rect -50650 81810 -50640 81880
rect -50860 81760 -50640 81810
rect -50360 81990 -50140 82040
rect -50360 81920 -50350 81990
rect -50150 81920 -50140 81990
rect -50360 81880 -50140 81920
rect -50360 81810 -50350 81880
rect -50150 81810 -50140 81880
rect -50360 81760 -50140 81810
rect -49860 81990 -49640 82040
rect -49860 81920 -49850 81990
rect -49650 81920 -49640 81990
rect -49860 81880 -49640 81920
rect -49860 81810 -49850 81880
rect -49650 81810 -49640 81880
rect -49860 81760 -49640 81810
rect -49360 81990 -49140 82040
rect -49360 81920 -49350 81990
rect -49150 81920 -49140 81990
rect -49360 81880 -49140 81920
rect -49360 81810 -49350 81880
rect -49150 81810 -49140 81880
rect -49360 81760 -49140 81810
rect -48860 81990 -48640 82040
rect -48860 81920 -48850 81990
rect -48650 81920 -48640 81990
rect -48860 81880 -48640 81920
rect -48860 81810 -48850 81880
rect -48650 81810 -48640 81880
rect -48860 81760 -48640 81810
rect -48360 81990 -48140 82040
rect -48360 81920 -48350 81990
rect -48150 81920 -48140 81990
rect -48360 81880 -48140 81920
rect -48360 81810 -48350 81880
rect -48150 81810 -48140 81880
rect -48360 81760 -48140 81810
rect -47860 81990 -47640 82040
rect -47860 81920 -47850 81990
rect -47650 81920 -47640 81990
rect -47860 81880 -47640 81920
rect -47860 81810 -47850 81880
rect -47650 81810 -47640 81880
rect -47860 81760 -47640 81810
rect -47360 81990 -47140 82040
rect -47360 81920 -47350 81990
rect -47150 81920 -47140 81990
rect -47360 81880 -47140 81920
rect -47360 81810 -47350 81880
rect -47150 81810 -47140 81880
rect -47360 81760 -47140 81810
rect -46860 81990 -46640 82040
rect -46860 81920 -46850 81990
rect -46650 81920 -46640 81990
rect -46860 81880 -46640 81920
rect -46860 81810 -46850 81880
rect -46650 81810 -46640 81880
rect -46860 81760 -46640 81810
rect -46360 81990 -46140 82040
rect -46360 81920 -46350 81990
rect -46150 81920 -46140 81990
rect -46360 81880 -46140 81920
rect -46360 81810 -46350 81880
rect -46150 81810 -46140 81880
rect -46360 81760 -46140 81810
rect -45860 81990 -45640 82040
rect -45860 81920 -45850 81990
rect -45650 81920 -45640 81990
rect -45860 81880 -45640 81920
rect -45860 81810 -45850 81880
rect -45650 81810 -45640 81880
rect -45860 81760 -45640 81810
rect -45360 81990 -45140 82040
rect -45360 81920 -45350 81990
rect -45150 81920 -45140 81990
rect -45360 81880 -45140 81920
rect -45360 81810 -45350 81880
rect -45150 81810 -45140 81880
rect -45360 81760 -45140 81810
rect -44860 81990 -44640 82040
rect -44860 81920 -44850 81990
rect -44650 81920 -44640 81990
rect -44860 81880 -44640 81920
rect -44860 81810 -44850 81880
rect -44650 81810 -44640 81880
rect -44860 81760 -44640 81810
rect -44360 81990 -44140 82040
rect -44360 81920 -44350 81990
rect -44150 81920 -44140 81990
rect -44360 81880 -44140 81920
rect -44360 81810 -44350 81880
rect -44150 81810 -44140 81880
rect -44360 81760 -44140 81810
rect -43860 81990 -43640 82040
rect -43860 81920 -43850 81990
rect -43650 81920 -43640 81990
rect -43860 81880 -43640 81920
rect -43860 81810 -43850 81880
rect -43650 81810 -43640 81880
rect -43860 81760 -43640 81810
rect -43360 81990 -43140 82040
rect -43360 81920 -43350 81990
rect -43150 81920 -43140 81990
rect -43360 81880 -43140 81920
rect -43360 81810 -43350 81880
rect -43150 81810 -43140 81880
rect -43360 81760 -43140 81810
rect -42860 81990 -42640 82040
rect -42860 81920 -42850 81990
rect -42650 81920 -42640 81990
rect -42860 81880 -42640 81920
rect -42860 81810 -42850 81880
rect -42650 81810 -42640 81880
rect -42860 81760 -42640 81810
rect -42360 81990 -42140 82040
rect -42360 81920 -42350 81990
rect -42150 81920 -42140 81990
rect -42360 81880 -42140 81920
rect -42360 81810 -42350 81880
rect -42150 81810 -42140 81880
rect -42360 81760 -42140 81810
rect -41860 81990 -41640 82040
rect -41860 81920 -41850 81990
rect -41650 81920 -41640 81990
rect -41860 81880 -41640 81920
rect -41860 81810 -41850 81880
rect -41650 81810 -41640 81880
rect -41860 81760 -41640 81810
rect -41360 81990 -41140 82040
rect -41360 81920 -41350 81990
rect -41150 81920 -41140 81990
rect -41360 81880 -41140 81920
rect -41360 81810 -41350 81880
rect -41150 81810 -41140 81880
rect -41360 81760 -41140 81810
rect -40860 81990 -40640 82040
rect -40860 81920 -40850 81990
rect -40650 81920 -40640 81990
rect -40860 81880 -40640 81920
rect -40860 81810 -40850 81880
rect -40650 81810 -40640 81880
rect -40860 81760 -40640 81810
rect -40360 81990 -40140 82040
rect -40360 81920 -40350 81990
rect -40150 81920 -40140 81990
rect -40360 81880 -40140 81920
rect -40360 81810 -40350 81880
rect -40150 81810 -40140 81880
rect -40360 81760 -40140 81810
rect -39860 81990 -39640 82040
rect -39860 81920 -39850 81990
rect -39650 81920 -39640 81990
rect -39860 81880 -39640 81920
rect -39860 81810 -39850 81880
rect -39650 81810 -39640 81880
rect -39860 81760 -39640 81810
rect -39360 81990 -39140 82040
rect -39360 81920 -39350 81990
rect -39150 81920 -39140 81990
rect -39360 81880 -39140 81920
rect -39360 81810 -39350 81880
rect -39150 81810 -39140 81880
rect -39360 81760 -39140 81810
rect -38860 81990 -38640 82040
rect -38860 81920 -38850 81990
rect -38650 81920 -38640 81990
rect -38860 81880 -38640 81920
rect -38860 81810 -38850 81880
rect -38650 81810 -38640 81880
rect -38860 81760 -38640 81810
rect -38360 81990 -38140 82040
rect -38360 81920 -38350 81990
rect -38150 81920 -38140 81990
rect -38360 81880 -38140 81920
rect -38360 81810 -38350 81880
rect -38150 81810 -38140 81880
rect -38360 81760 -38140 81810
rect -37860 81990 -37640 82040
rect -37860 81920 -37850 81990
rect -37650 81920 -37640 81990
rect -37860 81880 -37640 81920
rect -37860 81810 -37850 81880
rect -37650 81810 -37640 81880
rect -37860 81760 -37640 81810
rect -37360 81990 -37140 82040
rect -37360 81920 -37350 81990
rect -37150 81920 -37140 81990
rect -37360 81880 -37140 81920
rect -37360 81810 -37350 81880
rect -37150 81810 -37140 81880
rect -37360 81760 -37140 81810
rect -36860 81990 -36640 82040
rect -36860 81920 -36850 81990
rect -36650 81920 -36640 81990
rect -36860 81880 -36640 81920
rect -36860 81810 -36850 81880
rect -36650 81810 -36640 81880
rect -36860 81760 -36640 81810
rect -36360 81990 -36140 82040
rect -36360 81920 -36350 81990
rect -36150 81920 -36140 81990
rect -36360 81880 -36140 81920
rect -36360 81810 -36350 81880
rect -36150 81810 -36140 81880
rect -36360 81760 -36140 81810
rect -35860 81990 -35640 82040
rect -35860 81920 -35850 81990
rect -35650 81920 -35640 81990
rect -35860 81880 -35640 81920
rect -35860 81810 -35850 81880
rect -35650 81810 -35640 81880
rect -35860 81760 -35640 81810
rect -35360 81990 -35140 82040
rect -35360 81920 -35350 81990
rect -35150 81920 -35140 81990
rect -35360 81880 -35140 81920
rect -35360 81810 -35350 81880
rect -35150 81810 -35140 81880
rect -35360 81760 -35140 81810
rect -34860 81990 -34640 82040
rect -34860 81920 -34850 81990
rect -34650 81920 -34640 81990
rect -34860 81880 -34640 81920
rect -34860 81810 -34850 81880
rect -34650 81810 -34640 81880
rect -34860 81760 -34640 81810
rect -34360 81990 -34140 82040
rect -34360 81920 -34350 81990
rect -34150 81920 -34140 81990
rect -34360 81880 -34140 81920
rect -34360 81810 -34350 81880
rect -34150 81810 -34140 81880
rect -34360 81760 -34140 81810
rect -33860 81990 -33640 82040
rect -33860 81920 -33850 81990
rect -33650 81920 -33640 81990
rect -33860 81880 -33640 81920
rect -33860 81810 -33850 81880
rect -33650 81810 -33640 81880
rect -33860 81760 -33640 81810
rect -33360 81990 -33140 82040
rect -33360 81920 -33350 81990
rect -33150 81920 -33140 81990
rect -33360 81880 -33140 81920
rect -33360 81810 -33350 81880
rect -33150 81810 -33140 81880
rect -33360 81760 -33140 81810
rect -32860 81990 -32640 82040
rect -32860 81920 -32850 81990
rect -32650 81920 -32640 81990
rect -32860 81880 -32640 81920
rect -32860 81810 -32850 81880
rect -32650 81810 -32640 81880
rect -32860 81760 -32640 81810
rect -32360 81990 -32140 82040
rect -32360 81920 -32350 81990
rect -32150 81920 -32140 81990
rect -32360 81880 -32140 81920
rect -32360 81810 -32350 81880
rect -32150 81810 -32140 81880
rect -32360 81760 -32140 81810
rect -31860 81990 -31640 82040
rect -31860 81920 -31850 81990
rect -31650 81920 -31640 81990
rect -31860 81880 -31640 81920
rect -31860 81810 -31850 81880
rect -31650 81810 -31640 81880
rect -31860 81760 -31640 81810
rect -31360 81990 -31140 82040
rect -31360 81920 -31350 81990
rect -31150 81920 -31140 81990
rect -31360 81880 -31140 81920
rect -31360 81810 -31350 81880
rect -31150 81810 -31140 81880
rect -31360 81760 -31140 81810
rect -30860 81990 -30640 82040
rect -30860 81920 -30850 81990
rect -30650 81920 -30640 81990
rect -30860 81880 -30640 81920
rect -30860 81810 -30850 81880
rect -30650 81810 -30640 81880
rect -30860 81760 -30640 81810
rect -30360 81990 -30140 82040
rect -30360 81920 -30350 81990
rect -30150 81920 -30140 81990
rect -30360 81880 -30140 81920
rect -30360 81810 -30350 81880
rect -30150 81810 -30140 81880
rect -30360 81760 -30140 81810
rect -29860 81990 -29640 82040
rect -29860 81920 -29850 81990
rect -29650 81920 -29640 81990
rect -29860 81880 -29640 81920
rect -29860 81810 -29850 81880
rect -29650 81810 -29640 81880
rect -29860 81760 -29640 81810
rect -29360 81990 -29140 82040
rect -29360 81920 -29350 81990
rect -29150 81920 -29140 81990
rect -29360 81880 -29140 81920
rect -29360 81810 -29350 81880
rect -29150 81810 -29140 81880
rect -29360 81760 -29140 81810
rect -28860 81990 -28640 82040
rect -28860 81920 -28850 81990
rect -28650 81920 -28640 81990
rect -28860 81880 -28640 81920
rect -28860 81810 -28850 81880
rect -28650 81810 -28640 81880
rect -28860 81760 -28640 81810
rect -28360 81990 -28140 82040
rect -28360 81920 -28350 81990
rect -28150 81920 -28140 81990
rect -28360 81880 -28140 81920
rect -28360 81810 -28350 81880
rect -28150 81810 -28140 81880
rect -28360 81760 -28140 81810
rect -27860 81990 -27640 82040
rect -27860 81920 -27850 81990
rect -27650 81920 -27640 81990
rect -27860 81880 -27640 81920
rect -27860 81810 -27850 81880
rect -27650 81810 -27640 81880
rect -27860 81760 -27640 81810
rect -27360 81990 -27140 82040
rect -27360 81920 -27350 81990
rect -27150 81920 -27140 81990
rect -27360 81880 -27140 81920
rect -27360 81810 -27350 81880
rect -27150 81810 -27140 81880
rect -27360 81760 -27140 81810
rect -26860 81990 -26640 82040
rect -26860 81920 -26850 81990
rect -26650 81920 -26640 81990
rect -26860 81880 -26640 81920
rect -26860 81810 -26850 81880
rect -26650 81810 -26640 81880
rect -26860 81760 -26640 81810
rect -26360 81990 -26140 82040
rect -26360 81920 -26350 81990
rect -26150 81920 -26140 81990
rect -26360 81880 -26140 81920
rect -26360 81810 -26350 81880
rect -26150 81810 -26140 81880
rect -26360 81760 -26140 81810
rect -25860 81990 -25640 82040
rect -25860 81920 -25850 81990
rect -25650 81920 -25640 81990
rect -25860 81880 -25640 81920
rect -25860 81810 -25850 81880
rect -25650 81810 -25640 81880
rect -25860 81760 -25640 81810
rect -25360 81990 -25140 82040
rect -25360 81920 -25350 81990
rect -25150 81920 -25140 81990
rect -25360 81880 -25140 81920
rect -25360 81810 -25350 81880
rect -25150 81810 -25140 81880
rect -25360 81760 -25140 81810
rect -24860 81990 -24640 82040
rect -24860 81920 -24850 81990
rect -24650 81920 -24640 81990
rect -24860 81880 -24640 81920
rect -24860 81810 -24850 81880
rect -24650 81810 -24640 81880
rect -24860 81760 -24640 81810
rect -24360 81990 -24140 82040
rect -24360 81920 -24350 81990
rect -24150 81920 -24140 81990
rect -24360 81880 -24140 81920
rect -24360 81810 -24350 81880
rect -24150 81810 -24140 81880
rect -24360 81760 -24140 81810
rect -23860 81990 -23640 82040
rect -23860 81920 -23850 81990
rect -23650 81920 -23640 81990
rect -23860 81880 -23640 81920
rect -23860 81810 -23850 81880
rect -23650 81810 -23640 81880
rect -23860 81760 -23640 81810
rect -23360 81990 -23140 82040
rect -23360 81920 -23350 81990
rect -23150 81920 -23140 81990
rect -23360 81880 -23140 81920
rect -23360 81810 -23350 81880
rect -23150 81810 -23140 81880
rect -23360 81760 -23140 81810
rect -22860 81990 -22640 82040
rect -22860 81920 -22850 81990
rect -22650 81920 -22640 81990
rect -22860 81880 -22640 81920
rect -22860 81810 -22850 81880
rect -22650 81810 -22640 81880
rect -22860 81760 -22640 81810
rect -22360 81990 -22140 82040
rect -22360 81920 -22350 81990
rect -22150 81920 -22140 81990
rect -22360 81880 -22140 81920
rect -22360 81810 -22350 81880
rect -22150 81810 -22140 81880
rect -22360 81760 -22140 81810
rect -21860 81990 -21640 82040
rect -21860 81920 -21850 81990
rect -21650 81920 -21640 81990
rect -21860 81880 -21640 81920
rect -21860 81810 -21850 81880
rect -21650 81810 -21640 81880
rect -21860 81760 -21640 81810
rect -21360 81990 -21140 82040
rect -21360 81920 -21350 81990
rect -21150 81920 -21140 81990
rect -21360 81880 -21140 81920
rect -21360 81810 -21350 81880
rect -21150 81810 -21140 81880
rect -21360 81760 -21140 81810
rect -20860 81990 -20640 82040
rect -20860 81920 -20850 81990
rect -20650 81920 -20640 81990
rect -20860 81880 -20640 81920
rect -20860 81810 -20850 81880
rect -20650 81810 -20640 81880
rect -20860 81760 -20640 81810
rect -20360 81990 -20140 82040
rect -20360 81920 -20350 81990
rect -20150 81920 -20140 81990
rect -20360 81880 -20140 81920
rect -20360 81810 -20350 81880
rect -20150 81810 -20140 81880
rect -20360 81760 -20140 81810
rect -19860 81990 -19640 82040
rect -19860 81920 -19850 81990
rect -19650 81920 -19640 81990
rect -19860 81880 -19640 81920
rect -19860 81810 -19850 81880
rect -19650 81810 -19640 81880
rect -19860 81760 -19640 81810
rect -19360 81990 -19140 82040
rect -19360 81920 -19350 81990
rect -19150 81920 -19140 81990
rect -19360 81880 -19140 81920
rect -19360 81810 -19350 81880
rect -19150 81810 -19140 81880
rect -19360 81760 -19140 81810
rect -18860 81990 -18640 82040
rect -18860 81920 -18850 81990
rect -18650 81920 -18640 81990
rect -18860 81880 -18640 81920
rect -18860 81810 -18850 81880
rect -18650 81810 -18640 81880
rect -18860 81760 -18640 81810
rect -18360 81990 -18140 82040
rect -18360 81920 -18350 81990
rect -18150 81920 -18140 81990
rect -18360 81880 -18140 81920
rect -18360 81810 -18350 81880
rect -18150 81810 -18140 81880
rect -18360 81760 -18140 81810
rect -17860 81990 -17640 82040
rect -17860 81920 -17850 81990
rect -17650 81920 -17640 81990
rect -17860 81880 -17640 81920
rect -17860 81810 -17850 81880
rect -17650 81810 -17640 81880
rect -17860 81760 -17640 81810
rect -17360 81990 -17140 82040
rect -17360 81920 -17350 81990
rect -17150 81920 -17140 81990
rect -17360 81880 -17140 81920
rect -17360 81810 -17350 81880
rect -17150 81810 -17140 81880
rect -17360 81760 -17140 81810
rect -16860 81990 -16640 82040
rect -16860 81920 -16850 81990
rect -16650 81920 -16640 81990
rect -16860 81880 -16640 81920
rect -16860 81810 -16850 81880
rect -16650 81810 -16640 81880
rect -16860 81760 -16640 81810
rect -16360 81990 -16140 82040
rect -16360 81920 -16350 81990
rect -16150 81920 -16140 81990
rect -16360 81880 -16140 81920
rect -16360 81810 -16350 81880
rect -16150 81810 -16140 81880
rect -16360 81760 -16140 81810
rect -15860 81990 -15640 82040
rect -15860 81920 -15850 81990
rect -15650 81920 -15640 81990
rect -15860 81880 -15640 81920
rect -15860 81810 -15850 81880
rect -15650 81810 -15640 81880
rect -15860 81760 -15640 81810
rect -15360 81990 -15140 82040
rect -15360 81920 -15350 81990
rect -15150 81920 -15140 81990
rect -15360 81880 -15140 81920
rect -15360 81810 -15350 81880
rect -15150 81810 -15140 81880
rect -15360 81760 -15140 81810
rect -14860 81990 -14640 82040
rect -14860 81920 -14850 81990
rect -14650 81920 -14640 81990
rect -14860 81880 -14640 81920
rect -14860 81810 -14850 81880
rect -14650 81810 -14640 81880
rect -14860 81760 -14640 81810
rect -14360 81990 -14140 82040
rect -14360 81920 -14350 81990
rect -14150 81920 -14140 81990
rect -14360 81880 -14140 81920
rect -14360 81810 -14350 81880
rect -14150 81810 -14140 81880
rect -14360 81760 -14140 81810
rect -13860 81990 -13640 82040
rect -13860 81920 -13850 81990
rect -13650 81920 -13640 81990
rect -13860 81880 -13640 81920
rect -13860 81810 -13850 81880
rect -13650 81810 -13640 81880
rect -13860 81760 -13640 81810
rect -13360 81990 -13140 82040
rect -13360 81920 -13350 81990
rect -13150 81920 -13140 81990
rect -13360 81880 -13140 81920
rect -13360 81810 -13350 81880
rect -13150 81810 -13140 81880
rect -13360 81760 -13140 81810
rect -12860 81990 -12640 82040
rect -12860 81920 -12850 81990
rect -12650 81920 -12640 81990
rect -12860 81880 -12640 81920
rect -12860 81810 -12850 81880
rect -12650 81810 -12640 81880
rect -12860 81760 -12640 81810
rect -12360 81990 -12140 82040
rect -12360 81920 -12350 81990
rect -12150 81920 -12140 81990
rect -12360 81880 -12140 81920
rect -12360 81810 -12350 81880
rect -12150 81810 -12140 81880
rect -12360 81760 -12140 81810
rect -11860 81990 -11640 82040
rect -11860 81920 -11850 81990
rect -11650 81920 -11640 81990
rect -11860 81880 -11640 81920
rect -11860 81810 -11850 81880
rect -11650 81810 -11640 81880
rect -11860 81760 -11640 81810
rect -11360 81990 -11140 82040
rect -11360 81920 -11350 81990
rect -11150 81920 -11140 81990
rect -11360 81880 -11140 81920
rect -11360 81810 -11350 81880
rect -11150 81810 -11140 81880
rect -11360 81760 -11140 81810
rect -10860 81990 -10640 82040
rect -10860 81920 -10850 81990
rect -10650 81920 -10640 81990
rect -10860 81880 -10640 81920
rect -10860 81810 -10850 81880
rect -10650 81810 -10640 81880
rect -10860 81760 -10640 81810
rect -10360 81990 -10140 82040
rect -10360 81920 -10350 81990
rect -10150 81920 -10140 81990
rect -10360 81880 -10140 81920
rect -10360 81810 -10350 81880
rect -10150 81810 -10140 81880
rect -10360 81760 -10140 81810
rect -9860 81990 -9640 82040
rect -9860 81920 -9850 81990
rect -9650 81920 -9640 81990
rect -9860 81880 -9640 81920
rect -9860 81810 -9850 81880
rect -9650 81810 -9640 81880
rect -9860 81760 -9640 81810
rect -9360 81990 -9140 82040
rect -9360 81920 -9350 81990
rect -9150 81920 -9140 81990
rect -9360 81880 -9140 81920
rect -9360 81810 -9350 81880
rect -9150 81810 -9140 81880
rect -9360 81760 -9140 81810
rect -8860 81990 -8640 82040
rect -8860 81920 -8850 81990
rect -8650 81920 -8640 81990
rect -8860 81880 -8640 81920
rect -8860 81810 -8850 81880
rect -8650 81810 -8640 81880
rect -8860 81760 -8640 81810
rect -8360 81990 -8140 82040
rect -8360 81920 -8350 81990
rect -8150 81920 -8140 81990
rect -8360 81880 -8140 81920
rect -8360 81810 -8350 81880
rect -8150 81810 -8140 81880
rect -8360 81760 -8140 81810
rect -7860 81990 -7640 82040
rect -7860 81920 -7850 81990
rect -7650 81920 -7640 81990
rect -7860 81880 -7640 81920
rect -7860 81810 -7850 81880
rect -7650 81810 -7640 81880
rect -7860 81760 -7640 81810
rect -7360 81990 -7140 82040
rect -7360 81920 -7350 81990
rect -7150 81920 -7140 81990
rect -7360 81880 -7140 81920
rect -7360 81810 -7350 81880
rect -7150 81810 -7140 81880
rect -7360 81760 -7140 81810
rect -6860 81990 -6640 82040
rect -6860 81920 -6850 81990
rect -6650 81920 -6640 81990
rect -6860 81880 -6640 81920
rect -6860 81810 -6850 81880
rect -6650 81810 -6640 81880
rect -6860 81760 -6640 81810
rect -6360 81990 -6140 82040
rect -6360 81920 -6350 81990
rect -6150 81920 -6140 81990
rect -6360 81880 -6140 81920
rect -6360 81810 -6350 81880
rect -6150 81810 -6140 81880
rect -6360 81760 -6140 81810
rect -5860 81990 -5640 82040
rect -5860 81920 -5850 81990
rect -5650 81920 -5640 81990
rect -5860 81880 -5640 81920
rect -5860 81810 -5850 81880
rect -5650 81810 -5640 81880
rect -5860 81760 -5640 81810
rect -5360 81990 -5140 82040
rect -5360 81920 -5350 81990
rect -5150 81920 -5140 81990
rect -5360 81880 -5140 81920
rect -5360 81810 -5350 81880
rect -5150 81810 -5140 81880
rect -5360 81760 -5140 81810
rect -4860 81990 -4640 82040
rect -4860 81920 -4850 81990
rect -4650 81920 -4640 81990
rect -4860 81880 -4640 81920
rect -4860 81810 -4850 81880
rect -4650 81810 -4640 81880
rect -4860 81760 -4640 81810
rect -4360 81990 -4140 82040
rect -4360 81920 -4350 81990
rect -4150 81920 -4140 81990
rect -4360 81880 -4140 81920
rect -4360 81810 -4350 81880
rect -4150 81810 -4140 81880
rect -4360 81760 -4140 81810
rect -3860 81990 -3640 82040
rect -3860 81920 -3850 81990
rect -3650 81920 -3640 81990
rect -3860 81880 -3640 81920
rect -3860 81810 -3850 81880
rect -3650 81810 -3640 81880
rect -3860 81760 -3640 81810
rect -3360 81990 -3140 82040
rect -3360 81920 -3350 81990
rect -3150 81920 -3140 81990
rect -3360 81880 -3140 81920
rect -3360 81810 -3350 81880
rect -3150 81810 -3140 81880
rect -3360 81760 -3140 81810
rect -2860 81990 -2640 82040
rect -2860 81920 -2850 81990
rect -2650 81920 -2640 81990
rect -2860 81880 -2640 81920
rect -2860 81810 -2850 81880
rect -2650 81810 -2640 81880
rect -2860 81760 -2640 81810
rect -2360 81990 -2140 82040
rect -2360 81920 -2350 81990
rect -2150 81920 -2140 81990
rect -2360 81880 -2140 81920
rect -2360 81810 -2350 81880
rect -2150 81810 -2140 81880
rect -2360 81760 -2140 81810
rect -1860 81990 -1640 82040
rect -1860 81920 -1850 81990
rect -1650 81920 -1640 81990
rect -1860 81880 -1640 81920
rect -1860 81810 -1850 81880
rect -1650 81810 -1640 81880
rect -1860 81760 -1640 81810
rect -1360 81990 -1140 82040
rect -1360 81920 -1350 81990
rect -1150 81920 -1140 81990
rect -1360 81880 -1140 81920
rect -1360 81810 -1350 81880
rect -1150 81810 -1140 81880
rect -1360 81760 -1140 81810
rect -860 81990 -640 82040
rect -860 81920 -850 81990
rect -650 81920 -640 81990
rect -860 81880 -640 81920
rect -860 81810 -850 81880
rect -650 81810 -640 81880
rect -860 81760 -640 81810
rect -360 81990 -140 82040
rect -360 81920 -350 81990
rect -150 81920 -140 81990
rect -360 81880 -140 81920
rect -360 81810 -350 81880
rect -150 81810 -140 81880
rect -360 81760 -140 81810
rect 140 81990 360 82040
rect 140 81920 150 81990
rect 350 81920 360 81990
rect 140 81880 360 81920
rect 140 81810 150 81880
rect 350 81810 360 81880
rect 140 81760 360 81810
rect 640 81990 860 82040
rect 640 81920 650 81990
rect 850 81920 860 81990
rect 640 81880 860 81920
rect 640 81810 650 81880
rect 850 81810 860 81880
rect 640 81760 860 81810
rect 1140 81990 1360 82040
rect 1140 81920 1150 81990
rect 1350 81920 1360 81990
rect 1140 81880 1360 81920
rect 1140 81810 1150 81880
rect 1350 81810 1360 81880
rect 1140 81760 1360 81810
rect 1640 81990 1860 82040
rect 1640 81920 1650 81990
rect 1850 81920 1860 81990
rect 1640 81880 1860 81920
rect 1640 81810 1650 81880
rect 1850 81810 1860 81880
rect 1640 81760 1860 81810
rect 2140 81990 2360 82040
rect 2140 81920 2150 81990
rect 2350 81920 2360 81990
rect 2140 81880 2360 81920
rect 2140 81810 2150 81880
rect 2350 81810 2360 81880
rect 2140 81760 2360 81810
rect 2640 81990 2860 82040
rect 2640 81920 2650 81990
rect 2850 81920 2860 81990
rect 2640 81880 2860 81920
rect 2640 81810 2650 81880
rect 2850 81810 2860 81880
rect 2640 81760 2860 81810
rect 3140 81990 3360 82040
rect 3140 81920 3150 81990
rect 3350 81920 3360 81990
rect 3140 81880 3360 81920
rect 3140 81810 3150 81880
rect 3350 81810 3360 81880
rect 3140 81760 3360 81810
rect 3640 81990 3860 82040
rect 3640 81920 3650 81990
rect 3850 81920 3860 81990
rect 3640 81880 3860 81920
rect 3640 81810 3650 81880
rect 3850 81810 3860 81880
rect 3640 81760 3860 81810
rect 4140 81990 4360 82040
rect 4140 81920 4150 81990
rect 4350 81920 4360 81990
rect 4140 81880 4360 81920
rect 4140 81810 4150 81880
rect 4350 81810 4360 81880
rect 4140 81760 4360 81810
rect 4640 81990 4860 82040
rect 4640 81920 4650 81990
rect 4850 81920 4860 81990
rect 4640 81880 4860 81920
rect 4640 81810 4650 81880
rect 4850 81810 4860 81880
rect 4640 81760 4860 81810
rect 5140 81990 5360 82040
rect 5140 81920 5150 81990
rect 5350 81920 5360 81990
rect 5140 81880 5360 81920
rect 5140 81810 5150 81880
rect 5350 81810 5360 81880
rect 5140 81760 5360 81810
rect 5640 81990 5860 82040
rect 5640 81920 5650 81990
rect 5850 81920 5860 81990
rect 5640 81880 5860 81920
rect 5640 81810 5650 81880
rect 5850 81810 5860 81880
rect 5640 81760 5860 81810
rect 6140 81990 6360 82040
rect 6140 81920 6150 81990
rect 6350 81920 6360 81990
rect 6140 81880 6360 81920
rect 6140 81810 6150 81880
rect 6350 81810 6360 81880
rect 6140 81760 6360 81810
rect 6640 81990 6860 82040
rect 6640 81920 6650 81990
rect 6850 81920 6860 81990
rect 6640 81880 6860 81920
rect 6640 81810 6650 81880
rect 6850 81810 6860 81880
rect 6640 81760 6860 81810
rect 7140 81990 7360 82040
rect 7140 81920 7150 81990
rect 7350 81920 7360 81990
rect 7140 81880 7360 81920
rect 7140 81810 7150 81880
rect 7350 81810 7360 81880
rect 7140 81760 7360 81810
rect 7640 81990 7860 82040
rect 7640 81920 7650 81990
rect 7850 81920 7860 81990
rect 7640 81880 7860 81920
rect 7640 81810 7650 81880
rect 7850 81810 7860 81880
rect 7640 81760 7860 81810
rect 8140 81990 8360 82040
rect 8140 81920 8150 81990
rect 8350 81920 8360 81990
rect 8140 81880 8360 81920
rect 8140 81810 8150 81880
rect 8350 81810 8360 81880
rect 8140 81760 8360 81810
rect 8640 81990 8860 82040
rect 8640 81920 8650 81990
rect 8850 81920 8860 81990
rect 8640 81880 8860 81920
rect 8640 81810 8650 81880
rect 8850 81810 8860 81880
rect 8640 81760 8860 81810
rect 9140 81990 9360 82040
rect 9140 81920 9150 81990
rect 9350 81920 9360 81990
rect 9140 81880 9360 81920
rect 9140 81810 9150 81880
rect 9350 81810 9360 81880
rect 9140 81760 9360 81810
rect 9640 81990 9860 82040
rect 9640 81920 9650 81990
rect 9850 81920 9860 81990
rect 9640 81880 9860 81920
rect 9640 81810 9650 81880
rect 9850 81810 9860 81880
rect 9640 81760 9860 81810
rect 10140 81990 10360 82040
rect 10140 81920 10150 81990
rect 10350 81920 10360 81990
rect 10140 81880 10360 81920
rect 10140 81810 10150 81880
rect 10350 81810 10360 81880
rect 10140 81760 10360 81810
rect 10640 81990 10860 82040
rect 10640 81920 10650 81990
rect 10850 81920 10860 81990
rect 10640 81880 10860 81920
rect 10640 81810 10650 81880
rect 10850 81810 10860 81880
rect 10640 81760 10860 81810
rect 11140 81990 11360 82040
rect 11140 81920 11150 81990
rect 11350 81920 11360 81990
rect 11140 81880 11360 81920
rect 11140 81810 11150 81880
rect 11350 81810 11360 81880
rect 11140 81760 11360 81810
rect 11640 81990 11860 82040
rect 11640 81920 11650 81990
rect 11850 81920 11860 81990
rect 11640 81880 11860 81920
rect 11640 81810 11650 81880
rect 11850 81810 11860 81880
rect 11640 81760 11860 81810
rect 12140 81990 12360 82040
rect 12140 81920 12150 81990
rect 12350 81920 12360 81990
rect 12140 81880 12360 81920
rect 12140 81810 12150 81880
rect 12350 81810 12360 81880
rect 12140 81760 12360 81810
rect 12640 81990 12860 82040
rect 12640 81920 12650 81990
rect 12850 81920 12860 81990
rect 12640 81880 12860 81920
rect 12640 81810 12650 81880
rect 12850 81810 12860 81880
rect 12640 81760 12860 81810
rect 13140 81990 13360 82040
rect 13140 81920 13150 81990
rect 13350 81920 13360 81990
rect 13140 81880 13360 81920
rect 13140 81810 13150 81880
rect 13350 81810 13360 81880
rect 13140 81760 13360 81810
rect 13640 81990 13860 82040
rect 13640 81920 13650 81990
rect 13850 81920 13860 81990
rect 13640 81880 13860 81920
rect 13640 81810 13650 81880
rect 13850 81810 13860 81880
rect 13640 81760 13860 81810
rect 14140 81990 14360 82040
rect 14140 81920 14150 81990
rect 14350 81920 14360 81990
rect 14140 81880 14360 81920
rect 14140 81810 14150 81880
rect 14350 81810 14360 81880
rect 14140 81760 14360 81810
rect 14640 81990 14860 82040
rect 14640 81920 14650 81990
rect 14850 81920 14860 81990
rect 14640 81880 14860 81920
rect 14640 81810 14650 81880
rect 14850 81810 14860 81880
rect 14640 81760 14860 81810
rect 15140 81990 15360 82040
rect 15140 81920 15150 81990
rect 15350 81920 15360 81990
rect 15140 81880 15360 81920
rect 15140 81810 15150 81880
rect 15350 81810 15360 81880
rect 15140 81760 15360 81810
rect 15640 81990 15860 82040
rect 15640 81920 15650 81990
rect 15850 81920 15860 81990
rect 15640 81880 15860 81920
rect 15640 81810 15650 81880
rect 15850 81810 15860 81880
rect 15640 81760 15860 81810
rect 16140 81990 16360 82040
rect 16140 81920 16150 81990
rect 16350 81920 16360 81990
rect 16140 81880 16360 81920
rect 16140 81810 16150 81880
rect 16350 81810 16360 81880
rect 16140 81760 16360 81810
rect 16640 81990 16860 82040
rect 16640 81920 16650 81990
rect 16850 81920 16860 81990
rect 16640 81880 16860 81920
rect 16640 81810 16650 81880
rect 16850 81810 16860 81880
rect 16640 81760 16860 81810
rect 17140 81990 17360 82040
rect 17140 81920 17150 81990
rect 17350 81920 17360 81990
rect 17140 81880 17360 81920
rect 17140 81810 17150 81880
rect 17350 81810 17360 81880
rect 17140 81760 17360 81810
rect 17640 81990 17860 82040
rect 17640 81920 17650 81990
rect 17850 81920 17860 81990
rect 17640 81880 17860 81920
rect 17640 81810 17650 81880
rect 17850 81810 17860 81880
rect 17640 81760 17860 81810
rect 18140 81990 18360 82040
rect 18140 81920 18150 81990
rect 18350 81920 18360 81990
rect 18140 81880 18360 81920
rect 18140 81810 18150 81880
rect 18350 81810 18360 81880
rect 18140 81760 18360 81810
rect 18640 81990 18860 82040
rect 18640 81920 18650 81990
rect 18850 81920 18860 81990
rect 18640 81880 18860 81920
rect 18640 81810 18650 81880
rect 18850 81810 18860 81880
rect 18640 81760 18860 81810
rect 19140 81990 19360 82040
rect 19140 81920 19150 81990
rect 19350 81920 19360 81990
rect 19140 81880 19360 81920
rect 19140 81810 19150 81880
rect 19350 81810 19360 81880
rect 19140 81760 19360 81810
rect 19640 81990 19860 82040
rect 19640 81920 19650 81990
rect 19850 81920 19860 81990
rect 19640 81880 19860 81920
rect 19640 81810 19650 81880
rect 19850 81810 19860 81880
rect 19640 81760 19860 81810
rect 20140 81990 20360 82040
rect 20140 81920 20150 81990
rect 20350 81920 20360 81990
rect 20140 81880 20360 81920
rect 20140 81810 20150 81880
rect 20350 81810 20360 81880
rect 20140 81760 20360 81810
rect 20640 81990 20860 82040
rect 20640 81920 20650 81990
rect 20850 81920 20860 81990
rect 20640 81880 20860 81920
rect 20640 81810 20650 81880
rect 20850 81810 20860 81880
rect 20640 81760 20860 81810
rect 21140 81990 21360 82040
rect 21140 81920 21150 81990
rect 21350 81920 21360 81990
rect 21140 81880 21360 81920
rect 21140 81810 21150 81880
rect 21350 81810 21360 81880
rect 21140 81760 21360 81810
rect 21640 81990 21860 82040
rect 21640 81920 21650 81990
rect 21850 81920 21860 81990
rect 21640 81880 21860 81920
rect 21640 81810 21650 81880
rect 21850 81810 21860 81880
rect 21640 81760 21860 81810
rect 22140 81990 22360 82040
rect 22140 81920 22150 81990
rect 22350 81920 22360 81990
rect 22140 81880 22360 81920
rect 22140 81810 22150 81880
rect 22350 81810 22360 81880
rect 22140 81760 22360 81810
rect 22640 81990 22860 82040
rect 22640 81920 22650 81990
rect 22850 81920 22860 81990
rect 22640 81880 22860 81920
rect 22640 81810 22650 81880
rect 22850 81810 22860 81880
rect 22640 81760 22860 81810
rect 23140 81990 23360 82040
rect 23140 81920 23150 81990
rect 23350 81920 23360 81990
rect 23140 81880 23360 81920
rect 23140 81810 23150 81880
rect 23350 81810 23360 81880
rect 23140 81760 23360 81810
rect 23640 81990 23860 82040
rect 23640 81920 23650 81990
rect 23850 81920 23860 81990
rect 23640 81880 23860 81920
rect 23640 81810 23650 81880
rect 23850 81810 23860 81880
rect 23640 81760 23860 81810
rect 24140 81990 24360 82040
rect 24140 81920 24150 81990
rect 24350 81920 24360 81990
rect 24140 81880 24360 81920
rect 24140 81810 24150 81880
rect 24350 81810 24360 81880
rect 24140 81760 24360 81810
rect 24640 81990 24860 82040
rect 24640 81920 24650 81990
rect 24850 81920 24860 81990
rect 24640 81880 24860 81920
rect 24640 81810 24650 81880
rect 24850 81810 24860 81880
rect 24640 81760 24860 81810
rect 25140 81990 25360 82040
rect 25140 81920 25150 81990
rect 25350 81920 25360 81990
rect 25140 81880 25360 81920
rect 25140 81810 25150 81880
rect 25350 81810 25360 81880
rect 25140 81760 25360 81810
rect 25640 81990 25860 82040
rect 25640 81920 25650 81990
rect 25850 81920 25860 81990
rect 25640 81880 25860 81920
rect 25640 81810 25650 81880
rect 25850 81810 25860 81880
rect 25640 81760 25860 81810
rect 26140 81990 26360 82040
rect 26140 81920 26150 81990
rect 26350 81920 26360 81990
rect 26140 81880 26360 81920
rect 26140 81810 26150 81880
rect 26350 81810 26360 81880
rect 26140 81760 26360 81810
rect 26640 81990 26860 82040
rect 26640 81920 26650 81990
rect 26850 81920 26860 81990
rect 26640 81880 26860 81920
rect 26640 81810 26650 81880
rect 26850 81810 26860 81880
rect 26640 81760 26860 81810
rect 27140 81990 27360 82040
rect 27140 81920 27150 81990
rect 27350 81920 27360 81990
rect 27140 81880 27360 81920
rect 27140 81810 27150 81880
rect 27350 81810 27360 81880
rect 27140 81760 27360 81810
rect 27640 81990 27860 82040
rect 27640 81920 27650 81990
rect 27850 81920 27860 81990
rect 27640 81880 27860 81920
rect 27640 81810 27650 81880
rect 27850 81810 27860 81880
rect 27640 81760 27860 81810
rect 28140 81990 28360 82040
rect 28140 81920 28150 81990
rect 28350 81920 28360 81990
rect 28140 81880 28360 81920
rect 28140 81810 28150 81880
rect 28350 81810 28360 81880
rect 28140 81760 28360 81810
rect 28640 81990 28860 82040
rect 28640 81920 28650 81990
rect 28850 81920 28860 81990
rect 28640 81880 28860 81920
rect 28640 81810 28650 81880
rect 28850 81810 28860 81880
rect 28640 81760 28860 81810
rect 29140 81990 29360 82040
rect 29140 81920 29150 81990
rect 29350 81920 29360 81990
rect 29140 81880 29360 81920
rect 29140 81810 29150 81880
rect 29350 81810 29360 81880
rect 29140 81760 29360 81810
rect 29640 81990 29860 82040
rect 29640 81920 29650 81990
rect 29850 81920 29860 81990
rect 29640 81880 29860 81920
rect 29640 81810 29650 81880
rect 29850 81810 29860 81880
rect 29640 81760 29860 81810
rect 30140 81990 30360 82040
rect 30140 81920 30150 81990
rect 30350 81920 30360 81990
rect 30140 81880 30360 81920
rect 30140 81810 30150 81880
rect 30350 81810 30360 81880
rect 30140 81760 30360 81810
rect 30640 81990 30860 82040
rect 30640 81920 30650 81990
rect 30850 81920 30860 81990
rect 30640 81880 30860 81920
rect 30640 81810 30650 81880
rect 30850 81810 30860 81880
rect 30640 81760 30860 81810
rect 31140 81990 31360 82040
rect 31140 81920 31150 81990
rect 31350 81920 31360 81990
rect 31140 81880 31360 81920
rect 31140 81810 31150 81880
rect 31350 81810 31360 81880
rect 31140 81760 31360 81810
rect 31640 81990 31860 82040
rect 31640 81920 31650 81990
rect 31850 81920 31860 81990
rect 31640 81880 31860 81920
rect 31640 81810 31650 81880
rect 31850 81810 31860 81880
rect 31640 81760 31860 81810
rect 32140 81990 32360 82040
rect 32140 81920 32150 81990
rect 32350 81920 32360 81990
rect 32140 81880 32360 81920
rect 32140 81810 32150 81880
rect 32350 81810 32360 81880
rect 32140 81760 32360 81810
rect 32640 81990 32860 82040
rect 32640 81920 32650 81990
rect 32850 81920 32860 81990
rect 32640 81880 32860 81920
rect 32640 81810 32650 81880
rect 32850 81810 32860 81880
rect 32640 81760 32860 81810
rect 33140 81990 33360 82040
rect 33140 81920 33150 81990
rect 33350 81920 33360 81990
rect 33140 81880 33360 81920
rect 33140 81810 33150 81880
rect 33350 81810 33360 81880
rect 33140 81760 33360 81810
rect 33640 81990 33860 82040
rect 33640 81920 33650 81990
rect 33850 81920 33860 81990
rect 33640 81880 33860 81920
rect 33640 81810 33650 81880
rect 33850 81810 33860 81880
rect 33640 81760 33860 81810
rect 34140 81990 34360 82040
rect 34140 81920 34150 81990
rect 34350 81920 34360 81990
rect 34140 81880 34360 81920
rect 34140 81810 34150 81880
rect 34350 81810 34360 81880
rect 34140 81760 34360 81810
rect 34640 81990 34860 82040
rect 34640 81920 34650 81990
rect 34850 81920 34860 81990
rect 34640 81880 34860 81920
rect 34640 81810 34650 81880
rect 34850 81810 34860 81880
rect 34640 81760 34860 81810
rect 35140 81990 35360 82040
rect 35140 81920 35150 81990
rect 35350 81920 35360 81990
rect 35140 81880 35360 81920
rect 35140 81810 35150 81880
rect 35350 81810 35360 81880
rect 35140 81760 35360 81810
rect 35640 81990 35860 82040
rect 35640 81920 35650 81990
rect 35850 81920 35860 81990
rect 35640 81880 35860 81920
rect 35640 81810 35650 81880
rect 35850 81810 35860 81880
rect 35640 81760 35860 81810
rect 36140 81990 36360 82040
rect 36140 81920 36150 81990
rect 36350 81920 36360 81990
rect 36140 81880 36360 81920
rect 36140 81810 36150 81880
rect 36350 81810 36360 81880
rect 36140 81760 36360 81810
rect 36640 81990 36860 82040
rect 36640 81920 36650 81990
rect 36850 81920 36860 81990
rect 36640 81880 36860 81920
rect 36640 81810 36650 81880
rect 36850 81810 36860 81880
rect 36640 81760 36860 81810
rect 37140 81990 37360 82040
rect 37140 81920 37150 81990
rect 37350 81920 37360 81990
rect 37140 81880 37360 81920
rect 37140 81810 37150 81880
rect 37350 81810 37360 81880
rect 37140 81760 37360 81810
rect 37640 81990 37860 82040
rect 37640 81920 37650 81990
rect 37850 81920 37860 81990
rect 37640 81880 37860 81920
rect 37640 81810 37650 81880
rect 37850 81810 37860 81880
rect 37640 81760 37860 81810
rect 38140 81990 38360 82040
rect 38140 81920 38150 81990
rect 38350 81920 38360 81990
rect 38140 81880 38360 81920
rect 38140 81810 38150 81880
rect 38350 81810 38360 81880
rect 38140 81760 38360 81810
rect 38640 81990 38860 82040
rect 38640 81920 38650 81990
rect 38850 81920 38860 81990
rect 38640 81880 38860 81920
rect 38640 81810 38650 81880
rect 38850 81810 38860 81880
rect 38640 81760 38860 81810
rect 39140 81990 39360 82040
rect 39140 81920 39150 81990
rect 39350 81920 39360 81990
rect 39140 81880 39360 81920
rect 39140 81810 39150 81880
rect 39350 81810 39360 81880
rect 39140 81760 39360 81810
rect 39640 81990 39860 82040
rect 39640 81920 39650 81990
rect 39850 81920 39860 81990
rect 39640 81880 39860 81920
rect 39640 81810 39650 81880
rect 39850 81810 39860 81880
rect 39640 81760 39860 81810
rect 40140 81990 40360 82040
rect 40140 81920 40150 81990
rect 40350 81920 40360 81990
rect 40140 81880 40360 81920
rect 40140 81810 40150 81880
rect 40350 81810 40360 81880
rect 40140 81760 40360 81810
rect 40640 81990 40860 82040
rect 40640 81920 40650 81990
rect 40850 81920 40860 81990
rect 40640 81880 40860 81920
rect 40640 81810 40650 81880
rect 40850 81810 40860 81880
rect 40640 81760 40860 81810
rect 41140 81990 41360 82040
rect 41140 81920 41150 81990
rect 41350 81920 41360 81990
rect 41140 81880 41360 81920
rect 41140 81810 41150 81880
rect 41350 81810 41360 81880
rect 41140 81760 41360 81810
rect 41640 81990 41860 82040
rect 41640 81920 41650 81990
rect 41850 81920 41860 81990
rect 41640 81880 41860 81920
rect 41640 81810 41650 81880
rect 41850 81810 41860 81880
rect 41640 81760 41860 81810
rect 42140 81990 42360 82040
rect 42140 81920 42150 81990
rect 42350 81920 42360 81990
rect 42140 81880 42360 81920
rect 42140 81810 42150 81880
rect 42350 81810 42360 81880
rect 42140 81760 42360 81810
rect 42640 81990 42860 82040
rect 42640 81920 42650 81990
rect 42850 81920 42860 81990
rect 42640 81880 42860 81920
rect 42640 81810 42650 81880
rect 42850 81810 42860 81880
rect 42640 81760 42860 81810
rect 43140 81990 43360 82040
rect 43140 81920 43150 81990
rect 43350 81920 43360 81990
rect 43140 81880 43360 81920
rect 43140 81810 43150 81880
rect 43350 81810 43360 81880
rect 43140 81760 43360 81810
rect 43640 81990 43860 82040
rect 43640 81920 43650 81990
rect 43850 81920 43860 81990
rect 43640 81880 43860 81920
rect 43640 81810 43650 81880
rect 43850 81810 43860 81880
rect 43640 81760 43860 81810
rect 44140 81990 44360 82040
rect 44140 81920 44150 81990
rect 44350 81920 44360 81990
rect 44140 81880 44360 81920
rect 44140 81810 44150 81880
rect 44350 81810 44360 81880
rect 44140 81760 44360 81810
rect 44640 81990 44860 82040
rect 44640 81920 44650 81990
rect 44850 81920 44860 81990
rect 44640 81880 44860 81920
rect 44640 81810 44650 81880
rect 44850 81810 44860 81880
rect 44640 81760 44860 81810
rect 45140 81990 45360 82040
rect 45140 81920 45150 81990
rect 45350 81920 45360 81990
rect 45140 81880 45360 81920
rect 45140 81810 45150 81880
rect 45350 81810 45360 81880
rect 45140 81760 45360 81810
rect 45640 81990 45860 82040
rect 45640 81920 45650 81990
rect 45850 81920 45860 81990
rect 45640 81880 45860 81920
rect 45640 81810 45650 81880
rect 45850 81810 45860 81880
rect 45640 81760 45860 81810
rect 46140 81990 46360 82040
rect 46140 81920 46150 81990
rect 46350 81920 46360 81990
rect 46140 81880 46360 81920
rect 46140 81810 46150 81880
rect 46350 81810 46360 81880
rect 46140 81760 46360 81810
rect 46640 81990 46860 82040
rect 46640 81920 46650 81990
rect 46850 81920 46860 81990
rect 46640 81880 46860 81920
rect 46640 81810 46650 81880
rect 46850 81810 46860 81880
rect 46640 81760 46860 81810
rect 47140 81990 47360 82040
rect 47140 81920 47150 81990
rect 47350 81920 47360 81990
rect 47140 81880 47360 81920
rect 47140 81810 47150 81880
rect 47350 81810 47360 81880
rect 47140 81760 47360 81810
rect 47640 81990 47860 82040
rect 47640 81920 47650 81990
rect 47850 81920 47860 81990
rect 47640 81880 47860 81920
rect 47640 81810 47650 81880
rect 47850 81810 47860 81880
rect 47640 81760 47860 81810
rect 48140 81990 48360 82040
rect 48140 81920 48150 81990
rect 48350 81920 48360 81990
rect 48140 81880 48360 81920
rect 48140 81810 48150 81880
rect 48350 81810 48360 81880
rect 48140 81760 48360 81810
rect 48640 81990 48860 82040
rect 48640 81920 48650 81990
rect 48850 81920 48860 81990
rect 48640 81880 48860 81920
rect 48640 81810 48650 81880
rect 48850 81810 48860 81880
rect 48640 81760 48860 81810
rect 49140 81990 49360 82040
rect 49140 81920 49150 81990
rect 49350 81920 49360 81990
rect 49140 81880 49360 81920
rect 49140 81810 49150 81880
rect 49350 81810 49360 81880
rect 49140 81760 49360 81810
rect 49640 81990 49860 82040
rect 49640 81920 49650 81990
rect 49850 81920 49860 81990
rect 49640 81880 49860 81920
rect 49640 81810 49650 81880
rect 49850 81810 49860 81880
rect 49640 81760 49860 81810
rect 50140 81990 50360 82040
rect 50140 81920 50150 81990
rect 50350 81920 50360 81990
rect 50140 81880 50360 81920
rect 50140 81810 50150 81880
rect 50350 81810 50360 81880
rect 50140 81760 50360 81810
rect 50640 81990 50860 82040
rect 50640 81920 50650 81990
rect 50850 81920 50860 81990
rect 50640 81880 50860 81920
rect 50640 81810 50650 81880
rect 50850 81810 50860 81880
rect 50640 81760 50860 81810
rect 51140 81990 51360 82040
rect 51140 81920 51150 81990
rect 51350 81920 51360 81990
rect 51140 81880 51360 81920
rect 51140 81810 51150 81880
rect 51350 81810 51360 81880
rect 51140 81760 51360 81810
rect 51640 81990 51860 82040
rect 51640 81920 51650 81990
rect 51850 81920 51860 81990
rect 51640 81880 51860 81920
rect 51640 81810 51650 81880
rect 51850 81810 51860 81880
rect 51640 81760 51860 81810
rect 52140 81990 52360 82040
rect 52140 81920 52150 81990
rect 52350 81920 52360 81990
rect 52140 81880 52360 81920
rect 52140 81810 52150 81880
rect 52350 81810 52360 81880
rect 52140 81760 52360 81810
rect 52640 81990 52860 82040
rect 52640 81920 52650 81990
rect 52850 81920 52860 81990
rect 52640 81880 52860 81920
rect 52640 81810 52650 81880
rect 52850 81810 52860 81880
rect 52640 81760 52860 81810
rect 53140 81990 53360 82040
rect 53140 81920 53150 81990
rect 53350 81920 53360 81990
rect 53140 81880 53360 81920
rect 53140 81810 53150 81880
rect 53350 81810 53360 81880
rect 53140 81760 53360 81810
rect 53640 81990 53860 82040
rect 53640 81920 53650 81990
rect 53850 81920 53860 81990
rect 53640 81880 53860 81920
rect 53640 81810 53650 81880
rect 53850 81810 53860 81880
rect 53640 81760 53860 81810
rect 54140 81990 54360 82040
rect 54140 81920 54150 81990
rect 54350 81920 54360 81990
rect 54140 81880 54360 81920
rect 54140 81810 54150 81880
rect 54350 81810 54360 81880
rect 54140 81760 54360 81810
rect 54640 81990 54860 82040
rect 54640 81920 54650 81990
rect 54850 81920 54860 81990
rect 54640 81880 54860 81920
rect 54640 81810 54650 81880
rect 54850 81810 54860 81880
rect 54640 81760 54860 81810
rect 55140 81990 55360 82040
rect 55140 81920 55150 81990
rect 55350 81920 55360 81990
rect 55140 81880 55360 81920
rect 55140 81810 55150 81880
rect 55350 81810 55360 81880
rect 55140 81760 55360 81810
rect 55640 81990 55860 82040
rect 55640 81920 55650 81990
rect 55850 81920 55860 81990
rect 55640 81880 55860 81920
rect 55640 81810 55650 81880
rect 55850 81810 55860 81880
rect 55640 81760 55860 81810
rect 56140 81990 56360 82040
rect 56140 81920 56150 81990
rect 56350 81920 56360 81990
rect 56140 81880 56360 81920
rect 56140 81810 56150 81880
rect 56350 81810 56360 81880
rect 56140 81760 56360 81810
rect 56640 81990 56860 82040
rect 56640 81920 56650 81990
rect 56850 81920 56860 81990
rect 56640 81880 56860 81920
rect 56640 81810 56650 81880
rect 56850 81810 56860 81880
rect 56640 81760 56860 81810
rect 57140 81990 57360 82040
rect 57140 81920 57150 81990
rect 57350 81920 57360 81990
rect 57140 81880 57360 81920
rect 57140 81810 57150 81880
rect 57350 81810 57360 81880
rect 57140 81760 57360 81810
rect 57640 81990 57860 82040
rect 57640 81920 57650 81990
rect 57850 81920 57860 81990
rect 57640 81880 57860 81920
rect 57640 81810 57650 81880
rect 57850 81810 57860 81880
rect 57640 81760 57860 81810
rect 58140 81990 58360 82040
rect 58140 81920 58150 81990
rect 58350 81920 58360 81990
rect 58140 81880 58360 81920
rect 58140 81810 58150 81880
rect 58350 81810 58360 81880
rect 58140 81760 58360 81810
rect 58640 81990 58860 82040
rect 58640 81920 58650 81990
rect 58850 81920 58860 81990
rect 58640 81880 58860 81920
rect 58640 81810 58650 81880
rect 58850 81810 58860 81880
rect 58640 81760 58860 81810
rect 59140 81990 59360 82040
rect 59140 81920 59150 81990
rect 59350 81920 59360 81990
rect 59140 81880 59360 81920
rect 59140 81810 59150 81880
rect 59350 81810 59360 81880
rect 59140 81760 59360 81810
rect 59640 81990 59860 82040
rect 59640 81920 59650 81990
rect 59850 81920 59860 81990
rect 59640 81880 59860 81920
rect 59640 81810 59650 81880
rect 59850 81810 59860 81880
rect 59640 81760 59860 81810
rect 60140 81990 60360 82040
rect 60140 81920 60150 81990
rect 60350 81920 60360 81990
rect 60140 81880 60360 81920
rect 60140 81810 60150 81880
rect 60350 81810 60360 81880
rect 60140 81760 60360 81810
rect 60640 81990 60860 82040
rect 60640 81920 60650 81990
rect 60850 81920 60860 81990
rect 60640 81880 60860 81920
rect 60640 81810 60650 81880
rect 60850 81810 60860 81880
rect 60640 81760 60860 81810
rect 61140 81990 61360 82040
rect 61140 81920 61150 81990
rect 61350 81920 61360 81990
rect 61140 81880 61360 81920
rect 61140 81810 61150 81880
rect 61350 81810 61360 81880
rect 61140 81760 61360 81810
rect 61640 81990 61860 82040
rect 61640 81920 61650 81990
rect 61850 81920 61860 81990
rect 61640 81880 61860 81920
rect 61640 81810 61650 81880
rect 61850 81810 61860 81880
rect 61640 81760 61860 81810
rect 62140 81990 62360 82040
rect 62140 81920 62150 81990
rect 62350 81920 62360 81990
rect 62140 81880 62360 81920
rect 62140 81810 62150 81880
rect 62350 81810 62360 81880
rect 62140 81760 62360 81810
rect 62640 81990 62860 82040
rect 62640 81920 62650 81990
rect 62850 81920 62860 81990
rect 62640 81880 62860 81920
rect 62640 81810 62650 81880
rect 62850 81810 62860 81880
rect 62640 81760 62860 81810
rect 63140 81990 63360 82040
rect 63140 81920 63150 81990
rect 63350 81920 63360 81990
rect 63140 81880 63360 81920
rect 63140 81810 63150 81880
rect 63350 81810 63360 81880
rect 63140 81760 63360 81810
rect 63640 81990 63860 82040
rect 63640 81920 63650 81990
rect 63850 81920 63860 81990
rect 63640 81880 63860 81920
rect 63640 81810 63650 81880
rect 63850 81810 63860 81880
rect 63640 81760 63860 81810
rect 64140 81990 64360 82040
rect 64140 81920 64150 81990
rect 64350 81920 64360 81990
rect 64140 81880 64360 81920
rect 64140 81810 64150 81880
rect 64350 81810 64360 81880
rect 64140 81760 64360 81810
rect 64640 81990 64860 82040
rect 64640 81920 64650 81990
rect 64850 81920 64860 81990
rect 64640 81880 64860 81920
rect 64640 81810 64650 81880
rect 64850 81810 64860 81880
rect 64640 81760 64860 81810
rect 65140 81990 65360 82040
rect 65140 81920 65150 81990
rect 65350 81920 65360 81990
rect 65140 81880 65360 81920
rect 65140 81810 65150 81880
rect 65350 81810 65360 81880
rect 65140 81760 65360 81810
rect 65640 81990 65860 82040
rect 65640 81920 65650 81990
rect 65850 81920 65860 81990
rect 65640 81880 65860 81920
rect 65640 81810 65650 81880
rect 65850 81810 65860 81880
rect 65640 81760 65860 81810
rect 66140 81990 66360 82040
rect 66140 81920 66150 81990
rect 66350 81920 66360 81990
rect 66140 81880 66360 81920
rect 66140 81810 66150 81880
rect 66350 81810 66360 81880
rect 66140 81760 66360 81810
rect 66640 81990 66860 82040
rect 66640 81920 66650 81990
rect 66850 81920 66860 81990
rect 66640 81880 66860 81920
rect 66640 81810 66650 81880
rect 66850 81810 66860 81880
rect 66640 81760 66860 81810
rect 67140 81990 67360 82040
rect 67140 81920 67150 81990
rect 67350 81920 67360 81990
rect 67140 81880 67360 81920
rect 67140 81810 67150 81880
rect 67350 81810 67360 81880
rect 67140 81760 67360 81810
rect 67640 81990 67860 82040
rect 67640 81920 67650 81990
rect 67850 81920 67860 81990
rect 67640 81880 67860 81920
rect 67640 81810 67650 81880
rect 67850 81810 67860 81880
rect 67640 81760 67860 81810
rect 68140 81990 68360 82040
rect 68140 81920 68150 81990
rect 68350 81920 68360 81990
rect 68140 81880 68360 81920
rect 68140 81810 68150 81880
rect 68350 81810 68360 81880
rect 68140 81760 68360 81810
rect 68640 81990 68860 82040
rect 68640 81920 68650 81990
rect 68850 81920 68860 81990
rect 68640 81880 68860 81920
rect 68640 81810 68650 81880
rect 68850 81810 68860 81880
rect 68640 81760 68860 81810
rect 69140 81990 69360 82040
rect 69140 81920 69150 81990
rect 69350 81920 69360 81990
rect 69140 81880 69360 81920
rect 69140 81810 69150 81880
rect 69350 81810 69360 81880
rect 69140 81760 69360 81810
rect 69640 81990 69860 82040
rect 69640 81920 69650 81990
rect 69850 81920 69860 81990
rect 69640 81880 69860 81920
rect 69640 81810 69650 81880
rect 69850 81810 69860 81880
rect 69640 81760 69860 81810
rect 70140 81990 70360 82040
rect 70140 81920 70150 81990
rect 70350 81920 70360 81990
rect 70140 81880 70360 81920
rect 70140 81810 70150 81880
rect 70350 81810 70360 81880
rect 70140 81760 70360 81810
rect 70640 81990 70860 82040
rect 70640 81920 70650 81990
rect 70850 81920 70860 81990
rect 70640 81880 70860 81920
rect 70640 81810 70650 81880
rect 70850 81810 70860 81880
rect 70640 81760 70860 81810
rect 71140 81990 71360 82040
rect 71140 81920 71150 81990
rect 71350 81920 71360 81990
rect 71140 81880 71360 81920
rect 71140 81810 71150 81880
rect 71350 81810 71360 81880
rect 71140 81760 71360 81810
rect 71640 81990 71860 82040
rect 71640 81920 71650 81990
rect 71850 81920 71860 81990
rect 71640 81880 71860 81920
rect 71640 81810 71650 81880
rect 71850 81810 71860 81880
rect 71640 81760 71860 81810
rect 72140 81990 72360 82040
rect 72140 81920 72150 81990
rect 72350 81920 72360 81990
rect 72140 81880 72360 81920
rect 72140 81810 72150 81880
rect 72350 81810 72360 81880
rect 72140 81760 72360 81810
rect 72640 81990 72860 82040
rect 72640 81920 72650 81990
rect 72850 81920 72860 81990
rect 72640 81880 72860 81920
rect 72640 81810 72650 81880
rect 72850 81810 72860 81880
rect 72640 81760 72860 81810
rect 73140 81990 73360 82040
rect 73140 81920 73150 81990
rect 73350 81920 73360 81990
rect 73140 81880 73360 81920
rect 73140 81810 73150 81880
rect 73350 81810 73360 81880
rect 73140 81760 73360 81810
rect 73640 81990 73860 82040
rect 73640 81920 73650 81990
rect 73850 81920 73860 81990
rect 73640 81880 73860 81920
rect 73640 81810 73650 81880
rect 73850 81810 73860 81880
rect 73640 81760 73860 81810
rect 74140 81990 74360 82040
rect 74140 81920 74150 81990
rect 74350 81920 74360 81990
rect 74140 81880 74360 81920
rect 74140 81810 74150 81880
rect 74350 81810 74360 81880
rect 74140 81760 74360 81810
rect 74640 81990 74860 82040
rect 74640 81920 74650 81990
rect 74850 81920 74860 81990
rect 74640 81880 74860 81920
rect 74640 81810 74650 81880
rect 74850 81810 74860 81880
rect 74640 81760 74860 81810
rect 75140 81990 75360 82040
rect 75140 81920 75150 81990
rect 75350 81920 75360 81990
rect 75140 81880 75360 81920
rect 75140 81810 75150 81880
rect 75350 81810 75360 81880
rect 75140 81760 75360 81810
rect 75640 81990 75860 82040
rect 75640 81920 75650 81990
rect 75850 81920 75860 81990
rect 75640 81880 75860 81920
rect 75640 81810 75650 81880
rect 75850 81810 75860 81880
rect 75640 81760 75860 81810
rect 76140 81990 76360 82040
rect 76140 81920 76150 81990
rect 76350 81920 76360 81990
rect 76140 81880 76360 81920
rect 76140 81810 76150 81880
rect 76350 81810 76360 81880
rect 76140 81760 76360 81810
rect 76640 81990 76860 82040
rect 76640 81920 76650 81990
rect 76850 81920 76860 81990
rect 76640 81880 76860 81920
rect 76640 81810 76650 81880
rect 76850 81810 76860 81880
rect 76640 81760 76860 81810
rect 77140 81990 77360 82040
rect 77140 81920 77150 81990
rect 77350 81920 77360 81990
rect 77140 81880 77360 81920
rect 77140 81810 77150 81880
rect 77350 81810 77360 81880
rect 77140 81760 77360 81810
rect 77640 81990 77860 82040
rect 77640 81920 77650 81990
rect 77850 81920 77860 81990
rect 77640 81880 77860 81920
rect 77640 81810 77650 81880
rect 77850 81810 77860 81880
rect 77640 81760 77860 81810
rect 78140 81990 78360 82040
rect 78140 81920 78150 81990
rect 78350 81920 78360 81990
rect 78140 81880 78360 81920
rect 78140 81810 78150 81880
rect 78350 81810 78360 81880
rect 78140 81760 78360 81810
rect 78640 81990 78860 82040
rect 78640 81920 78650 81990
rect 78850 81920 78860 81990
rect 78640 81880 78860 81920
rect 78640 81810 78650 81880
rect 78850 81810 78860 81880
rect 78640 81760 78860 81810
rect 79140 81990 79360 82040
rect 79140 81920 79150 81990
rect 79350 81920 79360 81990
rect 79140 81880 79360 81920
rect 79140 81810 79150 81880
rect 79350 81810 79360 81880
rect 79140 81760 79360 81810
rect 79640 81990 79860 82040
rect 79640 81920 79650 81990
rect 79850 81920 79860 81990
rect 79640 81880 79860 81920
rect 79640 81810 79650 81880
rect 79850 81810 79860 81880
rect 79640 81760 79860 81810
rect 80140 81990 80360 82040
rect 80140 81920 80150 81990
rect 80350 81920 80360 81990
rect 80140 81880 80360 81920
rect 80140 81810 80150 81880
rect 80350 81810 80360 81880
rect 80140 81760 80360 81810
rect 80640 81990 80860 82040
rect 80640 81920 80650 81990
rect 80850 81920 80860 81990
rect 80640 81880 80860 81920
rect 80640 81810 80650 81880
rect 80850 81810 80860 81880
rect 80640 81760 80860 81810
rect 81140 81990 81360 82040
rect 81140 81920 81150 81990
rect 81350 81920 81360 81990
rect 81140 81880 81360 81920
rect 81140 81810 81150 81880
rect 81350 81810 81360 81880
rect 81140 81760 81360 81810
rect 81640 81990 81860 82040
rect 81640 81920 81650 81990
rect 81850 81920 81860 81990
rect 81640 81880 81860 81920
rect 81640 81810 81650 81880
rect 81850 81810 81860 81880
rect 81640 81760 81860 81810
rect 82140 81990 82360 82040
rect 82140 81920 82150 81990
rect 82350 81920 82360 81990
rect 82140 81880 82360 81920
rect 82140 81810 82150 81880
rect 82350 81810 82360 81880
rect 82140 81760 82360 81810
rect 82640 81990 82860 82040
rect 82640 81920 82650 81990
rect 82850 81920 82860 81990
rect 82640 81880 82860 81920
rect 82640 81810 82650 81880
rect 82850 81810 82860 81880
rect 82640 81760 82860 81810
rect 83140 81990 83360 82040
rect 83140 81920 83150 81990
rect 83350 81920 83360 81990
rect 83140 81880 83360 81920
rect 83140 81810 83150 81880
rect 83350 81810 83360 81880
rect 83140 81760 83360 81810
rect 83640 81990 83860 82040
rect 83640 81920 83650 81990
rect 83850 81920 83860 81990
rect 83640 81880 83860 81920
rect 83640 81810 83650 81880
rect 83850 81810 83860 81880
rect 83640 81760 83860 81810
rect 84140 81990 84360 82040
rect 84140 81920 84150 81990
rect 84350 81920 84360 81990
rect 84140 81880 84360 81920
rect 84140 81810 84150 81880
rect 84350 81810 84360 81880
rect 84140 81760 84360 81810
rect 84640 81990 84860 82040
rect 84640 81920 84650 81990
rect 84850 81920 84860 81990
rect 84640 81880 84860 81920
rect 84640 81810 84650 81880
rect 84850 81810 84860 81880
rect 84640 81760 84860 81810
rect 85140 81990 85360 82040
rect 85140 81920 85150 81990
rect 85350 81920 85360 81990
rect 85140 81880 85360 81920
rect 85140 81810 85150 81880
rect 85350 81810 85360 81880
rect 85140 81760 85360 81810
rect 85640 81990 85860 82040
rect 85640 81920 85650 81990
rect 85850 81920 85860 81990
rect 85640 81880 85860 81920
rect 85640 81810 85650 81880
rect 85850 81810 85860 81880
rect 85640 81760 85860 81810
rect 86140 81990 86360 82040
rect 86140 81920 86150 81990
rect 86350 81920 86360 81990
rect 86140 81880 86360 81920
rect 86140 81810 86150 81880
rect 86350 81810 86360 81880
rect 86140 81760 86360 81810
rect 86640 81990 86860 82040
rect 86640 81920 86650 81990
rect 86850 81920 86860 81990
rect 86640 81880 86860 81920
rect 86640 81810 86650 81880
rect 86850 81810 86860 81880
rect 86640 81760 86860 81810
rect 87140 81990 87360 82040
rect 87140 81920 87150 81990
rect 87350 81920 87360 81990
rect 87140 81880 87360 81920
rect 87140 81810 87150 81880
rect 87350 81810 87360 81880
rect 87140 81760 87360 81810
rect 87640 81990 87860 82040
rect 87640 81920 87650 81990
rect 87850 81920 87860 81990
rect 87640 81880 87860 81920
rect 87640 81810 87650 81880
rect 87850 81810 87860 81880
rect 87640 81760 87860 81810
rect 88140 81990 88360 82040
rect 88140 81920 88150 81990
rect 88350 81920 88360 81990
rect 88140 81880 88360 81920
rect 88140 81810 88150 81880
rect 88350 81810 88360 81880
rect 88140 81760 88360 81810
rect 88640 81990 88860 82040
rect 88640 81920 88650 81990
rect 88850 81920 88860 81990
rect 88640 81880 88860 81920
rect 88640 81810 88650 81880
rect 88850 81810 88860 81880
rect 88640 81760 88860 81810
rect 89140 81990 89360 82040
rect 89140 81920 89150 81990
rect 89350 81920 89360 81990
rect 89140 81880 89360 81920
rect 89140 81810 89150 81880
rect 89350 81810 89360 81880
rect 89140 81760 89360 81810
rect 89640 81990 89860 82040
rect 89640 81920 89650 81990
rect 89850 81920 89860 81990
rect 89640 81880 89860 81920
rect 89640 81810 89650 81880
rect 89850 81810 89860 81880
rect 89640 81760 89860 81810
rect 90140 81990 90360 82040
rect 90140 81920 90150 81990
rect 90350 81920 90360 81990
rect 90140 81880 90360 81920
rect 90140 81810 90150 81880
rect 90350 81810 90360 81880
rect 90140 81760 90360 81810
rect 90640 81990 90860 82040
rect 90640 81920 90650 81990
rect 90850 81920 90860 81990
rect 90640 81880 90860 81920
rect 90640 81810 90650 81880
rect 90850 81810 90860 81880
rect 90640 81760 90860 81810
rect 91140 81990 91360 82040
rect 91140 81920 91150 81990
rect 91350 81920 91360 81990
rect 91140 81880 91360 81920
rect 91140 81810 91150 81880
rect 91350 81810 91360 81880
rect 91140 81760 91360 81810
rect 91640 81990 91860 82040
rect 91640 81920 91650 81990
rect 91850 81920 91860 81990
rect 91640 81880 91860 81920
rect 91640 81810 91650 81880
rect 91850 81810 91860 81880
rect 91640 81760 91860 81810
rect 92140 81990 92360 82040
rect 92140 81920 92150 81990
rect 92350 81920 92360 81990
rect 92140 81880 92360 81920
rect 92140 81810 92150 81880
rect 92350 81810 92360 81880
rect 92140 81760 92360 81810
rect 92640 81990 92860 82040
rect 92640 81920 92650 81990
rect 92850 81920 92860 81990
rect 92640 81880 92860 81920
rect 92640 81810 92650 81880
rect 92850 81810 92860 81880
rect 92640 81760 92860 81810
rect 93140 81990 93360 82040
rect 93140 81920 93150 81990
rect 93350 81920 93360 81990
rect 93140 81880 93360 81920
rect 93140 81810 93150 81880
rect 93350 81810 93360 81880
rect 93140 81760 93360 81810
rect 93640 81990 93860 82040
rect 93640 81920 93650 81990
rect 93850 81920 93860 81990
rect 93640 81880 93860 81920
rect 93640 81810 93650 81880
rect 93850 81810 93860 81880
rect 93640 81760 93860 81810
rect 94140 81990 94360 82040
rect 94140 81920 94150 81990
rect 94350 81920 94360 81990
rect 94140 81880 94360 81920
rect 94140 81810 94150 81880
rect 94350 81810 94360 81880
rect 94140 81760 94360 81810
rect 94640 81990 94860 82040
rect 94640 81920 94650 81990
rect 94850 81920 94860 81990
rect 94640 81880 94860 81920
rect 94640 81810 94650 81880
rect 94850 81810 94860 81880
rect 94640 81760 94860 81810
rect 95140 81990 95360 82040
rect 95140 81920 95150 81990
rect 95350 81920 95360 81990
rect 95140 81880 95360 81920
rect 95140 81810 95150 81880
rect 95350 81810 95360 81880
rect 95140 81760 95360 81810
rect 95640 81990 95860 82040
rect 95640 81920 95650 81990
rect 95850 81920 95860 81990
rect 95640 81880 95860 81920
rect 95640 81810 95650 81880
rect 95850 81810 95860 81880
rect 95640 81760 95860 81810
rect 96140 81990 96360 82040
rect 96140 81920 96150 81990
rect 96350 81920 96360 81990
rect 96140 81880 96360 81920
rect 96140 81810 96150 81880
rect 96350 81810 96360 81880
rect 96140 81760 96360 81810
rect 96640 81990 96860 82040
rect 96640 81920 96650 81990
rect 96850 81920 96860 81990
rect 96640 81880 96860 81920
rect 96640 81810 96650 81880
rect 96850 81810 96860 81880
rect 96640 81760 96860 81810
rect 97140 81990 97360 82040
rect 97140 81920 97150 81990
rect 97350 81920 97360 81990
rect 97140 81880 97360 81920
rect 97140 81810 97150 81880
rect 97350 81810 97360 81880
rect 97140 81760 97360 81810
rect 97640 81990 97860 82040
rect 97640 81920 97650 81990
rect 97850 81920 97860 81990
rect 97640 81880 97860 81920
rect 97640 81810 97650 81880
rect 97850 81810 97860 81880
rect 97640 81760 97860 81810
rect 98140 81990 98360 82040
rect 98140 81920 98150 81990
rect 98350 81920 98360 81990
rect 98140 81880 98360 81920
rect 98140 81810 98150 81880
rect 98350 81810 98360 81880
rect 98140 81760 98360 81810
rect 98640 81990 98860 82040
rect 98640 81920 98650 81990
rect 98850 81920 98860 81990
rect 98640 81880 98860 81920
rect 98640 81810 98650 81880
rect 98850 81810 98860 81880
rect 98640 81760 98860 81810
rect 99140 81990 99360 82040
rect 99140 81920 99150 81990
rect 99350 81920 99360 81990
rect 99140 81880 99360 81920
rect 99140 81810 99150 81880
rect 99350 81810 99360 81880
rect 99140 81760 99360 81810
rect 99640 81990 99860 82040
rect 99640 81920 99650 81990
rect 99850 81920 99860 81990
rect 99640 81880 99860 81920
rect 99640 81810 99650 81880
rect 99850 81810 99860 81880
rect 99640 81760 99860 81810
rect 100140 81990 100360 82040
rect 100140 81920 100150 81990
rect 100350 81920 100360 81990
rect 100140 81880 100360 81920
rect 100140 81810 100150 81880
rect 100350 81810 100360 81880
rect 100140 81760 100360 81810
rect -83500 81750 100500 81760
rect -83500 81550 -83480 81750
rect -83410 81550 -83090 81750
rect -83020 81550 -82980 81750
rect -82910 81550 -82590 81750
rect -82520 81550 -82480 81750
rect -82410 81550 -82090 81750
rect -82020 81550 -81980 81750
rect -81910 81550 -81590 81750
rect -81520 81550 -81480 81750
rect -81410 81550 -81090 81750
rect -81020 81550 -80980 81750
rect -80910 81550 -80590 81750
rect -80520 81550 -80480 81750
rect -80410 81550 -80090 81750
rect -80020 81550 -79980 81750
rect -79910 81550 -79590 81750
rect -79520 81550 -79480 81750
rect -79410 81550 -79090 81750
rect -79020 81550 -78980 81750
rect -78910 81550 -78590 81750
rect -78520 81550 -78480 81750
rect -78410 81550 -78090 81750
rect -78020 81550 -77980 81750
rect -77910 81550 -77590 81750
rect -77520 81550 -77480 81750
rect -77410 81550 -77090 81750
rect -77020 81550 -76980 81750
rect -76910 81550 -76590 81750
rect -76520 81550 -76480 81750
rect -76410 81550 -76090 81750
rect -76020 81550 -75980 81750
rect -75910 81550 -75590 81750
rect -75520 81550 -75480 81750
rect -75410 81550 -75090 81750
rect -75020 81550 -74980 81750
rect -74910 81550 -74590 81750
rect -74520 81550 -74480 81750
rect -74410 81550 -74090 81750
rect -74020 81550 -73980 81750
rect -73910 81550 -73590 81750
rect -73520 81550 -73480 81750
rect -73410 81550 -73090 81750
rect -73020 81550 -72980 81750
rect -72910 81550 -72590 81750
rect -72520 81550 -72480 81750
rect -72410 81550 -72090 81750
rect -72020 81550 -71980 81750
rect -71910 81550 -71590 81750
rect -71520 81550 -71480 81750
rect -71410 81550 -71090 81750
rect -71020 81550 -70980 81750
rect -70910 81550 -70590 81750
rect -70520 81550 -70480 81750
rect -70410 81550 -70090 81750
rect -70020 81550 -69980 81750
rect -69910 81550 -69590 81750
rect -69520 81550 -69480 81750
rect -69410 81550 -69090 81750
rect -69020 81550 -68980 81750
rect -68910 81550 -68590 81750
rect -68520 81550 -68480 81750
rect -68410 81550 -68090 81750
rect -68020 81550 -67980 81750
rect -67910 81550 -67590 81750
rect -67520 81550 -67480 81750
rect -67410 81550 -67090 81750
rect -67020 81550 -66980 81750
rect -66910 81550 -66590 81750
rect -66520 81550 -66480 81750
rect -66410 81550 -66090 81750
rect -66020 81550 -65980 81750
rect -65910 81550 -65590 81750
rect -65520 81550 -65480 81750
rect -65410 81550 -65090 81750
rect -65020 81550 -64980 81750
rect -64910 81550 -64590 81750
rect -64520 81550 -64480 81750
rect -64410 81550 -64090 81750
rect -64020 81550 -63980 81750
rect -63910 81550 -63590 81750
rect -63520 81550 -63480 81750
rect -63410 81550 -63090 81750
rect -63020 81550 -62980 81750
rect -62910 81550 -62590 81750
rect -62520 81550 -62480 81750
rect -62410 81550 -62090 81750
rect -62020 81550 -61980 81750
rect -61910 81550 -61590 81750
rect -61520 81550 -61480 81750
rect -61410 81550 -61090 81750
rect -61020 81550 -60980 81750
rect -60910 81550 -60590 81750
rect -60520 81550 -60480 81750
rect -60410 81550 -60090 81750
rect -60020 81550 -59980 81750
rect -59910 81550 -59590 81750
rect -59520 81550 -59480 81750
rect -59410 81550 -59090 81750
rect -59020 81550 -58980 81750
rect -58910 81550 -58590 81750
rect -58520 81550 -58480 81750
rect -58410 81550 -58090 81750
rect -58020 81550 -57980 81750
rect -57910 81550 -57590 81750
rect -57520 81550 -57480 81750
rect -57410 81550 -57090 81750
rect -57020 81550 -56980 81750
rect -56910 81550 -56590 81750
rect -56520 81550 -56480 81750
rect -56410 81550 -56090 81750
rect -56020 81550 -55980 81750
rect -55910 81550 -55590 81750
rect -55520 81550 -55480 81750
rect -55410 81550 -55090 81750
rect -55020 81550 -54980 81750
rect -54910 81550 -54590 81750
rect -54520 81550 -54480 81750
rect -54410 81550 -54090 81750
rect -54020 81550 -53980 81750
rect -53910 81550 -53590 81750
rect -53520 81550 -53480 81750
rect -53410 81550 -53090 81750
rect -53020 81550 -52980 81750
rect -52910 81550 -52590 81750
rect -52520 81550 -52480 81750
rect -52410 81550 -52090 81750
rect -52020 81550 -51980 81750
rect -51910 81550 -51590 81750
rect -51520 81550 -51480 81750
rect -51410 81550 -51090 81750
rect -51020 81550 -50980 81750
rect -50910 81550 -50590 81750
rect -50520 81550 -50480 81750
rect -50410 81550 -50090 81750
rect -50020 81550 -49980 81750
rect -49910 81550 -49590 81750
rect -49520 81550 -49480 81750
rect -49410 81550 -49090 81750
rect -49020 81550 -48980 81750
rect -48910 81550 -48590 81750
rect -48520 81550 -48480 81750
rect -48410 81550 -48090 81750
rect -48020 81550 -47980 81750
rect -47910 81550 -47590 81750
rect -47520 81550 -47480 81750
rect -47410 81550 -47090 81750
rect -47020 81550 -46980 81750
rect -46910 81550 -46590 81750
rect -46520 81550 -46480 81750
rect -46410 81550 -46090 81750
rect -46020 81550 -45980 81750
rect -45910 81550 -45590 81750
rect -45520 81550 -45480 81750
rect -45410 81550 -45090 81750
rect -45020 81550 -44980 81750
rect -44910 81550 -44590 81750
rect -44520 81550 -44480 81750
rect -44410 81550 -44090 81750
rect -44020 81550 -43980 81750
rect -43910 81550 -43590 81750
rect -43520 81550 -43480 81750
rect -43410 81550 -43090 81750
rect -43020 81550 -42980 81750
rect -42910 81550 -42590 81750
rect -42520 81550 -42480 81750
rect -42410 81550 -42090 81750
rect -42020 81550 -41980 81750
rect -41910 81550 -41590 81750
rect -41520 81550 -41480 81750
rect -41410 81550 -41090 81750
rect -41020 81550 -40980 81750
rect -40910 81550 -40590 81750
rect -40520 81550 -40480 81750
rect -40410 81550 -40090 81750
rect -40020 81550 -39980 81750
rect -39910 81550 -39590 81750
rect -39520 81550 -39480 81750
rect -39410 81550 -39090 81750
rect -39020 81550 -38980 81750
rect -38910 81550 -38590 81750
rect -38520 81550 -38480 81750
rect -38410 81550 -38090 81750
rect -38020 81550 -37980 81750
rect -37910 81550 -37590 81750
rect -37520 81550 -37480 81750
rect -37410 81550 -37090 81750
rect -37020 81550 -36980 81750
rect -36910 81550 -36590 81750
rect -36520 81550 -36480 81750
rect -36410 81550 -36090 81750
rect -36020 81550 -35980 81750
rect -35910 81550 -35590 81750
rect -35520 81550 -35480 81750
rect -35410 81550 -35090 81750
rect -35020 81550 -34980 81750
rect -34910 81550 -34590 81750
rect -34520 81550 -34480 81750
rect -34410 81550 -34090 81750
rect -34020 81550 -33980 81750
rect -33910 81550 -33590 81750
rect -33520 81550 -33480 81750
rect -33410 81550 -33090 81750
rect -33020 81550 -32980 81750
rect -32910 81550 -32590 81750
rect -32520 81550 -32480 81750
rect -32410 81550 -32090 81750
rect -32020 81550 -31980 81750
rect -31910 81550 -31590 81750
rect -31520 81550 -31480 81750
rect -31410 81550 -31090 81750
rect -31020 81550 -30980 81750
rect -30910 81550 -30590 81750
rect -30520 81550 -30480 81750
rect -30410 81550 -30090 81750
rect -30020 81550 -29980 81750
rect -29910 81550 -29590 81750
rect -29520 81550 -29480 81750
rect -29410 81550 -29090 81750
rect -29020 81550 -28980 81750
rect -28910 81550 -28590 81750
rect -28520 81550 -28480 81750
rect -28410 81550 -28090 81750
rect -28020 81550 -27980 81750
rect -27910 81550 -27590 81750
rect -27520 81550 -27480 81750
rect -27410 81550 -27090 81750
rect -27020 81550 -26980 81750
rect -26910 81550 -26590 81750
rect -26520 81550 -26480 81750
rect -26410 81550 -26090 81750
rect -26020 81550 -25980 81750
rect -25910 81550 -25590 81750
rect -25520 81550 -25480 81750
rect -25410 81550 -25090 81750
rect -25020 81550 -24980 81750
rect -24910 81550 -24590 81750
rect -24520 81550 -24480 81750
rect -24410 81550 -24090 81750
rect -24020 81550 -23980 81750
rect -23910 81550 -23590 81750
rect -23520 81550 -23480 81750
rect -23410 81550 -23090 81750
rect -23020 81550 -22980 81750
rect -22910 81550 -22590 81750
rect -22520 81550 -22480 81750
rect -22410 81550 -22090 81750
rect -22020 81550 -21980 81750
rect -21910 81550 -21590 81750
rect -21520 81550 -21480 81750
rect -21410 81550 -21090 81750
rect -21020 81550 -20980 81750
rect -20910 81550 -20590 81750
rect -20520 81550 -20480 81750
rect -20410 81550 -20090 81750
rect -20020 81550 -19980 81750
rect -19910 81550 -19590 81750
rect -19520 81550 -19480 81750
rect -19410 81550 -19090 81750
rect -19020 81550 -18980 81750
rect -18910 81550 -18590 81750
rect -18520 81550 -18480 81750
rect -18410 81550 -18090 81750
rect -18020 81550 -17980 81750
rect -17910 81550 -17590 81750
rect -17520 81550 -17480 81750
rect -17410 81550 -17090 81750
rect -17020 81550 -16980 81750
rect -16910 81550 -16590 81750
rect -16520 81550 -16480 81750
rect -16410 81550 -16090 81750
rect -16020 81550 -15980 81750
rect -15910 81550 -15590 81750
rect -15520 81550 -15480 81750
rect -15410 81550 -15090 81750
rect -15020 81550 -14980 81750
rect -14910 81550 -14590 81750
rect -14520 81550 -14480 81750
rect -14410 81550 -14090 81750
rect -14020 81550 -13980 81750
rect -13910 81550 -13590 81750
rect -13520 81550 -13480 81750
rect -13410 81550 -13090 81750
rect -13020 81550 -12980 81750
rect -12910 81550 -12590 81750
rect -12520 81550 -12480 81750
rect -12410 81550 -12090 81750
rect -12020 81550 -11980 81750
rect -11910 81550 -11590 81750
rect -11520 81550 -11480 81750
rect -11410 81550 -11090 81750
rect -11020 81550 -10980 81750
rect -10910 81550 -10590 81750
rect -10520 81550 -10480 81750
rect -10410 81550 -10090 81750
rect -10020 81550 -9980 81750
rect -9910 81550 -9590 81750
rect -9520 81550 -9480 81750
rect -9410 81550 -9090 81750
rect -9020 81550 -8980 81750
rect -8910 81550 -8590 81750
rect -8520 81550 -8480 81750
rect -8410 81550 -8090 81750
rect -8020 81550 -7980 81750
rect -7910 81550 -7590 81750
rect -7520 81550 -7480 81750
rect -7410 81550 -7090 81750
rect -7020 81550 -6980 81750
rect -6910 81550 -6590 81750
rect -6520 81550 -6480 81750
rect -6410 81550 -6090 81750
rect -6020 81550 -5980 81750
rect -5910 81550 -5590 81750
rect -5520 81550 -5480 81750
rect -5410 81550 -5090 81750
rect -5020 81550 -4980 81750
rect -4910 81550 -4590 81750
rect -4520 81550 -4480 81750
rect -4410 81550 -4090 81750
rect -4020 81550 -3980 81750
rect -3910 81550 -3590 81750
rect -3520 81550 -3480 81750
rect -3410 81550 -3090 81750
rect -3020 81550 -2980 81750
rect -2910 81550 -2590 81750
rect -2520 81550 -2480 81750
rect -2410 81550 -2090 81750
rect -2020 81550 -1980 81750
rect -1910 81550 -1590 81750
rect -1520 81550 -1480 81750
rect -1410 81550 -1090 81750
rect -1020 81550 -980 81750
rect -910 81550 -590 81750
rect -520 81550 -480 81750
rect -410 81550 -90 81750
rect -20 81550 20 81750
rect 90 81550 410 81750
rect 480 81550 520 81750
rect 590 81550 910 81750
rect 980 81550 1020 81750
rect 1090 81550 1410 81750
rect 1480 81550 1520 81750
rect 1590 81550 1910 81750
rect 1980 81550 2020 81750
rect 2090 81550 2410 81750
rect 2480 81550 2520 81750
rect 2590 81550 2910 81750
rect 2980 81550 3020 81750
rect 3090 81550 3410 81750
rect 3480 81550 3520 81750
rect 3590 81550 3910 81750
rect 3980 81550 4020 81750
rect 4090 81550 4410 81750
rect 4480 81550 4520 81750
rect 4590 81550 4910 81750
rect 4980 81550 5020 81750
rect 5090 81550 5410 81750
rect 5480 81550 5520 81750
rect 5590 81550 5910 81750
rect 5980 81550 6020 81750
rect 6090 81550 6410 81750
rect 6480 81550 6520 81750
rect 6590 81550 6910 81750
rect 6980 81550 7020 81750
rect 7090 81550 7410 81750
rect 7480 81550 7520 81750
rect 7590 81550 7910 81750
rect 7980 81550 8020 81750
rect 8090 81550 8410 81750
rect 8480 81550 8520 81750
rect 8590 81550 8910 81750
rect 8980 81550 9020 81750
rect 9090 81550 9410 81750
rect 9480 81550 9520 81750
rect 9590 81550 9910 81750
rect 9980 81550 10020 81750
rect 10090 81550 10410 81750
rect 10480 81550 10520 81750
rect 10590 81550 10910 81750
rect 10980 81550 11020 81750
rect 11090 81550 11410 81750
rect 11480 81550 11520 81750
rect 11590 81550 11910 81750
rect 11980 81550 12020 81750
rect 12090 81550 12410 81750
rect 12480 81550 12520 81750
rect 12590 81550 12910 81750
rect 12980 81550 13020 81750
rect 13090 81550 13410 81750
rect 13480 81550 13520 81750
rect 13590 81550 13910 81750
rect 13980 81550 14020 81750
rect 14090 81550 14410 81750
rect 14480 81550 14520 81750
rect 14590 81550 14910 81750
rect 14980 81550 15020 81750
rect 15090 81550 15410 81750
rect 15480 81550 15520 81750
rect 15590 81550 15910 81750
rect 15980 81550 16020 81750
rect 16090 81550 16410 81750
rect 16480 81550 16520 81750
rect 16590 81550 16910 81750
rect 16980 81550 17020 81750
rect 17090 81550 17410 81750
rect 17480 81550 17520 81750
rect 17590 81550 17910 81750
rect 17980 81550 18020 81750
rect 18090 81550 18410 81750
rect 18480 81550 18520 81750
rect 18590 81550 18910 81750
rect 18980 81550 19020 81750
rect 19090 81550 19410 81750
rect 19480 81550 19520 81750
rect 19590 81550 19910 81750
rect 19980 81550 20020 81750
rect 20090 81550 20410 81750
rect 20480 81550 20520 81750
rect 20590 81550 20910 81750
rect 20980 81550 21020 81750
rect 21090 81550 21410 81750
rect 21480 81550 21520 81750
rect 21590 81550 21910 81750
rect 21980 81550 22020 81750
rect 22090 81550 22410 81750
rect 22480 81550 22520 81750
rect 22590 81550 22910 81750
rect 22980 81550 23020 81750
rect 23090 81550 23410 81750
rect 23480 81550 23520 81750
rect 23590 81550 23910 81750
rect 23980 81550 24020 81750
rect 24090 81550 24410 81750
rect 24480 81550 24520 81750
rect 24590 81550 24910 81750
rect 24980 81550 25020 81750
rect 25090 81550 25410 81750
rect 25480 81550 25520 81750
rect 25590 81550 25910 81750
rect 25980 81550 26020 81750
rect 26090 81550 26410 81750
rect 26480 81550 26520 81750
rect 26590 81550 26910 81750
rect 26980 81550 27020 81750
rect 27090 81550 27410 81750
rect 27480 81550 27520 81750
rect 27590 81550 27910 81750
rect 27980 81550 28020 81750
rect 28090 81550 28410 81750
rect 28480 81550 28520 81750
rect 28590 81550 28910 81750
rect 28980 81550 29020 81750
rect 29090 81550 29410 81750
rect 29480 81550 29520 81750
rect 29590 81550 29910 81750
rect 29980 81550 30020 81750
rect 30090 81550 30410 81750
rect 30480 81550 30520 81750
rect 30590 81550 30910 81750
rect 30980 81550 31020 81750
rect 31090 81550 31410 81750
rect 31480 81550 31520 81750
rect 31590 81550 31910 81750
rect 31980 81550 32020 81750
rect 32090 81550 32410 81750
rect 32480 81550 32520 81750
rect 32590 81550 32910 81750
rect 32980 81550 33020 81750
rect 33090 81550 33410 81750
rect 33480 81550 33520 81750
rect 33590 81550 33910 81750
rect 33980 81550 34020 81750
rect 34090 81550 34410 81750
rect 34480 81550 34520 81750
rect 34590 81550 34910 81750
rect 34980 81550 35020 81750
rect 35090 81550 35410 81750
rect 35480 81550 35520 81750
rect 35590 81550 35910 81750
rect 35980 81550 36020 81750
rect 36090 81550 36410 81750
rect 36480 81550 36520 81750
rect 36590 81550 36910 81750
rect 36980 81550 37020 81750
rect 37090 81550 37410 81750
rect 37480 81550 37520 81750
rect 37590 81550 37910 81750
rect 37980 81550 38020 81750
rect 38090 81550 38410 81750
rect 38480 81550 38520 81750
rect 38590 81550 38910 81750
rect 38980 81550 39020 81750
rect 39090 81550 39410 81750
rect 39480 81550 39520 81750
rect 39590 81550 39910 81750
rect 39980 81550 40020 81750
rect 40090 81550 40410 81750
rect 40480 81550 40520 81750
rect 40590 81550 40910 81750
rect 40980 81550 41020 81750
rect 41090 81550 41410 81750
rect 41480 81550 41520 81750
rect 41590 81550 41910 81750
rect 41980 81550 42020 81750
rect 42090 81550 42410 81750
rect 42480 81550 42520 81750
rect 42590 81550 42910 81750
rect 42980 81550 43020 81750
rect 43090 81550 43410 81750
rect 43480 81550 43520 81750
rect 43590 81550 43910 81750
rect 43980 81550 44020 81750
rect 44090 81550 44410 81750
rect 44480 81550 44520 81750
rect 44590 81550 44910 81750
rect 44980 81550 45020 81750
rect 45090 81550 45410 81750
rect 45480 81550 45520 81750
rect 45590 81550 45910 81750
rect 45980 81550 46020 81750
rect 46090 81550 46410 81750
rect 46480 81550 46520 81750
rect 46590 81550 46910 81750
rect 46980 81550 47020 81750
rect 47090 81550 47410 81750
rect 47480 81550 47520 81750
rect 47590 81550 47910 81750
rect 47980 81550 48020 81750
rect 48090 81550 48410 81750
rect 48480 81550 48520 81750
rect 48590 81550 48910 81750
rect 48980 81550 49020 81750
rect 49090 81550 49410 81750
rect 49480 81550 49520 81750
rect 49590 81550 49910 81750
rect 49980 81550 50020 81750
rect 50090 81550 50410 81750
rect 50480 81550 50520 81750
rect 50590 81550 50910 81750
rect 50980 81550 51020 81750
rect 51090 81550 51410 81750
rect 51480 81550 51520 81750
rect 51590 81550 51910 81750
rect 51980 81550 52020 81750
rect 52090 81550 52410 81750
rect 52480 81550 52520 81750
rect 52590 81550 52910 81750
rect 52980 81550 53020 81750
rect 53090 81550 53410 81750
rect 53480 81550 53520 81750
rect 53590 81550 53910 81750
rect 53980 81550 54020 81750
rect 54090 81550 54410 81750
rect 54480 81550 54520 81750
rect 54590 81550 54910 81750
rect 54980 81550 55020 81750
rect 55090 81550 55410 81750
rect 55480 81550 55520 81750
rect 55590 81550 55910 81750
rect 55980 81550 56020 81750
rect 56090 81550 56410 81750
rect 56480 81550 56520 81750
rect 56590 81550 56910 81750
rect 56980 81550 57020 81750
rect 57090 81550 57410 81750
rect 57480 81550 57520 81750
rect 57590 81550 57910 81750
rect 57980 81550 58020 81750
rect 58090 81550 58410 81750
rect 58480 81550 58520 81750
rect 58590 81550 58910 81750
rect 58980 81550 59020 81750
rect 59090 81550 59410 81750
rect 59480 81550 59520 81750
rect 59590 81550 59910 81750
rect 59980 81550 60020 81750
rect 60090 81550 60410 81750
rect 60480 81550 60520 81750
rect 60590 81550 60910 81750
rect 60980 81550 61020 81750
rect 61090 81550 61410 81750
rect 61480 81550 61520 81750
rect 61590 81550 61910 81750
rect 61980 81550 62020 81750
rect 62090 81550 62410 81750
rect 62480 81550 62520 81750
rect 62590 81550 62910 81750
rect 62980 81550 63020 81750
rect 63090 81550 63410 81750
rect 63480 81550 63520 81750
rect 63590 81550 63910 81750
rect 63980 81550 64020 81750
rect 64090 81550 64410 81750
rect 64480 81550 64520 81750
rect 64590 81550 64910 81750
rect 64980 81550 65020 81750
rect 65090 81550 65410 81750
rect 65480 81550 65520 81750
rect 65590 81550 65910 81750
rect 65980 81550 66020 81750
rect 66090 81550 66410 81750
rect 66480 81550 66520 81750
rect 66590 81550 66910 81750
rect 66980 81550 67020 81750
rect 67090 81550 67410 81750
rect 67480 81550 67520 81750
rect 67590 81550 67910 81750
rect 67980 81550 68020 81750
rect 68090 81550 68410 81750
rect 68480 81550 68520 81750
rect 68590 81550 68910 81750
rect 68980 81550 69020 81750
rect 69090 81550 69410 81750
rect 69480 81550 69520 81750
rect 69590 81550 69910 81750
rect 69980 81550 70020 81750
rect 70090 81550 70410 81750
rect 70480 81550 70520 81750
rect 70590 81550 70910 81750
rect 70980 81550 71020 81750
rect 71090 81550 71410 81750
rect 71480 81550 71520 81750
rect 71590 81550 71910 81750
rect 71980 81550 72020 81750
rect 72090 81550 72410 81750
rect 72480 81550 72520 81750
rect 72590 81550 72910 81750
rect 72980 81550 73020 81750
rect 73090 81550 73410 81750
rect 73480 81550 73520 81750
rect 73590 81550 73910 81750
rect 73980 81550 74020 81750
rect 74090 81550 74410 81750
rect 74480 81550 74520 81750
rect 74590 81550 74910 81750
rect 74980 81550 75020 81750
rect 75090 81550 75410 81750
rect 75480 81550 75520 81750
rect 75590 81550 75910 81750
rect 75980 81550 76020 81750
rect 76090 81550 76410 81750
rect 76480 81550 76520 81750
rect 76590 81550 76910 81750
rect 76980 81550 77020 81750
rect 77090 81550 77410 81750
rect 77480 81550 77520 81750
rect 77590 81550 77910 81750
rect 77980 81550 78020 81750
rect 78090 81550 78410 81750
rect 78480 81550 78520 81750
rect 78590 81550 78910 81750
rect 78980 81550 79020 81750
rect 79090 81550 79410 81750
rect 79480 81550 79520 81750
rect 79590 81550 79910 81750
rect 79980 81550 80020 81750
rect 80090 81550 80410 81750
rect 80480 81550 80520 81750
rect 80590 81550 80910 81750
rect 80980 81550 81020 81750
rect 81090 81550 81410 81750
rect 81480 81550 81520 81750
rect 81590 81550 81910 81750
rect 81980 81550 82020 81750
rect 82090 81550 82410 81750
rect 82480 81550 82520 81750
rect 82590 81550 82910 81750
rect 82980 81550 83020 81750
rect 83090 81550 83410 81750
rect 83480 81550 83520 81750
rect 83590 81550 83910 81750
rect 83980 81550 84020 81750
rect 84090 81550 84410 81750
rect 84480 81550 84520 81750
rect 84590 81550 84910 81750
rect 84980 81550 85020 81750
rect 85090 81550 85410 81750
rect 85480 81550 85520 81750
rect 85590 81550 85910 81750
rect 85980 81550 86020 81750
rect 86090 81550 86410 81750
rect 86480 81550 86520 81750
rect 86590 81550 86910 81750
rect 86980 81550 87020 81750
rect 87090 81550 87410 81750
rect 87480 81550 87520 81750
rect 87590 81550 87910 81750
rect 87980 81550 88020 81750
rect 88090 81550 88410 81750
rect 88480 81550 88520 81750
rect 88590 81550 88910 81750
rect 88980 81550 89020 81750
rect 89090 81550 89410 81750
rect 89480 81550 89520 81750
rect 89590 81550 89910 81750
rect 89980 81550 90020 81750
rect 90090 81550 90410 81750
rect 90480 81550 90520 81750
rect 90590 81550 90910 81750
rect 90980 81550 91020 81750
rect 91090 81550 91410 81750
rect 91480 81550 91520 81750
rect 91590 81550 91910 81750
rect 91980 81550 92020 81750
rect 92090 81550 92410 81750
rect 92480 81550 92520 81750
rect 92590 81550 92910 81750
rect 92980 81550 93020 81750
rect 93090 81550 93410 81750
rect 93480 81550 93520 81750
rect 93590 81550 93910 81750
rect 93980 81550 94020 81750
rect 94090 81550 94410 81750
rect 94480 81550 94520 81750
rect 94590 81550 94910 81750
rect 94980 81550 95020 81750
rect 95090 81550 95410 81750
rect 95480 81550 95520 81750
rect 95590 81550 95910 81750
rect 95980 81550 96020 81750
rect 96090 81550 96410 81750
rect 96480 81550 96520 81750
rect 96590 81550 96910 81750
rect 96980 81550 97020 81750
rect 97090 81550 97410 81750
rect 97480 81550 97520 81750
rect 97590 81550 97910 81750
rect 97980 81550 98020 81750
rect 98090 81550 98410 81750
rect 98480 81550 98520 81750
rect 98590 81550 98910 81750
rect 98980 81550 99020 81750
rect 99090 81550 99410 81750
rect 99480 81550 99520 81750
rect 99590 81550 99910 81750
rect 99980 81550 100020 81750
rect 100090 81550 100410 81750
rect 100480 81550 100500 81750
rect -83500 81540 100500 81550
rect -83360 81490 -83140 81540
rect -83360 81420 -83350 81490
rect -83150 81420 -83140 81490
rect -83360 81380 -83140 81420
rect -83360 81310 -83350 81380
rect -83150 81310 -83140 81380
rect -83360 81260 -83140 81310
rect -82860 81490 -82640 81540
rect -82860 81420 -82850 81490
rect -82650 81420 -82640 81490
rect -82860 81380 -82640 81420
rect -82860 81310 -82850 81380
rect -82650 81310 -82640 81380
rect -82860 81260 -82640 81310
rect -82360 81490 -82140 81540
rect -82360 81420 -82350 81490
rect -82150 81420 -82140 81490
rect -82360 81380 -82140 81420
rect -82360 81310 -82350 81380
rect -82150 81310 -82140 81380
rect -82360 81260 -82140 81310
rect -81860 81490 -81640 81540
rect -81860 81420 -81850 81490
rect -81650 81420 -81640 81490
rect -81860 81380 -81640 81420
rect -81860 81310 -81850 81380
rect -81650 81310 -81640 81380
rect -81860 81260 -81640 81310
rect -81360 81490 -81140 81540
rect -81360 81420 -81350 81490
rect -81150 81420 -81140 81490
rect -81360 81380 -81140 81420
rect -81360 81310 -81350 81380
rect -81150 81310 -81140 81380
rect -81360 81260 -81140 81310
rect -80860 81490 -80640 81540
rect -80860 81420 -80850 81490
rect -80650 81420 -80640 81490
rect -80860 81380 -80640 81420
rect -80860 81310 -80850 81380
rect -80650 81310 -80640 81380
rect -80860 81260 -80640 81310
rect -80360 81490 -80140 81540
rect -80360 81420 -80350 81490
rect -80150 81420 -80140 81490
rect -80360 81380 -80140 81420
rect -80360 81310 -80350 81380
rect -80150 81310 -80140 81380
rect -80360 81260 -80140 81310
rect -79860 81490 -79640 81540
rect -79860 81420 -79850 81490
rect -79650 81420 -79640 81490
rect -79860 81380 -79640 81420
rect -79860 81310 -79850 81380
rect -79650 81310 -79640 81380
rect -79860 81260 -79640 81310
rect -79360 81490 -79140 81540
rect -79360 81420 -79350 81490
rect -79150 81420 -79140 81490
rect -79360 81380 -79140 81420
rect -79360 81310 -79350 81380
rect -79150 81310 -79140 81380
rect -79360 81260 -79140 81310
rect -78860 81490 -78640 81540
rect -78860 81420 -78850 81490
rect -78650 81420 -78640 81490
rect -78860 81380 -78640 81420
rect -78860 81310 -78850 81380
rect -78650 81310 -78640 81380
rect -78860 81260 -78640 81310
rect -78360 81490 -78140 81540
rect -78360 81420 -78350 81490
rect -78150 81420 -78140 81490
rect -78360 81380 -78140 81420
rect -78360 81310 -78350 81380
rect -78150 81310 -78140 81380
rect -78360 81260 -78140 81310
rect -77860 81490 -77640 81540
rect -77860 81420 -77850 81490
rect -77650 81420 -77640 81490
rect -77860 81380 -77640 81420
rect -77860 81310 -77850 81380
rect -77650 81310 -77640 81380
rect -77860 81260 -77640 81310
rect -77360 81490 -77140 81540
rect -77360 81420 -77350 81490
rect -77150 81420 -77140 81490
rect -77360 81380 -77140 81420
rect -77360 81310 -77350 81380
rect -77150 81310 -77140 81380
rect -77360 81260 -77140 81310
rect -76860 81490 -76640 81540
rect -76860 81420 -76850 81490
rect -76650 81420 -76640 81490
rect -76860 81380 -76640 81420
rect -76860 81310 -76850 81380
rect -76650 81310 -76640 81380
rect -76860 81260 -76640 81310
rect -76360 81490 -76140 81540
rect -76360 81420 -76350 81490
rect -76150 81420 -76140 81490
rect -76360 81380 -76140 81420
rect -76360 81310 -76350 81380
rect -76150 81310 -76140 81380
rect -76360 81260 -76140 81310
rect -75860 81490 -75640 81540
rect -75860 81420 -75850 81490
rect -75650 81420 -75640 81490
rect -75860 81380 -75640 81420
rect -75860 81310 -75850 81380
rect -75650 81310 -75640 81380
rect -75860 81260 -75640 81310
rect -75360 81490 -75140 81540
rect -75360 81420 -75350 81490
rect -75150 81420 -75140 81490
rect -75360 81380 -75140 81420
rect -75360 81310 -75350 81380
rect -75150 81310 -75140 81380
rect -75360 81260 -75140 81310
rect -74860 81490 -74640 81540
rect -74860 81420 -74850 81490
rect -74650 81420 -74640 81490
rect -74860 81380 -74640 81420
rect -74860 81310 -74850 81380
rect -74650 81310 -74640 81380
rect -74860 81260 -74640 81310
rect -74360 81490 -74140 81540
rect -74360 81420 -74350 81490
rect -74150 81420 -74140 81490
rect -74360 81380 -74140 81420
rect -74360 81310 -74350 81380
rect -74150 81310 -74140 81380
rect -74360 81260 -74140 81310
rect -73860 81490 -73640 81540
rect -73860 81420 -73850 81490
rect -73650 81420 -73640 81490
rect -73860 81380 -73640 81420
rect -73860 81310 -73850 81380
rect -73650 81310 -73640 81380
rect -73860 81260 -73640 81310
rect -73360 81490 -73140 81540
rect -73360 81420 -73350 81490
rect -73150 81420 -73140 81490
rect -73360 81380 -73140 81420
rect -73360 81310 -73350 81380
rect -73150 81310 -73140 81380
rect -73360 81260 -73140 81310
rect -72860 81490 -72640 81540
rect -72860 81420 -72850 81490
rect -72650 81420 -72640 81490
rect -72860 81380 -72640 81420
rect -72860 81310 -72850 81380
rect -72650 81310 -72640 81380
rect -72860 81260 -72640 81310
rect -72360 81490 -72140 81540
rect -72360 81420 -72350 81490
rect -72150 81420 -72140 81490
rect -72360 81380 -72140 81420
rect -72360 81310 -72350 81380
rect -72150 81310 -72140 81380
rect -72360 81260 -72140 81310
rect -71860 81490 -71640 81540
rect -71860 81420 -71850 81490
rect -71650 81420 -71640 81490
rect -71860 81380 -71640 81420
rect -71860 81310 -71850 81380
rect -71650 81310 -71640 81380
rect -71860 81260 -71640 81310
rect -71360 81490 -71140 81540
rect -71360 81420 -71350 81490
rect -71150 81420 -71140 81490
rect -71360 81380 -71140 81420
rect -71360 81310 -71350 81380
rect -71150 81310 -71140 81380
rect -71360 81260 -71140 81310
rect -70860 81490 -70640 81540
rect -70860 81420 -70850 81490
rect -70650 81420 -70640 81490
rect -70860 81380 -70640 81420
rect -70860 81310 -70850 81380
rect -70650 81310 -70640 81380
rect -70860 81260 -70640 81310
rect -70360 81490 -70140 81540
rect -70360 81420 -70350 81490
rect -70150 81420 -70140 81490
rect -70360 81380 -70140 81420
rect -70360 81310 -70350 81380
rect -70150 81310 -70140 81380
rect -70360 81260 -70140 81310
rect -69860 81490 -69640 81540
rect -69860 81420 -69850 81490
rect -69650 81420 -69640 81490
rect -69860 81380 -69640 81420
rect -69860 81310 -69850 81380
rect -69650 81310 -69640 81380
rect -69860 81260 -69640 81310
rect -69360 81490 -69140 81540
rect -69360 81420 -69350 81490
rect -69150 81420 -69140 81490
rect -69360 81380 -69140 81420
rect -69360 81310 -69350 81380
rect -69150 81310 -69140 81380
rect -69360 81260 -69140 81310
rect -68860 81490 -68640 81540
rect -68860 81420 -68850 81490
rect -68650 81420 -68640 81490
rect -68860 81380 -68640 81420
rect -68860 81310 -68850 81380
rect -68650 81310 -68640 81380
rect -68860 81260 -68640 81310
rect -68360 81490 -68140 81540
rect -68360 81420 -68350 81490
rect -68150 81420 -68140 81490
rect -68360 81380 -68140 81420
rect -68360 81310 -68350 81380
rect -68150 81310 -68140 81380
rect -68360 81260 -68140 81310
rect -67860 81490 -67640 81540
rect -67860 81420 -67850 81490
rect -67650 81420 -67640 81490
rect -67860 81380 -67640 81420
rect -67860 81310 -67850 81380
rect -67650 81310 -67640 81380
rect -67860 81260 -67640 81310
rect -67360 81490 -67140 81540
rect -67360 81420 -67350 81490
rect -67150 81420 -67140 81490
rect -67360 81380 -67140 81420
rect -67360 81310 -67350 81380
rect -67150 81310 -67140 81380
rect -67360 81260 -67140 81310
rect -66860 81490 -66640 81540
rect -66860 81420 -66850 81490
rect -66650 81420 -66640 81490
rect -66860 81380 -66640 81420
rect -66860 81310 -66850 81380
rect -66650 81310 -66640 81380
rect -66860 81260 -66640 81310
rect -66360 81490 -66140 81540
rect -66360 81420 -66350 81490
rect -66150 81420 -66140 81490
rect -66360 81380 -66140 81420
rect -66360 81310 -66350 81380
rect -66150 81310 -66140 81380
rect -66360 81260 -66140 81310
rect -65860 81490 -65640 81540
rect -65860 81420 -65850 81490
rect -65650 81420 -65640 81490
rect -65860 81380 -65640 81420
rect -65860 81310 -65850 81380
rect -65650 81310 -65640 81380
rect -65860 81260 -65640 81310
rect -65360 81490 -65140 81540
rect -65360 81420 -65350 81490
rect -65150 81420 -65140 81490
rect -65360 81380 -65140 81420
rect -65360 81310 -65350 81380
rect -65150 81310 -65140 81380
rect -65360 81260 -65140 81310
rect -64860 81490 -64640 81540
rect -64860 81420 -64850 81490
rect -64650 81420 -64640 81490
rect -64860 81380 -64640 81420
rect -64860 81310 -64850 81380
rect -64650 81310 -64640 81380
rect -64860 81260 -64640 81310
rect -64360 81490 -64140 81540
rect -64360 81420 -64350 81490
rect -64150 81420 -64140 81490
rect -64360 81380 -64140 81420
rect -64360 81310 -64350 81380
rect -64150 81310 -64140 81380
rect -64360 81260 -64140 81310
rect -63860 81490 -63640 81540
rect -63860 81420 -63850 81490
rect -63650 81420 -63640 81490
rect -63860 81380 -63640 81420
rect -63860 81310 -63850 81380
rect -63650 81310 -63640 81380
rect -63860 81260 -63640 81310
rect -63360 81490 -63140 81540
rect -63360 81420 -63350 81490
rect -63150 81420 -63140 81490
rect -63360 81380 -63140 81420
rect -63360 81310 -63350 81380
rect -63150 81310 -63140 81380
rect -63360 81260 -63140 81310
rect -62860 81490 -62640 81540
rect -62860 81420 -62850 81490
rect -62650 81420 -62640 81490
rect -62860 81380 -62640 81420
rect -62860 81310 -62850 81380
rect -62650 81310 -62640 81380
rect -62860 81260 -62640 81310
rect -62360 81490 -62140 81540
rect -62360 81420 -62350 81490
rect -62150 81420 -62140 81490
rect -62360 81380 -62140 81420
rect -62360 81310 -62350 81380
rect -62150 81310 -62140 81380
rect -62360 81260 -62140 81310
rect -61860 81490 -61640 81540
rect -61860 81420 -61850 81490
rect -61650 81420 -61640 81490
rect -61860 81380 -61640 81420
rect -61860 81310 -61850 81380
rect -61650 81310 -61640 81380
rect -61860 81260 -61640 81310
rect -61360 81490 -61140 81540
rect -61360 81420 -61350 81490
rect -61150 81420 -61140 81490
rect -61360 81380 -61140 81420
rect -61360 81310 -61350 81380
rect -61150 81310 -61140 81380
rect -61360 81260 -61140 81310
rect -60860 81490 -60640 81540
rect -60860 81420 -60850 81490
rect -60650 81420 -60640 81490
rect -60860 81380 -60640 81420
rect -60860 81310 -60850 81380
rect -60650 81310 -60640 81380
rect -60860 81260 -60640 81310
rect -60360 81490 -60140 81540
rect -60360 81420 -60350 81490
rect -60150 81420 -60140 81490
rect -60360 81380 -60140 81420
rect -60360 81310 -60350 81380
rect -60150 81310 -60140 81380
rect -60360 81260 -60140 81310
rect -59860 81490 -59640 81540
rect -59860 81420 -59850 81490
rect -59650 81420 -59640 81490
rect -59860 81380 -59640 81420
rect -59860 81310 -59850 81380
rect -59650 81310 -59640 81380
rect -59860 81260 -59640 81310
rect -59360 81490 -59140 81540
rect -59360 81420 -59350 81490
rect -59150 81420 -59140 81490
rect -59360 81380 -59140 81420
rect -59360 81310 -59350 81380
rect -59150 81310 -59140 81380
rect -59360 81260 -59140 81310
rect -58860 81490 -58640 81540
rect -58860 81420 -58850 81490
rect -58650 81420 -58640 81490
rect -58860 81380 -58640 81420
rect -58860 81310 -58850 81380
rect -58650 81310 -58640 81380
rect -58860 81260 -58640 81310
rect -58360 81490 -58140 81540
rect -58360 81420 -58350 81490
rect -58150 81420 -58140 81490
rect -58360 81380 -58140 81420
rect -58360 81310 -58350 81380
rect -58150 81310 -58140 81380
rect -58360 81260 -58140 81310
rect -57860 81490 -57640 81540
rect -57860 81420 -57850 81490
rect -57650 81420 -57640 81490
rect -57860 81380 -57640 81420
rect -57860 81310 -57850 81380
rect -57650 81310 -57640 81380
rect -57860 81260 -57640 81310
rect -57360 81490 -57140 81540
rect -57360 81420 -57350 81490
rect -57150 81420 -57140 81490
rect -57360 81380 -57140 81420
rect -57360 81310 -57350 81380
rect -57150 81310 -57140 81380
rect -57360 81260 -57140 81310
rect -56860 81490 -56640 81540
rect -56860 81420 -56850 81490
rect -56650 81420 -56640 81490
rect -56860 81380 -56640 81420
rect -56860 81310 -56850 81380
rect -56650 81310 -56640 81380
rect -56860 81260 -56640 81310
rect -56360 81490 -56140 81540
rect -56360 81420 -56350 81490
rect -56150 81420 -56140 81490
rect -56360 81380 -56140 81420
rect -56360 81310 -56350 81380
rect -56150 81310 -56140 81380
rect -56360 81260 -56140 81310
rect -55860 81490 -55640 81540
rect -55860 81420 -55850 81490
rect -55650 81420 -55640 81490
rect -55860 81380 -55640 81420
rect -55860 81310 -55850 81380
rect -55650 81310 -55640 81380
rect -55860 81260 -55640 81310
rect -55360 81490 -55140 81540
rect -55360 81420 -55350 81490
rect -55150 81420 -55140 81490
rect -55360 81380 -55140 81420
rect -55360 81310 -55350 81380
rect -55150 81310 -55140 81380
rect -55360 81260 -55140 81310
rect -54860 81490 -54640 81540
rect -54860 81420 -54850 81490
rect -54650 81420 -54640 81490
rect -54860 81380 -54640 81420
rect -54860 81310 -54850 81380
rect -54650 81310 -54640 81380
rect -54860 81260 -54640 81310
rect -54360 81490 -54140 81540
rect -54360 81420 -54350 81490
rect -54150 81420 -54140 81490
rect -54360 81380 -54140 81420
rect -54360 81310 -54350 81380
rect -54150 81310 -54140 81380
rect -54360 81260 -54140 81310
rect -53860 81490 -53640 81540
rect -53860 81420 -53850 81490
rect -53650 81420 -53640 81490
rect -53860 81380 -53640 81420
rect -53860 81310 -53850 81380
rect -53650 81310 -53640 81380
rect -53860 81260 -53640 81310
rect -53360 81490 -53140 81540
rect -53360 81420 -53350 81490
rect -53150 81420 -53140 81490
rect -53360 81380 -53140 81420
rect -53360 81310 -53350 81380
rect -53150 81310 -53140 81380
rect -53360 81260 -53140 81310
rect -52860 81490 -52640 81540
rect -52860 81420 -52850 81490
rect -52650 81420 -52640 81490
rect -52860 81380 -52640 81420
rect -52860 81310 -52850 81380
rect -52650 81310 -52640 81380
rect -52860 81260 -52640 81310
rect -52360 81490 -52140 81540
rect -52360 81420 -52350 81490
rect -52150 81420 -52140 81490
rect -52360 81380 -52140 81420
rect -52360 81310 -52350 81380
rect -52150 81310 -52140 81380
rect -52360 81260 -52140 81310
rect -51860 81490 -51640 81540
rect -51860 81420 -51850 81490
rect -51650 81420 -51640 81490
rect -51860 81380 -51640 81420
rect -51860 81310 -51850 81380
rect -51650 81310 -51640 81380
rect -51860 81260 -51640 81310
rect -51360 81490 -51140 81540
rect -51360 81420 -51350 81490
rect -51150 81420 -51140 81490
rect -51360 81380 -51140 81420
rect -51360 81310 -51350 81380
rect -51150 81310 -51140 81380
rect -51360 81260 -51140 81310
rect -50860 81490 -50640 81540
rect -50860 81420 -50850 81490
rect -50650 81420 -50640 81490
rect -50860 81380 -50640 81420
rect -50860 81310 -50850 81380
rect -50650 81310 -50640 81380
rect -50860 81260 -50640 81310
rect -50360 81490 -50140 81540
rect -50360 81420 -50350 81490
rect -50150 81420 -50140 81490
rect -50360 81380 -50140 81420
rect -50360 81310 -50350 81380
rect -50150 81310 -50140 81380
rect -50360 81260 -50140 81310
rect -49860 81490 -49640 81540
rect -49860 81420 -49850 81490
rect -49650 81420 -49640 81490
rect -49860 81380 -49640 81420
rect -49860 81310 -49850 81380
rect -49650 81310 -49640 81380
rect -49860 81260 -49640 81310
rect -49360 81490 -49140 81540
rect -49360 81420 -49350 81490
rect -49150 81420 -49140 81490
rect -49360 81380 -49140 81420
rect -49360 81310 -49350 81380
rect -49150 81310 -49140 81380
rect -49360 81260 -49140 81310
rect -48860 81490 -48640 81540
rect -48860 81420 -48850 81490
rect -48650 81420 -48640 81490
rect -48860 81380 -48640 81420
rect -48860 81310 -48850 81380
rect -48650 81310 -48640 81380
rect -48860 81260 -48640 81310
rect -48360 81490 -48140 81540
rect -48360 81420 -48350 81490
rect -48150 81420 -48140 81490
rect -48360 81380 -48140 81420
rect -48360 81310 -48350 81380
rect -48150 81310 -48140 81380
rect -48360 81260 -48140 81310
rect -47860 81490 -47640 81540
rect -47860 81420 -47850 81490
rect -47650 81420 -47640 81490
rect -47860 81380 -47640 81420
rect -47860 81310 -47850 81380
rect -47650 81310 -47640 81380
rect -47860 81260 -47640 81310
rect -47360 81490 -47140 81540
rect -47360 81420 -47350 81490
rect -47150 81420 -47140 81490
rect -47360 81380 -47140 81420
rect -47360 81310 -47350 81380
rect -47150 81310 -47140 81380
rect -47360 81260 -47140 81310
rect -46860 81490 -46640 81540
rect -46860 81420 -46850 81490
rect -46650 81420 -46640 81490
rect -46860 81380 -46640 81420
rect -46860 81310 -46850 81380
rect -46650 81310 -46640 81380
rect -46860 81260 -46640 81310
rect -46360 81490 -46140 81540
rect -46360 81420 -46350 81490
rect -46150 81420 -46140 81490
rect -46360 81380 -46140 81420
rect -46360 81310 -46350 81380
rect -46150 81310 -46140 81380
rect -46360 81260 -46140 81310
rect -45860 81490 -45640 81540
rect -45860 81420 -45850 81490
rect -45650 81420 -45640 81490
rect -45860 81380 -45640 81420
rect -45860 81310 -45850 81380
rect -45650 81310 -45640 81380
rect -45860 81260 -45640 81310
rect -45360 81490 -45140 81540
rect -45360 81420 -45350 81490
rect -45150 81420 -45140 81490
rect -45360 81380 -45140 81420
rect -45360 81310 -45350 81380
rect -45150 81310 -45140 81380
rect -45360 81260 -45140 81310
rect -44860 81490 -44640 81540
rect -44860 81420 -44850 81490
rect -44650 81420 -44640 81490
rect -44860 81380 -44640 81420
rect -44860 81310 -44850 81380
rect -44650 81310 -44640 81380
rect -44860 81260 -44640 81310
rect -44360 81490 -44140 81540
rect -44360 81420 -44350 81490
rect -44150 81420 -44140 81490
rect -44360 81380 -44140 81420
rect -44360 81310 -44350 81380
rect -44150 81310 -44140 81380
rect -44360 81260 -44140 81310
rect -43860 81490 -43640 81540
rect -43860 81420 -43850 81490
rect -43650 81420 -43640 81490
rect -43860 81380 -43640 81420
rect -43860 81310 -43850 81380
rect -43650 81310 -43640 81380
rect -43860 81260 -43640 81310
rect -43360 81490 -43140 81540
rect -43360 81420 -43350 81490
rect -43150 81420 -43140 81490
rect -43360 81380 -43140 81420
rect -43360 81310 -43350 81380
rect -43150 81310 -43140 81380
rect -43360 81260 -43140 81310
rect -42860 81490 -42640 81540
rect -42860 81420 -42850 81490
rect -42650 81420 -42640 81490
rect -42860 81380 -42640 81420
rect -42860 81310 -42850 81380
rect -42650 81310 -42640 81380
rect -42860 81260 -42640 81310
rect -42360 81490 -42140 81540
rect -42360 81420 -42350 81490
rect -42150 81420 -42140 81490
rect -42360 81380 -42140 81420
rect -42360 81310 -42350 81380
rect -42150 81310 -42140 81380
rect -42360 81260 -42140 81310
rect -41860 81490 -41640 81540
rect -41860 81420 -41850 81490
rect -41650 81420 -41640 81490
rect -41860 81380 -41640 81420
rect -41860 81310 -41850 81380
rect -41650 81310 -41640 81380
rect -41860 81260 -41640 81310
rect -41360 81490 -41140 81540
rect -41360 81420 -41350 81490
rect -41150 81420 -41140 81490
rect -41360 81380 -41140 81420
rect -41360 81310 -41350 81380
rect -41150 81310 -41140 81380
rect -41360 81260 -41140 81310
rect -40860 81490 -40640 81540
rect -40860 81420 -40850 81490
rect -40650 81420 -40640 81490
rect -40860 81380 -40640 81420
rect -40860 81310 -40850 81380
rect -40650 81310 -40640 81380
rect -40860 81260 -40640 81310
rect -40360 81490 -40140 81540
rect -40360 81420 -40350 81490
rect -40150 81420 -40140 81490
rect -40360 81380 -40140 81420
rect -40360 81310 -40350 81380
rect -40150 81310 -40140 81380
rect -40360 81260 -40140 81310
rect -39860 81490 -39640 81540
rect -39860 81420 -39850 81490
rect -39650 81420 -39640 81490
rect -39860 81380 -39640 81420
rect -39860 81310 -39850 81380
rect -39650 81310 -39640 81380
rect -39860 81260 -39640 81310
rect -39360 81490 -39140 81540
rect -39360 81420 -39350 81490
rect -39150 81420 -39140 81490
rect -39360 81380 -39140 81420
rect -39360 81310 -39350 81380
rect -39150 81310 -39140 81380
rect -39360 81260 -39140 81310
rect -38860 81490 -38640 81540
rect -38860 81420 -38850 81490
rect -38650 81420 -38640 81490
rect -38860 81380 -38640 81420
rect -38860 81310 -38850 81380
rect -38650 81310 -38640 81380
rect -38860 81260 -38640 81310
rect -38360 81490 -38140 81540
rect -38360 81420 -38350 81490
rect -38150 81420 -38140 81490
rect -38360 81380 -38140 81420
rect -38360 81310 -38350 81380
rect -38150 81310 -38140 81380
rect -38360 81260 -38140 81310
rect -37860 81490 -37640 81540
rect -37860 81420 -37850 81490
rect -37650 81420 -37640 81490
rect -37860 81380 -37640 81420
rect -37860 81310 -37850 81380
rect -37650 81310 -37640 81380
rect -37860 81260 -37640 81310
rect -37360 81490 -37140 81540
rect -37360 81420 -37350 81490
rect -37150 81420 -37140 81490
rect -37360 81380 -37140 81420
rect -37360 81310 -37350 81380
rect -37150 81310 -37140 81380
rect -37360 81260 -37140 81310
rect -36860 81490 -36640 81540
rect -36860 81420 -36850 81490
rect -36650 81420 -36640 81490
rect -36860 81380 -36640 81420
rect -36860 81310 -36850 81380
rect -36650 81310 -36640 81380
rect -36860 81260 -36640 81310
rect -36360 81490 -36140 81540
rect -36360 81420 -36350 81490
rect -36150 81420 -36140 81490
rect -36360 81380 -36140 81420
rect -36360 81310 -36350 81380
rect -36150 81310 -36140 81380
rect -36360 81260 -36140 81310
rect -35860 81490 -35640 81540
rect -35860 81420 -35850 81490
rect -35650 81420 -35640 81490
rect -35860 81380 -35640 81420
rect -35860 81310 -35850 81380
rect -35650 81310 -35640 81380
rect -35860 81260 -35640 81310
rect -35360 81490 -35140 81540
rect -35360 81420 -35350 81490
rect -35150 81420 -35140 81490
rect -35360 81380 -35140 81420
rect -35360 81310 -35350 81380
rect -35150 81310 -35140 81380
rect -35360 81260 -35140 81310
rect -34860 81490 -34640 81540
rect -34860 81420 -34850 81490
rect -34650 81420 -34640 81490
rect -34860 81380 -34640 81420
rect -34860 81310 -34850 81380
rect -34650 81310 -34640 81380
rect -34860 81260 -34640 81310
rect -34360 81490 -34140 81540
rect -34360 81420 -34350 81490
rect -34150 81420 -34140 81490
rect -34360 81380 -34140 81420
rect -34360 81310 -34350 81380
rect -34150 81310 -34140 81380
rect -34360 81260 -34140 81310
rect -33860 81490 -33640 81540
rect -33860 81420 -33850 81490
rect -33650 81420 -33640 81490
rect -33860 81380 -33640 81420
rect -33860 81310 -33850 81380
rect -33650 81310 -33640 81380
rect -33860 81260 -33640 81310
rect -33360 81490 -33140 81540
rect -33360 81420 -33350 81490
rect -33150 81420 -33140 81490
rect -33360 81380 -33140 81420
rect -33360 81310 -33350 81380
rect -33150 81310 -33140 81380
rect -33360 81260 -33140 81310
rect -32860 81490 -32640 81540
rect -32860 81420 -32850 81490
rect -32650 81420 -32640 81490
rect -32860 81380 -32640 81420
rect -32860 81310 -32850 81380
rect -32650 81310 -32640 81380
rect -32860 81260 -32640 81310
rect -32360 81490 -32140 81540
rect -32360 81420 -32350 81490
rect -32150 81420 -32140 81490
rect -32360 81380 -32140 81420
rect -32360 81310 -32350 81380
rect -32150 81310 -32140 81380
rect -32360 81260 -32140 81310
rect -31860 81490 -31640 81540
rect -31860 81420 -31850 81490
rect -31650 81420 -31640 81490
rect -31860 81380 -31640 81420
rect -31860 81310 -31850 81380
rect -31650 81310 -31640 81380
rect -31860 81260 -31640 81310
rect -31360 81490 -31140 81540
rect -31360 81420 -31350 81490
rect -31150 81420 -31140 81490
rect -31360 81380 -31140 81420
rect -31360 81310 -31350 81380
rect -31150 81310 -31140 81380
rect -31360 81260 -31140 81310
rect -30860 81490 -30640 81540
rect -30860 81420 -30850 81490
rect -30650 81420 -30640 81490
rect -30860 81380 -30640 81420
rect -30860 81310 -30850 81380
rect -30650 81310 -30640 81380
rect -30860 81260 -30640 81310
rect -30360 81490 -30140 81540
rect -30360 81420 -30350 81490
rect -30150 81420 -30140 81490
rect -30360 81380 -30140 81420
rect -30360 81310 -30350 81380
rect -30150 81310 -30140 81380
rect -30360 81260 -30140 81310
rect -29860 81490 -29640 81540
rect -29860 81420 -29850 81490
rect -29650 81420 -29640 81490
rect -29860 81380 -29640 81420
rect -29860 81310 -29850 81380
rect -29650 81310 -29640 81380
rect -29860 81260 -29640 81310
rect -29360 81490 -29140 81540
rect -29360 81420 -29350 81490
rect -29150 81420 -29140 81490
rect -29360 81380 -29140 81420
rect -29360 81310 -29350 81380
rect -29150 81310 -29140 81380
rect -29360 81260 -29140 81310
rect -28860 81490 -28640 81540
rect -28860 81420 -28850 81490
rect -28650 81420 -28640 81490
rect -28860 81380 -28640 81420
rect -28860 81310 -28850 81380
rect -28650 81310 -28640 81380
rect -28860 81260 -28640 81310
rect -28360 81490 -28140 81540
rect -28360 81420 -28350 81490
rect -28150 81420 -28140 81490
rect -28360 81380 -28140 81420
rect -28360 81310 -28350 81380
rect -28150 81310 -28140 81380
rect -28360 81260 -28140 81310
rect -27860 81490 -27640 81540
rect -27860 81420 -27850 81490
rect -27650 81420 -27640 81490
rect -27860 81380 -27640 81420
rect -27860 81310 -27850 81380
rect -27650 81310 -27640 81380
rect -27860 81260 -27640 81310
rect -27360 81490 -27140 81540
rect -27360 81420 -27350 81490
rect -27150 81420 -27140 81490
rect -27360 81380 -27140 81420
rect -27360 81310 -27350 81380
rect -27150 81310 -27140 81380
rect -27360 81260 -27140 81310
rect -26860 81490 -26640 81540
rect -26860 81420 -26850 81490
rect -26650 81420 -26640 81490
rect -26860 81380 -26640 81420
rect -26860 81310 -26850 81380
rect -26650 81310 -26640 81380
rect -26860 81260 -26640 81310
rect -26360 81490 -26140 81540
rect -26360 81420 -26350 81490
rect -26150 81420 -26140 81490
rect -26360 81380 -26140 81420
rect -26360 81310 -26350 81380
rect -26150 81310 -26140 81380
rect -26360 81260 -26140 81310
rect -25860 81490 -25640 81540
rect -25860 81420 -25850 81490
rect -25650 81420 -25640 81490
rect -25860 81380 -25640 81420
rect -25860 81310 -25850 81380
rect -25650 81310 -25640 81380
rect -25860 81260 -25640 81310
rect -25360 81490 -25140 81540
rect -25360 81420 -25350 81490
rect -25150 81420 -25140 81490
rect -25360 81380 -25140 81420
rect -25360 81310 -25350 81380
rect -25150 81310 -25140 81380
rect -25360 81260 -25140 81310
rect -24860 81490 -24640 81540
rect -24860 81420 -24850 81490
rect -24650 81420 -24640 81490
rect -24860 81380 -24640 81420
rect -24860 81310 -24850 81380
rect -24650 81310 -24640 81380
rect -24860 81260 -24640 81310
rect -24360 81490 -24140 81540
rect -24360 81420 -24350 81490
rect -24150 81420 -24140 81490
rect -24360 81380 -24140 81420
rect -24360 81310 -24350 81380
rect -24150 81310 -24140 81380
rect -24360 81260 -24140 81310
rect -23860 81490 -23640 81540
rect -23860 81420 -23850 81490
rect -23650 81420 -23640 81490
rect -23860 81380 -23640 81420
rect -23860 81310 -23850 81380
rect -23650 81310 -23640 81380
rect -23860 81260 -23640 81310
rect -23360 81490 -23140 81540
rect -23360 81420 -23350 81490
rect -23150 81420 -23140 81490
rect -23360 81380 -23140 81420
rect -23360 81310 -23350 81380
rect -23150 81310 -23140 81380
rect -23360 81260 -23140 81310
rect -22860 81490 -22640 81540
rect -22860 81420 -22850 81490
rect -22650 81420 -22640 81490
rect -22860 81380 -22640 81420
rect -22860 81310 -22850 81380
rect -22650 81310 -22640 81380
rect -22860 81260 -22640 81310
rect -22360 81490 -22140 81540
rect -22360 81420 -22350 81490
rect -22150 81420 -22140 81490
rect -22360 81380 -22140 81420
rect -22360 81310 -22350 81380
rect -22150 81310 -22140 81380
rect -22360 81260 -22140 81310
rect -21860 81490 -21640 81540
rect -21860 81420 -21850 81490
rect -21650 81420 -21640 81490
rect -21860 81380 -21640 81420
rect -21860 81310 -21850 81380
rect -21650 81310 -21640 81380
rect -21860 81260 -21640 81310
rect -21360 81490 -21140 81540
rect -21360 81420 -21350 81490
rect -21150 81420 -21140 81490
rect -21360 81380 -21140 81420
rect -21360 81310 -21350 81380
rect -21150 81310 -21140 81380
rect -21360 81260 -21140 81310
rect -20860 81490 -20640 81540
rect -20860 81420 -20850 81490
rect -20650 81420 -20640 81490
rect -20860 81380 -20640 81420
rect -20860 81310 -20850 81380
rect -20650 81310 -20640 81380
rect -20860 81260 -20640 81310
rect -20360 81490 -20140 81540
rect -20360 81420 -20350 81490
rect -20150 81420 -20140 81490
rect -20360 81380 -20140 81420
rect -20360 81310 -20350 81380
rect -20150 81310 -20140 81380
rect -20360 81260 -20140 81310
rect -19860 81490 -19640 81540
rect -19860 81420 -19850 81490
rect -19650 81420 -19640 81490
rect -19860 81380 -19640 81420
rect -19860 81310 -19850 81380
rect -19650 81310 -19640 81380
rect -19860 81260 -19640 81310
rect -19360 81490 -19140 81540
rect -19360 81420 -19350 81490
rect -19150 81420 -19140 81490
rect -19360 81380 -19140 81420
rect -19360 81310 -19350 81380
rect -19150 81310 -19140 81380
rect -19360 81260 -19140 81310
rect -18860 81490 -18640 81540
rect -18860 81420 -18850 81490
rect -18650 81420 -18640 81490
rect -18860 81380 -18640 81420
rect -18860 81310 -18850 81380
rect -18650 81310 -18640 81380
rect -18860 81260 -18640 81310
rect -18360 81490 -18140 81540
rect -18360 81420 -18350 81490
rect -18150 81420 -18140 81490
rect -18360 81380 -18140 81420
rect -18360 81310 -18350 81380
rect -18150 81310 -18140 81380
rect -18360 81260 -18140 81310
rect -17860 81490 -17640 81540
rect -17860 81420 -17850 81490
rect -17650 81420 -17640 81490
rect -17860 81380 -17640 81420
rect -17860 81310 -17850 81380
rect -17650 81310 -17640 81380
rect -17860 81260 -17640 81310
rect -17360 81490 -17140 81540
rect -17360 81420 -17350 81490
rect -17150 81420 -17140 81490
rect -17360 81380 -17140 81420
rect -17360 81310 -17350 81380
rect -17150 81310 -17140 81380
rect -17360 81260 -17140 81310
rect -16860 81490 -16640 81540
rect -16860 81420 -16850 81490
rect -16650 81420 -16640 81490
rect -16860 81380 -16640 81420
rect -16860 81310 -16850 81380
rect -16650 81310 -16640 81380
rect -16860 81260 -16640 81310
rect -16360 81490 -16140 81540
rect -16360 81420 -16350 81490
rect -16150 81420 -16140 81490
rect -16360 81380 -16140 81420
rect -16360 81310 -16350 81380
rect -16150 81310 -16140 81380
rect -16360 81260 -16140 81310
rect -15860 81490 -15640 81540
rect -15860 81420 -15850 81490
rect -15650 81420 -15640 81490
rect -15860 81380 -15640 81420
rect -15860 81310 -15850 81380
rect -15650 81310 -15640 81380
rect -15860 81260 -15640 81310
rect -15360 81490 -15140 81540
rect -15360 81420 -15350 81490
rect -15150 81420 -15140 81490
rect -15360 81380 -15140 81420
rect -15360 81310 -15350 81380
rect -15150 81310 -15140 81380
rect -15360 81260 -15140 81310
rect -14860 81490 -14640 81540
rect -14860 81420 -14850 81490
rect -14650 81420 -14640 81490
rect -14860 81380 -14640 81420
rect -14860 81310 -14850 81380
rect -14650 81310 -14640 81380
rect -14860 81260 -14640 81310
rect -14360 81490 -14140 81540
rect -14360 81420 -14350 81490
rect -14150 81420 -14140 81490
rect -14360 81380 -14140 81420
rect -14360 81310 -14350 81380
rect -14150 81310 -14140 81380
rect -14360 81260 -14140 81310
rect -13860 81490 -13640 81540
rect -13860 81420 -13850 81490
rect -13650 81420 -13640 81490
rect -13860 81380 -13640 81420
rect -13860 81310 -13850 81380
rect -13650 81310 -13640 81380
rect -13860 81260 -13640 81310
rect -13360 81490 -13140 81540
rect -13360 81420 -13350 81490
rect -13150 81420 -13140 81490
rect -13360 81380 -13140 81420
rect -13360 81310 -13350 81380
rect -13150 81310 -13140 81380
rect -13360 81260 -13140 81310
rect -12860 81490 -12640 81540
rect -12860 81420 -12850 81490
rect -12650 81420 -12640 81490
rect -12860 81380 -12640 81420
rect -12860 81310 -12850 81380
rect -12650 81310 -12640 81380
rect -12860 81260 -12640 81310
rect -12360 81490 -12140 81540
rect -12360 81420 -12350 81490
rect -12150 81420 -12140 81490
rect -12360 81380 -12140 81420
rect -12360 81310 -12350 81380
rect -12150 81310 -12140 81380
rect -12360 81260 -12140 81310
rect -11860 81490 -11640 81540
rect -11860 81420 -11850 81490
rect -11650 81420 -11640 81490
rect -11860 81380 -11640 81420
rect -11860 81310 -11850 81380
rect -11650 81310 -11640 81380
rect -11860 81260 -11640 81310
rect -11360 81490 -11140 81540
rect -11360 81420 -11350 81490
rect -11150 81420 -11140 81490
rect -11360 81380 -11140 81420
rect -11360 81310 -11350 81380
rect -11150 81310 -11140 81380
rect -11360 81260 -11140 81310
rect -10860 81490 -10640 81540
rect -10860 81420 -10850 81490
rect -10650 81420 -10640 81490
rect -10860 81380 -10640 81420
rect -10860 81310 -10850 81380
rect -10650 81310 -10640 81380
rect -10860 81260 -10640 81310
rect -10360 81490 -10140 81540
rect -10360 81420 -10350 81490
rect -10150 81420 -10140 81490
rect -10360 81380 -10140 81420
rect -10360 81310 -10350 81380
rect -10150 81310 -10140 81380
rect -10360 81260 -10140 81310
rect -9860 81490 -9640 81540
rect -9860 81420 -9850 81490
rect -9650 81420 -9640 81490
rect -9860 81380 -9640 81420
rect -9860 81310 -9850 81380
rect -9650 81310 -9640 81380
rect -9860 81260 -9640 81310
rect -9360 81490 -9140 81540
rect -9360 81420 -9350 81490
rect -9150 81420 -9140 81490
rect -9360 81380 -9140 81420
rect -9360 81310 -9350 81380
rect -9150 81310 -9140 81380
rect -9360 81260 -9140 81310
rect -8860 81490 -8640 81540
rect -8860 81420 -8850 81490
rect -8650 81420 -8640 81490
rect -8860 81380 -8640 81420
rect -8860 81310 -8850 81380
rect -8650 81310 -8640 81380
rect -8860 81260 -8640 81310
rect -8360 81490 -8140 81540
rect -8360 81420 -8350 81490
rect -8150 81420 -8140 81490
rect -8360 81380 -8140 81420
rect -8360 81310 -8350 81380
rect -8150 81310 -8140 81380
rect -8360 81260 -8140 81310
rect -7860 81490 -7640 81540
rect -7860 81420 -7850 81490
rect -7650 81420 -7640 81490
rect -7860 81380 -7640 81420
rect -7860 81310 -7850 81380
rect -7650 81310 -7640 81380
rect -7860 81260 -7640 81310
rect -7360 81490 -7140 81540
rect -7360 81420 -7350 81490
rect -7150 81420 -7140 81490
rect -7360 81380 -7140 81420
rect -7360 81310 -7350 81380
rect -7150 81310 -7140 81380
rect -7360 81260 -7140 81310
rect -6860 81490 -6640 81540
rect -6860 81420 -6850 81490
rect -6650 81420 -6640 81490
rect -6860 81380 -6640 81420
rect -6860 81310 -6850 81380
rect -6650 81310 -6640 81380
rect -6860 81260 -6640 81310
rect -6360 81490 -6140 81540
rect -6360 81420 -6350 81490
rect -6150 81420 -6140 81490
rect -6360 81380 -6140 81420
rect -6360 81310 -6350 81380
rect -6150 81310 -6140 81380
rect -6360 81260 -6140 81310
rect -5860 81490 -5640 81540
rect -5860 81420 -5850 81490
rect -5650 81420 -5640 81490
rect -5860 81380 -5640 81420
rect -5860 81310 -5850 81380
rect -5650 81310 -5640 81380
rect -5860 81260 -5640 81310
rect -5360 81490 -5140 81540
rect -5360 81420 -5350 81490
rect -5150 81420 -5140 81490
rect -5360 81380 -5140 81420
rect -5360 81310 -5350 81380
rect -5150 81310 -5140 81380
rect -5360 81260 -5140 81310
rect -4860 81490 -4640 81540
rect -4860 81420 -4850 81490
rect -4650 81420 -4640 81490
rect -4860 81380 -4640 81420
rect -4860 81310 -4850 81380
rect -4650 81310 -4640 81380
rect -4860 81260 -4640 81310
rect -4360 81490 -4140 81540
rect -4360 81420 -4350 81490
rect -4150 81420 -4140 81490
rect -4360 81380 -4140 81420
rect -4360 81310 -4350 81380
rect -4150 81310 -4140 81380
rect -4360 81260 -4140 81310
rect -3860 81490 -3640 81540
rect -3860 81420 -3850 81490
rect -3650 81420 -3640 81490
rect -3860 81380 -3640 81420
rect -3860 81310 -3850 81380
rect -3650 81310 -3640 81380
rect -3860 81260 -3640 81310
rect -3360 81490 -3140 81540
rect -3360 81420 -3350 81490
rect -3150 81420 -3140 81490
rect -3360 81380 -3140 81420
rect -3360 81310 -3350 81380
rect -3150 81310 -3140 81380
rect -3360 81260 -3140 81310
rect -2860 81490 -2640 81540
rect -2860 81420 -2850 81490
rect -2650 81420 -2640 81490
rect -2860 81380 -2640 81420
rect -2860 81310 -2850 81380
rect -2650 81310 -2640 81380
rect -2860 81260 -2640 81310
rect -2360 81490 -2140 81540
rect -2360 81420 -2350 81490
rect -2150 81420 -2140 81490
rect -2360 81380 -2140 81420
rect -2360 81310 -2350 81380
rect -2150 81310 -2140 81380
rect -2360 81260 -2140 81310
rect -1860 81490 -1640 81540
rect -1860 81420 -1850 81490
rect -1650 81420 -1640 81490
rect -1860 81380 -1640 81420
rect -1860 81310 -1850 81380
rect -1650 81310 -1640 81380
rect -1860 81260 -1640 81310
rect -1360 81490 -1140 81540
rect -1360 81420 -1350 81490
rect -1150 81420 -1140 81490
rect -1360 81380 -1140 81420
rect -1360 81310 -1350 81380
rect -1150 81310 -1140 81380
rect -1360 81260 -1140 81310
rect -860 81490 -640 81540
rect -860 81420 -850 81490
rect -650 81420 -640 81490
rect -860 81380 -640 81420
rect -860 81310 -850 81380
rect -650 81310 -640 81380
rect -860 81260 -640 81310
rect -360 81490 -140 81540
rect -360 81420 -350 81490
rect -150 81420 -140 81490
rect -360 81380 -140 81420
rect -360 81310 -350 81380
rect -150 81310 -140 81380
rect -360 81260 -140 81310
rect 140 81490 360 81540
rect 140 81420 150 81490
rect 350 81420 360 81490
rect 140 81380 360 81420
rect 140 81310 150 81380
rect 350 81310 360 81380
rect 140 81260 360 81310
rect 640 81490 860 81540
rect 640 81420 650 81490
rect 850 81420 860 81490
rect 640 81380 860 81420
rect 640 81310 650 81380
rect 850 81310 860 81380
rect 640 81260 860 81310
rect 1140 81490 1360 81540
rect 1140 81420 1150 81490
rect 1350 81420 1360 81490
rect 1140 81380 1360 81420
rect 1140 81310 1150 81380
rect 1350 81310 1360 81380
rect 1140 81260 1360 81310
rect 1640 81490 1860 81540
rect 1640 81420 1650 81490
rect 1850 81420 1860 81490
rect 1640 81380 1860 81420
rect 1640 81310 1650 81380
rect 1850 81310 1860 81380
rect 1640 81260 1860 81310
rect 2140 81490 2360 81540
rect 2140 81420 2150 81490
rect 2350 81420 2360 81490
rect 2140 81380 2360 81420
rect 2140 81310 2150 81380
rect 2350 81310 2360 81380
rect 2140 81260 2360 81310
rect 2640 81490 2860 81540
rect 2640 81420 2650 81490
rect 2850 81420 2860 81490
rect 2640 81380 2860 81420
rect 2640 81310 2650 81380
rect 2850 81310 2860 81380
rect 2640 81260 2860 81310
rect 3140 81490 3360 81540
rect 3140 81420 3150 81490
rect 3350 81420 3360 81490
rect 3140 81380 3360 81420
rect 3140 81310 3150 81380
rect 3350 81310 3360 81380
rect 3140 81260 3360 81310
rect 3640 81490 3860 81540
rect 3640 81420 3650 81490
rect 3850 81420 3860 81490
rect 3640 81380 3860 81420
rect 3640 81310 3650 81380
rect 3850 81310 3860 81380
rect 3640 81260 3860 81310
rect 4140 81490 4360 81540
rect 4140 81420 4150 81490
rect 4350 81420 4360 81490
rect 4140 81380 4360 81420
rect 4140 81310 4150 81380
rect 4350 81310 4360 81380
rect 4140 81260 4360 81310
rect 4640 81490 4860 81540
rect 4640 81420 4650 81490
rect 4850 81420 4860 81490
rect 4640 81380 4860 81420
rect 4640 81310 4650 81380
rect 4850 81310 4860 81380
rect 4640 81260 4860 81310
rect 5140 81490 5360 81540
rect 5140 81420 5150 81490
rect 5350 81420 5360 81490
rect 5140 81380 5360 81420
rect 5140 81310 5150 81380
rect 5350 81310 5360 81380
rect 5140 81260 5360 81310
rect 5640 81490 5860 81540
rect 5640 81420 5650 81490
rect 5850 81420 5860 81490
rect 5640 81380 5860 81420
rect 5640 81310 5650 81380
rect 5850 81310 5860 81380
rect 5640 81260 5860 81310
rect 6140 81490 6360 81540
rect 6140 81420 6150 81490
rect 6350 81420 6360 81490
rect 6140 81380 6360 81420
rect 6140 81310 6150 81380
rect 6350 81310 6360 81380
rect 6140 81260 6360 81310
rect 6640 81490 6860 81540
rect 6640 81420 6650 81490
rect 6850 81420 6860 81490
rect 6640 81380 6860 81420
rect 6640 81310 6650 81380
rect 6850 81310 6860 81380
rect 6640 81260 6860 81310
rect 7140 81490 7360 81540
rect 7140 81420 7150 81490
rect 7350 81420 7360 81490
rect 7140 81380 7360 81420
rect 7140 81310 7150 81380
rect 7350 81310 7360 81380
rect 7140 81260 7360 81310
rect 7640 81490 7860 81540
rect 7640 81420 7650 81490
rect 7850 81420 7860 81490
rect 7640 81380 7860 81420
rect 7640 81310 7650 81380
rect 7850 81310 7860 81380
rect 7640 81260 7860 81310
rect 8140 81490 8360 81540
rect 8140 81420 8150 81490
rect 8350 81420 8360 81490
rect 8140 81380 8360 81420
rect 8140 81310 8150 81380
rect 8350 81310 8360 81380
rect 8140 81260 8360 81310
rect 8640 81490 8860 81540
rect 8640 81420 8650 81490
rect 8850 81420 8860 81490
rect 8640 81380 8860 81420
rect 8640 81310 8650 81380
rect 8850 81310 8860 81380
rect 8640 81260 8860 81310
rect 9140 81490 9360 81540
rect 9140 81420 9150 81490
rect 9350 81420 9360 81490
rect 9140 81380 9360 81420
rect 9140 81310 9150 81380
rect 9350 81310 9360 81380
rect 9140 81260 9360 81310
rect 9640 81490 9860 81540
rect 9640 81420 9650 81490
rect 9850 81420 9860 81490
rect 9640 81380 9860 81420
rect 9640 81310 9650 81380
rect 9850 81310 9860 81380
rect 9640 81260 9860 81310
rect 10140 81490 10360 81540
rect 10140 81420 10150 81490
rect 10350 81420 10360 81490
rect 10140 81380 10360 81420
rect 10140 81310 10150 81380
rect 10350 81310 10360 81380
rect 10140 81260 10360 81310
rect 10640 81490 10860 81540
rect 10640 81420 10650 81490
rect 10850 81420 10860 81490
rect 10640 81380 10860 81420
rect 10640 81310 10650 81380
rect 10850 81310 10860 81380
rect 10640 81260 10860 81310
rect 11140 81490 11360 81540
rect 11140 81420 11150 81490
rect 11350 81420 11360 81490
rect 11140 81380 11360 81420
rect 11140 81310 11150 81380
rect 11350 81310 11360 81380
rect 11140 81260 11360 81310
rect 11640 81490 11860 81540
rect 11640 81420 11650 81490
rect 11850 81420 11860 81490
rect 11640 81380 11860 81420
rect 11640 81310 11650 81380
rect 11850 81310 11860 81380
rect 11640 81260 11860 81310
rect 12140 81490 12360 81540
rect 12140 81420 12150 81490
rect 12350 81420 12360 81490
rect 12140 81380 12360 81420
rect 12140 81310 12150 81380
rect 12350 81310 12360 81380
rect 12140 81260 12360 81310
rect 12640 81490 12860 81540
rect 12640 81420 12650 81490
rect 12850 81420 12860 81490
rect 12640 81380 12860 81420
rect 12640 81310 12650 81380
rect 12850 81310 12860 81380
rect 12640 81260 12860 81310
rect 13140 81490 13360 81540
rect 13140 81420 13150 81490
rect 13350 81420 13360 81490
rect 13140 81380 13360 81420
rect 13140 81310 13150 81380
rect 13350 81310 13360 81380
rect 13140 81260 13360 81310
rect 13640 81490 13860 81540
rect 13640 81420 13650 81490
rect 13850 81420 13860 81490
rect 13640 81380 13860 81420
rect 13640 81310 13650 81380
rect 13850 81310 13860 81380
rect 13640 81260 13860 81310
rect 14140 81490 14360 81540
rect 14140 81420 14150 81490
rect 14350 81420 14360 81490
rect 14140 81380 14360 81420
rect 14140 81310 14150 81380
rect 14350 81310 14360 81380
rect 14140 81260 14360 81310
rect 14640 81490 14860 81540
rect 14640 81420 14650 81490
rect 14850 81420 14860 81490
rect 14640 81380 14860 81420
rect 14640 81310 14650 81380
rect 14850 81310 14860 81380
rect 14640 81260 14860 81310
rect 15140 81490 15360 81540
rect 15140 81420 15150 81490
rect 15350 81420 15360 81490
rect 15140 81380 15360 81420
rect 15140 81310 15150 81380
rect 15350 81310 15360 81380
rect 15140 81260 15360 81310
rect 15640 81490 15860 81540
rect 15640 81420 15650 81490
rect 15850 81420 15860 81490
rect 15640 81380 15860 81420
rect 15640 81310 15650 81380
rect 15850 81310 15860 81380
rect 15640 81260 15860 81310
rect 16140 81490 16360 81540
rect 16140 81420 16150 81490
rect 16350 81420 16360 81490
rect 16140 81380 16360 81420
rect 16140 81310 16150 81380
rect 16350 81310 16360 81380
rect 16140 81260 16360 81310
rect 16640 81490 16860 81540
rect 16640 81420 16650 81490
rect 16850 81420 16860 81490
rect 16640 81380 16860 81420
rect 16640 81310 16650 81380
rect 16850 81310 16860 81380
rect 16640 81260 16860 81310
rect 17140 81490 17360 81540
rect 17140 81420 17150 81490
rect 17350 81420 17360 81490
rect 17140 81380 17360 81420
rect 17140 81310 17150 81380
rect 17350 81310 17360 81380
rect 17140 81260 17360 81310
rect 17640 81490 17860 81540
rect 17640 81420 17650 81490
rect 17850 81420 17860 81490
rect 17640 81380 17860 81420
rect 17640 81310 17650 81380
rect 17850 81310 17860 81380
rect 17640 81260 17860 81310
rect 18140 81490 18360 81540
rect 18140 81420 18150 81490
rect 18350 81420 18360 81490
rect 18140 81380 18360 81420
rect 18140 81310 18150 81380
rect 18350 81310 18360 81380
rect 18140 81260 18360 81310
rect 18640 81490 18860 81540
rect 18640 81420 18650 81490
rect 18850 81420 18860 81490
rect 18640 81380 18860 81420
rect 18640 81310 18650 81380
rect 18850 81310 18860 81380
rect 18640 81260 18860 81310
rect 19140 81490 19360 81540
rect 19140 81420 19150 81490
rect 19350 81420 19360 81490
rect 19140 81380 19360 81420
rect 19140 81310 19150 81380
rect 19350 81310 19360 81380
rect 19140 81260 19360 81310
rect 19640 81490 19860 81540
rect 19640 81420 19650 81490
rect 19850 81420 19860 81490
rect 19640 81380 19860 81420
rect 19640 81310 19650 81380
rect 19850 81310 19860 81380
rect 19640 81260 19860 81310
rect 20140 81490 20360 81540
rect 20140 81420 20150 81490
rect 20350 81420 20360 81490
rect 20140 81380 20360 81420
rect 20140 81310 20150 81380
rect 20350 81310 20360 81380
rect 20140 81260 20360 81310
rect 20640 81490 20860 81540
rect 20640 81420 20650 81490
rect 20850 81420 20860 81490
rect 20640 81380 20860 81420
rect 20640 81310 20650 81380
rect 20850 81310 20860 81380
rect 20640 81260 20860 81310
rect 21140 81490 21360 81540
rect 21140 81420 21150 81490
rect 21350 81420 21360 81490
rect 21140 81380 21360 81420
rect 21140 81310 21150 81380
rect 21350 81310 21360 81380
rect 21140 81260 21360 81310
rect 21640 81490 21860 81540
rect 21640 81420 21650 81490
rect 21850 81420 21860 81490
rect 21640 81380 21860 81420
rect 21640 81310 21650 81380
rect 21850 81310 21860 81380
rect 21640 81260 21860 81310
rect 22140 81490 22360 81540
rect 22140 81420 22150 81490
rect 22350 81420 22360 81490
rect 22140 81380 22360 81420
rect 22140 81310 22150 81380
rect 22350 81310 22360 81380
rect 22140 81260 22360 81310
rect 22640 81490 22860 81540
rect 22640 81420 22650 81490
rect 22850 81420 22860 81490
rect 22640 81380 22860 81420
rect 22640 81310 22650 81380
rect 22850 81310 22860 81380
rect 22640 81260 22860 81310
rect 23140 81490 23360 81540
rect 23140 81420 23150 81490
rect 23350 81420 23360 81490
rect 23140 81380 23360 81420
rect 23140 81310 23150 81380
rect 23350 81310 23360 81380
rect 23140 81260 23360 81310
rect 23640 81490 23860 81540
rect 23640 81420 23650 81490
rect 23850 81420 23860 81490
rect 23640 81380 23860 81420
rect 23640 81310 23650 81380
rect 23850 81310 23860 81380
rect 23640 81260 23860 81310
rect 24140 81490 24360 81540
rect 24140 81420 24150 81490
rect 24350 81420 24360 81490
rect 24140 81380 24360 81420
rect 24140 81310 24150 81380
rect 24350 81310 24360 81380
rect 24140 81260 24360 81310
rect 24640 81490 24860 81540
rect 24640 81420 24650 81490
rect 24850 81420 24860 81490
rect 24640 81380 24860 81420
rect 24640 81310 24650 81380
rect 24850 81310 24860 81380
rect 24640 81260 24860 81310
rect 25140 81490 25360 81540
rect 25140 81420 25150 81490
rect 25350 81420 25360 81490
rect 25140 81380 25360 81420
rect 25140 81310 25150 81380
rect 25350 81310 25360 81380
rect 25140 81260 25360 81310
rect 25640 81490 25860 81540
rect 25640 81420 25650 81490
rect 25850 81420 25860 81490
rect 25640 81380 25860 81420
rect 25640 81310 25650 81380
rect 25850 81310 25860 81380
rect 25640 81260 25860 81310
rect 26140 81490 26360 81540
rect 26140 81420 26150 81490
rect 26350 81420 26360 81490
rect 26140 81380 26360 81420
rect 26140 81310 26150 81380
rect 26350 81310 26360 81380
rect 26140 81260 26360 81310
rect 26640 81490 26860 81540
rect 26640 81420 26650 81490
rect 26850 81420 26860 81490
rect 26640 81380 26860 81420
rect 26640 81310 26650 81380
rect 26850 81310 26860 81380
rect 26640 81260 26860 81310
rect 27140 81490 27360 81540
rect 27140 81420 27150 81490
rect 27350 81420 27360 81490
rect 27140 81380 27360 81420
rect 27140 81310 27150 81380
rect 27350 81310 27360 81380
rect 27140 81260 27360 81310
rect 27640 81490 27860 81540
rect 27640 81420 27650 81490
rect 27850 81420 27860 81490
rect 27640 81380 27860 81420
rect 27640 81310 27650 81380
rect 27850 81310 27860 81380
rect 27640 81260 27860 81310
rect 28140 81490 28360 81540
rect 28140 81420 28150 81490
rect 28350 81420 28360 81490
rect 28140 81380 28360 81420
rect 28140 81310 28150 81380
rect 28350 81310 28360 81380
rect 28140 81260 28360 81310
rect 28640 81490 28860 81540
rect 28640 81420 28650 81490
rect 28850 81420 28860 81490
rect 28640 81380 28860 81420
rect 28640 81310 28650 81380
rect 28850 81310 28860 81380
rect 28640 81260 28860 81310
rect 29140 81490 29360 81540
rect 29140 81420 29150 81490
rect 29350 81420 29360 81490
rect 29140 81380 29360 81420
rect 29140 81310 29150 81380
rect 29350 81310 29360 81380
rect 29140 81260 29360 81310
rect 29640 81490 29860 81540
rect 29640 81420 29650 81490
rect 29850 81420 29860 81490
rect 29640 81380 29860 81420
rect 29640 81310 29650 81380
rect 29850 81310 29860 81380
rect 29640 81260 29860 81310
rect 30140 81490 30360 81540
rect 30140 81420 30150 81490
rect 30350 81420 30360 81490
rect 30140 81380 30360 81420
rect 30140 81310 30150 81380
rect 30350 81310 30360 81380
rect 30140 81260 30360 81310
rect 30640 81490 30860 81540
rect 30640 81420 30650 81490
rect 30850 81420 30860 81490
rect 30640 81380 30860 81420
rect 30640 81310 30650 81380
rect 30850 81310 30860 81380
rect 30640 81260 30860 81310
rect 31140 81490 31360 81540
rect 31140 81420 31150 81490
rect 31350 81420 31360 81490
rect 31140 81380 31360 81420
rect 31140 81310 31150 81380
rect 31350 81310 31360 81380
rect 31140 81260 31360 81310
rect 31640 81490 31860 81540
rect 31640 81420 31650 81490
rect 31850 81420 31860 81490
rect 31640 81380 31860 81420
rect 31640 81310 31650 81380
rect 31850 81310 31860 81380
rect 31640 81260 31860 81310
rect 32140 81490 32360 81540
rect 32140 81420 32150 81490
rect 32350 81420 32360 81490
rect 32140 81380 32360 81420
rect 32140 81310 32150 81380
rect 32350 81310 32360 81380
rect 32140 81260 32360 81310
rect 32640 81490 32860 81540
rect 32640 81420 32650 81490
rect 32850 81420 32860 81490
rect 32640 81380 32860 81420
rect 32640 81310 32650 81380
rect 32850 81310 32860 81380
rect 32640 81260 32860 81310
rect 33140 81490 33360 81540
rect 33140 81420 33150 81490
rect 33350 81420 33360 81490
rect 33140 81380 33360 81420
rect 33140 81310 33150 81380
rect 33350 81310 33360 81380
rect 33140 81260 33360 81310
rect 33640 81490 33860 81540
rect 33640 81420 33650 81490
rect 33850 81420 33860 81490
rect 33640 81380 33860 81420
rect 33640 81310 33650 81380
rect 33850 81310 33860 81380
rect 33640 81260 33860 81310
rect 34140 81490 34360 81540
rect 34140 81420 34150 81490
rect 34350 81420 34360 81490
rect 34140 81380 34360 81420
rect 34140 81310 34150 81380
rect 34350 81310 34360 81380
rect 34140 81260 34360 81310
rect 34640 81490 34860 81540
rect 34640 81420 34650 81490
rect 34850 81420 34860 81490
rect 34640 81380 34860 81420
rect 34640 81310 34650 81380
rect 34850 81310 34860 81380
rect 34640 81260 34860 81310
rect 35140 81490 35360 81540
rect 35140 81420 35150 81490
rect 35350 81420 35360 81490
rect 35140 81380 35360 81420
rect 35140 81310 35150 81380
rect 35350 81310 35360 81380
rect 35140 81260 35360 81310
rect 35640 81490 35860 81540
rect 35640 81420 35650 81490
rect 35850 81420 35860 81490
rect 35640 81380 35860 81420
rect 35640 81310 35650 81380
rect 35850 81310 35860 81380
rect 35640 81260 35860 81310
rect 36140 81490 36360 81540
rect 36140 81420 36150 81490
rect 36350 81420 36360 81490
rect 36140 81380 36360 81420
rect 36140 81310 36150 81380
rect 36350 81310 36360 81380
rect 36140 81260 36360 81310
rect 36640 81490 36860 81540
rect 36640 81420 36650 81490
rect 36850 81420 36860 81490
rect 36640 81380 36860 81420
rect 36640 81310 36650 81380
rect 36850 81310 36860 81380
rect 36640 81260 36860 81310
rect 37140 81490 37360 81540
rect 37140 81420 37150 81490
rect 37350 81420 37360 81490
rect 37140 81380 37360 81420
rect 37140 81310 37150 81380
rect 37350 81310 37360 81380
rect 37140 81260 37360 81310
rect 37640 81490 37860 81540
rect 37640 81420 37650 81490
rect 37850 81420 37860 81490
rect 37640 81380 37860 81420
rect 37640 81310 37650 81380
rect 37850 81310 37860 81380
rect 37640 81260 37860 81310
rect 38140 81490 38360 81540
rect 38140 81420 38150 81490
rect 38350 81420 38360 81490
rect 38140 81380 38360 81420
rect 38140 81310 38150 81380
rect 38350 81310 38360 81380
rect 38140 81260 38360 81310
rect 38640 81490 38860 81540
rect 38640 81420 38650 81490
rect 38850 81420 38860 81490
rect 38640 81380 38860 81420
rect 38640 81310 38650 81380
rect 38850 81310 38860 81380
rect 38640 81260 38860 81310
rect 39140 81490 39360 81540
rect 39140 81420 39150 81490
rect 39350 81420 39360 81490
rect 39140 81380 39360 81420
rect 39140 81310 39150 81380
rect 39350 81310 39360 81380
rect 39140 81260 39360 81310
rect 39640 81490 39860 81540
rect 39640 81420 39650 81490
rect 39850 81420 39860 81490
rect 39640 81380 39860 81420
rect 39640 81310 39650 81380
rect 39850 81310 39860 81380
rect 39640 81260 39860 81310
rect 40140 81490 40360 81540
rect 40140 81420 40150 81490
rect 40350 81420 40360 81490
rect 40140 81380 40360 81420
rect 40140 81310 40150 81380
rect 40350 81310 40360 81380
rect 40140 81260 40360 81310
rect 40640 81490 40860 81540
rect 40640 81420 40650 81490
rect 40850 81420 40860 81490
rect 40640 81380 40860 81420
rect 40640 81310 40650 81380
rect 40850 81310 40860 81380
rect 40640 81260 40860 81310
rect 41140 81490 41360 81540
rect 41140 81420 41150 81490
rect 41350 81420 41360 81490
rect 41140 81380 41360 81420
rect 41140 81310 41150 81380
rect 41350 81310 41360 81380
rect 41140 81260 41360 81310
rect 41640 81490 41860 81540
rect 41640 81420 41650 81490
rect 41850 81420 41860 81490
rect 41640 81380 41860 81420
rect 41640 81310 41650 81380
rect 41850 81310 41860 81380
rect 41640 81260 41860 81310
rect 42140 81490 42360 81540
rect 42140 81420 42150 81490
rect 42350 81420 42360 81490
rect 42140 81380 42360 81420
rect 42140 81310 42150 81380
rect 42350 81310 42360 81380
rect 42140 81260 42360 81310
rect 42640 81490 42860 81540
rect 42640 81420 42650 81490
rect 42850 81420 42860 81490
rect 42640 81380 42860 81420
rect 42640 81310 42650 81380
rect 42850 81310 42860 81380
rect 42640 81260 42860 81310
rect 43140 81490 43360 81540
rect 43140 81420 43150 81490
rect 43350 81420 43360 81490
rect 43140 81380 43360 81420
rect 43140 81310 43150 81380
rect 43350 81310 43360 81380
rect 43140 81260 43360 81310
rect 43640 81490 43860 81540
rect 43640 81420 43650 81490
rect 43850 81420 43860 81490
rect 43640 81380 43860 81420
rect 43640 81310 43650 81380
rect 43850 81310 43860 81380
rect 43640 81260 43860 81310
rect 44140 81490 44360 81540
rect 44140 81420 44150 81490
rect 44350 81420 44360 81490
rect 44140 81380 44360 81420
rect 44140 81310 44150 81380
rect 44350 81310 44360 81380
rect 44140 81260 44360 81310
rect 44640 81490 44860 81540
rect 44640 81420 44650 81490
rect 44850 81420 44860 81490
rect 44640 81380 44860 81420
rect 44640 81310 44650 81380
rect 44850 81310 44860 81380
rect 44640 81260 44860 81310
rect 45140 81490 45360 81540
rect 45140 81420 45150 81490
rect 45350 81420 45360 81490
rect 45140 81380 45360 81420
rect 45140 81310 45150 81380
rect 45350 81310 45360 81380
rect 45140 81260 45360 81310
rect 45640 81490 45860 81540
rect 45640 81420 45650 81490
rect 45850 81420 45860 81490
rect 45640 81380 45860 81420
rect 45640 81310 45650 81380
rect 45850 81310 45860 81380
rect 45640 81260 45860 81310
rect 46140 81490 46360 81540
rect 46140 81420 46150 81490
rect 46350 81420 46360 81490
rect 46140 81380 46360 81420
rect 46140 81310 46150 81380
rect 46350 81310 46360 81380
rect 46140 81260 46360 81310
rect 46640 81490 46860 81540
rect 46640 81420 46650 81490
rect 46850 81420 46860 81490
rect 46640 81380 46860 81420
rect 46640 81310 46650 81380
rect 46850 81310 46860 81380
rect 46640 81260 46860 81310
rect 47140 81490 47360 81540
rect 47140 81420 47150 81490
rect 47350 81420 47360 81490
rect 47140 81380 47360 81420
rect 47140 81310 47150 81380
rect 47350 81310 47360 81380
rect 47140 81260 47360 81310
rect 47640 81490 47860 81540
rect 47640 81420 47650 81490
rect 47850 81420 47860 81490
rect 47640 81380 47860 81420
rect 47640 81310 47650 81380
rect 47850 81310 47860 81380
rect 47640 81260 47860 81310
rect 48140 81490 48360 81540
rect 48140 81420 48150 81490
rect 48350 81420 48360 81490
rect 48140 81380 48360 81420
rect 48140 81310 48150 81380
rect 48350 81310 48360 81380
rect 48140 81260 48360 81310
rect 48640 81490 48860 81540
rect 48640 81420 48650 81490
rect 48850 81420 48860 81490
rect 48640 81380 48860 81420
rect 48640 81310 48650 81380
rect 48850 81310 48860 81380
rect 48640 81260 48860 81310
rect 49140 81490 49360 81540
rect 49140 81420 49150 81490
rect 49350 81420 49360 81490
rect 49140 81380 49360 81420
rect 49140 81310 49150 81380
rect 49350 81310 49360 81380
rect 49140 81260 49360 81310
rect 49640 81490 49860 81540
rect 49640 81420 49650 81490
rect 49850 81420 49860 81490
rect 49640 81380 49860 81420
rect 49640 81310 49650 81380
rect 49850 81310 49860 81380
rect 49640 81260 49860 81310
rect 50140 81490 50360 81540
rect 50140 81420 50150 81490
rect 50350 81420 50360 81490
rect 50140 81380 50360 81420
rect 50140 81310 50150 81380
rect 50350 81310 50360 81380
rect 50140 81260 50360 81310
rect 50640 81490 50860 81540
rect 50640 81420 50650 81490
rect 50850 81420 50860 81490
rect 50640 81380 50860 81420
rect 50640 81310 50650 81380
rect 50850 81310 50860 81380
rect 50640 81260 50860 81310
rect 51140 81490 51360 81540
rect 51140 81420 51150 81490
rect 51350 81420 51360 81490
rect 51140 81380 51360 81420
rect 51140 81310 51150 81380
rect 51350 81310 51360 81380
rect 51140 81260 51360 81310
rect 51640 81490 51860 81540
rect 51640 81420 51650 81490
rect 51850 81420 51860 81490
rect 51640 81380 51860 81420
rect 51640 81310 51650 81380
rect 51850 81310 51860 81380
rect 51640 81260 51860 81310
rect 52140 81490 52360 81540
rect 52140 81420 52150 81490
rect 52350 81420 52360 81490
rect 52140 81380 52360 81420
rect 52140 81310 52150 81380
rect 52350 81310 52360 81380
rect 52140 81260 52360 81310
rect 52640 81490 52860 81540
rect 52640 81420 52650 81490
rect 52850 81420 52860 81490
rect 52640 81380 52860 81420
rect 52640 81310 52650 81380
rect 52850 81310 52860 81380
rect 52640 81260 52860 81310
rect 53140 81490 53360 81540
rect 53140 81420 53150 81490
rect 53350 81420 53360 81490
rect 53140 81380 53360 81420
rect 53140 81310 53150 81380
rect 53350 81310 53360 81380
rect 53140 81260 53360 81310
rect 53640 81490 53860 81540
rect 53640 81420 53650 81490
rect 53850 81420 53860 81490
rect 53640 81380 53860 81420
rect 53640 81310 53650 81380
rect 53850 81310 53860 81380
rect 53640 81260 53860 81310
rect 54140 81490 54360 81540
rect 54140 81420 54150 81490
rect 54350 81420 54360 81490
rect 54140 81380 54360 81420
rect 54140 81310 54150 81380
rect 54350 81310 54360 81380
rect 54140 81260 54360 81310
rect 54640 81490 54860 81540
rect 54640 81420 54650 81490
rect 54850 81420 54860 81490
rect 54640 81380 54860 81420
rect 54640 81310 54650 81380
rect 54850 81310 54860 81380
rect 54640 81260 54860 81310
rect 55140 81490 55360 81540
rect 55140 81420 55150 81490
rect 55350 81420 55360 81490
rect 55140 81380 55360 81420
rect 55140 81310 55150 81380
rect 55350 81310 55360 81380
rect 55140 81260 55360 81310
rect 55640 81490 55860 81540
rect 55640 81420 55650 81490
rect 55850 81420 55860 81490
rect 55640 81380 55860 81420
rect 55640 81310 55650 81380
rect 55850 81310 55860 81380
rect 55640 81260 55860 81310
rect 56140 81490 56360 81540
rect 56140 81420 56150 81490
rect 56350 81420 56360 81490
rect 56140 81380 56360 81420
rect 56140 81310 56150 81380
rect 56350 81310 56360 81380
rect 56140 81260 56360 81310
rect 56640 81490 56860 81540
rect 56640 81420 56650 81490
rect 56850 81420 56860 81490
rect 56640 81380 56860 81420
rect 56640 81310 56650 81380
rect 56850 81310 56860 81380
rect 56640 81260 56860 81310
rect 57140 81490 57360 81540
rect 57140 81420 57150 81490
rect 57350 81420 57360 81490
rect 57140 81380 57360 81420
rect 57140 81310 57150 81380
rect 57350 81310 57360 81380
rect 57140 81260 57360 81310
rect 57640 81490 57860 81540
rect 57640 81420 57650 81490
rect 57850 81420 57860 81490
rect 57640 81380 57860 81420
rect 57640 81310 57650 81380
rect 57850 81310 57860 81380
rect 57640 81260 57860 81310
rect 58140 81490 58360 81540
rect 58140 81420 58150 81490
rect 58350 81420 58360 81490
rect 58140 81380 58360 81420
rect 58140 81310 58150 81380
rect 58350 81310 58360 81380
rect 58140 81260 58360 81310
rect 58640 81490 58860 81540
rect 58640 81420 58650 81490
rect 58850 81420 58860 81490
rect 58640 81380 58860 81420
rect 58640 81310 58650 81380
rect 58850 81310 58860 81380
rect 58640 81260 58860 81310
rect 59140 81490 59360 81540
rect 59140 81420 59150 81490
rect 59350 81420 59360 81490
rect 59140 81380 59360 81420
rect 59140 81310 59150 81380
rect 59350 81310 59360 81380
rect 59140 81260 59360 81310
rect 59640 81490 59860 81540
rect 59640 81420 59650 81490
rect 59850 81420 59860 81490
rect 59640 81380 59860 81420
rect 59640 81310 59650 81380
rect 59850 81310 59860 81380
rect 59640 81260 59860 81310
rect 60140 81490 60360 81540
rect 60140 81420 60150 81490
rect 60350 81420 60360 81490
rect 60140 81380 60360 81420
rect 60140 81310 60150 81380
rect 60350 81310 60360 81380
rect 60140 81260 60360 81310
rect 60640 81490 60860 81540
rect 60640 81420 60650 81490
rect 60850 81420 60860 81490
rect 60640 81380 60860 81420
rect 60640 81310 60650 81380
rect 60850 81310 60860 81380
rect 60640 81260 60860 81310
rect 61140 81490 61360 81540
rect 61140 81420 61150 81490
rect 61350 81420 61360 81490
rect 61140 81380 61360 81420
rect 61140 81310 61150 81380
rect 61350 81310 61360 81380
rect 61140 81260 61360 81310
rect 61640 81490 61860 81540
rect 61640 81420 61650 81490
rect 61850 81420 61860 81490
rect 61640 81380 61860 81420
rect 61640 81310 61650 81380
rect 61850 81310 61860 81380
rect 61640 81260 61860 81310
rect 62140 81490 62360 81540
rect 62140 81420 62150 81490
rect 62350 81420 62360 81490
rect 62140 81380 62360 81420
rect 62140 81310 62150 81380
rect 62350 81310 62360 81380
rect 62140 81260 62360 81310
rect 62640 81490 62860 81540
rect 62640 81420 62650 81490
rect 62850 81420 62860 81490
rect 62640 81380 62860 81420
rect 62640 81310 62650 81380
rect 62850 81310 62860 81380
rect 62640 81260 62860 81310
rect 63140 81490 63360 81540
rect 63140 81420 63150 81490
rect 63350 81420 63360 81490
rect 63140 81380 63360 81420
rect 63140 81310 63150 81380
rect 63350 81310 63360 81380
rect 63140 81260 63360 81310
rect 63640 81490 63860 81540
rect 63640 81420 63650 81490
rect 63850 81420 63860 81490
rect 63640 81380 63860 81420
rect 63640 81310 63650 81380
rect 63850 81310 63860 81380
rect 63640 81260 63860 81310
rect 64140 81490 64360 81540
rect 64140 81420 64150 81490
rect 64350 81420 64360 81490
rect 64140 81380 64360 81420
rect 64140 81310 64150 81380
rect 64350 81310 64360 81380
rect 64140 81260 64360 81310
rect 64640 81490 64860 81540
rect 64640 81420 64650 81490
rect 64850 81420 64860 81490
rect 64640 81380 64860 81420
rect 64640 81310 64650 81380
rect 64850 81310 64860 81380
rect 64640 81260 64860 81310
rect 65140 81490 65360 81540
rect 65140 81420 65150 81490
rect 65350 81420 65360 81490
rect 65140 81380 65360 81420
rect 65140 81310 65150 81380
rect 65350 81310 65360 81380
rect 65140 81260 65360 81310
rect 65640 81490 65860 81540
rect 65640 81420 65650 81490
rect 65850 81420 65860 81490
rect 65640 81380 65860 81420
rect 65640 81310 65650 81380
rect 65850 81310 65860 81380
rect 65640 81260 65860 81310
rect 66140 81490 66360 81540
rect 66140 81420 66150 81490
rect 66350 81420 66360 81490
rect 66140 81380 66360 81420
rect 66140 81310 66150 81380
rect 66350 81310 66360 81380
rect 66140 81260 66360 81310
rect 66640 81490 66860 81540
rect 66640 81420 66650 81490
rect 66850 81420 66860 81490
rect 66640 81380 66860 81420
rect 66640 81310 66650 81380
rect 66850 81310 66860 81380
rect 66640 81260 66860 81310
rect 67140 81490 67360 81540
rect 67140 81420 67150 81490
rect 67350 81420 67360 81490
rect 67140 81380 67360 81420
rect 67140 81310 67150 81380
rect 67350 81310 67360 81380
rect 67140 81260 67360 81310
rect 67640 81490 67860 81540
rect 67640 81420 67650 81490
rect 67850 81420 67860 81490
rect 67640 81380 67860 81420
rect 67640 81310 67650 81380
rect 67850 81310 67860 81380
rect 67640 81260 67860 81310
rect 68140 81490 68360 81540
rect 68140 81420 68150 81490
rect 68350 81420 68360 81490
rect 68140 81380 68360 81420
rect 68140 81310 68150 81380
rect 68350 81310 68360 81380
rect 68140 81260 68360 81310
rect 68640 81490 68860 81540
rect 68640 81420 68650 81490
rect 68850 81420 68860 81490
rect 68640 81380 68860 81420
rect 68640 81310 68650 81380
rect 68850 81310 68860 81380
rect 68640 81260 68860 81310
rect 69140 81490 69360 81540
rect 69140 81420 69150 81490
rect 69350 81420 69360 81490
rect 69140 81380 69360 81420
rect 69140 81310 69150 81380
rect 69350 81310 69360 81380
rect 69140 81260 69360 81310
rect 69640 81490 69860 81540
rect 69640 81420 69650 81490
rect 69850 81420 69860 81490
rect 69640 81380 69860 81420
rect 69640 81310 69650 81380
rect 69850 81310 69860 81380
rect 69640 81260 69860 81310
rect 70140 81490 70360 81540
rect 70140 81420 70150 81490
rect 70350 81420 70360 81490
rect 70140 81380 70360 81420
rect 70140 81310 70150 81380
rect 70350 81310 70360 81380
rect 70140 81260 70360 81310
rect 70640 81490 70860 81540
rect 70640 81420 70650 81490
rect 70850 81420 70860 81490
rect 70640 81380 70860 81420
rect 70640 81310 70650 81380
rect 70850 81310 70860 81380
rect 70640 81260 70860 81310
rect 71140 81490 71360 81540
rect 71140 81420 71150 81490
rect 71350 81420 71360 81490
rect 71140 81380 71360 81420
rect 71140 81310 71150 81380
rect 71350 81310 71360 81380
rect 71140 81260 71360 81310
rect 71640 81490 71860 81540
rect 71640 81420 71650 81490
rect 71850 81420 71860 81490
rect 71640 81380 71860 81420
rect 71640 81310 71650 81380
rect 71850 81310 71860 81380
rect 71640 81260 71860 81310
rect 72140 81490 72360 81540
rect 72140 81420 72150 81490
rect 72350 81420 72360 81490
rect 72140 81380 72360 81420
rect 72140 81310 72150 81380
rect 72350 81310 72360 81380
rect 72140 81260 72360 81310
rect 72640 81490 72860 81540
rect 72640 81420 72650 81490
rect 72850 81420 72860 81490
rect 72640 81380 72860 81420
rect 72640 81310 72650 81380
rect 72850 81310 72860 81380
rect 72640 81260 72860 81310
rect 73140 81490 73360 81540
rect 73140 81420 73150 81490
rect 73350 81420 73360 81490
rect 73140 81380 73360 81420
rect 73140 81310 73150 81380
rect 73350 81310 73360 81380
rect 73140 81260 73360 81310
rect 73640 81490 73860 81540
rect 73640 81420 73650 81490
rect 73850 81420 73860 81490
rect 73640 81380 73860 81420
rect 73640 81310 73650 81380
rect 73850 81310 73860 81380
rect 73640 81260 73860 81310
rect 74140 81490 74360 81540
rect 74140 81420 74150 81490
rect 74350 81420 74360 81490
rect 74140 81380 74360 81420
rect 74140 81310 74150 81380
rect 74350 81310 74360 81380
rect 74140 81260 74360 81310
rect 74640 81490 74860 81540
rect 74640 81420 74650 81490
rect 74850 81420 74860 81490
rect 74640 81380 74860 81420
rect 74640 81310 74650 81380
rect 74850 81310 74860 81380
rect 74640 81260 74860 81310
rect 75140 81490 75360 81540
rect 75140 81420 75150 81490
rect 75350 81420 75360 81490
rect 75140 81380 75360 81420
rect 75140 81310 75150 81380
rect 75350 81310 75360 81380
rect 75140 81260 75360 81310
rect 75640 81490 75860 81540
rect 75640 81420 75650 81490
rect 75850 81420 75860 81490
rect 75640 81380 75860 81420
rect 75640 81310 75650 81380
rect 75850 81310 75860 81380
rect 75640 81260 75860 81310
rect 76140 81490 76360 81540
rect 76140 81420 76150 81490
rect 76350 81420 76360 81490
rect 76140 81380 76360 81420
rect 76140 81310 76150 81380
rect 76350 81310 76360 81380
rect 76140 81260 76360 81310
rect 76640 81490 76860 81540
rect 76640 81420 76650 81490
rect 76850 81420 76860 81490
rect 76640 81380 76860 81420
rect 76640 81310 76650 81380
rect 76850 81310 76860 81380
rect 76640 81260 76860 81310
rect 77140 81490 77360 81540
rect 77140 81420 77150 81490
rect 77350 81420 77360 81490
rect 77140 81380 77360 81420
rect 77140 81310 77150 81380
rect 77350 81310 77360 81380
rect 77140 81260 77360 81310
rect 77640 81490 77860 81540
rect 77640 81420 77650 81490
rect 77850 81420 77860 81490
rect 77640 81380 77860 81420
rect 77640 81310 77650 81380
rect 77850 81310 77860 81380
rect 77640 81260 77860 81310
rect 78140 81490 78360 81540
rect 78140 81420 78150 81490
rect 78350 81420 78360 81490
rect 78140 81380 78360 81420
rect 78140 81310 78150 81380
rect 78350 81310 78360 81380
rect 78140 81260 78360 81310
rect 78640 81490 78860 81540
rect 78640 81420 78650 81490
rect 78850 81420 78860 81490
rect 78640 81380 78860 81420
rect 78640 81310 78650 81380
rect 78850 81310 78860 81380
rect 78640 81260 78860 81310
rect 79140 81490 79360 81540
rect 79140 81420 79150 81490
rect 79350 81420 79360 81490
rect 79140 81380 79360 81420
rect 79140 81310 79150 81380
rect 79350 81310 79360 81380
rect 79140 81260 79360 81310
rect 79640 81490 79860 81540
rect 79640 81420 79650 81490
rect 79850 81420 79860 81490
rect 79640 81380 79860 81420
rect 79640 81310 79650 81380
rect 79850 81310 79860 81380
rect 79640 81260 79860 81310
rect 80140 81490 80360 81540
rect 80140 81420 80150 81490
rect 80350 81420 80360 81490
rect 80140 81380 80360 81420
rect 80140 81310 80150 81380
rect 80350 81310 80360 81380
rect 80140 81260 80360 81310
rect 80640 81490 80860 81540
rect 80640 81420 80650 81490
rect 80850 81420 80860 81490
rect 80640 81380 80860 81420
rect 80640 81310 80650 81380
rect 80850 81310 80860 81380
rect 80640 81260 80860 81310
rect 81140 81490 81360 81540
rect 81140 81420 81150 81490
rect 81350 81420 81360 81490
rect 81140 81380 81360 81420
rect 81140 81310 81150 81380
rect 81350 81310 81360 81380
rect 81140 81260 81360 81310
rect 81640 81490 81860 81540
rect 81640 81420 81650 81490
rect 81850 81420 81860 81490
rect 81640 81380 81860 81420
rect 81640 81310 81650 81380
rect 81850 81310 81860 81380
rect 81640 81260 81860 81310
rect 82140 81490 82360 81540
rect 82140 81420 82150 81490
rect 82350 81420 82360 81490
rect 82140 81380 82360 81420
rect 82140 81310 82150 81380
rect 82350 81310 82360 81380
rect 82140 81260 82360 81310
rect 82640 81490 82860 81540
rect 82640 81420 82650 81490
rect 82850 81420 82860 81490
rect 82640 81380 82860 81420
rect 82640 81310 82650 81380
rect 82850 81310 82860 81380
rect 82640 81260 82860 81310
rect 83140 81490 83360 81540
rect 83140 81420 83150 81490
rect 83350 81420 83360 81490
rect 83140 81380 83360 81420
rect 83140 81310 83150 81380
rect 83350 81310 83360 81380
rect 83140 81260 83360 81310
rect 83640 81490 83860 81540
rect 83640 81420 83650 81490
rect 83850 81420 83860 81490
rect 83640 81380 83860 81420
rect 83640 81310 83650 81380
rect 83850 81310 83860 81380
rect 83640 81260 83860 81310
rect 84140 81490 84360 81540
rect 84140 81420 84150 81490
rect 84350 81420 84360 81490
rect 84140 81380 84360 81420
rect 84140 81310 84150 81380
rect 84350 81310 84360 81380
rect 84140 81260 84360 81310
rect 84640 81490 84860 81540
rect 84640 81420 84650 81490
rect 84850 81420 84860 81490
rect 84640 81380 84860 81420
rect 84640 81310 84650 81380
rect 84850 81310 84860 81380
rect 84640 81260 84860 81310
rect 85140 81490 85360 81540
rect 85140 81420 85150 81490
rect 85350 81420 85360 81490
rect 85140 81380 85360 81420
rect 85140 81310 85150 81380
rect 85350 81310 85360 81380
rect 85140 81260 85360 81310
rect 85640 81490 85860 81540
rect 85640 81420 85650 81490
rect 85850 81420 85860 81490
rect 85640 81380 85860 81420
rect 85640 81310 85650 81380
rect 85850 81310 85860 81380
rect 85640 81260 85860 81310
rect 86140 81490 86360 81540
rect 86140 81420 86150 81490
rect 86350 81420 86360 81490
rect 86140 81380 86360 81420
rect 86140 81310 86150 81380
rect 86350 81310 86360 81380
rect 86140 81260 86360 81310
rect 86640 81490 86860 81540
rect 86640 81420 86650 81490
rect 86850 81420 86860 81490
rect 86640 81380 86860 81420
rect 86640 81310 86650 81380
rect 86850 81310 86860 81380
rect 86640 81260 86860 81310
rect 87140 81490 87360 81540
rect 87140 81420 87150 81490
rect 87350 81420 87360 81490
rect 87140 81380 87360 81420
rect 87140 81310 87150 81380
rect 87350 81310 87360 81380
rect 87140 81260 87360 81310
rect 87640 81490 87860 81540
rect 87640 81420 87650 81490
rect 87850 81420 87860 81490
rect 87640 81380 87860 81420
rect 87640 81310 87650 81380
rect 87850 81310 87860 81380
rect 87640 81260 87860 81310
rect 88140 81490 88360 81540
rect 88140 81420 88150 81490
rect 88350 81420 88360 81490
rect 88140 81380 88360 81420
rect 88140 81310 88150 81380
rect 88350 81310 88360 81380
rect 88140 81260 88360 81310
rect 88640 81490 88860 81540
rect 88640 81420 88650 81490
rect 88850 81420 88860 81490
rect 88640 81380 88860 81420
rect 88640 81310 88650 81380
rect 88850 81310 88860 81380
rect 88640 81260 88860 81310
rect 89140 81490 89360 81540
rect 89140 81420 89150 81490
rect 89350 81420 89360 81490
rect 89140 81380 89360 81420
rect 89140 81310 89150 81380
rect 89350 81310 89360 81380
rect 89140 81260 89360 81310
rect 89640 81490 89860 81540
rect 89640 81420 89650 81490
rect 89850 81420 89860 81490
rect 89640 81380 89860 81420
rect 89640 81310 89650 81380
rect 89850 81310 89860 81380
rect 89640 81260 89860 81310
rect 90140 81490 90360 81540
rect 90140 81420 90150 81490
rect 90350 81420 90360 81490
rect 90140 81380 90360 81420
rect 90140 81310 90150 81380
rect 90350 81310 90360 81380
rect 90140 81260 90360 81310
rect 90640 81490 90860 81540
rect 90640 81420 90650 81490
rect 90850 81420 90860 81490
rect 90640 81380 90860 81420
rect 90640 81310 90650 81380
rect 90850 81310 90860 81380
rect 90640 81260 90860 81310
rect 91140 81490 91360 81540
rect 91140 81420 91150 81490
rect 91350 81420 91360 81490
rect 91140 81380 91360 81420
rect 91140 81310 91150 81380
rect 91350 81310 91360 81380
rect 91140 81260 91360 81310
rect 91640 81490 91860 81540
rect 91640 81420 91650 81490
rect 91850 81420 91860 81490
rect 91640 81380 91860 81420
rect 91640 81310 91650 81380
rect 91850 81310 91860 81380
rect 91640 81260 91860 81310
rect 92140 81490 92360 81540
rect 92140 81420 92150 81490
rect 92350 81420 92360 81490
rect 92140 81380 92360 81420
rect 92140 81310 92150 81380
rect 92350 81310 92360 81380
rect 92140 81260 92360 81310
rect 92640 81490 92860 81540
rect 92640 81420 92650 81490
rect 92850 81420 92860 81490
rect 92640 81380 92860 81420
rect 92640 81310 92650 81380
rect 92850 81310 92860 81380
rect 92640 81260 92860 81310
rect 93140 81490 93360 81540
rect 93140 81420 93150 81490
rect 93350 81420 93360 81490
rect 93140 81380 93360 81420
rect 93140 81310 93150 81380
rect 93350 81310 93360 81380
rect 93140 81260 93360 81310
rect 93640 81490 93860 81540
rect 93640 81420 93650 81490
rect 93850 81420 93860 81490
rect 93640 81380 93860 81420
rect 93640 81310 93650 81380
rect 93850 81310 93860 81380
rect 93640 81260 93860 81310
rect 94140 81490 94360 81540
rect 94140 81420 94150 81490
rect 94350 81420 94360 81490
rect 94140 81380 94360 81420
rect 94140 81310 94150 81380
rect 94350 81310 94360 81380
rect 94140 81260 94360 81310
rect 94640 81490 94860 81540
rect 94640 81420 94650 81490
rect 94850 81420 94860 81490
rect 94640 81380 94860 81420
rect 94640 81310 94650 81380
rect 94850 81310 94860 81380
rect 94640 81260 94860 81310
rect 95140 81490 95360 81540
rect 95140 81420 95150 81490
rect 95350 81420 95360 81490
rect 95140 81380 95360 81420
rect 95140 81310 95150 81380
rect 95350 81310 95360 81380
rect 95140 81260 95360 81310
rect 95640 81490 95860 81540
rect 95640 81420 95650 81490
rect 95850 81420 95860 81490
rect 95640 81380 95860 81420
rect 95640 81310 95650 81380
rect 95850 81310 95860 81380
rect 95640 81260 95860 81310
rect 96140 81490 96360 81540
rect 96140 81420 96150 81490
rect 96350 81420 96360 81490
rect 96140 81380 96360 81420
rect 96140 81310 96150 81380
rect 96350 81310 96360 81380
rect 96140 81260 96360 81310
rect 96640 81490 96860 81540
rect 96640 81420 96650 81490
rect 96850 81420 96860 81490
rect 96640 81380 96860 81420
rect 96640 81310 96650 81380
rect 96850 81310 96860 81380
rect 96640 81260 96860 81310
rect 97140 81490 97360 81540
rect 97140 81420 97150 81490
rect 97350 81420 97360 81490
rect 97140 81380 97360 81420
rect 97140 81310 97150 81380
rect 97350 81310 97360 81380
rect 97140 81260 97360 81310
rect 97640 81490 97860 81540
rect 97640 81420 97650 81490
rect 97850 81420 97860 81490
rect 97640 81380 97860 81420
rect 97640 81310 97650 81380
rect 97850 81310 97860 81380
rect 97640 81260 97860 81310
rect 98140 81490 98360 81540
rect 98140 81420 98150 81490
rect 98350 81420 98360 81490
rect 98140 81380 98360 81420
rect 98140 81310 98150 81380
rect 98350 81310 98360 81380
rect 98140 81260 98360 81310
rect 98640 81490 98860 81540
rect 98640 81420 98650 81490
rect 98850 81420 98860 81490
rect 98640 81380 98860 81420
rect 98640 81310 98650 81380
rect 98850 81310 98860 81380
rect 98640 81260 98860 81310
rect 99140 81490 99360 81540
rect 99140 81420 99150 81490
rect 99350 81420 99360 81490
rect 99140 81380 99360 81420
rect 99140 81310 99150 81380
rect 99350 81310 99360 81380
rect 99140 81260 99360 81310
rect 99640 81490 99860 81540
rect 99640 81420 99650 81490
rect 99850 81420 99860 81490
rect 99640 81380 99860 81420
rect 99640 81310 99650 81380
rect 99850 81310 99860 81380
rect 99640 81260 99860 81310
rect 100140 81490 100360 81540
rect 100140 81420 100150 81490
rect 100350 81420 100360 81490
rect 100140 81380 100360 81420
rect 100140 81310 100150 81380
rect 100350 81310 100360 81380
rect 100140 81260 100360 81310
rect -83500 81250 100500 81260
rect -83500 81050 -83480 81250
rect -83410 81050 -83090 81250
rect -83020 81050 -82980 81250
rect -82910 81050 -82590 81250
rect -82520 81050 -82480 81250
rect -82410 81050 -82090 81250
rect -82020 81050 -81980 81250
rect -81910 81050 -81590 81250
rect -81520 81050 -81480 81250
rect -81410 81050 -81090 81250
rect -81020 81050 -80980 81250
rect -80910 81050 -80590 81250
rect -80520 81050 -80480 81250
rect -80410 81050 -80090 81250
rect -80020 81050 -79980 81250
rect -79910 81050 -79590 81250
rect -79520 81050 -79480 81250
rect -79410 81050 -79090 81250
rect -79020 81050 -78980 81250
rect -78910 81050 -78590 81250
rect -78520 81050 -78480 81250
rect -78410 81050 -78090 81250
rect -78020 81050 -77980 81250
rect -77910 81050 -77590 81250
rect -77520 81050 -77480 81250
rect -77410 81050 -77090 81250
rect -77020 81050 -76980 81250
rect -76910 81050 -76590 81250
rect -76520 81050 -76480 81250
rect -76410 81050 -76090 81250
rect -76020 81050 -75980 81250
rect -75910 81050 -75590 81250
rect -75520 81050 -75480 81250
rect -75410 81050 -75090 81250
rect -75020 81050 -74980 81250
rect -74910 81050 -74590 81250
rect -74520 81050 -74480 81250
rect -74410 81050 -74090 81250
rect -74020 81050 -73980 81250
rect -73910 81050 -73590 81250
rect -73520 81050 -73480 81250
rect -73410 81050 -73090 81250
rect -73020 81050 -72980 81250
rect -72910 81050 -72590 81250
rect -72520 81050 -72480 81250
rect -72410 81050 -72090 81250
rect -72020 81050 -71980 81250
rect -71910 81050 -71590 81250
rect -71520 81050 -71480 81250
rect -71410 81050 -71090 81250
rect -71020 81050 -70980 81250
rect -70910 81050 -70590 81250
rect -70520 81050 -70480 81250
rect -70410 81050 -70090 81250
rect -70020 81050 -69980 81250
rect -69910 81050 -69590 81250
rect -69520 81050 -69480 81250
rect -69410 81050 -69090 81250
rect -69020 81050 -68980 81250
rect -68910 81050 -68590 81250
rect -68520 81050 -68480 81250
rect -68410 81050 -68090 81250
rect -68020 81050 -67980 81250
rect -67910 81050 -67590 81250
rect -67520 81050 -67480 81250
rect -67410 81050 -67090 81250
rect -67020 81050 -66980 81250
rect -66910 81050 -66590 81250
rect -66520 81050 -66480 81250
rect -66410 81050 -66090 81250
rect -66020 81050 -65980 81250
rect -65910 81050 -65590 81250
rect -65520 81050 -65480 81250
rect -65410 81050 -65090 81250
rect -65020 81050 -64980 81250
rect -64910 81050 -64590 81250
rect -64520 81050 -64480 81250
rect -64410 81050 -64090 81250
rect -64020 81050 -63980 81250
rect -63910 81050 -63590 81250
rect -63520 81050 -63480 81250
rect -63410 81050 -63090 81250
rect -63020 81050 -62980 81250
rect -62910 81050 -62590 81250
rect -62520 81050 -62480 81250
rect -62410 81050 -62090 81250
rect -62020 81050 -61980 81250
rect -61910 81050 -61590 81250
rect -61520 81050 -61480 81250
rect -61410 81050 -61090 81250
rect -61020 81050 -60980 81250
rect -60910 81050 -60590 81250
rect -60520 81050 -60480 81250
rect -60410 81050 -60090 81250
rect -60020 81050 -59980 81250
rect -59910 81050 -59590 81250
rect -59520 81050 -59480 81250
rect -59410 81050 -59090 81250
rect -59020 81050 -58980 81250
rect -58910 81050 -58590 81250
rect -58520 81050 -58480 81250
rect -58410 81050 -58090 81250
rect -58020 81050 -57980 81250
rect -57910 81050 -57590 81250
rect -57520 81050 -57480 81250
rect -57410 81050 -57090 81250
rect -57020 81050 -56980 81250
rect -56910 81050 -56590 81250
rect -56520 81050 -56480 81250
rect -56410 81050 -56090 81250
rect -56020 81050 -55980 81250
rect -55910 81050 -55590 81250
rect -55520 81050 -55480 81250
rect -55410 81050 -55090 81250
rect -55020 81050 -54980 81250
rect -54910 81050 -54590 81250
rect -54520 81050 -54480 81250
rect -54410 81050 -54090 81250
rect -54020 81050 -53980 81250
rect -53910 81050 -53590 81250
rect -53520 81050 -53480 81250
rect -53410 81050 -53090 81250
rect -53020 81050 -52980 81250
rect -52910 81050 -52590 81250
rect -52520 81050 -52480 81250
rect -52410 81050 -52090 81250
rect -52020 81050 -51980 81250
rect -51910 81050 -51590 81250
rect -51520 81050 -51480 81250
rect -51410 81050 -51090 81250
rect -51020 81050 -50980 81250
rect -50910 81050 -50590 81250
rect -50520 81050 -50480 81250
rect -50410 81050 -50090 81250
rect -50020 81050 -49980 81250
rect -49910 81050 -49590 81250
rect -49520 81050 -49480 81250
rect -49410 81050 -49090 81250
rect -49020 81050 -48980 81250
rect -48910 81050 -48590 81250
rect -48520 81050 -48480 81250
rect -48410 81050 -48090 81250
rect -48020 81050 -47980 81250
rect -47910 81050 -47590 81250
rect -47520 81050 -47480 81250
rect -47410 81050 -47090 81250
rect -47020 81050 -46980 81250
rect -46910 81050 -46590 81250
rect -46520 81050 -46480 81250
rect -46410 81050 -46090 81250
rect -46020 81050 -45980 81250
rect -45910 81050 -45590 81250
rect -45520 81050 -45480 81250
rect -45410 81050 -45090 81250
rect -45020 81050 -44980 81250
rect -44910 81050 -44590 81250
rect -44520 81050 -44480 81250
rect -44410 81050 -44090 81250
rect -44020 81050 -43980 81250
rect -43910 81050 -43590 81250
rect -43520 81050 -43480 81250
rect -43410 81050 -43090 81250
rect -43020 81050 -42980 81250
rect -42910 81050 -42590 81250
rect -42520 81050 -42480 81250
rect -42410 81050 -42090 81250
rect -42020 81050 -41980 81250
rect -41910 81050 -41590 81250
rect -41520 81050 -41480 81250
rect -41410 81050 -41090 81250
rect -41020 81050 -40980 81250
rect -40910 81050 -40590 81250
rect -40520 81050 -40480 81250
rect -40410 81050 -40090 81250
rect -40020 81050 -39980 81250
rect -39910 81050 -39590 81250
rect -39520 81050 -39480 81250
rect -39410 81050 -39090 81250
rect -39020 81050 -38980 81250
rect -38910 81050 -38590 81250
rect -38520 81050 -38480 81250
rect -38410 81050 -38090 81250
rect -38020 81050 -37980 81250
rect -37910 81050 -37590 81250
rect -37520 81050 -37480 81250
rect -37410 81050 -37090 81250
rect -37020 81050 -36980 81250
rect -36910 81050 -36590 81250
rect -36520 81050 -36480 81250
rect -36410 81050 -36090 81250
rect -36020 81050 -35980 81250
rect -35910 81050 -35590 81250
rect -35520 81050 -35480 81250
rect -35410 81050 -35090 81250
rect -35020 81050 -34980 81250
rect -34910 81050 -34590 81250
rect -34520 81050 -34480 81250
rect -34410 81050 -34090 81250
rect -34020 81050 -33980 81250
rect -33910 81050 -33590 81250
rect -33520 81050 -33480 81250
rect -33410 81050 -33090 81250
rect -33020 81050 -32980 81250
rect -32910 81050 -32590 81250
rect -32520 81050 -32480 81250
rect -32410 81050 -32090 81250
rect -32020 81050 -31980 81250
rect -31910 81050 -31590 81250
rect -31520 81050 -31480 81250
rect -31410 81050 -31090 81250
rect -31020 81050 -30980 81250
rect -30910 81050 -30590 81250
rect -30520 81050 -30480 81250
rect -30410 81050 -30090 81250
rect -30020 81050 -29980 81250
rect -29910 81050 -29590 81250
rect -29520 81050 -29480 81250
rect -29410 81050 -29090 81250
rect -29020 81050 -28980 81250
rect -28910 81050 -28590 81250
rect -28520 81050 -28480 81250
rect -28410 81050 -28090 81250
rect -28020 81050 -27980 81250
rect -27910 81050 -27590 81250
rect -27520 81050 -27480 81250
rect -27410 81050 -27090 81250
rect -27020 81050 -26980 81250
rect -26910 81050 -26590 81250
rect -26520 81050 -26480 81250
rect -26410 81050 -26090 81250
rect -26020 81050 -25980 81250
rect -25910 81050 -25590 81250
rect -25520 81050 -25480 81250
rect -25410 81050 -25090 81250
rect -25020 81050 -24980 81250
rect -24910 81050 -24590 81250
rect -24520 81050 -24480 81250
rect -24410 81050 -24090 81250
rect -24020 81050 -23980 81250
rect -23910 81050 -23590 81250
rect -23520 81050 -23480 81250
rect -23410 81050 -23090 81250
rect -23020 81050 -22980 81250
rect -22910 81050 -22590 81250
rect -22520 81050 -22480 81250
rect -22410 81050 -22090 81250
rect -22020 81050 -21980 81250
rect -21910 81050 -21590 81250
rect -21520 81050 -21480 81250
rect -21410 81050 -21090 81250
rect -21020 81050 -20980 81250
rect -20910 81050 -20590 81250
rect -20520 81050 -20480 81250
rect -20410 81050 -20090 81250
rect -20020 81050 -19980 81250
rect -19910 81050 -19590 81250
rect -19520 81050 -19480 81250
rect -19410 81050 -19090 81250
rect -19020 81050 -18980 81250
rect -18910 81050 -18590 81250
rect -18520 81050 -18480 81250
rect -18410 81050 -18090 81250
rect -18020 81050 -17980 81250
rect -17910 81050 -17590 81250
rect -17520 81050 -17480 81250
rect -17410 81050 -17090 81250
rect -17020 81050 -16980 81250
rect -16910 81050 -16590 81250
rect -16520 81050 -16480 81250
rect -16410 81050 -16090 81250
rect -16020 81050 -15980 81250
rect -15910 81050 -15590 81250
rect -15520 81050 -15480 81250
rect -15410 81050 -15090 81250
rect -15020 81050 -14980 81250
rect -14910 81050 -14590 81250
rect -14520 81050 -14480 81250
rect -14410 81050 -14090 81250
rect -14020 81050 -13980 81250
rect -13910 81050 -13590 81250
rect -13520 81050 -13480 81250
rect -13410 81050 -13090 81250
rect -13020 81050 -12980 81250
rect -12910 81050 -12590 81250
rect -12520 81050 -12480 81250
rect -12410 81050 -12090 81250
rect -12020 81050 -11980 81250
rect -11910 81050 -11590 81250
rect -11520 81050 -11480 81250
rect -11410 81050 -11090 81250
rect -11020 81050 -10980 81250
rect -10910 81050 -10590 81250
rect -10520 81050 -10480 81250
rect -10410 81050 -10090 81250
rect -10020 81050 -9980 81250
rect -9910 81050 -9590 81250
rect -9520 81050 -9480 81250
rect -9410 81050 -9090 81250
rect -9020 81050 -8980 81250
rect -8910 81050 -8590 81250
rect -8520 81050 -8480 81250
rect -8410 81050 -8090 81250
rect -8020 81050 -7980 81250
rect -7910 81050 -7590 81250
rect -7520 81050 -7480 81250
rect -7410 81050 -7090 81250
rect -7020 81050 -6980 81250
rect -6910 81050 -6590 81250
rect -6520 81050 -6480 81250
rect -6410 81050 -6090 81250
rect -6020 81050 -5980 81250
rect -5910 81050 -5590 81250
rect -5520 81050 -5480 81250
rect -5410 81050 -5090 81250
rect -5020 81050 -4980 81250
rect -4910 81050 -4590 81250
rect -4520 81050 -4480 81250
rect -4410 81050 -4090 81250
rect -4020 81050 -3980 81250
rect -3910 81050 -3590 81250
rect -3520 81050 -3480 81250
rect -3410 81050 -3090 81250
rect -3020 81050 -2980 81250
rect -2910 81050 -2590 81250
rect -2520 81050 -2480 81250
rect -2410 81050 -2090 81250
rect -2020 81050 -1980 81250
rect -1910 81050 -1590 81250
rect -1520 81050 -1480 81250
rect -1410 81050 -1090 81250
rect -1020 81050 -980 81250
rect -910 81050 -590 81250
rect -520 81050 -480 81250
rect -410 81050 -90 81250
rect -20 81050 20 81250
rect 90 81050 410 81250
rect 480 81050 520 81250
rect 590 81050 910 81250
rect 980 81050 1020 81250
rect 1090 81050 1410 81250
rect 1480 81050 1520 81250
rect 1590 81050 1910 81250
rect 1980 81050 2020 81250
rect 2090 81050 2410 81250
rect 2480 81050 2520 81250
rect 2590 81050 2910 81250
rect 2980 81050 3020 81250
rect 3090 81050 3410 81250
rect 3480 81050 3520 81250
rect 3590 81050 3910 81250
rect 3980 81050 4020 81250
rect 4090 81050 4410 81250
rect 4480 81050 4520 81250
rect 4590 81050 4910 81250
rect 4980 81050 5020 81250
rect 5090 81050 5410 81250
rect 5480 81050 5520 81250
rect 5590 81050 5910 81250
rect 5980 81050 6020 81250
rect 6090 81050 6410 81250
rect 6480 81050 6520 81250
rect 6590 81050 6910 81250
rect 6980 81050 7020 81250
rect 7090 81050 7410 81250
rect 7480 81050 7520 81250
rect 7590 81050 7910 81250
rect 7980 81050 8020 81250
rect 8090 81050 8410 81250
rect 8480 81050 8520 81250
rect 8590 81050 8910 81250
rect 8980 81050 9020 81250
rect 9090 81050 9410 81250
rect 9480 81050 9520 81250
rect 9590 81050 9910 81250
rect 9980 81050 10020 81250
rect 10090 81050 10410 81250
rect 10480 81050 10520 81250
rect 10590 81050 10910 81250
rect 10980 81050 11020 81250
rect 11090 81050 11410 81250
rect 11480 81050 11520 81250
rect 11590 81050 11910 81250
rect 11980 81050 12020 81250
rect 12090 81050 12410 81250
rect 12480 81050 12520 81250
rect 12590 81050 12910 81250
rect 12980 81050 13020 81250
rect 13090 81050 13410 81250
rect 13480 81050 13520 81250
rect 13590 81050 13910 81250
rect 13980 81050 14020 81250
rect 14090 81050 14410 81250
rect 14480 81050 14520 81250
rect 14590 81050 14910 81250
rect 14980 81050 15020 81250
rect 15090 81050 15410 81250
rect 15480 81050 15520 81250
rect 15590 81050 15910 81250
rect 15980 81050 16020 81250
rect 16090 81050 16410 81250
rect 16480 81050 16520 81250
rect 16590 81050 16910 81250
rect 16980 81050 17020 81250
rect 17090 81050 17410 81250
rect 17480 81050 17520 81250
rect 17590 81050 17910 81250
rect 17980 81050 18020 81250
rect 18090 81050 18410 81250
rect 18480 81050 18520 81250
rect 18590 81050 18910 81250
rect 18980 81050 19020 81250
rect 19090 81050 19410 81250
rect 19480 81050 19520 81250
rect 19590 81050 19910 81250
rect 19980 81050 20020 81250
rect 20090 81050 20410 81250
rect 20480 81050 20520 81250
rect 20590 81050 20910 81250
rect 20980 81050 21020 81250
rect 21090 81050 21410 81250
rect 21480 81050 21520 81250
rect 21590 81050 21910 81250
rect 21980 81050 22020 81250
rect 22090 81050 22410 81250
rect 22480 81050 22520 81250
rect 22590 81050 22910 81250
rect 22980 81050 23020 81250
rect 23090 81050 23410 81250
rect 23480 81050 23520 81250
rect 23590 81050 23910 81250
rect 23980 81050 24020 81250
rect 24090 81050 24410 81250
rect 24480 81050 24520 81250
rect 24590 81050 24910 81250
rect 24980 81050 25020 81250
rect 25090 81050 25410 81250
rect 25480 81050 25520 81250
rect 25590 81050 25910 81250
rect 25980 81050 26020 81250
rect 26090 81050 26410 81250
rect 26480 81050 26520 81250
rect 26590 81050 26910 81250
rect 26980 81050 27020 81250
rect 27090 81050 27410 81250
rect 27480 81050 27520 81250
rect 27590 81050 27910 81250
rect 27980 81050 28020 81250
rect 28090 81050 28410 81250
rect 28480 81050 28520 81250
rect 28590 81050 28910 81250
rect 28980 81050 29020 81250
rect 29090 81050 29410 81250
rect 29480 81050 29520 81250
rect 29590 81050 29910 81250
rect 29980 81050 30020 81250
rect 30090 81050 30410 81250
rect 30480 81050 30520 81250
rect 30590 81050 30910 81250
rect 30980 81050 31020 81250
rect 31090 81050 31410 81250
rect 31480 81050 31520 81250
rect 31590 81050 31910 81250
rect 31980 81050 32020 81250
rect 32090 81050 32410 81250
rect 32480 81050 32520 81250
rect 32590 81050 32910 81250
rect 32980 81050 33020 81250
rect 33090 81050 33410 81250
rect 33480 81050 33520 81250
rect 33590 81050 33910 81250
rect 33980 81050 34020 81250
rect 34090 81050 34410 81250
rect 34480 81050 34520 81250
rect 34590 81050 34910 81250
rect 34980 81050 35020 81250
rect 35090 81050 35410 81250
rect 35480 81050 35520 81250
rect 35590 81050 35910 81250
rect 35980 81050 36020 81250
rect 36090 81050 36410 81250
rect 36480 81050 36520 81250
rect 36590 81050 36910 81250
rect 36980 81050 37020 81250
rect 37090 81050 37410 81250
rect 37480 81050 37520 81250
rect 37590 81050 37910 81250
rect 37980 81050 38020 81250
rect 38090 81050 38410 81250
rect 38480 81050 38520 81250
rect 38590 81050 38910 81250
rect 38980 81050 39020 81250
rect 39090 81050 39410 81250
rect 39480 81050 39520 81250
rect 39590 81050 39910 81250
rect 39980 81050 40020 81250
rect 40090 81050 40410 81250
rect 40480 81050 40520 81250
rect 40590 81050 40910 81250
rect 40980 81050 41020 81250
rect 41090 81050 41410 81250
rect 41480 81050 41520 81250
rect 41590 81050 41910 81250
rect 41980 81050 42020 81250
rect 42090 81050 42410 81250
rect 42480 81050 42520 81250
rect 42590 81050 42910 81250
rect 42980 81050 43020 81250
rect 43090 81050 43410 81250
rect 43480 81050 43520 81250
rect 43590 81050 43910 81250
rect 43980 81050 44020 81250
rect 44090 81050 44410 81250
rect 44480 81050 44520 81250
rect 44590 81050 44910 81250
rect 44980 81050 45020 81250
rect 45090 81050 45410 81250
rect 45480 81050 45520 81250
rect 45590 81050 45910 81250
rect 45980 81050 46020 81250
rect 46090 81050 46410 81250
rect 46480 81050 46520 81250
rect 46590 81050 46910 81250
rect 46980 81050 47020 81250
rect 47090 81050 47410 81250
rect 47480 81050 47520 81250
rect 47590 81050 47910 81250
rect 47980 81050 48020 81250
rect 48090 81050 48410 81250
rect 48480 81050 48520 81250
rect 48590 81050 48910 81250
rect 48980 81050 49020 81250
rect 49090 81050 49410 81250
rect 49480 81050 49520 81250
rect 49590 81050 49910 81250
rect 49980 81050 50020 81250
rect 50090 81050 50410 81250
rect 50480 81050 50520 81250
rect 50590 81050 50910 81250
rect 50980 81050 51020 81250
rect 51090 81050 51410 81250
rect 51480 81050 51520 81250
rect 51590 81050 51910 81250
rect 51980 81050 52020 81250
rect 52090 81050 52410 81250
rect 52480 81050 52520 81250
rect 52590 81050 52910 81250
rect 52980 81050 53020 81250
rect 53090 81050 53410 81250
rect 53480 81050 53520 81250
rect 53590 81050 53910 81250
rect 53980 81050 54020 81250
rect 54090 81050 54410 81250
rect 54480 81050 54520 81250
rect 54590 81050 54910 81250
rect 54980 81050 55020 81250
rect 55090 81050 55410 81250
rect 55480 81050 55520 81250
rect 55590 81050 55910 81250
rect 55980 81050 56020 81250
rect 56090 81050 56410 81250
rect 56480 81050 56520 81250
rect 56590 81050 56910 81250
rect 56980 81050 57020 81250
rect 57090 81050 57410 81250
rect 57480 81050 57520 81250
rect 57590 81050 57910 81250
rect 57980 81050 58020 81250
rect 58090 81050 58410 81250
rect 58480 81050 58520 81250
rect 58590 81050 58910 81250
rect 58980 81050 59020 81250
rect 59090 81050 59410 81250
rect 59480 81050 59520 81250
rect 59590 81050 59910 81250
rect 59980 81050 60020 81250
rect 60090 81050 60410 81250
rect 60480 81050 60520 81250
rect 60590 81050 60910 81250
rect 60980 81050 61020 81250
rect 61090 81050 61410 81250
rect 61480 81050 61520 81250
rect 61590 81050 61910 81250
rect 61980 81050 62020 81250
rect 62090 81050 62410 81250
rect 62480 81050 62520 81250
rect 62590 81050 62910 81250
rect 62980 81050 63020 81250
rect 63090 81050 63410 81250
rect 63480 81050 63520 81250
rect 63590 81050 63910 81250
rect 63980 81050 64020 81250
rect 64090 81050 64410 81250
rect 64480 81050 64520 81250
rect 64590 81050 64910 81250
rect 64980 81050 65020 81250
rect 65090 81050 65410 81250
rect 65480 81050 65520 81250
rect 65590 81050 65910 81250
rect 65980 81050 66020 81250
rect 66090 81050 66410 81250
rect 66480 81050 66520 81250
rect 66590 81050 66910 81250
rect 66980 81050 67020 81250
rect 67090 81050 67410 81250
rect 67480 81050 67520 81250
rect 67590 81050 67910 81250
rect 67980 81050 68020 81250
rect 68090 81050 68410 81250
rect 68480 81050 68520 81250
rect 68590 81050 68910 81250
rect 68980 81050 69020 81250
rect 69090 81050 69410 81250
rect 69480 81050 69520 81250
rect 69590 81050 69910 81250
rect 69980 81050 70020 81250
rect 70090 81050 70410 81250
rect 70480 81050 70520 81250
rect 70590 81050 70910 81250
rect 70980 81050 71020 81250
rect 71090 81050 71410 81250
rect 71480 81050 71520 81250
rect 71590 81050 71910 81250
rect 71980 81050 72020 81250
rect 72090 81050 72410 81250
rect 72480 81050 72520 81250
rect 72590 81050 72910 81250
rect 72980 81050 73020 81250
rect 73090 81050 73410 81250
rect 73480 81050 73520 81250
rect 73590 81050 73910 81250
rect 73980 81050 74020 81250
rect 74090 81050 74410 81250
rect 74480 81050 74520 81250
rect 74590 81050 74910 81250
rect 74980 81050 75020 81250
rect 75090 81050 75410 81250
rect 75480 81050 75520 81250
rect 75590 81050 75910 81250
rect 75980 81050 76020 81250
rect 76090 81050 76410 81250
rect 76480 81050 76520 81250
rect 76590 81050 76910 81250
rect 76980 81050 77020 81250
rect 77090 81050 77410 81250
rect 77480 81050 77520 81250
rect 77590 81050 77910 81250
rect 77980 81050 78020 81250
rect 78090 81050 78410 81250
rect 78480 81050 78520 81250
rect 78590 81050 78910 81250
rect 78980 81050 79020 81250
rect 79090 81050 79410 81250
rect 79480 81050 79520 81250
rect 79590 81050 79910 81250
rect 79980 81050 80020 81250
rect 80090 81050 80410 81250
rect 80480 81050 80520 81250
rect 80590 81050 80910 81250
rect 80980 81050 81020 81250
rect 81090 81050 81410 81250
rect 81480 81050 81520 81250
rect 81590 81050 81910 81250
rect 81980 81050 82020 81250
rect 82090 81050 82410 81250
rect 82480 81050 82520 81250
rect 82590 81050 82910 81250
rect 82980 81050 83020 81250
rect 83090 81050 83410 81250
rect 83480 81050 83520 81250
rect 83590 81050 83910 81250
rect 83980 81050 84020 81250
rect 84090 81050 84410 81250
rect 84480 81050 84520 81250
rect 84590 81050 84910 81250
rect 84980 81050 85020 81250
rect 85090 81050 85410 81250
rect 85480 81050 85520 81250
rect 85590 81050 85910 81250
rect 85980 81050 86020 81250
rect 86090 81050 86410 81250
rect 86480 81050 86520 81250
rect 86590 81050 86910 81250
rect 86980 81050 87020 81250
rect 87090 81050 87410 81250
rect 87480 81050 87520 81250
rect 87590 81050 87910 81250
rect 87980 81050 88020 81250
rect 88090 81050 88410 81250
rect 88480 81050 88520 81250
rect 88590 81050 88910 81250
rect 88980 81050 89020 81250
rect 89090 81050 89410 81250
rect 89480 81050 89520 81250
rect 89590 81050 89910 81250
rect 89980 81050 90020 81250
rect 90090 81050 90410 81250
rect 90480 81050 90520 81250
rect 90590 81050 90910 81250
rect 90980 81050 91020 81250
rect 91090 81050 91410 81250
rect 91480 81050 91520 81250
rect 91590 81050 91910 81250
rect 91980 81050 92020 81250
rect 92090 81050 92410 81250
rect 92480 81050 92520 81250
rect 92590 81050 92910 81250
rect 92980 81050 93020 81250
rect 93090 81050 93410 81250
rect 93480 81050 93520 81250
rect 93590 81050 93910 81250
rect 93980 81050 94020 81250
rect 94090 81050 94410 81250
rect 94480 81050 94520 81250
rect 94590 81050 94910 81250
rect 94980 81050 95020 81250
rect 95090 81050 95410 81250
rect 95480 81050 95520 81250
rect 95590 81050 95910 81250
rect 95980 81050 96020 81250
rect 96090 81050 96410 81250
rect 96480 81050 96520 81250
rect 96590 81050 96910 81250
rect 96980 81050 97020 81250
rect 97090 81050 97410 81250
rect 97480 81050 97520 81250
rect 97590 81050 97910 81250
rect 97980 81050 98020 81250
rect 98090 81050 98410 81250
rect 98480 81050 98520 81250
rect 98590 81050 98910 81250
rect 98980 81050 99020 81250
rect 99090 81050 99410 81250
rect 99480 81050 99520 81250
rect 99590 81050 99910 81250
rect 99980 81050 100020 81250
rect 100090 81050 100410 81250
rect 100480 81050 100500 81250
rect -83500 81040 100500 81050
rect -83360 80990 -83140 81040
rect -83360 80920 -83350 80990
rect -83150 80920 -83140 80990
rect -83360 80880 -83140 80920
rect -83360 80810 -83350 80880
rect -83150 80810 -83140 80880
rect -83360 80760 -83140 80810
rect -82860 80990 -82640 81040
rect -82860 80920 -82850 80990
rect -82650 80920 -82640 80990
rect -82860 80880 -82640 80920
rect -82860 80810 -82850 80880
rect -82650 80810 -82640 80880
rect -82860 80760 -82640 80810
rect -82360 80990 -82140 81040
rect -82360 80920 -82350 80990
rect -82150 80920 -82140 80990
rect -82360 80880 -82140 80920
rect -82360 80810 -82350 80880
rect -82150 80810 -82140 80880
rect -82360 80760 -82140 80810
rect -81860 80990 -81640 81040
rect -81860 80920 -81850 80990
rect -81650 80920 -81640 80990
rect -81860 80880 -81640 80920
rect -81860 80810 -81850 80880
rect -81650 80810 -81640 80880
rect -81860 80760 -81640 80810
rect -81360 80990 -81140 81040
rect -81360 80920 -81350 80990
rect -81150 80920 -81140 80990
rect -81360 80880 -81140 80920
rect -81360 80810 -81350 80880
rect -81150 80810 -81140 80880
rect -81360 80760 -81140 80810
rect -80860 80990 -80640 81040
rect -80860 80920 -80850 80990
rect -80650 80920 -80640 80990
rect -80860 80880 -80640 80920
rect -80860 80810 -80850 80880
rect -80650 80810 -80640 80880
rect -80860 80760 -80640 80810
rect -80360 80990 -80140 81040
rect -80360 80920 -80350 80990
rect -80150 80920 -80140 80990
rect -80360 80880 -80140 80920
rect -80360 80810 -80350 80880
rect -80150 80810 -80140 80880
rect -80360 80760 -80140 80810
rect -79860 80990 -79640 81040
rect -79860 80920 -79850 80990
rect -79650 80920 -79640 80990
rect -79860 80880 -79640 80920
rect -79860 80810 -79850 80880
rect -79650 80810 -79640 80880
rect -79860 80760 -79640 80810
rect -79360 80990 -79140 81040
rect -79360 80920 -79350 80990
rect -79150 80920 -79140 80990
rect -79360 80880 -79140 80920
rect -79360 80810 -79350 80880
rect -79150 80810 -79140 80880
rect -79360 80760 -79140 80810
rect -78860 80990 -78640 81040
rect -78860 80920 -78850 80990
rect -78650 80920 -78640 80990
rect -78860 80880 -78640 80920
rect -78860 80810 -78850 80880
rect -78650 80810 -78640 80880
rect -78860 80760 -78640 80810
rect -78360 80990 -78140 81040
rect -78360 80920 -78350 80990
rect -78150 80920 -78140 80990
rect -78360 80880 -78140 80920
rect -78360 80810 -78350 80880
rect -78150 80810 -78140 80880
rect -78360 80760 -78140 80810
rect -77860 80990 -77640 81040
rect -77860 80920 -77850 80990
rect -77650 80920 -77640 80990
rect -77860 80880 -77640 80920
rect -77860 80810 -77850 80880
rect -77650 80810 -77640 80880
rect -77860 80760 -77640 80810
rect -77360 80990 -77140 81040
rect -77360 80920 -77350 80990
rect -77150 80920 -77140 80990
rect -77360 80880 -77140 80920
rect -77360 80810 -77350 80880
rect -77150 80810 -77140 80880
rect -77360 80760 -77140 80810
rect -76860 80990 -76640 81040
rect -76860 80920 -76850 80990
rect -76650 80920 -76640 80990
rect -76860 80880 -76640 80920
rect -76860 80810 -76850 80880
rect -76650 80810 -76640 80880
rect -76860 80760 -76640 80810
rect -76360 80990 -76140 81040
rect -76360 80920 -76350 80990
rect -76150 80920 -76140 80990
rect -76360 80880 -76140 80920
rect -76360 80810 -76350 80880
rect -76150 80810 -76140 80880
rect -76360 80760 -76140 80810
rect -75860 80990 -75640 81040
rect -75860 80920 -75850 80990
rect -75650 80920 -75640 80990
rect -75860 80880 -75640 80920
rect -75860 80810 -75850 80880
rect -75650 80810 -75640 80880
rect -75860 80760 -75640 80810
rect -75360 80990 -75140 81040
rect -75360 80920 -75350 80990
rect -75150 80920 -75140 80990
rect -75360 80880 -75140 80920
rect -75360 80810 -75350 80880
rect -75150 80810 -75140 80880
rect -75360 80760 -75140 80810
rect -74860 80990 -74640 81040
rect -74860 80920 -74850 80990
rect -74650 80920 -74640 80990
rect -74860 80880 -74640 80920
rect -74860 80810 -74850 80880
rect -74650 80810 -74640 80880
rect -74860 80760 -74640 80810
rect -74360 80990 -74140 81040
rect -74360 80920 -74350 80990
rect -74150 80920 -74140 80990
rect -74360 80880 -74140 80920
rect -74360 80810 -74350 80880
rect -74150 80810 -74140 80880
rect -74360 80760 -74140 80810
rect -73860 80990 -73640 81040
rect -73860 80920 -73850 80990
rect -73650 80920 -73640 80990
rect -73860 80880 -73640 80920
rect -73860 80810 -73850 80880
rect -73650 80810 -73640 80880
rect -73860 80760 -73640 80810
rect -73360 80990 -73140 81040
rect -73360 80920 -73350 80990
rect -73150 80920 -73140 80990
rect -73360 80880 -73140 80920
rect -73360 80810 -73350 80880
rect -73150 80810 -73140 80880
rect -73360 80760 -73140 80810
rect -72860 80990 -72640 81040
rect -72860 80920 -72850 80990
rect -72650 80920 -72640 80990
rect -72860 80880 -72640 80920
rect -72860 80810 -72850 80880
rect -72650 80810 -72640 80880
rect -72860 80760 -72640 80810
rect -72360 80990 -72140 81040
rect -72360 80920 -72350 80990
rect -72150 80920 -72140 80990
rect -72360 80880 -72140 80920
rect -72360 80810 -72350 80880
rect -72150 80810 -72140 80880
rect -72360 80760 -72140 80810
rect -71860 80990 -71640 81040
rect -71860 80920 -71850 80990
rect -71650 80920 -71640 80990
rect -71860 80880 -71640 80920
rect -71860 80810 -71850 80880
rect -71650 80810 -71640 80880
rect -71860 80760 -71640 80810
rect -71360 80990 -71140 81040
rect -71360 80920 -71350 80990
rect -71150 80920 -71140 80990
rect -71360 80880 -71140 80920
rect -71360 80810 -71350 80880
rect -71150 80810 -71140 80880
rect -71360 80760 -71140 80810
rect -70860 80990 -70640 81040
rect -70860 80920 -70850 80990
rect -70650 80920 -70640 80990
rect -70860 80880 -70640 80920
rect -70860 80810 -70850 80880
rect -70650 80810 -70640 80880
rect -70860 80760 -70640 80810
rect -70360 80990 -70140 81040
rect -70360 80920 -70350 80990
rect -70150 80920 -70140 80990
rect -70360 80880 -70140 80920
rect -70360 80810 -70350 80880
rect -70150 80810 -70140 80880
rect -70360 80760 -70140 80810
rect -69860 80990 -69640 81040
rect -69860 80920 -69850 80990
rect -69650 80920 -69640 80990
rect -69860 80880 -69640 80920
rect -69860 80810 -69850 80880
rect -69650 80810 -69640 80880
rect -69860 80760 -69640 80810
rect -69360 80990 -69140 81040
rect -69360 80920 -69350 80990
rect -69150 80920 -69140 80990
rect -69360 80880 -69140 80920
rect -69360 80810 -69350 80880
rect -69150 80810 -69140 80880
rect -69360 80760 -69140 80810
rect -68860 80990 -68640 81040
rect -68860 80920 -68850 80990
rect -68650 80920 -68640 80990
rect -68860 80880 -68640 80920
rect -68860 80810 -68850 80880
rect -68650 80810 -68640 80880
rect -68860 80760 -68640 80810
rect -68360 80990 -68140 81040
rect -68360 80920 -68350 80990
rect -68150 80920 -68140 80990
rect -68360 80880 -68140 80920
rect -68360 80810 -68350 80880
rect -68150 80810 -68140 80880
rect -68360 80760 -68140 80810
rect -67860 80990 -67640 81040
rect -67860 80920 -67850 80990
rect -67650 80920 -67640 80990
rect -67860 80880 -67640 80920
rect -67860 80810 -67850 80880
rect -67650 80810 -67640 80880
rect -67860 80760 -67640 80810
rect -67360 80990 -67140 81040
rect -67360 80920 -67350 80990
rect -67150 80920 -67140 80990
rect -67360 80880 -67140 80920
rect -67360 80810 -67350 80880
rect -67150 80810 -67140 80880
rect -67360 80760 -67140 80810
rect -66860 80990 -66640 81040
rect -66860 80920 -66850 80990
rect -66650 80920 -66640 80990
rect -66860 80880 -66640 80920
rect -66860 80810 -66850 80880
rect -66650 80810 -66640 80880
rect -66860 80760 -66640 80810
rect -66360 80990 -66140 81040
rect -66360 80920 -66350 80990
rect -66150 80920 -66140 80990
rect -66360 80880 -66140 80920
rect -66360 80810 -66350 80880
rect -66150 80810 -66140 80880
rect -66360 80760 -66140 80810
rect -65860 80990 -65640 81040
rect -65860 80920 -65850 80990
rect -65650 80920 -65640 80990
rect -65860 80880 -65640 80920
rect -65860 80810 -65850 80880
rect -65650 80810 -65640 80880
rect -65860 80760 -65640 80810
rect -65360 80990 -65140 81040
rect -65360 80920 -65350 80990
rect -65150 80920 -65140 80990
rect -65360 80880 -65140 80920
rect -65360 80810 -65350 80880
rect -65150 80810 -65140 80880
rect -65360 80760 -65140 80810
rect -64860 80990 -64640 81040
rect -64860 80920 -64850 80990
rect -64650 80920 -64640 80990
rect -64860 80880 -64640 80920
rect -64860 80810 -64850 80880
rect -64650 80810 -64640 80880
rect -64860 80760 -64640 80810
rect -64360 80990 -64140 81040
rect -64360 80920 -64350 80990
rect -64150 80920 -64140 80990
rect -64360 80880 -64140 80920
rect -64360 80810 -64350 80880
rect -64150 80810 -64140 80880
rect -64360 80760 -64140 80810
rect -63860 80990 -63640 81040
rect -63860 80920 -63850 80990
rect -63650 80920 -63640 80990
rect -63860 80880 -63640 80920
rect -63860 80810 -63850 80880
rect -63650 80810 -63640 80880
rect -63860 80760 -63640 80810
rect -63360 80990 -63140 81040
rect -63360 80920 -63350 80990
rect -63150 80920 -63140 80990
rect -63360 80880 -63140 80920
rect -63360 80810 -63350 80880
rect -63150 80810 -63140 80880
rect -63360 80760 -63140 80810
rect -62860 80990 -62640 81040
rect -62860 80920 -62850 80990
rect -62650 80920 -62640 80990
rect -62860 80880 -62640 80920
rect -62860 80810 -62850 80880
rect -62650 80810 -62640 80880
rect -62860 80760 -62640 80810
rect -62360 80990 -62140 81040
rect -62360 80920 -62350 80990
rect -62150 80920 -62140 80990
rect -62360 80880 -62140 80920
rect -62360 80810 -62350 80880
rect -62150 80810 -62140 80880
rect -62360 80760 -62140 80810
rect -61860 80990 -61640 81040
rect -61860 80920 -61850 80990
rect -61650 80920 -61640 80990
rect -61860 80880 -61640 80920
rect -61860 80810 -61850 80880
rect -61650 80810 -61640 80880
rect -61860 80760 -61640 80810
rect -61360 80990 -61140 81040
rect -61360 80920 -61350 80990
rect -61150 80920 -61140 80990
rect -61360 80880 -61140 80920
rect -61360 80810 -61350 80880
rect -61150 80810 -61140 80880
rect -61360 80760 -61140 80810
rect -60860 80990 -60640 81040
rect -60860 80920 -60850 80990
rect -60650 80920 -60640 80990
rect -60860 80880 -60640 80920
rect -60860 80810 -60850 80880
rect -60650 80810 -60640 80880
rect -60860 80760 -60640 80810
rect -60360 80990 -60140 81040
rect -60360 80920 -60350 80990
rect -60150 80920 -60140 80990
rect -60360 80880 -60140 80920
rect -60360 80810 -60350 80880
rect -60150 80810 -60140 80880
rect -60360 80760 -60140 80810
rect -59860 80990 -59640 81040
rect -59860 80920 -59850 80990
rect -59650 80920 -59640 80990
rect -59860 80880 -59640 80920
rect -59860 80810 -59850 80880
rect -59650 80810 -59640 80880
rect -59860 80760 -59640 80810
rect -59360 80990 -59140 81040
rect -59360 80920 -59350 80990
rect -59150 80920 -59140 80990
rect -59360 80880 -59140 80920
rect -59360 80810 -59350 80880
rect -59150 80810 -59140 80880
rect -59360 80760 -59140 80810
rect -58860 80990 -58640 81040
rect -58860 80920 -58850 80990
rect -58650 80920 -58640 80990
rect -58860 80880 -58640 80920
rect -58860 80810 -58850 80880
rect -58650 80810 -58640 80880
rect -58860 80760 -58640 80810
rect -58360 80990 -58140 81040
rect -58360 80920 -58350 80990
rect -58150 80920 -58140 80990
rect -58360 80880 -58140 80920
rect -58360 80810 -58350 80880
rect -58150 80810 -58140 80880
rect -58360 80760 -58140 80810
rect -57860 80990 -57640 81040
rect -57860 80920 -57850 80990
rect -57650 80920 -57640 80990
rect -57860 80880 -57640 80920
rect -57860 80810 -57850 80880
rect -57650 80810 -57640 80880
rect -57860 80760 -57640 80810
rect -57360 80990 -57140 81040
rect -57360 80920 -57350 80990
rect -57150 80920 -57140 80990
rect -57360 80880 -57140 80920
rect -57360 80810 -57350 80880
rect -57150 80810 -57140 80880
rect -57360 80760 -57140 80810
rect -56860 80990 -56640 81040
rect -56860 80920 -56850 80990
rect -56650 80920 -56640 80990
rect -56860 80880 -56640 80920
rect -56860 80810 -56850 80880
rect -56650 80810 -56640 80880
rect -56860 80760 -56640 80810
rect -56360 80990 -56140 81040
rect -56360 80920 -56350 80990
rect -56150 80920 -56140 80990
rect -56360 80880 -56140 80920
rect -56360 80810 -56350 80880
rect -56150 80810 -56140 80880
rect -56360 80760 -56140 80810
rect -55860 80990 -55640 81040
rect -55860 80920 -55850 80990
rect -55650 80920 -55640 80990
rect -55860 80880 -55640 80920
rect -55860 80810 -55850 80880
rect -55650 80810 -55640 80880
rect -55860 80760 -55640 80810
rect -55360 80990 -55140 81040
rect -55360 80920 -55350 80990
rect -55150 80920 -55140 80990
rect -55360 80880 -55140 80920
rect -55360 80810 -55350 80880
rect -55150 80810 -55140 80880
rect -55360 80760 -55140 80810
rect -54860 80990 -54640 81040
rect -54860 80920 -54850 80990
rect -54650 80920 -54640 80990
rect -54860 80880 -54640 80920
rect -54860 80810 -54850 80880
rect -54650 80810 -54640 80880
rect -54860 80760 -54640 80810
rect -54360 80990 -54140 81040
rect -54360 80920 -54350 80990
rect -54150 80920 -54140 80990
rect -54360 80880 -54140 80920
rect -54360 80810 -54350 80880
rect -54150 80810 -54140 80880
rect -54360 80760 -54140 80810
rect -53860 80990 -53640 81040
rect -53860 80920 -53850 80990
rect -53650 80920 -53640 80990
rect -53860 80880 -53640 80920
rect -53860 80810 -53850 80880
rect -53650 80810 -53640 80880
rect -53860 80760 -53640 80810
rect -53360 80990 -53140 81040
rect -53360 80920 -53350 80990
rect -53150 80920 -53140 80990
rect -53360 80880 -53140 80920
rect -53360 80810 -53350 80880
rect -53150 80810 -53140 80880
rect -53360 80760 -53140 80810
rect -52860 80990 -52640 81040
rect -52860 80920 -52850 80990
rect -52650 80920 -52640 80990
rect -52860 80880 -52640 80920
rect -52860 80810 -52850 80880
rect -52650 80810 -52640 80880
rect -52860 80760 -52640 80810
rect -52360 80990 -52140 81040
rect -52360 80920 -52350 80990
rect -52150 80920 -52140 80990
rect -52360 80880 -52140 80920
rect -52360 80810 -52350 80880
rect -52150 80810 -52140 80880
rect -52360 80760 -52140 80810
rect -51860 80990 -51640 81040
rect -51860 80920 -51850 80990
rect -51650 80920 -51640 80990
rect -51860 80880 -51640 80920
rect -51860 80810 -51850 80880
rect -51650 80810 -51640 80880
rect -51860 80760 -51640 80810
rect -51360 80990 -51140 81040
rect -51360 80920 -51350 80990
rect -51150 80920 -51140 80990
rect -51360 80880 -51140 80920
rect -51360 80810 -51350 80880
rect -51150 80810 -51140 80880
rect -51360 80760 -51140 80810
rect -50860 80990 -50640 81040
rect -50860 80920 -50850 80990
rect -50650 80920 -50640 80990
rect -50860 80880 -50640 80920
rect -50860 80810 -50850 80880
rect -50650 80810 -50640 80880
rect -50860 80760 -50640 80810
rect -50360 80990 -50140 81040
rect -50360 80920 -50350 80990
rect -50150 80920 -50140 80990
rect -50360 80880 -50140 80920
rect -50360 80810 -50350 80880
rect -50150 80810 -50140 80880
rect -50360 80760 -50140 80810
rect -49860 80990 -49640 81040
rect -49860 80920 -49850 80990
rect -49650 80920 -49640 80990
rect -49860 80880 -49640 80920
rect -49860 80810 -49850 80880
rect -49650 80810 -49640 80880
rect -49860 80760 -49640 80810
rect -49360 80990 -49140 81040
rect -49360 80920 -49350 80990
rect -49150 80920 -49140 80990
rect -49360 80880 -49140 80920
rect -49360 80810 -49350 80880
rect -49150 80810 -49140 80880
rect -49360 80760 -49140 80810
rect -48860 80990 -48640 81040
rect -48860 80920 -48850 80990
rect -48650 80920 -48640 80990
rect -48860 80880 -48640 80920
rect -48860 80810 -48850 80880
rect -48650 80810 -48640 80880
rect -48860 80760 -48640 80810
rect -48360 80990 -48140 81040
rect -48360 80920 -48350 80990
rect -48150 80920 -48140 80990
rect -48360 80880 -48140 80920
rect -48360 80810 -48350 80880
rect -48150 80810 -48140 80880
rect -48360 80760 -48140 80810
rect -47860 80990 -47640 81040
rect -47860 80920 -47850 80990
rect -47650 80920 -47640 80990
rect -47860 80880 -47640 80920
rect -47860 80810 -47850 80880
rect -47650 80810 -47640 80880
rect -47860 80760 -47640 80810
rect -47360 80990 -47140 81040
rect -47360 80920 -47350 80990
rect -47150 80920 -47140 80990
rect -47360 80880 -47140 80920
rect -47360 80810 -47350 80880
rect -47150 80810 -47140 80880
rect -47360 80760 -47140 80810
rect -46860 80990 -46640 81040
rect -46860 80920 -46850 80990
rect -46650 80920 -46640 80990
rect -46860 80880 -46640 80920
rect -46860 80810 -46850 80880
rect -46650 80810 -46640 80880
rect -46860 80760 -46640 80810
rect -46360 80990 -46140 81040
rect -46360 80920 -46350 80990
rect -46150 80920 -46140 80990
rect -46360 80880 -46140 80920
rect -46360 80810 -46350 80880
rect -46150 80810 -46140 80880
rect -46360 80760 -46140 80810
rect -45860 80990 -45640 81040
rect -45860 80920 -45850 80990
rect -45650 80920 -45640 80990
rect -45860 80880 -45640 80920
rect -45860 80810 -45850 80880
rect -45650 80810 -45640 80880
rect -45860 80760 -45640 80810
rect -45360 80990 -45140 81040
rect -45360 80920 -45350 80990
rect -45150 80920 -45140 80990
rect -45360 80880 -45140 80920
rect -45360 80810 -45350 80880
rect -45150 80810 -45140 80880
rect -45360 80760 -45140 80810
rect -44860 80990 -44640 81040
rect -44860 80920 -44850 80990
rect -44650 80920 -44640 80990
rect -44860 80880 -44640 80920
rect -44860 80810 -44850 80880
rect -44650 80810 -44640 80880
rect -44860 80760 -44640 80810
rect -44360 80990 -44140 81040
rect -44360 80920 -44350 80990
rect -44150 80920 -44140 80990
rect -44360 80880 -44140 80920
rect -44360 80810 -44350 80880
rect -44150 80810 -44140 80880
rect -44360 80760 -44140 80810
rect -43860 80990 -43640 81040
rect -43860 80920 -43850 80990
rect -43650 80920 -43640 80990
rect -43860 80880 -43640 80920
rect -43860 80810 -43850 80880
rect -43650 80810 -43640 80880
rect -43860 80760 -43640 80810
rect -43360 80990 -43140 81040
rect -43360 80920 -43350 80990
rect -43150 80920 -43140 80990
rect -43360 80880 -43140 80920
rect -43360 80810 -43350 80880
rect -43150 80810 -43140 80880
rect -43360 80760 -43140 80810
rect -42860 80990 -42640 81040
rect -42860 80920 -42850 80990
rect -42650 80920 -42640 80990
rect -42860 80880 -42640 80920
rect -42860 80810 -42850 80880
rect -42650 80810 -42640 80880
rect -42860 80760 -42640 80810
rect -42360 80990 -42140 81040
rect -42360 80920 -42350 80990
rect -42150 80920 -42140 80990
rect -42360 80880 -42140 80920
rect -42360 80810 -42350 80880
rect -42150 80810 -42140 80880
rect -42360 80760 -42140 80810
rect -41860 80990 -41640 81040
rect -41860 80920 -41850 80990
rect -41650 80920 -41640 80990
rect -41860 80880 -41640 80920
rect -41860 80810 -41850 80880
rect -41650 80810 -41640 80880
rect -41860 80760 -41640 80810
rect -41360 80990 -41140 81040
rect -41360 80920 -41350 80990
rect -41150 80920 -41140 80990
rect -41360 80880 -41140 80920
rect -41360 80810 -41350 80880
rect -41150 80810 -41140 80880
rect -41360 80760 -41140 80810
rect -40860 80990 -40640 81040
rect -40860 80920 -40850 80990
rect -40650 80920 -40640 80990
rect -40860 80880 -40640 80920
rect -40860 80810 -40850 80880
rect -40650 80810 -40640 80880
rect -40860 80760 -40640 80810
rect -40360 80990 -40140 81040
rect -40360 80920 -40350 80990
rect -40150 80920 -40140 80990
rect -40360 80880 -40140 80920
rect -40360 80810 -40350 80880
rect -40150 80810 -40140 80880
rect -40360 80760 -40140 80810
rect -39860 80990 -39640 81040
rect -39860 80920 -39850 80990
rect -39650 80920 -39640 80990
rect -39860 80880 -39640 80920
rect -39860 80810 -39850 80880
rect -39650 80810 -39640 80880
rect -39860 80760 -39640 80810
rect -39360 80990 -39140 81040
rect -39360 80920 -39350 80990
rect -39150 80920 -39140 80990
rect -39360 80880 -39140 80920
rect -39360 80810 -39350 80880
rect -39150 80810 -39140 80880
rect -39360 80760 -39140 80810
rect -38860 80990 -38640 81040
rect -38860 80920 -38850 80990
rect -38650 80920 -38640 80990
rect -38860 80880 -38640 80920
rect -38860 80810 -38850 80880
rect -38650 80810 -38640 80880
rect -38860 80760 -38640 80810
rect -38360 80990 -38140 81040
rect -38360 80920 -38350 80990
rect -38150 80920 -38140 80990
rect -38360 80880 -38140 80920
rect -38360 80810 -38350 80880
rect -38150 80810 -38140 80880
rect -38360 80760 -38140 80810
rect -37860 80990 -37640 81040
rect -37860 80920 -37850 80990
rect -37650 80920 -37640 80990
rect -37860 80880 -37640 80920
rect -37860 80810 -37850 80880
rect -37650 80810 -37640 80880
rect -37860 80760 -37640 80810
rect -37360 80990 -37140 81040
rect -37360 80920 -37350 80990
rect -37150 80920 -37140 80990
rect -37360 80880 -37140 80920
rect -37360 80810 -37350 80880
rect -37150 80810 -37140 80880
rect -37360 80760 -37140 80810
rect -36860 80990 -36640 81040
rect -36860 80920 -36850 80990
rect -36650 80920 -36640 80990
rect -36860 80880 -36640 80920
rect -36860 80810 -36850 80880
rect -36650 80810 -36640 80880
rect -36860 80760 -36640 80810
rect -36360 80990 -36140 81040
rect -36360 80920 -36350 80990
rect -36150 80920 -36140 80990
rect -36360 80880 -36140 80920
rect -36360 80810 -36350 80880
rect -36150 80810 -36140 80880
rect -36360 80760 -36140 80810
rect -35860 80990 -35640 81040
rect -35860 80920 -35850 80990
rect -35650 80920 -35640 80990
rect -35860 80880 -35640 80920
rect -35860 80810 -35850 80880
rect -35650 80810 -35640 80880
rect -35860 80760 -35640 80810
rect -35360 80990 -35140 81040
rect -35360 80920 -35350 80990
rect -35150 80920 -35140 80990
rect -35360 80880 -35140 80920
rect -35360 80810 -35350 80880
rect -35150 80810 -35140 80880
rect -35360 80760 -35140 80810
rect -34860 80990 -34640 81040
rect -34860 80920 -34850 80990
rect -34650 80920 -34640 80990
rect -34860 80880 -34640 80920
rect -34860 80810 -34850 80880
rect -34650 80810 -34640 80880
rect -34860 80760 -34640 80810
rect -34360 80990 -34140 81040
rect -34360 80920 -34350 80990
rect -34150 80920 -34140 80990
rect -34360 80880 -34140 80920
rect -34360 80810 -34350 80880
rect -34150 80810 -34140 80880
rect -34360 80760 -34140 80810
rect -33860 80990 -33640 81040
rect -33860 80920 -33850 80990
rect -33650 80920 -33640 80990
rect -33860 80880 -33640 80920
rect -33860 80810 -33850 80880
rect -33650 80810 -33640 80880
rect -33860 80760 -33640 80810
rect -33360 80990 -33140 81040
rect -33360 80920 -33350 80990
rect -33150 80920 -33140 80990
rect -33360 80880 -33140 80920
rect -33360 80810 -33350 80880
rect -33150 80810 -33140 80880
rect -33360 80760 -33140 80810
rect -32860 80990 -32640 81040
rect -32860 80920 -32850 80990
rect -32650 80920 -32640 80990
rect -32860 80880 -32640 80920
rect -32860 80810 -32850 80880
rect -32650 80810 -32640 80880
rect -32860 80760 -32640 80810
rect -32360 80990 -32140 81040
rect -32360 80920 -32350 80990
rect -32150 80920 -32140 80990
rect -32360 80880 -32140 80920
rect -32360 80810 -32350 80880
rect -32150 80810 -32140 80880
rect -32360 80760 -32140 80810
rect -31860 80990 -31640 81040
rect -31860 80920 -31850 80990
rect -31650 80920 -31640 80990
rect -31860 80880 -31640 80920
rect -31860 80810 -31850 80880
rect -31650 80810 -31640 80880
rect -31860 80760 -31640 80810
rect -31360 80990 -31140 81040
rect -31360 80920 -31350 80990
rect -31150 80920 -31140 80990
rect -31360 80880 -31140 80920
rect -31360 80810 -31350 80880
rect -31150 80810 -31140 80880
rect -31360 80760 -31140 80810
rect -30860 80990 -30640 81040
rect -30860 80920 -30850 80990
rect -30650 80920 -30640 80990
rect -30860 80880 -30640 80920
rect -30860 80810 -30850 80880
rect -30650 80810 -30640 80880
rect -30860 80760 -30640 80810
rect -30360 80990 -30140 81040
rect -30360 80920 -30350 80990
rect -30150 80920 -30140 80990
rect -30360 80880 -30140 80920
rect -30360 80810 -30350 80880
rect -30150 80810 -30140 80880
rect -30360 80760 -30140 80810
rect -29860 80990 -29640 81040
rect -29860 80920 -29850 80990
rect -29650 80920 -29640 80990
rect -29860 80880 -29640 80920
rect -29860 80810 -29850 80880
rect -29650 80810 -29640 80880
rect -29860 80760 -29640 80810
rect -29360 80990 -29140 81040
rect -29360 80920 -29350 80990
rect -29150 80920 -29140 80990
rect -29360 80880 -29140 80920
rect -29360 80810 -29350 80880
rect -29150 80810 -29140 80880
rect -29360 80760 -29140 80810
rect -28860 80990 -28640 81040
rect -28860 80920 -28850 80990
rect -28650 80920 -28640 80990
rect -28860 80880 -28640 80920
rect -28860 80810 -28850 80880
rect -28650 80810 -28640 80880
rect -28860 80760 -28640 80810
rect -28360 80990 -28140 81040
rect -28360 80920 -28350 80990
rect -28150 80920 -28140 80990
rect -28360 80880 -28140 80920
rect -28360 80810 -28350 80880
rect -28150 80810 -28140 80880
rect -28360 80760 -28140 80810
rect -27860 80990 -27640 81040
rect -27860 80920 -27850 80990
rect -27650 80920 -27640 80990
rect -27860 80880 -27640 80920
rect -27860 80810 -27850 80880
rect -27650 80810 -27640 80880
rect -27860 80760 -27640 80810
rect -27360 80990 -27140 81040
rect -27360 80920 -27350 80990
rect -27150 80920 -27140 80990
rect -27360 80880 -27140 80920
rect -27360 80810 -27350 80880
rect -27150 80810 -27140 80880
rect -27360 80760 -27140 80810
rect -26860 80990 -26640 81040
rect -26860 80920 -26850 80990
rect -26650 80920 -26640 80990
rect -26860 80880 -26640 80920
rect -26860 80810 -26850 80880
rect -26650 80810 -26640 80880
rect -26860 80760 -26640 80810
rect -26360 80990 -26140 81040
rect -26360 80920 -26350 80990
rect -26150 80920 -26140 80990
rect -26360 80880 -26140 80920
rect -26360 80810 -26350 80880
rect -26150 80810 -26140 80880
rect -26360 80760 -26140 80810
rect -25860 80990 -25640 81040
rect -25860 80920 -25850 80990
rect -25650 80920 -25640 80990
rect -25860 80880 -25640 80920
rect -25860 80810 -25850 80880
rect -25650 80810 -25640 80880
rect -25860 80760 -25640 80810
rect -25360 80990 -25140 81040
rect -25360 80920 -25350 80990
rect -25150 80920 -25140 80990
rect -25360 80880 -25140 80920
rect -25360 80810 -25350 80880
rect -25150 80810 -25140 80880
rect -25360 80760 -25140 80810
rect -24860 80990 -24640 81040
rect -24860 80920 -24850 80990
rect -24650 80920 -24640 80990
rect -24860 80880 -24640 80920
rect -24860 80810 -24850 80880
rect -24650 80810 -24640 80880
rect -24860 80760 -24640 80810
rect -24360 80990 -24140 81040
rect -24360 80920 -24350 80990
rect -24150 80920 -24140 80990
rect -24360 80880 -24140 80920
rect -24360 80810 -24350 80880
rect -24150 80810 -24140 80880
rect -24360 80760 -24140 80810
rect -23860 80990 -23640 81040
rect -23860 80920 -23850 80990
rect -23650 80920 -23640 80990
rect -23860 80880 -23640 80920
rect -23860 80810 -23850 80880
rect -23650 80810 -23640 80880
rect -23860 80760 -23640 80810
rect -23360 80990 -23140 81040
rect -23360 80920 -23350 80990
rect -23150 80920 -23140 80990
rect -23360 80880 -23140 80920
rect -23360 80810 -23350 80880
rect -23150 80810 -23140 80880
rect -23360 80760 -23140 80810
rect -22860 80990 -22640 81040
rect -22860 80920 -22850 80990
rect -22650 80920 -22640 80990
rect -22860 80880 -22640 80920
rect -22860 80810 -22850 80880
rect -22650 80810 -22640 80880
rect -22860 80760 -22640 80810
rect -22360 80990 -22140 81040
rect -22360 80920 -22350 80990
rect -22150 80920 -22140 80990
rect -22360 80880 -22140 80920
rect -22360 80810 -22350 80880
rect -22150 80810 -22140 80880
rect -22360 80760 -22140 80810
rect -21860 80990 -21640 81040
rect -21860 80920 -21850 80990
rect -21650 80920 -21640 80990
rect -21860 80880 -21640 80920
rect -21860 80810 -21850 80880
rect -21650 80810 -21640 80880
rect -21860 80760 -21640 80810
rect -21360 80990 -21140 81040
rect -21360 80920 -21350 80990
rect -21150 80920 -21140 80990
rect -21360 80880 -21140 80920
rect -21360 80810 -21350 80880
rect -21150 80810 -21140 80880
rect -21360 80760 -21140 80810
rect -20860 80990 -20640 81040
rect -20860 80920 -20850 80990
rect -20650 80920 -20640 80990
rect -20860 80880 -20640 80920
rect -20860 80810 -20850 80880
rect -20650 80810 -20640 80880
rect -20860 80760 -20640 80810
rect -20360 80990 -20140 81040
rect -20360 80920 -20350 80990
rect -20150 80920 -20140 80990
rect -20360 80880 -20140 80920
rect -20360 80810 -20350 80880
rect -20150 80810 -20140 80880
rect -20360 80760 -20140 80810
rect -19860 80990 -19640 81040
rect -19860 80920 -19850 80990
rect -19650 80920 -19640 80990
rect -19860 80880 -19640 80920
rect -19860 80810 -19850 80880
rect -19650 80810 -19640 80880
rect -19860 80760 -19640 80810
rect -19360 80990 -19140 81040
rect -19360 80920 -19350 80990
rect -19150 80920 -19140 80990
rect -19360 80880 -19140 80920
rect -19360 80810 -19350 80880
rect -19150 80810 -19140 80880
rect -19360 80760 -19140 80810
rect -18860 80990 -18640 81040
rect -18860 80920 -18850 80990
rect -18650 80920 -18640 80990
rect -18860 80880 -18640 80920
rect -18860 80810 -18850 80880
rect -18650 80810 -18640 80880
rect -18860 80760 -18640 80810
rect -18360 80990 -18140 81040
rect -18360 80920 -18350 80990
rect -18150 80920 -18140 80990
rect -18360 80880 -18140 80920
rect -18360 80810 -18350 80880
rect -18150 80810 -18140 80880
rect -18360 80760 -18140 80810
rect -17860 80990 -17640 81040
rect -17860 80920 -17850 80990
rect -17650 80920 -17640 80990
rect -17860 80880 -17640 80920
rect -17860 80810 -17850 80880
rect -17650 80810 -17640 80880
rect -17860 80760 -17640 80810
rect -17360 80990 -17140 81040
rect -17360 80920 -17350 80990
rect -17150 80920 -17140 80990
rect -17360 80880 -17140 80920
rect -17360 80810 -17350 80880
rect -17150 80810 -17140 80880
rect -17360 80760 -17140 80810
rect -16860 80990 -16640 81040
rect -16860 80920 -16850 80990
rect -16650 80920 -16640 80990
rect -16860 80880 -16640 80920
rect -16860 80810 -16850 80880
rect -16650 80810 -16640 80880
rect -16860 80760 -16640 80810
rect -16360 80990 -16140 81040
rect -16360 80920 -16350 80990
rect -16150 80920 -16140 80990
rect -16360 80880 -16140 80920
rect -16360 80810 -16350 80880
rect -16150 80810 -16140 80880
rect -16360 80760 -16140 80810
rect -15860 80990 -15640 81040
rect -15860 80920 -15850 80990
rect -15650 80920 -15640 80990
rect -15860 80880 -15640 80920
rect -15860 80810 -15850 80880
rect -15650 80810 -15640 80880
rect -15860 80760 -15640 80810
rect -15360 80990 -15140 81040
rect -15360 80920 -15350 80990
rect -15150 80920 -15140 80990
rect -15360 80880 -15140 80920
rect -15360 80810 -15350 80880
rect -15150 80810 -15140 80880
rect -15360 80760 -15140 80810
rect -14860 80990 -14640 81040
rect -14860 80920 -14850 80990
rect -14650 80920 -14640 80990
rect -14860 80880 -14640 80920
rect -14860 80810 -14850 80880
rect -14650 80810 -14640 80880
rect -14860 80760 -14640 80810
rect -14360 80990 -14140 81040
rect -14360 80920 -14350 80990
rect -14150 80920 -14140 80990
rect -14360 80880 -14140 80920
rect -14360 80810 -14350 80880
rect -14150 80810 -14140 80880
rect -14360 80760 -14140 80810
rect -13860 80990 -13640 81040
rect -13860 80920 -13850 80990
rect -13650 80920 -13640 80990
rect -13860 80880 -13640 80920
rect -13860 80810 -13850 80880
rect -13650 80810 -13640 80880
rect -13860 80760 -13640 80810
rect -13360 80990 -13140 81040
rect -13360 80920 -13350 80990
rect -13150 80920 -13140 80990
rect -13360 80880 -13140 80920
rect -13360 80810 -13350 80880
rect -13150 80810 -13140 80880
rect -13360 80760 -13140 80810
rect -12860 80990 -12640 81040
rect -12860 80920 -12850 80990
rect -12650 80920 -12640 80990
rect -12860 80880 -12640 80920
rect -12860 80810 -12850 80880
rect -12650 80810 -12640 80880
rect -12860 80760 -12640 80810
rect -12360 80990 -12140 81040
rect -12360 80920 -12350 80990
rect -12150 80920 -12140 80990
rect -12360 80880 -12140 80920
rect -12360 80810 -12350 80880
rect -12150 80810 -12140 80880
rect -12360 80760 -12140 80810
rect -11860 80990 -11640 81040
rect -11860 80920 -11850 80990
rect -11650 80920 -11640 80990
rect -11860 80880 -11640 80920
rect -11860 80810 -11850 80880
rect -11650 80810 -11640 80880
rect -11860 80760 -11640 80810
rect -11360 80990 -11140 81040
rect -11360 80920 -11350 80990
rect -11150 80920 -11140 80990
rect -11360 80880 -11140 80920
rect -11360 80810 -11350 80880
rect -11150 80810 -11140 80880
rect -11360 80760 -11140 80810
rect -10860 80990 -10640 81040
rect -10860 80920 -10850 80990
rect -10650 80920 -10640 80990
rect -10860 80880 -10640 80920
rect -10860 80810 -10850 80880
rect -10650 80810 -10640 80880
rect -10860 80760 -10640 80810
rect -10360 80990 -10140 81040
rect -10360 80920 -10350 80990
rect -10150 80920 -10140 80990
rect -10360 80880 -10140 80920
rect -10360 80810 -10350 80880
rect -10150 80810 -10140 80880
rect -10360 80760 -10140 80810
rect -9860 80990 -9640 81040
rect -9860 80920 -9850 80990
rect -9650 80920 -9640 80990
rect -9860 80880 -9640 80920
rect -9860 80810 -9850 80880
rect -9650 80810 -9640 80880
rect -9860 80760 -9640 80810
rect -9360 80990 -9140 81040
rect -9360 80920 -9350 80990
rect -9150 80920 -9140 80990
rect -9360 80880 -9140 80920
rect -9360 80810 -9350 80880
rect -9150 80810 -9140 80880
rect -9360 80760 -9140 80810
rect -8860 80990 -8640 81040
rect -8860 80920 -8850 80990
rect -8650 80920 -8640 80990
rect -8860 80880 -8640 80920
rect -8860 80810 -8850 80880
rect -8650 80810 -8640 80880
rect -8860 80760 -8640 80810
rect -8360 80990 -8140 81040
rect -8360 80920 -8350 80990
rect -8150 80920 -8140 80990
rect -8360 80880 -8140 80920
rect -8360 80810 -8350 80880
rect -8150 80810 -8140 80880
rect -8360 80760 -8140 80810
rect -7860 80990 -7640 81040
rect -7860 80920 -7850 80990
rect -7650 80920 -7640 80990
rect -7860 80880 -7640 80920
rect -7860 80810 -7850 80880
rect -7650 80810 -7640 80880
rect -7860 80760 -7640 80810
rect -7360 80990 -7140 81040
rect -7360 80920 -7350 80990
rect -7150 80920 -7140 80990
rect -7360 80880 -7140 80920
rect -7360 80810 -7350 80880
rect -7150 80810 -7140 80880
rect -7360 80760 -7140 80810
rect -6860 80990 -6640 81040
rect -6860 80920 -6850 80990
rect -6650 80920 -6640 80990
rect -6860 80880 -6640 80920
rect -6860 80810 -6850 80880
rect -6650 80810 -6640 80880
rect -6860 80760 -6640 80810
rect -6360 80990 -6140 81040
rect -6360 80920 -6350 80990
rect -6150 80920 -6140 80990
rect -6360 80880 -6140 80920
rect -6360 80810 -6350 80880
rect -6150 80810 -6140 80880
rect -6360 80760 -6140 80810
rect -5860 80990 -5640 81040
rect -5860 80920 -5850 80990
rect -5650 80920 -5640 80990
rect -5860 80880 -5640 80920
rect -5860 80810 -5850 80880
rect -5650 80810 -5640 80880
rect -5860 80760 -5640 80810
rect -5360 80990 -5140 81040
rect -5360 80920 -5350 80990
rect -5150 80920 -5140 80990
rect -5360 80880 -5140 80920
rect -5360 80810 -5350 80880
rect -5150 80810 -5140 80880
rect -5360 80760 -5140 80810
rect -4860 80990 -4640 81040
rect -4860 80920 -4850 80990
rect -4650 80920 -4640 80990
rect -4860 80880 -4640 80920
rect -4860 80810 -4850 80880
rect -4650 80810 -4640 80880
rect -4860 80760 -4640 80810
rect -4360 80990 -4140 81040
rect -4360 80920 -4350 80990
rect -4150 80920 -4140 80990
rect -4360 80880 -4140 80920
rect -4360 80810 -4350 80880
rect -4150 80810 -4140 80880
rect -4360 80760 -4140 80810
rect -3860 80990 -3640 81040
rect -3860 80920 -3850 80990
rect -3650 80920 -3640 80990
rect -3860 80880 -3640 80920
rect -3860 80810 -3850 80880
rect -3650 80810 -3640 80880
rect -3860 80760 -3640 80810
rect -3360 80990 -3140 81040
rect -3360 80920 -3350 80990
rect -3150 80920 -3140 80990
rect -3360 80880 -3140 80920
rect -3360 80810 -3350 80880
rect -3150 80810 -3140 80880
rect -3360 80760 -3140 80810
rect -2860 80990 -2640 81040
rect -2860 80920 -2850 80990
rect -2650 80920 -2640 80990
rect -2860 80880 -2640 80920
rect -2860 80810 -2850 80880
rect -2650 80810 -2640 80880
rect -2860 80760 -2640 80810
rect -2360 80990 -2140 81040
rect -2360 80920 -2350 80990
rect -2150 80920 -2140 80990
rect -2360 80880 -2140 80920
rect -2360 80810 -2350 80880
rect -2150 80810 -2140 80880
rect -2360 80760 -2140 80810
rect -1860 80990 -1640 81040
rect -1860 80920 -1850 80990
rect -1650 80920 -1640 80990
rect -1860 80880 -1640 80920
rect -1860 80810 -1850 80880
rect -1650 80810 -1640 80880
rect -1860 80760 -1640 80810
rect -1360 80990 -1140 81040
rect -1360 80920 -1350 80990
rect -1150 80920 -1140 80990
rect -1360 80880 -1140 80920
rect -1360 80810 -1350 80880
rect -1150 80810 -1140 80880
rect -1360 80760 -1140 80810
rect -860 80990 -640 81040
rect -860 80920 -850 80990
rect -650 80920 -640 80990
rect -860 80880 -640 80920
rect -860 80810 -850 80880
rect -650 80810 -640 80880
rect -860 80760 -640 80810
rect -360 80990 -140 81040
rect -360 80920 -350 80990
rect -150 80920 -140 80990
rect -360 80880 -140 80920
rect -360 80810 -350 80880
rect -150 80810 -140 80880
rect -360 80760 -140 80810
rect 140 80990 360 81040
rect 140 80920 150 80990
rect 350 80920 360 80990
rect 140 80880 360 80920
rect 140 80810 150 80880
rect 350 80810 360 80880
rect 140 80760 360 80810
rect 640 80990 860 81040
rect 640 80920 650 80990
rect 850 80920 860 80990
rect 640 80880 860 80920
rect 640 80810 650 80880
rect 850 80810 860 80880
rect 640 80760 860 80810
rect 1140 80990 1360 81040
rect 1140 80920 1150 80990
rect 1350 80920 1360 80990
rect 1140 80880 1360 80920
rect 1140 80810 1150 80880
rect 1350 80810 1360 80880
rect 1140 80760 1360 80810
rect 1640 80990 1860 81040
rect 1640 80920 1650 80990
rect 1850 80920 1860 80990
rect 1640 80880 1860 80920
rect 1640 80810 1650 80880
rect 1850 80810 1860 80880
rect 1640 80760 1860 80810
rect 2140 80990 2360 81040
rect 2140 80920 2150 80990
rect 2350 80920 2360 80990
rect 2140 80880 2360 80920
rect 2140 80810 2150 80880
rect 2350 80810 2360 80880
rect 2140 80760 2360 80810
rect 2640 80990 2860 81040
rect 2640 80920 2650 80990
rect 2850 80920 2860 80990
rect 2640 80880 2860 80920
rect 2640 80810 2650 80880
rect 2850 80810 2860 80880
rect 2640 80760 2860 80810
rect 3140 80990 3360 81040
rect 3140 80920 3150 80990
rect 3350 80920 3360 80990
rect 3140 80880 3360 80920
rect 3140 80810 3150 80880
rect 3350 80810 3360 80880
rect 3140 80760 3360 80810
rect 3640 80990 3860 81040
rect 3640 80920 3650 80990
rect 3850 80920 3860 80990
rect 3640 80880 3860 80920
rect 3640 80810 3650 80880
rect 3850 80810 3860 80880
rect 3640 80760 3860 80810
rect 4140 80990 4360 81040
rect 4140 80920 4150 80990
rect 4350 80920 4360 80990
rect 4140 80880 4360 80920
rect 4140 80810 4150 80880
rect 4350 80810 4360 80880
rect 4140 80760 4360 80810
rect 4640 80990 4860 81040
rect 4640 80920 4650 80990
rect 4850 80920 4860 80990
rect 4640 80880 4860 80920
rect 4640 80810 4650 80880
rect 4850 80810 4860 80880
rect 4640 80760 4860 80810
rect 5140 80990 5360 81040
rect 5140 80920 5150 80990
rect 5350 80920 5360 80990
rect 5140 80880 5360 80920
rect 5140 80810 5150 80880
rect 5350 80810 5360 80880
rect 5140 80760 5360 80810
rect 5640 80990 5860 81040
rect 5640 80920 5650 80990
rect 5850 80920 5860 80990
rect 5640 80880 5860 80920
rect 5640 80810 5650 80880
rect 5850 80810 5860 80880
rect 5640 80760 5860 80810
rect 6140 80990 6360 81040
rect 6140 80920 6150 80990
rect 6350 80920 6360 80990
rect 6140 80880 6360 80920
rect 6140 80810 6150 80880
rect 6350 80810 6360 80880
rect 6140 80760 6360 80810
rect 6640 80990 6860 81040
rect 6640 80920 6650 80990
rect 6850 80920 6860 80990
rect 6640 80880 6860 80920
rect 6640 80810 6650 80880
rect 6850 80810 6860 80880
rect 6640 80760 6860 80810
rect 7140 80990 7360 81040
rect 7140 80920 7150 80990
rect 7350 80920 7360 80990
rect 7140 80880 7360 80920
rect 7140 80810 7150 80880
rect 7350 80810 7360 80880
rect 7140 80760 7360 80810
rect 7640 80990 7860 81040
rect 7640 80920 7650 80990
rect 7850 80920 7860 80990
rect 7640 80880 7860 80920
rect 7640 80810 7650 80880
rect 7850 80810 7860 80880
rect 7640 80760 7860 80810
rect 8140 80990 8360 81040
rect 8140 80920 8150 80990
rect 8350 80920 8360 80990
rect 8140 80880 8360 80920
rect 8140 80810 8150 80880
rect 8350 80810 8360 80880
rect 8140 80760 8360 80810
rect 8640 80990 8860 81040
rect 8640 80920 8650 80990
rect 8850 80920 8860 80990
rect 8640 80880 8860 80920
rect 8640 80810 8650 80880
rect 8850 80810 8860 80880
rect 8640 80760 8860 80810
rect 9140 80990 9360 81040
rect 9140 80920 9150 80990
rect 9350 80920 9360 80990
rect 9140 80880 9360 80920
rect 9140 80810 9150 80880
rect 9350 80810 9360 80880
rect 9140 80760 9360 80810
rect 9640 80990 9860 81040
rect 9640 80920 9650 80990
rect 9850 80920 9860 80990
rect 9640 80880 9860 80920
rect 9640 80810 9650 80880
rect 9850 80810 9860 80880
rect 9640 80760 9860 80810
rect 10140 80990 10360 81040
rect 10140 80920 10150 80990
rect 10350 80920 10360 80990
rect 10140 80880 10360 80920
rect 10140 80810 10150 80880
rect 10350 80810 10360 80880
rect 10140 80760 10360 80810
rect 10640 80990 10860 81040
rect 10640 80920 10650 80990
rect 10850 80920 10860 80990
rect 10640 80880 10860 80920
rect 10640 80810 10650 80880
rect 10850 80810 10860 80880
rect 10640 80760 10860 80810
rect 11140 80990 11360 81040
rect 11140 80920 11150 80990
rect 11350 80920 11360 80990
rect 11140 80880 11360 80920
rect 11140 80810 11150 80880
rect 11350 80810 11360 80880
rect 11140 80760 11360 80810
rect 11640 80990 11860 81040
rect 11640 80920 11650 80990
rect 11850 80920 11860 80990
rect 11640 80880 11860 80920
rect 11640 80810 11650 80880
rect 11850 80810 11860 80880
rect 11640 80760 11860 80810
rect 12140 80990 12360 81040
rect 12140 80920 12150 80990
rect 12350 80920 12360 80990
rect 12140 80880 12360 80920
rect 12140 80810 12150 80880
rect 12350 80810 12360 80880
rect 12140 80760 12360 80810
rect 12640 80990 12860 81040
rect 12640 80920 12650 80990
rect 12850 80920 12860 80990
rect 12640 80880 12860 80920
rect 12640 80810 12650 80880
rect 12850 80810 12860 80880
rect 12640 80760 12860 80810
rect 13140 80990 13360 81040
rect 13140 80920 13150 80990
rect 13350 80920 13360 80990
rect 13140 80880 13360 80920
rect 13140 80810 13150 80880
rect 13350 80810 13360 80880
rect 13140 80760 13360 80810
rect 13640 80990 13860 81040
rect 13640 80920 13650 80990
rect 13850 80920 13860 80990
rect 13640 80880 13860 80920
rect 13640 80810 13650 80880
rect 13850 80810 13860 80880
rect 13640 80760 13860 80810
rect 14140 80990 14360 81040
rect 14140 80920 14150 80990
rect 14350 80920 14360 80990
rect 14140 80880 14360 80920
rect 14140 80810 14150 80880
rect 14350 80810 14360 80880
rect 14140 80760 14360 80810
rect 14640 80990 14860 81040
rect 14640 80920 14650 80990
rect 14850 80920 14860 80990
rect 14640 80880 14860 80920
rect 14640 80810 14650 80880
rect 14850 80810 14860 80880
rect 14640 80760 14860 80810
rect 15140 80990 15360 81040
rect 15140 80920 15150 80990
rect 15350 80920 15360 80990
rect 15140 80880 15360 80920
rect 15140 80810 15150 80880
rect 15350 80810 15360 80880
rect 15140 80760 15360 80810
rect 15640 80990 15860 81040
rect 15640 80920 15650 80990
rect 15850 80920 15860 80990
rect 15640 80880 15860 80920
rect 15640 80810 15650 80880
rect 15850 80810 15860 80880
rect 15640 80760 15860 80810
rect 16140 80990 16360 81040
rect 16140 80920 16150 80990
rect 16350 80920 16360 80990
rect 16140 80880 16360 80920
rect 16140 80810 16150 80880
rect 16350 80810 16360 80880
rect 16140 80760 16360 80810
rect 16640 80990 16860 81040
rect 16640 80920 16650 80990
rect 16850 80920 16860 80990
rect 16640 80880 16860 80920
rect 16640 80810 16650 80880
rect 16850 80810 16860 80880
rect 16640 80760 16860 80810
rect 17140 80990 17360 81040
rect 17140 80920 17150 80990
rect 17350 80920 17360 80990
rect 17140 80880 17360 80920
rect 17140 80810 17150 80880
rect 17350 80810 17360 80880
rect 17140 80760 17360 80810
rect 17640 80990 17860 81040
rect 17640 80920 17650 80990
rect 17850 80920 17860 80990
rect 17640 80880 17860 80920
rect 17640 80810 17650 80880
rect 17850 80810 17860 80880
rect 17640 80760 17860 80810
rect 18140 80990 18360 81040
rect 18140 80920 18150 80990
rect 18350 80920 18360 80990
rect 18140 80880 18360 80920
rect 18140 80810 18150 80880
rect 18350 80810 18360 80880
rect 18140 80760 18360 80810
rect 18640 80990 18860 81040
rect 18640 80920 18650 80990
rect 18850 80920 18860 80990
rect 18640 80880 18860 80920
rect 18640 80810 18650 80880
rect 18850 80810 18860 80880
rect 18640 80760 18860 80810
rect 19140 80990 19360 81040
rect 19140 80920 19150 80990
rect 19350 80920 19360 80990
rect 19140 80880 19360 80920
rect 19140 80810 19150 80880
rect 19350 80810 19360 80880
rect 19140 80760 19360 80810
rect 19640 80990 19860 81040
rect 19640 80920 19650 80990
rect 19850 80920 19860 80990
rect 19640 80880 19860 80920
rect 19640 80810 19650 80880
rect 19850 80810 19860 80880
rect 19640 80760 19860 80810
rect 20140 80990 20360 81040
rect 20140 80920 20150 80990
rect 20350 80920 20360 80990
rect 20140 80880 20360 80920
rect 20140 80810 20150 80880
rect 20350 80810 20360 80880
rect 20140 80760 20360 80810
rect 20640 80990 20860 81040
rect 20640 80920 20650 80990
rect 20850 80920 20860 80990
rect 20640 80880 20860 80920
rect 20640 80810 20650 80880
rect 20850 80810 20860 80880
rect 20640 80760 20860 80810
rect 21140 80990 21360 81040
rect 21140 80920 21150 80990
rect 21350 80920 21360 80990
rect 21140 80880 21360 80920
rect 21140 80810 21150 80880
rect 21350 80810 21360 80880
rect 21140 80760 21360 80810
rect 21640 80990 21860 81040
rect 21640 80920 21650 80990
rect 21850 80920 21860 80990
rect 21640 80880 21860 80920
rect 21640 80810 21650 80880
rect 21850 80810 21860 80880
rect 21640 80760 21860 80810
rect 22140 80990 22360 81040
rect 22140 80920 22150 80990
rect 22350 80920 22360 80990
rect 22140 80880 22360 80920
rect 22140 80810 22150 80880
rect 22350 80810 22360 80880
rect 22140 80760 22360 80810
rect 22640 80990 22860 81040
rect 22640 80920 22650 80990
rect 22850 80920 22860 80990
rect 22640 80880 22860 80920
rect 22640 80810 22650 80880
rect 22850 80810 22860 80880
rect 22640 80760 22860 80810
rect 23140 80990 23360 81040
rect 23140 80920 23150 80990
rect 23350 80920 23360 80990
rect 23140 80880 23360 80920
rect 23140 80810 23150 80880
rect 23350 80810 23360 80880
rect 23140 80760 23360 80810
rect 23640 80990 23860 81040
rect 23640 80920 23650 80990
rect 23850 80920 23860 80990
rect 23640 80880 23860 80920
rect 23640 80810 23650 80880
rect 23850 80810 23860 80880
rect 23640 80760 23860 80810
rect 24140 80990 24360 81040
rect 24140 80920 24150 80990
rect 24350 80920 24360 80990
rect 24140 80880 24360 80920
rect 24140 80810 24150 80880
rect 24350 80810 24360 80880
rect 24140 80760 24360 80810
rect 24640 80990 24860 81040
rect 24640 80920 24650 80990
rect 24850 80920 24860 80990
rect 24640 80880 24860 80920
rect 24640 80810 24650 80880
rect 24850 80810 24860 80880
rect 24640 80760 24860 80810
rect 25140 80990 25360 81040
rect 25140 80920 25150 80990
rect 25350 80920 25360 80990
rect 25140 80880 25360 80920
rect 25140 80810 25150 80880
rect 25350 80810 25360 80880
rect 25140 80760 25360 80810
rect 25640 80990 25860 81040
rect 25640 80920 25650 80990
rect 25850 80920 25860 80990
rect 25640 80880 25860 80920
rect 25640 80810 25650 80880
rect 25850 80810 25860 80880
rect 25640 80760 25860 80810
rect 26140 80990 26360 81040
rect 26140 80920 26150 80990
rect 26350 80920 26360 80990
rect 26140 80880 26360 80920
rect 26140 80810 26150 80880
rect 26350 80810 26360 80880
rect 26140 80760 26360 80810
rect 26640 80990 26860 81040
rect 26640 80920 26650 80990
rect 26850 80920 26860 80990
rect 26640 80880 26860 80920
rect 26640 80810 26650 80880
rect 26850 80810 26860 80880
rect 26640 80760 26860 80810
rect 27140 80990 27360 81040
rect 27140 80920 27150 80990
rect 27350 80920 27360 80990
rect 27140 80880 27360 80920
rect 27140 80810 27150 80880
rect 27350 80810 27360 80880
rect 27140 80760 27360 80810
rect 27640 80990 27860 81040
rect 27640 80920 27650 80990
rect 27850 80920 27860 80990
rect 27640 80880 27860 80920
rect 27640 80810 27650 80880
rect 27850 80810 27860 80880
rect 27640 80760 27860 80810
rect 28140 80990 28360 81040
rect 28140 80920 28150 80990
rect 28350 80920 28360 80990
rect 28140 80880 28360 80920
rect 28140 80810 28150 80880
rect 28350 80810 28360 80880
rect 28140 80760 28360 80810
rect 28640 80990 28860 81040
rect 28640 80920 28650 80990
rect 28850 80920 28860 80990
rect 28640 80880 28860 80920
rect 28640 80810 28650 80880
rect 28850 80810 28860 80880
rect 28640 80760 28860 80810
rect 29140 80990 29360 81040
rect 29140 80920 29150 80990
rect 29350 80920 29360 80990
rect 29140 80880 29360 80920
rect 29140 80810 29150 80880
rect 29350 80810 29360 80880
rect 29140 80760 29360 80810
rect 29640 80990 29860 81040
rect 29640 80920 29650 80990
rect 29850 80920 29860 80990
rect 29640 80880 29860 80920
rect 29640 80810 29650 80880
rect 29850 80810 29860 80880
rect 29640 80760 29860 80810
rect 30140 80990 30360 81040
rect 30140 80920 30150 80990
rect 30350 80920 30360 80990
rect 30140 80880 30360 80920
rect 30140 80810 30150 80880
rect 30350 80810 30360 80880
rect 30140 80760 30360 80810
rect 30640 80990 30860 81040
rect 30640 80920 30650 80990
rect 30850 80920 30860 80990
rect 30640 80880 30860 80920
rect 30640 80810 30650 80880
rect 30850 80810 30860 80880
rect 30640 80760 30860 80810
rect 31140 80990 31360 81040
rect 31140 80920 31150 80990
rect 31350 80920 31360 80990
rect 31140 80880 31360 80920
rect 31140 80810 31150 80880
rect 31350 80810 31360 80880
rect 31140 80760 31360 80810
rect 31640 80990 31860 81040
rect 31640 80920 31650 80990
rect 31850 80920 31860 80990
rect 31640 80880 31860 80920
rect 31640 80810 31650 80880
rect 31850 80810 31860 80880
rect 31640 80760 31860 80810
rect 32140 80990 32360 81040
rect 32140 80920 32150 80990
rect 32350 80920 32360 80990
rect 32140 80880 32360 80920
rect 32140 80810 32150 80880
rect 32350 80810 32360 80880
rect 32140 80760 32360 80810
rect 32640 80990 32860 81040
rect 32640 80920 32650 80990
rect 32850 80920 32860 80990
rect 32640 80880 32860 80920
rect 32640 80810 32650 80880
rect 32850 80810 32860 80880
rect 32640 80760 32860 80810
rect 33140 80990 33360 81040
rect 33140 80920 33150 80990
rect 33350 80920 33360 80990
rect 33140 80880 33360 80920
rect 33140 80810 33150 80880
rect 33350 80810 33360 80880
rect 33140 80760 33360 80810
rect 33640 80990 33860 81040
rect 33640 80920 33650 80990
rect 33850 80920 33860 80990
rect 33640 80880 33860 80920
rect 33640 80810 33650 80880
rect 33850 80810 33860 80880
rect 33640 80760 33860 80810
rect 34140 80990 34360 81040
rect 34140 80920 34150 80990
rect 34350 80920 34360 80990
rect 34140 80880 34360 80920
rect 34140 80810 34150 80880
rect 34350 80810 34360 80880
rect 34140 80760 34360 80810
rect 34640 80990 34860 81040
rect 34640 80920 34650 80990
rect 34850 80920 34860 80990
rect 34640 80880 34860 80920
rect 34640 80810 34650 80880
rect 34850 80810 34860 80880
rect 34640 80760 34860 80810
rect 35140 80990 35360 81040
rect 35140 80920 35150 80990
rect 35350 80920 35360 80990
rect 35140 80880 35360 80920
rect 35140 80810 35150 80880
rect 35350 80810 35360 80880
rect 35140 80760 35360 80810
rect 35640 80990 35860 81040
rect 35640 80920 35650 80990
rect 35850 80920 35860 80990
rect 35640 80880 35860 80920
rect 35640 80810 35650 80880
rect 35850 80810 35860 80880
rect 35640 80760 35860 80810
rect 36140 80990 36360 81040
rect 36140 80920 36150 80990
rect 36350 80920 36360 80990
rect 36140 80880 36360 80920
rect 36140 80810 36150 80880
rect 36350 80810 36360 80880
rect 36140 80760 36360 80810
rect 36640 80990 36860 81040
rect 36640 80920 36650 80990
rect 36850 80920 36860 80990
rect 36640 80880 36860 80920
rect 36640 80810 36650 80880
rect 36850 80810 36860 80880
rect 36640 80760 36860 80810
rect 37140 80990 37360 81040
rect 37140 80920 37150 80990
rect 37350 80920 37360 80990
rect 37140 80880 37360 80920
rect 37140 80810 37150 80880
rect 37350 80810 37360 80880
rect 37140 80760 37360 80810
rect 37640 80990 37860 81040
rect 37640 80920 37650 80990
rect 37850 80920 37860 80990
rect 37640 80880 37860 80920
rect 37640 80810 37650 80880
rect 37850 80810 37860 80880
rect 37640 80760 37860 80810
rect 38140 80990 38360 81040
rect 38140 80920 38150 80990
rect 38350 80920 38360 80990
rect 38140 80880 38360 80920
rect 38140 80810 38150 80880
rect 38350 80810 38360 80880
rect 38140 80760 38360 80810
rect 38640 80990 38860 81040
rect 38640 80920 38650 80990
rect 38850 80920 38860 80990
rect 38640 80880 38860 80920
rect 38640 80810 38650 80880
rect 38850 80810 38860 80880
rect 38640 80760 38860 80810
rect 39140 80990 39360 81040
rect 39140 80920 39150 80990
rect 39350 80920 39360 80990
rect 39140 80880 39360 80920
rect 39140 80810 39150 80880
rect 39350 80810 39360 80880
rect 39140 80760 39360 80810
rect 39640 80990 39860 81040
rect 39640 80920 39650 80990
rect 39850 80920 39860 80990
rect 39640 80880 39860 80920
rect 39640 80810 39650 80880
rect 39850 80810 39860 80880
rect 39640 80760 39860 80810
rect 40140 80990 40360 81040
rect 40140 80920 40150 80990
rect 40350 80920 40360 80990
rect 40140 80880 40360 80920
rect 40140 80810 40150 80880
rect 40350 80810 40360 80880
rect 40140 80760 40360 80810
rect 40640 80990 40860 81040
rect 40640 80920 40650 80990
rect 40850 80920 40860 80990
rect 40640 80880 40860 80920
rect 40640 80810 40650 80880
rect 40850 80810 40860 80880
rect 40640 80760 40860 80810
rect 41140 80990 41360 81040
rect 41140 80920 41150 80990
rect 41350 80920 41360 80990
rect 41140 80880 41360 80920
rect 41140 80810 41150 80880
rect 41350 80810 41360 80880
rect 41140 80760 41360 80810
rect 41640 80990 41860 81040
rect 41640 80920 41650 80990
rect 41850 80920 41860 80990
rect 41640 80880 41860 80920
rect 41640 80810 41650 80880
rect 41850 80810 41860 80880
rect 41640 80760 41860 80810
rect 42140 80990 42360 81040
rect 42140 80920 42150 80990
rect 42350 80920 42360 80990
rect 42140 80880 42360 80920
rect 42140 80810 42150 80880
rect 42350 80810 42360 80880
rect 42140 80760 42360 80810
rect 42640 80990 42860 81040
rect 42640 80920 42650 80990
rect 42850 80920 42860 80990
rect 42640 80880 42860 80920
rect 42640 80810 42650 80880
rect 42850 80810 42860 80880
rect 42640 80760 42860 80810
rect 43140 80990 43360 81040
rect 43140 80920 43150 80990
rect 43350 80920 43360 80990
rect 43140 80880 43360 80920
rect 43140 80810 43150 80880
rect 43350 80810 43360 80880
rect 43140 80760 43360 80810
rect 43640 80990 43860 81040
rect 43640 80920 43650 80990
rect 43850 80920 43860 80990
rect 43640 80880 43860 80920
rect 43640 80810 43650 80880
rect 43850 80810 43860 80880
rect 43640 80760 43860 80810
rect 44140 80990 44360 81040
rect 44140 80920 44150 80990
rect 44350 80920 44360 80990
rect 44140 80880 44360 80920
rect 44140 80810 44150 80880
rect 44350 80810 44360 80880
rect 44140 80760 44360 80810
rect 44640 80990 44860 81040
rect 44640 80920 44650 80990
rect 44850 80920 44860 80990
rect 44640 80880 44860 80920
rect 44640 80810 44650 80880
rect 44850 80810 44860 80880
rect 44640 80760 44860 80810
rect 45140 80990 45360 81040
rect 45140 80920 45150 80990
rect 45350 80920 45360 80990
rect 45140 80880 45360 80920
rect 45140 80810 45150 80880
rect 45350 80810 45360 80880
rect 45140 80760 45360 80810
rect 45640 80990 45860 81040
rect 45640 80920 45650 80990
rect 45850 80920 45860 80990
rect 45640 80880 45860 80920
rect 45640 80810 45650 80880
rect 45850 80810 45860 80880
rect 45640 80760 45860 80810
rect 46140 80990 46360 81040
rect 46140 80920 46150 80990
rect 46350 80920 46360 80990
rect 46140 80880 46360 80920
rect 46140 80810 46150 80880
rect 46350 80810 46360 80880
rect 46140 80760 46360 80810
rect 46640 80990 46860 81040
rect 46640 80920 46650 80990
rect 46850 80920 46860 80990
rect 46640 80880 46860 80920
rect 46640 80810 46650 80880
rect 46850 80810 46860 80880
rect 46640 80760 46860 80810
rect 47140 80990 47360 81040
rect 47140 80920 47150 80990
rect 47350 80920 47360 80990
rect 47140 80880 47360 80920
rect 47140 80810 47150 80880
rect 47350 80810 47360 80880
rect 47140 80760 47360 80810
rect 47640 80990 47860 81040
rect 47640 80920 47650 80990
rect 47850 80920 47860 80990
rect 47640 80880 47860 80920
rect 47640 80810 47650 80880
rect 47850 80810 47860 80880
rect 47640 80760 47860 80810
rect 48140 80990 48360 81040
rect 48140 80920 48150 80990
rect 48350 80920 48360 80990
rect 48140 80880 48360 80920
rect 48140 80810 48150 80880
rect 48350 80810 48360 80880
rect 48140 80760 48360 80810
rect 48640 80990 48860 81040
rect 48640 80920 48650 80990
rect 48850 80920 48860 80990
rect 48640 80880 48860 80920
rect 48640 80810 48650 80880
rect 48850 80810 48860 80880
rect 48640 80760 48860 80810
rect 49140 80990 49360 81040
rect 49140 80920 49150 80990
rect 49350 80920 49360 80990
rect 49140 80880 49360 80920
rect 49140 80810 49150 80880
rect 49350 80810 49360 80880
rect 49140 80760 49360 80810
rect 49640 80990 49860 81040
rect 49640 80920 49650 80990
rect 49850 80920 49860 80990
rect 49640 80880 49860 80920
rect 49640 80810 49650 80880
rect 49850 80810 49860 80880
rect 49640 80760 49860 80810
rect 50140 80990 50360 81040
rect 50140 80920 50150 80990
rect 50350 80920 50360 80990
rect 50140 80880 50360 80920
rect 50140 80810 50150 80880
rect 50350 80810 50360 80880
rect 50140 80760 50360 80810
rect 50640 80990 50860 81040
rect 50640 80920 50650 80990
rect 50850 80920 50860 80990
rect 50640 80880 50860 80920
rect 50640 80810 50650 80880
rect 50850 80810 50860 80880
rect 50640 80760 50860 80810
rect 51140 80990 51360 81040
rect 51140 80920 51150 80990
rect 51350 80920 51360 80990
rect 51140 80880 51360 80920
rect 51140 80810 51150 80880
rect 51350 80810 51360 80880
rect 51140 80760 51360 80810
rect 51640 80990 51860 81040
rect 51640 80920 51650 80990
rect 51850 80920 51860 80990
rect 51640 80880 51860 80920
rect 51640 80810 51650 80880
rect 51850 80810 51860 80880
rect 51640 80760 51860 80810
rect 52140 80990 52360 81040
rect 52140 80920 52150 80990
rect 52350 80920 52360 80990
rect 52140 80880 52360 80920
rect 52140 80810 52150 80880
rect 52350 80810 52360 80880
rect 52140 80760 52360 80810
rect 52640 80990 52860 81040
rect 52640 80920 52650 80990
rect 52850 80920 52860 80990
rect 52640 80880 52860 80920
rect 52640 80810 52650 80880
rect 52850 80810 52860 80880
rect 52640 80760 52860 80810
rect 53140 80990 53360 81040
rect 53140 80920 53150 80990
rect 53350 80920 53360 80990
rect 53140 80880 53360 80920
rect 53140 80810 53150 80880
rect 53350 80810 53360 80880
rect 53140 80760 53360 80810
rect 53640 80990 53860 81040
rect 53640 80920 53650 80990
rect 53850 80920 53860 80990
rect 53640 80880 53860 80920
rect 53640 80810 53650 80880
rect 53850 80810 53860 80880
rect 53640 80760 53860 80810
rect 54140 80990 54360 81040
rect 54140 80920 54150 80990
rect 54350 80920 54360 80990
rect 54140 80880 54360 80920
rect 54140 80810 54150 80880
rect 54350 80810 54360 80880
rect 54140 80760 54360 80810
rect 54640 80990 54860 81040
rect 54640 80920 54650 80990
rect 54850 80920 54860 80990
rect 54640 80880 54860 80920
rect 54640 80810 54650 80880
rect 54850 80810 54860 80880
rect 54640 80760 54860 80810
rect 55140 80990 55360 81040
rect 55140 80920 55150 80990
rect 55350 80920 55360 80990
rect 55140 80880 55360 80920
rect 55140 80810 55150 80880
rect 55350 80810 55360 80880
rect 55140 80760 55360 80810
rect 55640 80990 55860 81040
rect 55640 80920 55650 80990
rect 55850 80920 55860 80990
rect 55640 80880 55860 80920
rect 55640 80810 55650 80880
rect 55850 80810 55860 80880
rect 55640 80760 55860 80810
rect 56140 80990 56360 81040
rect 56140 80920 56150 80990
rect 56350 80920 56360 80990
rect 56140 80880 56360 80920
rect 56140 80810 56150 80880
rect 56350 80810 56360 80880
rect 56140 80760 56360 80810
rect 56640 80990 56860 81040
rect 56640 80920 56650 80990
rect 56850 80920 56860 80990
rect 56640 80880 56860 80920
rect 56640 80810 56650 80880
rect 56850 80810 56860 80880
rect 56640 80760 56860 80810
rect 57140 80990 57360 81040
rect 57140 80920 57150 80990
rect 57350 80920 57360 80990
rect 57140 80880 57360 80920
rect 57140 80810 57150 80880
rect 57350 80810 57360 80880
rect 57140 80760 57360 80810
rect 57640 80990 57860 81040
rect 57640 80920 57650 80990
rect 57850 80920 57860 80990
rect 57640 80880 57860 80920
rect 57640 80810 57650 80880
rect 57850 80810 57860 80880
rect 57640 80760 57860 80810
rect 58140 80990 58360 81040
rect 58140 80920 58150 80990
rect 58350 80920 58360 80990
rect 58140 80880 58360 80920
rect 58140 80810 58150 80880
rect 58350 80810 58360 80880
rect 58140 80760 58360 80810
rect 58640 80990 58860 81040
rect 58640 80920 58650 80990
rect 58850 80920 58860 80990
rect 58640 80880 58860 80920
rect 58640 80810 58650 80880
rect 58850 80810 58860 80880
rect 58640 80760 58860 80810
rect 59140 80990 59360 81040
rect 59140 80920 59150 80990
rect 59350 80920 59360 80990
rect 59140 80880 59360 80920
rect 59140 80810 59150 80880
rect 59350 80810 59360 80880
rect 59140 80760 59360 80810
rect 59640 80990 59860 81040
rect 59640 80920 59650 80990
rect 59850 80920 59860 80990
rect 59640 80880 59860 80920
rect 59640 80810 59650 80880
rect 59850 80810 59860 80880
rect 59640 80760 59860 80810
rect 60140 80990 60360 81040
rect 60140 80920 60150 80990
rect 60350 80920 60360 80990
rect 60140 80880 60360 80920
rect 60140 80810 60150 80880
rect 60350 80810 60360 80880
rect 60140 80760 60360 80810
rect 60640 80990 60860 81040
rect 60640 80920 60650 80990
rect 60850 80920 60860 80990
rect 60640 80880 60860 80920
rect 60640 80810 60650 80880
rect 60850 80810 60860 80880
rect 60640 80760 60860 80810
rect 61140 80990 61360 81040
rect 61140 80920 61150 80990
rect 61350 80920 61360 80990
rect 61140 80880 61360 80920
rect 61140 80810 61150 80880
rect 61350 80810 61360 80880
rect 61140 80760 61360 80810
rect 61640 80990 61860 81040
rect 61640 80920 61650 80990
rect 61850 80920 61860 80990
rect 61640 80880 61860 80920
rect 61640 80810 61650 80880
rect 61850 80810 61860 80880
rect 61640 80760 61860 80810
rect 62140 80990 62360 81040
rect 62140 80920 62150 80990
rect 62350 80920 62360 80990
rect 62140 80880 62360 80920
rect 62140 80810 62150 80880
rect 62350 80810 62360 80880
rect 62140 80760 62360 80810
rect 62640 80990 62860 81040
rect 62640 80920 62650 80990
rect 62850 80920 62860 80990
rect 62640 80880 62860 80920
rect 62640 80810 62650 80880
rect 62850 80810 62860 80880
rect 62640 80760 62860 80810
rect 63140 80990 63360 81040
rect 63140 80920 63150 80990
rect 63350 80920 63360 80990
rect 63140 80880 63360 80920
rect 63140 80810 63150 80880
rect 63350 80810 63360 80880
rect 63140 80760 63360 80810
rect 63640 80990 63860 81040
rect 63640 80920 63650 80990
rect 63850 80920 63860 80990
rect 63640 80880 63860 80920
rect 63640 80810 63650 80880
rect 63850 80810 63860 80880
rect 63640 80760 63860 80810
rect 64140 80990 64360 81040
rect 64140 80920 64150 80990
rect 64350 80920 64360 80990
rect 64140 80880 64360 80920
rect 64140 80810 64150 80880
rect 64350 80810 64360 80880
rect 64140 80760 64360 80810
rect 64640 80990 64860 81040
rect 64640 80920 64650 80990
rect 64850 80920 64860 80990
rect 64640 80880 64860 80920
rect 64640 80810 64650 80880
rect 64850 80810 64860 80880
rect 64640 80760 64860 80810
rect 65140 80990 65360 81040
rect 65140 80920 65150 80990
rect 65350 80920 65360 80990
rect 65140 80880 65360 80920
rect 65140 80810 65150 80880
rect 65350 80810 65360 80880
rect 65140 80760 65360 80810
rect 65640 80990 65860 81040
rect 65640 80920 65650 80990
rect 65850 80920 65860 80990
rect 65640 80880 65860 80920
rect 65640 80810 65650 80880
rect 65850 80810 65860 80880
rect 65640 80760 65860 80810
rect 66140 80990 66360 81040
rect 66140 80920 66150 80990
rect 66350 80920 66360 80990
rect 66140 80880 66360 80920
rect 66140 80810 66150 80880
rect 66350 80810 66360 80880
rect 66140 80760 66360 80810
rect 66640 80990 66860 81040
rect 66640 80920 66650 80990
rect 66850 80920 66860 80990
rect 66640 80880 66860 80920
rect 66640 80810 66650 80880
rect 66850 80810 66860 80880
rect 66640 80760 66860 80810
rect 67140 80990 67360 81040
rect 67140 80920 67150 80990
rect 67350 80920 67360 80990
rect 67140 80880 67360 80920
rect 67140 80810 67150 80880
rect 67350 80810 67360 80880
rect 67140 80760 67360 80810
rect 67640 80990 67860 81040
rect 67640 80920 67650 80990
rect 67850 80920 67860 80990
rect 67640 80880 67860 80920
rect 67640 80810 67650 80880
rect 67850 80810 67860 80880
rect 67640 80760 67860 80810
rect 68140 80990 68360 81040
rect 68140 80920 68150 80990
rect 68350 80920 68360 80990
rect 68140 80880 68360 80920
rect 68140 80810 68150 80880
rect 68350 80810 68360 80880
rect 68140 80760 68360 80810
rect 68640 80990 68860 81040
rect 68640 80920 68650 80990
rect 68850 80920 68860 80990
rect 68640 80880 68860 80920
rect 68640 80810 68650 80880
rect 68850 80810 68860 80880
rect 68640 80760 68860 80810
rect 69140 80990 69360 81040
rect 69140 80920 69150 80990
rect 69350 80920 69360 80990
rect 69140 80880 69360 80920
rect 69140 80810 69150 80880
rect 69350 80810 69360 80880
rect 69140 80760 69360 80810
rect 69640 80990 69860 81040
rect 69640 80920 69650 80990
rect 69850 80920 69860 80990
rect 69640 80880 69860 80920
rect 69640 80810 69650 80880
rect 69850 80810 69860 80880
rect 69640 80760 69860 80810
rect 70140 80990 70360 81040
rect 70140 80920 70150 80990
rect 70350 80920 70360 80990
rect 70140 80880 70360 80920
rect 70140 80810 70150 80880
rect 70350 80810 70360 80880
rect 70140 80760 70360 80810
rect 70640 80990 70860 81040
rect 70640 80920 70650 80990
rect 70850 80920 70860 80990
rect 70640 80880 70860 80920
rect 70640 80810 70650 80880
rect 70850 80810 70860 80880
rect 70640 80760 70860 80810
rect 71140 80990 71360 81040
rect 71140 80920 71150 80990
rect 71350 80920 71360 80990
rect 71140 80880 71360 80920
rect 71140 80810 71150 80880
rect 71350 80810 71360 80880
rect 71140 80760 71360 80810
rect 71640 80990 71860 81040
rect 71640 80920 71650 80990
rect 71850 80920 71860 80990
rect 71640 80880 71860 80920
rect 71640 80810 71650 80880
rect 71850 80810 71860 80880
rect 71640 80760 71860 80810
rect 72140 80990 72360 81040
rect 72140 80920 72150 80990
rect 72350 80920 72360 80990
rect 72140 80880 72360 80920
rect 72140 80810 72150 80880
rect 72350 80810 72360 80880
rect 72140 80760 72360 80810
rect 72640 80990 72860 81040
rect 72640 80920 72650 80990
rect 72850 80920 72860 80990
rect 72640 80880 72860 80920
rect 72640 80810 72650 80880
rect 72850 80810 72860 80880
rect 72640 80760 72860 80810
rect 73140 80990 73360 81040
rect 73140 80920 73150 80990
rect 73350 80920 73360 80990
rect 73140 80880 73360 80920
rect 73140 80810 73150 80880
rect 73350 80810 73360 80880
rect 73140 80760 73360 80810
rect 73640 80990 73860 81040
rect 73640 80920 73650 80990
rect 73850 80920 73860 80990
rect 73640 80880 73860 80920
rect 73640 80810 73650 80880
rect 73850 80810 73860 80880
rect 73640 80760 73860 80810
rect 74140 80990 74360 81040
rect 74140 80920 74150 80990
rect 74350 80920 74360 80990
rect 74140 80880 74360 80920
rect 74140 80810 74150 80880
rect 74350 80810 74360 80880
rect 74140 80760 74360 80810
rect 74640 80990 74860 81040
rect 74640 80920 74650 80990
rect 74850 80920 74860 80990
rect 74640 80880 74860 80920
rect 74640 80810 74650 80880
rect 74850 80810 74860 80880
rect 74640 80760 74860 80810
rect 75140 80990 75360 81040
rect 75140 80920 75150 80990
rect 75350 80920 75360 80990
rect 75140 80880 75360 80920
rect 75140 80810 75150 80880
rect 75350 80810 75360 80880
rect 75140 80760 75360 80810
rect 75640 80990 75860 81040
rect 75640 80920 75650 80990
rect 75850 80920 75860 80990
rect 75640 80880 75860 80920
rect 75640 80810 75650 80880
rect 75850 80810 75860 80880
rect 75640 80760 75860 80810
rect 76140 80990 76360 81040
rect 76140 80920 76150 80990
rect 76350 80920 76360 80990
rect 76140 80880 76360 80920
rect 76140 80810 76150 80880
rect 76350 80810 76360 80880
rect 76140 80760 76360 80810
rect 76640 80990 76860 81040
rect 76640 80920 76650 80990
rect 76850 80920 76860 80990
rect 76640 80880 76860 80920
rect 76640 80810 76650 80880
rect 76850 80810 76860 80880
rect 76640 80760 76860 80810
rect 77140 80990 77360 81040
rect 77140 80920 77150 80990
rect 77350 80920 77360 80990
rect 77140 80880 77360 80920
rect 77140 80810 77150 80880
rect 77350 80810 77360 80880
rect 77140 80760 77360 80810
rect 77640 80990 77860 81040
rect 77640 80920 77650 80990
rect 77850 80920 77860 80990
rect 77640 80880 77860 80920
rect 77640 80810 77650 80880
rect 77850 80810 77860 80880
rect 77640 80760 77860 80810
rect 78140 80990 78360 81040
rect 78140 80920 78150 80990
rect 78350 80920 78360 80990
rect 78140 80880 78360 80920
rect 78140 80810 78150 80880
rect 78350 80810 78360 80880
rect 78140 80760 78360 80810
rect 78640 80990 78860 81040
rect 78640 80920 78650 80990
rect 78850 80920 78860 80990
rect 78640 80880 78860 80920
rect 78640 80810 78650 80880
rect 78850 80810 78860 80880
rect 78640 80760 78860 80810
rect 79140 80990 79360 81040
rect 79140 80920 79150 80990
rect 79350 80920 79360 80990
rect 79140 80880 79360 80920
rect 79140 80810 79150 80880
rect 79350 80810 79360 80880
rect 79140 80760 79360 80810
rect 79640 80990 79860 81040
rect 79640 80920 79650 80990
rect 79850 80920 79860 80990
rect 79640 80880 79860 80920
rect 79640 80810 79650 80880
rect 79850 80810 79860 80880
rect 79640 80760 79860 80810
rect 80140 80990 80360 81040
rect 80140 80920 80150 80990
rect 80350 80920 80360 80990
rect 80140 80880 80360 80920
rect 80140 80810 80150 80880
rect 80350 80810 80360 80880
rect 80140 80760 80360 80810
rect 80640 80990 80860 81040
rect 80640 80920 80650 80990
rect 80850 80920 80860 80990
rect 80640 80880 80860 80920
rect 80640 80810 80650 80880
rect 80850 80810 80860 80880
rect 80640 80760 80860 80810
rect 81140 80990 81360 81040
rect 81140 80920 81150 80990
rect 81350 80920 81360 80990
rect 81140 80880 81360 80920
rect 81140 80810 81150 80880
rect 81350 80810 81360 80880
rect 81140 80760 81360 80810
rect 81640 80990 81860 81040
rect 81640 80920 81650 80990
rect 81850 80920 81860 80990
rect 81640 80880 81860 80920
rect 81640 80810 81650 80880
rect 81850 80810 81860 80880
rect 81640 80760 81860 80810
rect 82140 80990 82360 81040
rect 82140 80920 82150 80990
rect 82350 80920 82360 80990
rect 82140 80880 82360 80920
rect 82140 80810 82150 80880
rect 82350 80810 82360 80880
rect 82140 80760 82360 80810
rect 82640 80990 82860 81040
rect 82640 80920 82650 80990
rect 82850 80920 82860 80990
rect 82640 80880 82860 80920
rect 82640 80810 82650 80880
rect 82850 80810 82860 80880
rect 82640 80760 82860 80810
rect 83140 80990 83360 81040
rect 83140 80920 83150 80990
rect 83350 80920 83360 80990
rect 83140 80880 83360 80920
rect 83140 80810 83150 80880
rect 83350 80810 83360 80880
rect 83140 80760 83360 80810
rect 83640 80990 83860 81040
rect 83640 80920 83650 80990
rect 83850 80920 83860 80990
rect 83640 80880 83860 80920
rect 83640 80810 83650 80880
rect 83850 80810 83860 80880
rect 83640 80760 83860 80810
rect 84140 80990 84360 81040
rect 84140 80920 84150 80990
rect 84350 80920 84360 80990
rect 84140 80880 84360 80920
rect 84140 80810 84150 80880
rect 84350 80810 84360 80880
rect 84140 80760 84360 80810
rect 84640 80990 84860 81040
rect 84640 80920 84650 80990
rect 84850 80920 84860 80990
rect 84640 80880 84860 80920
rect 84640 80810 84650 80880
rect 84850 80810 84860 80880
rect 84640 80760 84860 80810
rect 85140 80990 85360 81040
rect 85140 80920 85150 80990
rect 85350 80920 85360 80990
rect 85140 80880 85360 80920
rect 85140 80810 85150 80880
rect 85350 80810 85360 80880
rect 85140 80760 85360 80810
rect 85640 80990 85860 81040
rect 85640 80920 85650 80990
rect 85850 80920 85860 80990
rect 85640 80880 85860 80920
rect 85640 80810 85650 80880
rect 85850 80810 85860 80880
rect 85640 80760 85860 80810
rect 86140 80990 86360 81040
rect 86140 80920 86150 80990
rect 86350 80920 86360 80990
rect 86140 80880 86360 80920
rect 86140 80810 86150 80880
rect 86350 80810 86360 80880
rect 86140 80760 86360 80810
rect 86640 80990 86860 81040
rect 86640 80920 86650 80990
rect 86850 80920 86860 80990
rect 86640 80880 86860 80920
rect 86640 80810 86650 80880
rect 86850 80810 86860 80880
rect 86640 80760 86860 80810
rect 87140 80990 87360 81040
rect 87140 80920 87150 80990
rect 87350 80920 87360 80990
rect 87140 80880 87360 80920
rect 87140 80810 87150 80880
rect 87350 80810 87360 80880
rect 87140 80760 87360 80810
rect 87640 80990 87860 81040
rect 87640 80920 87650 80990
rect 87850 80920 87860 80990
rect 87640 80880 87860 80920
rect 87640 80810 87650 80880
rect 87850 80810 87860 80880
rect 87640 80760 87860 80810
rect 88140 80990 88360 81040
rect 88140 80920 88150 80990
rect 88350 80920 88360 80990
rect 88140 80880 88360 80920
rect 88140 80810 88150 80880
rect 88350 80810 88360 80880
rect 88140 80760 88360 80810
rect 88640 80990 88860 81040
rect 88640 80920 88650 80990
rect 88850 80920 88860 80990
rect 88640 80880 88860 80920
rect 88640 80810 88650 80880
rect 88850 80810 88860 80880
rect 88640 80760 88860 80810
rect 89140 80990 89360 81040
rect 89140 80920 89150 80990
rect 89350 80920 89360 80990
rect 89140 80880 89360 80920
rect 89140 80810 89150 80880
rect 89350 80810 89360 80880
rect 89140 80760 89360 80810
rect 89640 80990 89860 81040
rect 89640 80920 89650 80990
rect 89850 80920 89860 80990
rect 89640 80880 89860 80920
rect 89640 80810 89650 80880
rect 89850 80810 89860 80880
rect 89640 80760 89860 80810
rect 90140 80990 90360 81040
rect 90140 80920 90150 80990
rect 90350 80920 90360 80990
rect 90140 80880 90360 80920
rect 90140 80810 90150 80880
rect 90350 80810 90360 80880
rect 90140 80760 90360 80810
rect 90640 80990 90860 81040
rect 90640 80920 90650 80990
rect 90850 80920 90860 80990
rect 90640 80880 90860 80920
rect 90640 80810 90650 80880
rect 90850 80810 90860 80880
rect 90640 80760 90860 80810
rect 91140 80990 91360 81040
rect 91140 80920 91150 80990
rect 91350 80920 91360 80990
rect 91140 80880 91360 80920
rect 91140 80810 91150 80880
rect 91350 80810 91360 80880
rect 91140 80760 91360 80810
rect 91640 80990 91860 81040
rect 91640 80920 91650 80990
rect 91850 80920 91860 80990
rect 91640 80880 91860 80920
rect 91640 80810 91650 80880
rect 91850 80810 91860 80880
rect 91640 80760 91860 80810
rect 92140 80990 92360 81040
rect 92140 80920 92150 80990
rect 92350 80920 92360 80990
rect 92140 80880 92360 80920
rect 92140 80810 92150 80880
rect 92350 80810 92360 80880
rect 92140 80760 92360 80810
rect 92640 80990 92860 81040
rect 92640 80920 92650 80990
rect 92850 80920 92860 80990
rect 92640 80880 92860 80920
rect 92640 80810 92650 80880
rect 92850 80810 92860 80880
rect 92640 80760 92860 80810
rect 93140 80990 93360 81040
rect 93140 80920 93150 80990
rect 93350 80920 93360 80990
rect 93140 80880 93360 80920
rect 93140 80810 93150 80880
rect 93350 80810 93360 80880
rect 93140 80760 93360 80810
rect 93640 80990 93860 81040
rect 93640 80920 93650 80990
rect 93850 80920 93860 80990
rect 93640 80880 93860 80920
rect 93640 80810 93650 80880
rect 93850 80810 93860 80880
rect 93640 80760 93860 80810
rect 94140 80990 94360 81040
rect 94140 80920 94150 80990
rect 94350 80920 94360 80990
rect 94140 80880 94360 80920
rect 94140 80810 94150 80880
rect 94350 80810 94360 80880
rect 94140 80760 94360 80810
rect 94640 80990 94860 81040
rect 94640 80920 94650 80990
rect 94850 80920 94860 80990
rect 94640 80880 94860 80920
rect 94640 80810 94650 80880
rect 94850 80810 94860 80880
rect 94640 80760 94860 80810
rect 95140 80990 95360 81040
rect 95140 80920 95150 80990
rect 95350 80920 95360 80990
rect 95140 80880 95360 80920
rect 95140 80810 95150 80880
rect 95350 80810 95360 80880
rect 95140 80760 95360 80810
rect 95640 80990 95860 81040
rect 95640 80920 95650 80990
rect 95850 80920 95860 80990
rect 95640 80880 95860 80920
rect 95640 80810 95650 80880
rect 95850 80810 95860 80880
rect 95640 80760 95860 80810
rect 96140 80990 96360 81040
rect 96140 80920 96150 80990
rect 96350 80920 96360 80990
rect 96140 80880 96360 80920
rect 96140 80810 96150 80880
rect 96350 80810 96360 80880
rect 96140 80760 96360 80810
rect 96640 80990 96860 81040
rect 96640 80920 96650 80990
rect 96850 80920 96860 80990
rect 96640 80880 96860 80920
rect 96640 80810 96650 80880
rect 96850 80810 96860 80880
rect 96640 80760 96860 80810
rect 97140 80990 97360 81040
rect 97140 80920 97150 80990
rect 97350 80920 97360 80990
rect 97140 80880 97360 80920
rect 97140 80810 97150 80880
rect 97350 80810 97360 80880
rect 97140 80760 97360 80810
rect 97640 80990 97860 81040
rect 97640 80920 97650 80990
rect 97850 80920 97860 80990
rect 97640 80880 97860 80920
rect 97640 80810 97650 80880
rect 97850 80810 97860 80880
rect 97640 80760 97860 80810
rect 98140 80990 98360 81040
rect 98140 80920 98150 80990
rect 98350 80920 98360 80990
rect 98140 80880 98360 80920
rect 98140 80810 98150 80880
rect 98350 80810 98360 80880
rect 98140 80760 98360 80810
rect 98640 80990 98860 81040
rect 98640 80920 98650 80990
rect 98850 80920 98860 80990
rect 98640 80880 98860 80920
rect 98640 80810 98650 80880
rect 98850 80810 98860 80880
rect 98640 80760 98860 80810
rect 99140 80990 99360 81040
rect 99140 80920 99150 80990
rect 99350 80920 99360 80990
rect 99140 80880 99360 80920
rect 99140 80810 99150 80880
rect 99350 80810 99360 80880
rect 99140 80760 99360 80810
rect 99640 80990 99860 81040
rect 99640 80920 99650 80990
rect 99850 80920 99860 80990
rect 99640 80880 99860 80920
rect 99640 80810 99650 80880
rect 99850 80810 99860 80880
rect 99640 80760 99860 80810
rect 100140 80990 100360 81040
rect 100140 80920 100150 80990
rect 100350 80920 100360 80990
rect 100140 80880 100360 80920
rect 100140 80810 100150 80880
rect 100350 80810 100360 80880
rect 100140 80760 100360 80810
rect -83500 80750 100500 80760
rect -83500 80550 -83480 80750
rect -83410 80550 -83090 80750
rect -83020 80550 -82980 80750
rect -82910 80550 -82590 80750
rect -82520 80550 -82480 80750
rect -82410 80550 -82090 80750
rect -82020 80550 -81980 80750
rect -81910 80550 -81590 80750
rect -81520 80550 -81480 80750
rect -81410 80550 -81090 80750
rect -81020 80550 -80980 80750
rect -80910 80550 -80590 80750
rect -80520 80550 -80480 80750
rect -80410 80550 -80090 80750
rect -80020 80550 -79980 80750
rect -79910 80550 -79590 80750
rect -79520 80550 -79480 80750
rect -79410 80550 -79090 80750
rect -79020 80550 -78980 80750
rect -78910 80550 -78590 80750
rect -78520 80550 -78480 80750
rect -78410 80550 -78090 80750
rect -78020 80550 -77980 80750
rect -77910 80550 -77590 80750
rect -77520 80550 -77480 80750
rect -77410 80550 -77090 80750
rect -77020 80550 -76980 80750
rect -76910 80550 -76590 80750
rect -76520 80550 -76480 80750
rect -76410 80550 -76090 80750
rect -76020 80550 -75980 80750
rect -75910 80550 -75590 80750
rect -75520 80550 -75480 80750
rect -75410 80550 -75090 80750
rect -75020 80550 -74980 80750
rect -74910 80550 -74590 80750
rect -74520 80550 -74480 80750
rect -74410 80550 -74090 80750
rect -74020 80550 -73980 80750
rect -73910 80550 -73590 80750
rect -73520 80550 -73480 80750
rect -73410 80550 -73090 80750
rect -73020 80550 -72980 80750
rect -72910 80550 -72590 80750
rect -72520 80550 -72480 80750
rect -72410 80550 -72090 80750
rect -72020 80550 -71980 80750
rect -71910 80550 -71590 80750
rect -71520 80550 -71480 80750
rect -71410 80550 -71090 80750
rect -71020 80550 -70980 80750
rect -70910 80550 -70590 80750
rect -70520 80550 -70480 80750
rect -70410 80550 -70090 80750
rect -70020 80550 -69980 80750
rect -69910 80550 -69590 80750
rect -69520 80550 -69480 80750
rect -69410 80550 -69090 80750
rect -69020 80550 -68980 80750
rect -68910 80550 -68590 80750
rect -68520 80550 -68480 80750
rect -68410 80550 -68090 80750
rect -68020 80550 -67980 80750
rect -67910 80550 -67590 80750
rect -67520 80550 -67480 80750
rect -67410 80550 -67090 80750
rect -67020 80550 -66980 80750
rect -66910 80550 -66590 80750
rect -66520 80550 -66480 80750
rect -66410 80550 -66090 80750
rect -66020 80550 -65980 80750
rect -65910 80550 -65590 80750
rect -65520 80550 -65480 80750
rect -65410 80550 -65090 80750
rect -65020 80550 -64980 80750
rect -64910 80550 -64590 80750
rect -64520 80550 -64480 80750
rect -64410 80550 -64090 80750
rect -64020 80550 -63980 80750
rect -63910 80550 -63590 80750
rect -63520 80550 -63480 80750
rect -63410 80550 -63090 80750
rect -63020 80550 -62980 80750
rect -62910 80550 -62590 80750
rect -62520 80550 -62480 80750
rect -62410 80550 -62090 80750
rect -62020 80550 -61980 80750
rect -61910 80550 -61590 80750
rect -61520 80550 -61480 80750
rect -61410 80550 -61090 80750
rect -61020 80550 -60980 80750
rect -60910 80550 -60590 80750
rect -60520 80550 -60480 80750
rect -60410 80550 -60090 80750
rect -60020 80550 -59980 80750
rect -59910 80550 -59590 80750
rect -59520 80550 -59480 80750
rect -59410 80550 -59090 80750
rect -59020 80550 -58980 80750
rect -58910 80550 -58590 80750
rect -58520 80550 -58480 80750
rect -58410 80550 -58090 80750
rect -58020 80550 -57980 80750
rect -57910 80550 -57590 80750
rect -57520 80550 -57480 80750
rect -57410 80550 -57090 80750
rect -57020 80550 -56980 80750
rect -56910 80550 -56590 80750
rect -56520 80550 -56480 80750
rect -56410 80550 -56090 80750
rect -56020 80550 -55980 80750
rect -55910 80550 -55590 80750
rect -55520 80550 -55480 80750
rect -55410 80550 -55090 80750
rect -55020 80550 -54980 80750
rect -54910 80550 -54590 80750
rect -54520 80550 -54480 80750
rect -54410 80550 -54090 80750
rect -54020 80550 -53980 80750
rect -53910 80550 -53590 80750
rect -53520 80550 -53480 80750
rect -53410 80550 -53090 80750
rect -53020 80550 -52980 80750
rect -52910 80550 -52590 80750
rect -52520 80550 -52480 80750
rect -52410 80550 -52090 80750
rect -52020 80550 -51980 80750
rect -51910 80550 -51590 80750
rect -51520 80550 -51480 80750
rect -51410 80550 -51090 80750
rect -51020 80550 -50980 80750
rect -50910 80550 -50590 80750
rect -50520 80550 -50480 80750
rect -50410 80550 -50090 80750
rect -50020 80550 -49980 80750
rect -49910 80550 -49590 80750
rect -49520 80550 -49480 80750
rect -49410 80550 -49090 80750
rect -49020 80550 -48980 80750
rect -48910 80550 -48590 80750
rect -48520 80550 -48480 80750
rect -48410 80550 -48090 80750
rect -48020 80550 -47980 80750
rect -47910 80550 -47590 80750
rect -47520 80550 -47480 80750
rect -47410 80550 -47090 80750
rect -47020 80550 -46980 80750
rect -46910 80550 -46590 80750
rect -46520 80550 -46480 80750
rect -46410 80550 -46090 80750
rect -46020 80550 -45980 80750
rect -45910 80550 -45590 80750
rect -45520 80550 -45480 80750
rect -45410 80550 -45090 80750
rect -45020 80550 -44980 80750
rect -44910 80550 -44590 80750
rect -44520 80550 -44480 80750
rect -44410 80550 -44090 80750
rect -44020 80550 -43980 80750
rect -43910 80550 -43590 80750
rect -43520 80550 -43480 80750
rect -43410 80550 -43090 80750
rect -43020 80550 -42980 80750
rect -42910 80550 -42590 80750
rect -42520 80550 -42480 80750
rect -42410 80550 -42090 80750
rect -42020 80550 -41980 80750
rect -41910 80550 -41590 80750
rect -41520 80550 -41480 80750
rect -41410 80550 -41090 80750
rect -41020 80550 -40980 80750
rect -40910 80550 -40590 80750
rect -40520 80550 -40480 80750
rect -40410 80550 -40090 80750
rect -40020 80550 -39980 80750
rect -39910 80550 -39590 80750
rect -39520 80550 -39480 80750
rect -39410 80550 -39090 80750
rect -39020 80550 -38980 80750
rect -38910 80550 -38590 80750
rect -38520 80550 -38480 80750
rect -38410 80550 -38090 80750
rect -38020 80550 -37980 80750
rect -37910 80550 -37590 80750
rect -37520 80550 -37480 80750
rect -37410 80550 -37090 80750
rect -37020 80550 -36980 80750
rect -36910 80550 -36590 80750
rect -36520 80550 -36480 80750
rect -36410 80550 -36090 80750
rect -36020 80550 -35980 80750
rect -35910 80550 -35590 80750
rect -35520 80550 -35480 80750
rect -35410 80550 -35090 80750
rect -35020 80550 -34980 80750
rect -34910 80550 -34590 80750
rect -34520 80550 -34480 80750
rect -34410 80550 -34090 80750
rect -34020 80550 -33980 80750
rect -33910 80550 -33590 80750
rect -33520 80550 -33480 80750
rect -33410 80550 -33090 80750
rect -33020 80550 -32980 80750
rect -32910 80550 -32590 80750
rect -32520 80550 -32480 80750
rect -32410 80550 -32090 80750
rect -32020 80550 -31980 80750
rect -31910 80550 -31590 80750
rect -31520 80550 -31480 80750
rect -31410 80550 -31090 80750
rect -31020 80550 -30980 80750
rect -30910 80550 -30590 80750
rect -30520 80550 -30480 80750
rect -30410 80550 -30090 80750
rect -30020 80550 -29980 80750
rect -29910 80550 -29590 80750
rect -29520 80550 -29480 80750
rect -29410 80550 -29090 80750
rect -29020 80550 -28980 80750
rect -28910 80550 -28590 80750
rect -28520 80550 -28480 80750
rect -28410 80550 -28090 80750
rect -28020 80550 -27980 80750
rect -27910 80550 -27590 80750
rect -27520 80550 -27480 80750
rect -27410 80550 -27090 80750
rect -27020 80550 -26980 80750
rect -26910 80550 -26590 80750
rect -26520 80550 -26480 80750
rect -26410 80550 -26090 80750
rect -26020 80550 -25980 80750
rect -25910 80550 -25590 80750
rect -25520 80550 -25480 80750
rect -25410 80550 -25090 80750
rect -25020 80550 -24980 80750
rect -24910 80550 -24590 80750
rect -24520 80550 -24480 80750
rect -24410 80550 -24090 80750
rect -24020 80550 -23980 80750
rect -23910 80550 -23590 80750
rect -23520 80550 -23480 80750
rect -23410 80550 -23090 80750
rect -23020 80550 -22980 80750
rect -22910 80550 -22590 80750
rect -22520 80550 -22480 80750
rect -22410 80550 -22090 80750
rect -22020 80550 -21980 80750
rect -21910 80550 -21590 80750
rect -21520 80550 -21480 80750
rect -21410 80550 -21090 80750
rect -21020 80550 -20980 80750
rect -20910 80550 -20590 80750
rect -20520 80550 -20480 80750
rect -20410 80550 -20090 80750
rect -20020 80550 -19980 80750
rect -19910 80550 -19590 80750
rect -19520 80550 -19480 80750
rect -19410 80550 -19090 80750
rect -19020 80550 -18980 80750
rect -18910 80550 -18590 80750
rect -18520 80550 -18480 80750
rect -18410 80550 -18090 80750
rect -18020 80550 -17980 80750
rect -17910 80550 -17590 80750
rect -17520 80550 -17480 80750
rect -17410 80550 -17090 80750
rect -17020 80550 -16980 80750
rect -16910 80550 -16590 80750
rect -16520 80550 -16480 80750
rect -16410 80550 -16090 80750
rect -16020 80550 -15980 80750
rect -15910 80550 -15590 80750
rect -15520 80550 -15480 80750
rect -15410 80550 -15090 80750
rect -15020 80550 -14980 80750
rect -14910 80550 -14590 80750
rect -14520 80550 -14480 80750
rect -14410 80550 -14090 80750
rect -14020 80550 -13980 80750
rect -13910 80550 -13590 80750
rect -13520 80550 -13480 80750
rect -13410 80550 -13090 80750
rect -13020 80550 -12980 80750
rect -12910 80550 -12590 80750
rect -12520 80550 -12480 80750
rect -12410 80550 -12090 80750
rect -12020 80550 -11980 80750
rect -11910 80550 -11590 80750
rect -11520 80550 -11480 80750
rect -11410 80550 -11090 80750
rect -11020 80550 -10980 80750
rect -10910 80550 -10590 80750
rect -10520 80550 -10480 80750
rect -10410 80550 -10090 80750
rect -10020 80550 -9980 80750
rect -9910 80550 -9590 80750
rect -9520 80550 -9480 80750
rect -9410 80550 -9090 80750
rect -9020 80550 -8980 80750
rect -8910 80550 -8590 80750
rect -8520 80550 -8480 80750
rect -8410 80550 -8090 80750
rect -8020 80550 -7980 80750
rect -7910 80550 -7590 80750
rect -7520 80550 -7480 80750
rect -7410 80550 -7090 80750
rect -7020 80550 -6980 80750
rect -6910 80550 -6590 80750
rect -6520 80550 -6480 80750
rect -6410 80550 -6090 80750
rect -6020 80550 -5980 80750
rect -5910 80550 -5590 80750
rect -5520 80550 -5480 80750
rect -5410 80550 -5090 80750
rect -5020 80550 -4980 80750
rect -4910 80550 -4590 80750
rect -4520 80550 -4480 80750
rect -4410 80550 -4090 80750
rect -4020 80550 -3980 80750
rect -3910 80550 -3590 80750
rect -3520 80550 -3480 80750
rect -3410 80550 -3090 80750
rect -3020 80550 -2980 80750
rect -2910 80550 -2590 80750
rect -2520 80550 -2480 80750
rect -2410 80550 -2090 80750
rect -2020 80550 -1980 80750
rect -1910 80550 -1590 80750
rect -1520 80550 -1480 80750
rect -1410 80550 -1090 80750
rect -1020 80550 -980 80750
rect -910 80550 -590 80750
rect -520 80550 -480 80750
rect -410 80550 -90 80750
rect -20 80550 20 80750
rect 90 80550 410 80750
rect 480 80550 520 80750
rect 590 80550 910 80750
rect 980 80550 1020 80750
rect 1090 80550 1410 80750
rect 1480 80550 1520 80750
rect 1590 80550 1910 80750
rect 1980 80550 2020 80750
rect 2090 80550 2410 80750
rect 2480 80550 2520 80750
rect 2590 80550 2910 80750
rect 2980 80550 3020 80750
rect 3090 80550 3410 80750
rect 3480 80550 3520 80750
rect 3590 80550 3910 80750
rect 3980 80550 4020 80750
rect 4090 80550 4410 80750
rect 4480 80550 4520 80750
rect 4590 80550 4910 80750
rect 4980 80550 5020 80750
rect 5090 80550 5410 80750
rect 5480 80550 5520 80750
rect 5590 80550 5910 80750
rect 5980 80550 6020 80750
rect 6090 80550 6410 80750
rect 6480 80550 6520 80750
rect 6590 80550 6910 80750
rect 6980 80550 7020 80750
rect 7090 80550 7410 80750
rect 7480 80550 7520 80750
rect 7590 80550 7910 80750
rect 7980 80550 8020 80750
rect 8090 80550 8410 80750
rect 8480 80550 8520 80750
rect 8590 80550 8910 80750
rect 8980 80550 9020 80750
rect 9090 80550 9410 80750
rect 9480 80550 9520 80750
rect 9590 80550 9910 80750
rect 9980 80550 10020 80750
rect 10090 80550 10410 80750
rect 10480 80550 10520 80750
rect 10590 80550 10910 80750
rect 10980 80550 11020 80750
rect 11090 80550 11410 80750
rect 11480 80550 11520 80750
rect 11590 80550 11910 80750
rect 11980 80550 12020 80750
rect 12090 80550 12410 80750
rect 12480 80550 12520 80750
rect 12590 80550 12910 80750
rect 12980 80550 13020 80750
rect 13090 80550 13410 80750
rect 13480 80550 13520 80750
rect 13590 80550 13910 80750
rect 13980 80550 14020 80750
rect 14090 80550 14410 80750
rect 14480 80550 14520 80750
rect 14590 80550 14910 80750
rect 14980 80550 15020 80750
rect 15090 80550 15410 80750
rect 15480 80550 15520 80750
rect 15590 80550 15910 80750
rect 15980 80550 16020 80750
rect 16090 80550 16410 80750
rect 16480 80550 16520 80750
rect 16590 80550 16910 80750
rect 16980 80550 17020 80750
rect 17090 80550 17410 80750
rect 17480 80550 17520 80750
rect 17590 80550 17910 80750
rect 17980 80550 18020 80750
rect 18090 80550 18410 80750
rect 18480 80550 18520 80750
rect 18590 80550 18910 80750
rect 18980 80550 19020 80750
rect 19090 80550 19410 80750
rect 19480 80550 19520 80750
rect 19590 80550 19910 80750
rect 19980 80550 20020 80750
rect 20090 80550 20410 80750
rect 20480 80550 20520 80750
rect 20590 80550 20910 80750
rect 20980 80550 21020 80750
rect 21090 80550 21410 80750
rect 21480 80550 21520 80750
rect 21590 80550 21910 80750
rect 21980 80550 22020 80750
rect 22090 80550 22410 80750
rect 22480 80550 22520 80750
rect 22590 80550 22910 80750
rect 22980 80550 23020 80750
rect 23090 80550 23410 80750
rect 23480 80550 23520 80750
rect 23590 80550 23910 80750
rect 23980 80550 24020 80750
rect 24090 80550 24410 80750
rect 24480 80550 24520 80750
rect 24590 80550 24910 80750
rect 24980 80550 25020 80750
rect 25090 80550 25410 80750
rect 25480 80550 25520 80750
rect 25590 80550 25910 80750
rect 25980 80550 26020 80750
rect 26090 80550 26410 80750
rect 26480 80550 26520 80750
rect 26590 80550 26910 80750
rect 26980 80550 27020 80750
rect 27090 80550 27410 80750
rect 27480 80550 27520 80750
rect 27590 80550 27910 80750
rect 27980 80550 28020 80750
rect 28090 80550 28410 80750
rect 28480 80550 28520 80750
rect 28590 80550 28910 80750
rect 28980 80550 29020 80750
rect 29090 80550 29410 80750
rect 29480 80550 29520 80750
rect 29590 80550 29910 80750
rect 29980 80550 30020 80750
rect 30090 80550 30410 80750
rect 30480 80550 30520 80750
rect 30590 80550 30910 80750
rect 30980 80550 31020 80750
rect 31090 80550 31410 80750
rect 31480 80550 31520 80750
rect 31590 80550 31910 80750
rect 31980 80550 32020 80750
rect 32090 80550 32410 80750
rect 32480 80550 32520 80750
rect 32590 80550 32910 80750
rect 32980 80550 33020 80750
rect 33090 80550 33410 80750
rect 33480 80550 33520 80750
rect 33590 80550 33910 80750
rect 33980 80550 34020 80750
rect 34090 80550 34410 80750
rect 34480 80550 34520 80750
rect 34590 80550 34910 80750
rect 34980 80550 35020 80750
rect 35090 80550 35410 80750
rect 35480 80550 35520 80750
rect 35590 80550 35910 80750
rect 35980 80550 36020 80750
rect 36090 80550 36410 80750
rect 36480 80550 36520 80750
rect 36590 80550 36910 80750
rect 36980 80550 37020 80750
rect 37090 80550 37410 80750
rect 37480 80550 37520 80750
rect 37590 80550 37910 80750
rect 37980 80550 38020 80750
rect 38090 80550 38410 80750
rect 38480 80550 38520 80750
rect 38590 80550 38910 80750
rect 38980 80550 39020 80750
rect 39090 80550 39410 80750
rect 39480 80550 39520 80750
rect 39590 80550 39910 80750
rect 39980 80550 40020 80750
rect 40090 80550 40410 80750
rect 40480 80550 40520 80750
rect 40590 80550 40910 80750
rect 40980 80550 41020 80750
rect 41090 80550 41410 80750
rect 41480 80550 41520 80750
rect 41590 80550 41910 80750
rect 41980 80550 42020 80750
rect 42090 80550 42410 80750
rect 42480 80550 42520 80750
rect 42590 80550 42910 80750
rect 42980 80550 43020 80750
rect 43090 80550 43410 80750
rect 43480 80550 43520 80750
rect 43590 80550 43910 80750
rect 43980 80550 44020 80750
rect 44090 80550 44410 80750
rect 44480 80550 44520 80750
rect 44590 80550 44910 80750
rect 44980 80550 45020 80750
rect 45090 80550 45410 80750
rect 45480 80550 45520 80750
rect 45590 80550 45910 80750
rect 45980 80550 46020 80750
rect 46090 80550 46410 80750
rect 46480 80550 46520 80750
rect 46590 80550 46910 80750
rect 46980 80550 47020 80750
rect 47090 80550 47410 80750
rect 47480 80550 47520 80750
rect 47590 80550 47910 80750
rect 47980 80550 48020 80750
rect 48090 80550 48410 80750
rect 48480 80550 48520 80750
rect 48590 80550 48910 80750
rect 48980 80550 49020 80750
rect 49090 80550 49410 80750
rect 49480 80550 49520 80750
rect 49590 80550 49910 80750
rect 49980 80550 50020 80750
rect 50090 80550 50410 80750
rect 50480 80550 50520 80750
rect 50590 80550 50910 80750
rect 50980 80550 51020 80750
rect 51090 80550 51410 80750
rect 51480 80550 51520 80750
rect 51590 80550 51910 80750
rect 51980 80550 52020 80750
rect 52090 80550 52410 80750
rect 52480 80550 52520 80750
rect 52590 80550 52910 80750
rect 52980 80550 53020 80750
rect 53090 80550 53410 80750
rect 53480 80550 53520 80750
rect 53590 80550 53910 80750
rect 53980 80550 54020 80750
rect 54090 80550 54410 80750
rect 54480 80550 54520 80750
rect 54590 80550 54910 80750
rect 54980 80550 55020 80750
rect 55090 80550 55410 80750
rect 55480 80550 55520 80750
rect 55590 80550 55910 80750
rect 55980 80550 56020 80750
rect 56090 80550 56410 80750
rect 56480 80550 56520 80750
rect 56590 80550 56910 80750
rect 56980 80550 57020 80750
rect 57090 80550 57410 80750
rect 57480 80550 57520 80750
rect 57590 80550 57910 80750
rect 57980 80550 58020 80750
rect 58090 80550 58410 80750
rect 58480 80550 58520 80750
rect 58590 80550 58910 80750
rect 58980 80550 59020 80750
rect 59090 80550 59410 80750
rect 59480 80550 59520 80750
rect 59590 80550 59910 80750
rect 59980 80550 60020 80750
rect 60090 80550 60410 80750
rect 60480 80550 60520 80750
rect 60590 80550 60910 80750
rect 60980 80550 61020 80750
rect 61090 80550 61410 80750
rect 61480 80550 61520 80750
rect 61590 80550 61910 80750
rect 61980 80550 62020 80750
rect 62090 80550 62410 80750
rect 62480 80550 62520 80750
rect 62590 80550 62910 80750
rect 62980 80550 63020 80750
rect 63090 80550 63410 80750
rect 63480 80550 63520 80750
rect 63590 80550 63910 80750
rect 63980 80550 64020 80750
rect 64090 80550 64410 80750
rect 64480 80550 64520 80750
rect 64590 80550 64910 80750
rect 64980 80550 65020 80750
rect 65090 80550 65410 80750
rect 65480 80550 65520 80750
rect 65590 80550 65910 80750
rect 65980 80550 66020 80750
rect 66090 80550 66410 80750
rect 66480 80550 66520 80750
rect 66590 80550 66910 80750
rect 66980 80550 67020 80750
rect 67090 80550 67410 80750
rect 67480 80550 67520 80750
rect 67590 80550 67910 80750
rect 67980 80550 68020 80750
rect 68090 80550 68410 80750
rect 68480 80550 68520 80750
rect 68590 80550 68910 80750
rect 68980 80550 69020 80750
rect 69090 80550 69410 80750
rect 69480 80550 69520 80750
rect 69590 80550 69910 80750
rect 69980 80550 70020 80750
rect 70090 80550 70410 80750
rect 70480 80550 70520 80750
rect 70590 80550 70910 80750
rect 70980 80550 71020 80750
rect 71090 80550 71410 80750
rect 71480 80550 71520 80750
rect 71590 80550 71910 80750
rect 71980 80550 72020 80750
rect 72090 80550 72410 80750
rect 72480 80550 72520 80750
rect 72590 80550 72910 80750
rect 72980 80550 73020 80750
rect 73090 80550 73410 80750
rect 73480 80550 73520 80750
rect 73590 80550 73910 80750
rect 73980 80550 74020 80750
rect 74090 80550 74410 80750
rect 74480 80550 74520 80750
rect 74590 80550 74910 80750
rect 74980 80550 75020 80750
rect 75090 80550 75410 80750
rect 75480 80550 75520 80750
rect 75590 80550 75910 80750
rect 75980 80550 76020 80750
rect 76090 80550 76410 80750
rect 76480 80550 76520 80750
rect 76590 80550 76910 80750
rect 76980 80550 77020 80750
rect 77090 80550 77410 80750
rect 77480 80550 77520 80750
rect 77590 80550 77910 80750
rect 77980 80550 78020 80750
rect 78090 80550 78410 80750
rect 78480 80550 78520 80750
rect 78590 80550 78910 80750
rect 78980 80550 79020 80750
rect 79090 80550 79410 80750
rect 79480 80550 79520 80750
rect 79590 80550 79910 80750
rect 79980 80550 80020 80750
rect 80090 80550 80410 80750
rect 80480 80550 80520 80750
rect 80590 80550 80910 80750
rect 80980 80550 81020 80750
rect 81090 80550 81410 80750
rect 81480 80550 81520 80750
rect 81590 80550 81910 80750
rect 81980 80550 82020 80750
rect 82090 80550 82410 80750
rect 82480 80550 82520 80750
rect 82590 80550 82910 80750
rect 82980 80550 83020 80750
rect 83090 80550 83410 80750
rect 83480 80550 83520 80750
rect 83590 80550 83910 80750
rect 83980 80550 84020 80750
rect 84090 80550 84410 80750
rect 84480 80550 84520 80750
rect 84590 80550 84910 80750
rect 84980 80550 85020 80750
rect 85090 80550 85410 80750
rect 85480 80550 85520 80750
rect 85590 80550 85910 80750
rect 85980 80550 86020 80750
rect 86090 80550 86410 80750
rect 86480 80550 86520 80750
rect 86590 80550 86910 80750
rect 86980 80550 87020 80750
rect 87090 80550 87410 80750
rect 87480 80550 87520 80750
rect 87590 80550 87910 80750
rect 87980 80550 88020 80750
rect 88090 80550 88410 80750
rect 88480 80550 88520 80750
rect 88590 80550 88910 80750
rect 88980 80550 89020 80750
rect 89090 80550 89410 80750
rect 89480 80550 89520 80750
rect 89590 80550 89910 80750
rect 89980 80550 90020 80750
rect 90090 80550 90410 80750
rect 90480 80550 90520 80750
rect 90590 80550 90910 80750
rect 90980 80550 91020 80750
rect 91090 80550 91410 80750
rect 91480 80550 91520 80750
rect 91590 80550 91910 80750
rect 91980 80550 92020 80750
rect 92090 80550 92410 80750
rect 92480 80550 92520 80750
rect 92590 80550 92910 80750
rect 92980 80550 93020 80750
rect 93090 80550 93410 80750
rect 93480 80550 93520 80750
rect 93590 80550 93910 80750
rect 93980 80550 94020 80750
rect 94090 80550 94410 80750
rect 94480 80550 94520 80750
rect 94590 80550 94910 80750
rect 94980 80550 95020 80750
rect 95090 80550 95410 80750
rect 95480 80550 95520 80750
rect 95590 80550 95910 80750
rect 95980 80550 96020 80750
rect 96090 80550 96410 80750
rect 96480 80550 96520 80750
rect 96590 80550 96910 80750
rect 96980 80550 97020 80750
rect 97090 80550 97410 80750
rect 97480 80550 97520 80750
rect 97590 80550 97910 80750
rect 97980 80550 98020 80750
rect 98090 80550 98410 80750
rect 98480 80550 98520 80750
rect 98590 80550 98910 80750
rect 98980 80550 99020 80750
rect 99090 80550 99410 80750
rect 99480 80550 99520 80750
rect 99590 80550 99910 80750
rect 99980 80550 100020 80750
rect 100090 80550 100410 80750
rect 100480 80550 100500 80750
rect -83500 80540 100500 80550
rect -83360 80490 -83140 80540
rect -83360 80420 -83350 80490
rect -83150 80420 -83140 80490
rect -83360 80380 -83140 80420
rect -83360 80310 -83350 80380
rect -83150 80310 -83140 80380
rect -83360 80260 -83140 80310
rect -82860 80490 -82640 80540
rect -82860 80420 -82850 80490
rect -82650 80420 -82640 80490
rect -82860 80380 -82640 80420
rect -82860 80310 -82850 80380
rect -82650 80310 -82640 80380
rect -82860 80260 -82640 80310
rect -82360 80490 -82140 80540
rect -82360 80420 -82350 80490
rect -82150 80420 -82140 80490
rect -82360 80380 -82140 80420
rect -82360 80310 -82350 80380
rect -82150 80310 -82140 80380
rect -82360 80260 -82140 80310
rect -81860 80490 -81640 80540
rect -81860 80420 -81850 80490
rect -81650 80420 -81640 80490
rect -81860 80380 -81640 80420
rect -81860 80310 -81850 80380
rect -81650 80310 -81640 80380
rect -81860 80260 -81640 80310
rect -81360 80490 -81140 80540
rect -81360 80420 -81350 80490
rect -81150 80420 -81140 80490
rect -81360 80380 -81140 80420
rect -81360 80310 -81350 80380
rect -81150 80310 -81140 80380
rect -81360 80260 -81140 80310
rect -80860 80490 -80640 80540
rect -80860 80420 -80850 80490
rect -80650 80420 -80640 80490
rect -80860 80380 -80640 80420
rect -80860 80310 -80850 80380
rect -80650 80310 -80640 80380
rect -80860 80260 -80640 80310
rect -80360 80490 -80140 80540
rect -80360 80420 -80350 80490
rect -80150 80420 -80140 80490
rect -80360 80380 -80140 80420
rect -80360 80310 -80350 80380
rect -80150 80310 -80140 80380
rect -80360 80260 -80140 80310
rect -79860 80490 -79640 80540
rect -79860 80420 -79850 80490
rect -79650 80420 -79640 80490
rect -79860 80380 -79640 80420
rect -79860 80310 -79850 80380
rect -79650 80310 -79640 80380
rect -79860 80260 -79640 80310
rect -79360 80490 -79140 80540
rect -79360 80420 -79350 80490
rect -79150 80420 -79140 80490
rect -79360 80380 -79140 80420
rect -79360 80310 -79350 80380
rect -79150 80310 -79140 80380
rect -79360 80260 -79140 80310
rect -78860 80490 -78640 80540
rect -78860 80420 -78850 80490
rect -78650 80420 -78640 80490
rect -78860 80380 -78640 80420
rect -78860 80310 -78850 80380
rect -78650 80310 -78640 80380
rect -78860 80260 -78640 80310
rect -78360 80490 -78140 80540
rect -78360 80420 -78350 80490
rect -78150 80420 -78140 80490
rect -78360 80380 -78140 80420
rect -78360 80310 -78350 80380
rect -78150 80310 -78140 80380
rect -78360 80260 -78140 80310
rect -77860 80490 -77640 80540
rect -77860 80420 -77850 80490
rect -77650 80420 -77640 80490
rect -77860 80380 -77640 80420
rect -77860 80310 -77850 80380
rect -77650 80310 -77640 80380
rect -77860 80260 -77640 80310
rect -77360 80490 -77140 80540
rect -77360 80420 -77350 80490
rect -77150 80420 -77140 80490
rect -77360 80380 -77140 80420
rect -77360 80310 -77350 80380
rect -77150 80310 -77140 80380
rect -77360 80260 -77140 80310
rect -76860 80490 -76640 80540
rect -76860 80420 -76850 80490
rect -76650 80420 -76640 80490
rect -76860 80380 -76640 80420
rect -76860 80310 -76850 80380
rect -76650 80310 -76640 80380
rect -76860 80260 -76640 80310
rect -76360 80490 -76140 80540
rect -76360 80420 -76350 80490
rect -76150 80420 -76140 80490
rect -76360 80380 -76140 80420
rect -76360 80310 -76350 80380
rect -76150 80310 -76140 80380
rect -76360 80260 -76140 80310
rect -75860 80490 -75640 80540
rect -75860 80420 -75850 80490
rect -75650 80420 -75640 80490
rect -75860 80380 -75640 80420
rect -75860 80310 -75850 80380
rect -75650 80310 -75640 80380
rect -75860 80260 -75640 80310
rect -75360 80490 -75140 80540
rect -75360 80420 -75350 80490
rect -75150 80420 -75140 80490
rect -75360 80380 -75140 80420
rect -75360 80310 -75350 80380
rect -75150 80310 -75140 80380
rect -75360 80260 -75140 80310
rect -74860 80490 -74640 80540
rect -74860 80420 -74850 80490
rect -74650 80420 -74640 80490
rect -74860 80380 -74640 80420
rect -74860 80310 -74850 80380
rect -74650 80310 -74640 80380
rect -74860 80260 -74640 80310
rect -74360 80490 -74140 80540
rect -74360 80420 -74350 80490
rect -74150 80420 -74140 80490
rect -74360 80380 -74140 80420
rect -74360 80310 -74350 80380
rect -74150 80310 -74140 80380
rect -74360 80260 -74140 80310
rect -73860 80490 -73640 80540
rect -73860 80420 -73850 80490
rect -73650 80420 -73640 80490
rect -73860 80380 -73640 80420
rect -73860 80310 -73850 80380
rect -73650 80310 -73640 80380
rect -73860 80260 -73640 80310
rect -73360 80490 -73140 80540
rect -73360 80420 -73350 80490
rect -73150 80420 -73140 80490
rect -73360 80380 -73140 80420
rect -73360 80310 -73350 80380
rect -73150 80310 -73140 80380
rect -73360 80260 -73140 80310
rect -72860 80490 -72640 80540
rect -72860 80420 -72850 80490
rect -72650 80420 -72640 80490
rect -72860 80380 -72640 80420
rect -72860 80310 -72850 80380
rect -72650 80310 -72640 80380
rect -72860 80260 -72640 80310
rect -72360 80490 -72140 80540
rect -72360 80420 -72350 80490
rect -72150 80420 -72140 80490
rect -72360 80380 -72140 80420
rect -72360 80310 -72350 80380
rect -72150 80310 -72140 80380
rect -72360 80260 -72140 80310
rect -71860 80490 -71640 80540
rect -71860 80420 -71850 80490
rect -71650 80420 -71640 80490
rect -71860 80380 -71640 80420
rect -71860 80310 -71850 80380
rect -71650 80310 -71640 80380
rect -71860 80260 -71640 80310
rect -71360 80490 -71140 80540
rect -71360 80420 -71350 80490
rect -71150 80420 -71140 80490
rect -71360 80380 -71140 80420
rect -71360 80310 -71350 80380
rect -71150 80310 -71140 80380
rect -71360 80260 -71140 80310
rect -70860 80490 -70640 80540
rect -70860 80420 -70850 80490
rect -70650 80420 -70640 80490
rect -70860 80380 -70640 80420
rect -70860 80310 -70850 80380
rect -70650 80310 -70640 80380
rect -70860 80260 -70640 80310
rect -70360 80490 -70140 80540
rect -70360 80420 -70350 80490
rect -70150 80420 -70140 80490
rect -70360 80380 -70140 80420
rect -70360 80310 -70350 80380
rect -70150 80310 -70140 80380
rect -70360 80260 -70140 80310
rect -69860 80490 -69640 80540
rect -69860 80420 -69850 80490
rect -69650 80420 -69640 80490
rect -69860 80380 -69640 80420
rect -69860 80310 -69850 80380
rect -69650 80310 -69640 80380
rect -69860 80260 -69640 80310
rect -69360 80490 -69140 80540
rect -69360 80420 -69350 80490
rect -69150 80420 -69140 80490
rect -69360 80380 -69140 80420
rect -69360 80310 -69350 80380
rect -69150 80310 -69140 80380
rect -69360 80260 -69140 80310
rect -68860 80490 -68640 80540
rect -68860 80420 -68850 80490
rect -68650 80420 -68640 80490
rect -68860 80380 -68640 80420
rect -68860 80310 -68850 80380
rect -68650 80310 -68640 80380
rect -68860 80260 -68640 80310
rect -68360 80490 -68140 80540
rect -68360 80420 -68350 80490
rect -68150 80420 -68140 80490
rect -68360 80380 -68140 80420
rect -68360 80310 -68350 80380
rect -68150 80310 -68140 80380
rect -68360 80260 -68140 80310
rect -67860 80490 -67640 80540
rect -67860 80420 -67850 80490
rect -67650 80420 -67640 80490
rect -67860 80380 -67640 80420
rect -67860 80310 -67850 80380
rect -67650 80310 -67640 80380
rect -67860 80260 -67640 80310
rect -67360 80490 -67140 80540
rect -67360 80420 -67350 80490
rect -67150 80420 -67140 80490
rect -67360 80380 -67140 80420
rect -67360 80310 -67350 80380
rect -67150 80310 -67140 80380
rect -67360 80260 -67140 80310
rect -66860 80490 -66640 80540
rect -66860 80420 -66850 80490
rect -66650 80420 -66640 80490
rect -66860 80380 -66640 80420
rect -66860 80310 -66850 80380
rect -66650 80310 -66640 80380
rect -66860 80260 -66640 80310
rect -66360 80490 -66140 80540
rect -66360 80420 -66350 80490
rect -66150 80420 -66140 80490
rect -66360 80380 -66140 80420
rect -66360 80310 -66350 80380
rect -66150 80310 -66140 80380
rect -66360 80260 -66140 80310
rect -65860 80490 -65640 80540
rect -65860 80420 -65850 80490
rect -65650 80420 -65640 80490
rect -65860 80380 -65640 80420
rect -65860 80310 -65850 80380
rect -65650 80310 -65640 80380
rect -65860 80260 -65640 80310
rect -65360 80490 -65140 80540
rect -65360 80420 -65350 80490
rect -65150 80420 -65140 80490
rect -65360 80380 -65140 80420
rect -65360 80310 -65350 80380
rect -65150 80310 -65140 80380
rect -65360 80260 -65140 80310
rect -64860 80490 -64640 80540
rect -64860 80420 -64850 80490
rect -64650 80420 -64640 80490
rect -64860 80380 -64640 80420
rect -64860 80310 -64850 80380
rect -64650 80310 -64640 80380
rect -64860 80260 -64640 80310
rect -64360 80490 -64140 80540
rect -64360 80420 -64350 80490
rect -64150 80420 -64140 80490
rect -64360 80380 -64140 80420
rect -64360 80310 -64350 80380
rect -64150 80310 -64140 80380
rect -64360 80260 -64140 80310
rect -63860 80490 -63640 80540
rect -63860 80420 -63850 80490
rect -63650 80420 -63640 80490
rect -63860 80380 -63640 80420
rect -63860 80310 -63850 80380
rect -63650 80310 -63640 80380
rect -63860 80260 -63640 80310
rect -63360 80490 -63140 80540
rect -63360 80420 -63350 80490
rect -63150 80420 -63140 80490
rect -63360 80380 -63140 80420
rect -63360 80310 -63350 80380
rect -63150 80310 -63140 80380
rect -63360 80260 -63140 80310
rect -62860 80490 -62640 80540
rect -62860 80420 -62850 80490
rect -62650 80420 -62640 80490
rect -62860 80380 -62640 80420
rect -62860 80310 -62850 80380
rect -62650 80310 -62640 80380
rect -62860 80260 -62640 80310
rect -62360 80490 -62140 80540
rect -62360 80420 -62350 80490
rect -62150 80420 -62140 80490
rect -62360 80380 -62140 80420
rect -62360 80310 -62350 80380
rect -62150 80310 -62140 80380
rect -62360 80260 -62140 80310
rect -61860 80490 -61640 80540
rect -61860 80420 -61850 80490
rect -61650 80420 -61640 80490
rect -61860 80380 -61640 80420
rect -61860 80310 -61850 80380
rect -61650 80310 -61640 80380
rect -61860 80260 -61640 80310
rect -61360 80490 -61140 80540
rect -61360 80420 -61350 80490
rect -61150 80420 -61140 80490
rect -61360 80380 -61140 80420
rect -61360 80310 -61350 80380
rect -61150 80310 -61140 80380
rect -61360 80260 -61140 80310
rect -60860 80490 -60640 80540
rect -60860 80420 -60850 80490
rect -60650 80420 -60640 80490
rect -60860 80380 -60640 80420
rect -60860 80310 -60850 80380
rect -60650 80310 -60640 80380
rect -60860 80260 -60640 80310
rect -60360 80490 -60140 80540
rect -60360 80420 -60350 80490
rect -60150 80420 -60140 80490
rect -60360 80380 -60140 80420
rect -60360 80310 -60350 80380
rect -60150 80310 -60140 80380
rect -60360 80260 -60140 80310
rect -59860 80490 -59640 80540
rect -59860 80420 -59850 80490
rect -59650 80420 -59640 80490
rect -59860 80380 -59640 80420
rect -59860 80310 -59850 80380
rect -59650 80310 -59640 80380
rect -59860 80260 -59640 80310
rect -59360 80490 -59140 80540
rect -59360 80420 -59350 80490
rect -59150 80420 -59140 80490
rect -59360 80380 -59140 80420
rect -59360 80310 -59350 80380
rect -59150 80310 -59140 80380
rect -59360 80260 -59140 80310
rect -58860 80490 -58640 80540
rect -58860 80420 -58850 80490
rect -58650 80420 -58640 80490
rect -58860 80380 -58640 80420
rect -58860 80310 -58850 80380
rect -58650 80310 -58640 80380
rect -58860 80260 -58640 80310
rect -58360 80490 -58140 80540
rect -58360 80420 -58350 80490
rect -58150 80420 -58140 80490
rect -58360 80380 -58140 80420
rect -58360 80310 -58350 80380
rect -58150 80310 -58140 80380
rect -58360 80260 -58140 80310
rect -57860 80490 -57640 80540
rect -57860 80420 -57850 80490
rect -57650 80420 -57640 80490
rect -57860 80380 -57640 80420
rect -57860 80310 -57850 80380
rect -57650 80310 -57640 80380
rect -57860 80260 -57640 80310
rect -57360 80490 -57140 80540
rect -57360 80420 -57350 80490
rect -57150 80420 -57140 80490
rect -57360 80380 -57140 80420
rect -57360 80310 -57350 80380
rect -57150 80310 -57140 80380
rect -57360 80260 -57140 80310
rect -56860 80490 -56640 80540
rect -56860 80420 -56850 80490
rect -56650 80420 -56640 80490
rect -56860 80380 -56640 80420
rect -56860 80310 -56850 80380
rect -56650 80310 -56640 80380
rect -56860 80260 -56640 80310
rect -56360 80490 -56140 80540
rect -56360 80420 -56350 80490
rect -56150 80420 -56140 80490
rect -56360 80380 -56140 80420
rect -56360 80310 -56350 80380
rect -56150 80310 -56140 80380
rect -56360 80260 -56140 80310
rect -55860 80490 -55640 80540
rect -55860 80420 -55850 80490
rect -55650 80420 -55640 80490
rect -55860 80380 -55640 80420
rect -55860 80310 -55850 80380
rect -55650 80310 -55640 80380
rect -55860 80260 -55640 80310
rect -55360 80490 -55140 80540
rect -55360 80420 -55350 80490
rect -55150 80420 -55140 80490
rect -55360 80380 -55140 80420
rect -55360 80310 -55350 80380
rect -55150 80310 -55140 80380
rect -55360 80260 -55140 80310
rect -54860 80490 -54640 80540
rect -54860 80420 -54850 80490
rect -54650 80420 -54640 80490
rect -54860 80380 -54640 80420
rect -54860 80310 -54850 80380
rect -54650 80310 -54640 80380
rect -54860 80260 -54640 80310
rect -54360 80490 -54140 80540
rect -54360 80420 -54350 80490
rect -54150 80420 -54140 80490
rect -54360 80380 -54140 80420
rect -54360 80310 -54350 80380
rect -54150 80310 -54140 80380
rect -54360 80260 -54140 80310
rect -53860 80490 -53640 80540
rect -53860 80420 -53850 80490
rect -53650 80420 -53640 80490
rect -53860 80380 -53640 80420
rect -53860 80310 -53850 80380
rect -53650 80310 -53640 80380
rect -53860 80260 -53640 80310
rect -53360 80490 -53140 80540
rect -53360 80420 -53350 80490
rect -53150 80420 -53140 80490
rect -53360 80380 -53140 80420
rect -53360 80310 -53350 80380
rect -53150 80310 -53140 80380
rect -53360 80260 -53140 80310
rect -52860 80490 -52640 80540
rect -52860 80420 -52850 80490
rect -52650 80420 -52640 80490
rect -52860 80380 -52640 80420
rect -52860 80310 -52850 80380
rect -52650 80310 -52640 80380
rect -52860 80260 -52640 80310
rect -52360 80490 -52140 80540
rect -52360 80420 -52350 80490
rect -52150 80420 -52140 80490
rect -52360 80380 -52140 80420
rect -52360 80310 -52350 80380
rect -52150 80310 -52140 80380
rect -52360 80260 -52140 80310
rect -51860 80490 -51640 80540
rect -51860 80420 -51850 80490
rect -51650 80420 -51640 80490
rect -51860 80380 -51640 80420
rect -51860 80310 -51850 80380
rect -51650 80310 -51640 80380
rect -51860 80260 -51640 80310
rect -51360 80490 -51140 80540
rect -51360 80420 -51350 80490
rect -51150 80420 -51140 80490
rect -51360 80380 -51140 80420
rect -51360 80310 -51350 80380
rect -51150 80310 -51140 80380
rect -51360 80260 -51140 80310
rect -50860 80490 -50640 80540
rect -50860 80420 -50850 80490
rect -50650 80420 -50640 80490
rect -50860 80380 -50640 80420
rect -50860 80310 -50850 80380
rect -50650 80310 -50640 80380
rect -50860 80260 -50640 80310
rect -50360 80490 -50140 80540
rect -50360 80420 -50350 80490
rect -50150 80420 -50140 80490
rect -50360 80380 -50140 80420
rect -50360 80310 -50350 80380
rect -50150 80310 -50140 80380
rect -50360 80260 -50140 80310
rect -49860 80490 -49640 80540
rect -49860 80420 -49850 80490
rect -49650 80420 -49640 80490
rect -49860 80380 -49640 80420
rect -49860 80310 -49850 80380
rect -49650 80310 -49640 80380
rect -49860 80260 -49640 80310
rect -49360 80490 -49140 80540
rect -49360 80420 -49350 80490
rect -49150 80420 -49140 80490
rect -49360 80380 -49140 80420
rect -49360 80310 -49350 80380
rect -49150 80310 -49140 80380
rect -49360 80260 -49140 80310
rect -48860 80490 -48640 80540
rect -48860 80420 -48850 80490
rect -48650 80420 -48640 80490
rect -48860 80380 -48640 80420
rect -48860 80310 -48850 80380
rect -48650 80310 -48640 80380
rect -48860 80260 -48640 80310
rect -48360 80490 -48140 80540
rect -48360 80420 -48350 80490
rect -48150 80420 -48140 80490
rect -48360 80380 -48140 80420
rect -48360 80310 -48350 80380
rect -48150 80310 -48140 80380
rect -48360 80260 -48140 80310
rect -47860 80490 -47640 80540
rect -47860 80420 -47850 80490
rect -47650 80420 -47640 80490
rect -47860 80380 -47640 80420
rect -47860 80310 -47850 80380
rect -47650 80310 -47640 80380
rect -47860 80260 -47640 80310
rect -47360 80490 -47140 80540
rect -47360 80420 -47350 80490
rect -47150 80420 -47140 80490
rect -47360 80380 -47140 80420
rect -47360 80310 -47350 80380
rect -47150 80310 -47140 80380
rect -47360 80260 -47140 80310
rect -46860 80490 -46640 80540
rect -46860 80420 -46850 80490
rect -46650 80420 -46640 80490
rect -46860 80380 -46640 80420
rect -46860 80310 -46850 80380
rect -46650 80310 -46640 80380
rect -46860 80260 -46640 80310
rect -46360 80490 -46140 80540
rect -46360 80420 -46350 80490
rect -46150 80420 -46140 80490
rect -46360 80380 -46140 80420
rect -46360 80310 -46350 80380
rect -46150 80310 -46140 80380
rect -46360 80260 -46140 80310
rect -45860 80490 -45640 80540
rect -45860 80420 -45850 80490
rect -45650 80420 -45640 80490
rect -45860 80380 -45640 80420
rect -45860 80310 -45850 80380
rect -45650 80310 -45640 80380
rect -45860 80260 -45640 80310
rect -45360 80490 -45140 80540
rect -45360 80420 -45350 80490
rect -45150 80420 -45140 80490
rect -45360 80380 -45140 80420
rect -45360 80310 -45350 80380
rect -45150 80310 -45140 80380
rect -45360 80260 -45140 80310
rect -44860 80490 -44640 80540
rect -44860 80420 -44850 80490
rect -44650 80420 -44640 80490
rect -44860 80380 -44640 80420
rect -44860 80310 -44850 80380
rect -44650 80310 -44640 80380
rect -44860 80260 -44640 80310
rect -44360 80490 -44140 80540
rect -44360 80420 -44350 80490
rect -44150 80420 -44140 80490
rect -44360 80380 -44140 80420
rect -44360 80310 -44350 80380
rect -44150 80310 -44140 80380
rect -44360 80260 -44140 80310
rect -43860 80490 -43640 80540
rect -43860 80420 -43850 80490
rect -43650 80420 -43640 80490
rect -43860 80380 -43640 80420
rect -43860 80310 -43850 80380
rect -43650 80310 -43640 80380
rect -43860 80260 -43640 80310
rect -43360 80490 -43140 80540
rect -43360 80420 -43350 80490
rect -43150 80420 -43140 80490
rect -43360 80380 -43140 80420
rect -43360 80310 -43350 80380
rect -43150 80310 -43140 80380
rect -43360 80260 -43140 80310
rect -42860 80490 -42640 80540
rect -42860 80420 -42850 80490
rect -42650 80420 -42640 80490
rect -42860 80380 -42640 80420
rect -42860 80310 -42850 80380
rect -42650 80310 -42640 80380
rect -42860 80260 -42640 80310
rect -42360 80490 -42140 80540
rect -42360 80420 -42350 80490
rect -42150 80420 -42140 80490
rect -42360 80380 -42140 80420
rect -42360 80310 -42350 80380
rect -42150 80310 -42140 80380
rect -42360 80260 -42140 80310
rect -41860 80490 -41640 80540
rect -41860 80420 -41850 80490
rect -41650 80420 -41640 80490
rect -41860 80380 -41640 80420
rect -41860 80310 -41850 80380
rect -41650 80310 -41640 80380
rect -41860 80260 -41640 80310
rect -41360 80490 -41140 80540
rect -41360 80420 -41350 80490
rect -41150 80420 -41140 80490
rect -41360 80380 -41140 80420
rect -41360 80310 -41350 80380
rect -41150 80310 -41140 80380
rect -41360 80260 -41140 80310
rect -40860 80490 -40640 80540
rect -40860 80420 -40850 80490
rect -40650 80420 -40640 80490
rect -40860 80380 -40640 80420
rect -40860 80310 -40850 80380
rect -40650 80310 -40640 80380
rect -40860 80260 -40640 80310
rect -40360 80490 -40140 80540
rect -40360 80420 -40350 80490
rect -40150 80420 -40140 80490
rect -40360 80380 -40140 80420
rect -40360 80310 -40350 80380
rect -40150 80310 -40140 80380
rect -40360 80260 -40140 80310
rect -39860 80490 -39640 80540
rect -39860 80420 -39850 80490
rect -39650 80420 -39640 80490
rect -39860 80380 -39640 80420
rect -39860 80310 -39850 80380
rect -39650 80310 -39640 80380
rect -39860 80260 -39640 80310
rect -39360 80490 -39140 80540
rect -39360 80420 -39350 80490
rect -39150 80420 -39140 80490
rect -39360 80380 -39140 80420
rect -39360 80310 -39350 80380
rect -39150 80310 -39140 80380
rect -39360 80260 -39140 80310
rect -38860 80490 -38640 80540
rect -38860 80420 -38850 80490
rect -38650 80420 -38640 80490
rect -38860 80380 -38640 80420
rect -38860 80310 -38850 80380
rect -38650 80310 -38640 80380
rect -38860 80260 -38640 80310
rect -38360 80490 -38140 80540
rect -38360 80420 -38350 80490
rect -38150 80420 -38140 80490
rect -38360 80380 -38140 80420
rect -38360 80310 -38350 80380
rect -38150 80310 -38140 80380
rect -38360 80260 -38140 80310
rect -37860 80490 -37640 80540
rect -37860 80420 -37850 80490
rect -37650 80420 -37640 80490
rect -37860 80380 -37640 80420
rect -37860 80310 -37850 80380
rect -37650 80310 -37640 80380
rect -37860 80260 -37640 80310
rect -37360 80490 -37140 80540
rect -37360 80420 -37350 80490
rect -37150 80420 -37140 80490
rect -37360 80380 -37140 80420
rect -37360 80310 -37350 80380
rect -37150 80310 -37140 80380
rect -37360 80260 -37140 80310
rect -36860 80490 -36640 80540
rect -36860 80420 -36850 80490
rect -36650 80420 -36640 80490
rect -36860 80380 -36640 80420
rect -36860 80310 -36850 80380
rect -36650 80310 -36640 80380
rect -36860 80260 -36640 80310
rect -36360 80490 -36140 80540
rect -36360 80420 -36350 80490
rect -36150 80420 -36140 80490
rect -36360 80380 -36140 80420
rect -36360 80310 -36350 80380
rect -36150 80310 -36140 80380
rect -36360 80260 -36140 80310
rect -35860 80490 -35640 80540
rect -35860 80420 -35850 80490
rect -35650 80420 -35640 80490
rect -35860 80380 -35640 80420
rect -35860 80310 -35850 80380
rect -35650 80310 -35640 80380
rect -35860 80260 -35640 80310
rect -35360 80490 -35140 80540
rect -35360 80420 -35350 80490
rect -35150 80420 -35140 80490
rect -35360 80380 -35140 80420
rect -35360 80310 -35350 80380
rect -35150 80310 -35140 80380
rect -35360 80260 -35140 80310
rect -34860 80490 -34640 80540
rect -34860 80420 -34850 80490
rect -34650 80420 -34640 80490
rect -34860 80380 -34640 80420
rect -34860 80310 -34850 80380
rect -34650 80310 -34640 80380
rect -34860 80260 -34640 80310
rect -34360 80490 -34140 80540
rect -34360 80420 -34350 80490
rect -34150 80420 -34140 80490
rect -34360 80380 -34140 80420
rect -34360 80310 -34350 80380
rect -34150 80310 -34140 80380
rect -34360 80260 -34140 80310
rect -33860 80490 -33640 80540
rect -33860 80420 -33850 80490
rect -33650 80420 -33640 80490
rect -33860 80380 -33640 80420
rect -33860 80310 -33850 80380
rect -33650 80310 -33640 80380
rect -33860 80260 -33640 80310
rect -33360 80490 -33140 80540
rect -33360 80420 -33350 80490
rect -33150 80420 -33140 80490
rect -33360 80380 -33140 80420
rect -33360 80310 -33350 80380
rect -33150 80310 -33140 80380
rect -33360 80260 -33140 80310
rect -32860 80490 -32640 80540
rect -32860 80420 -32850 80490
rect -32650 80420 -32640 80490
rect -32860 80380 -32640 80420
rect -32860 80310 -32850 80380
rect -32650 80310 -32640 80380
rect -32860 80260 -32640 80310
rect -32360 80490 -32140 80540
rect -32360 80420 -32350 80490
rect -32150 80420 -32140 80490
rect -32360 80380 -32140 80420
rect -32360 80310 -32350 80380
rect -32150 80310 -32140 80380
rect -32360 80260 -32140 80310
rect -31860 80490 -31640 80540
rect -31860 80420 -31850 80490
rect -31650 80420 -31640 80490
rect -31860 80380 -31640 80420
rect -31860 80310 -31850 80380
rect -31650 80310 -31640 80380
rect -31860 80260 -31640 80310
rect -31360 80490 -31140 80540
rect -31360 80420 -31350 80490
rect -31150 80420 -31140 80490
rect -31360 80380 -31140 80420
rect -31360 80310 -31350 80380
rect -31150 80310 -31140 80380
rect -31360 80260 -31140 80310
rect -30860 80490 -30640 80540
rect -30860 80420 -30850 80490
rect -30650 80420 -30640 80490
rect -30860 80380 -30640 80420
rect -30860 80310 -30850 80380
rect -30650 80310 -30640 80380
rect -30860 80260 -30640 80310
rect -30360 80490 -30140 80540
rect -30360 80420 -30350 80490
rect -30150 80420 -30140 80490
rect -30360 80380 -30140 80420
rect -30360 80310 -30350 80380
rect -30150 80310 -30140 80380
rect -30360 80260 -30140 80310
rect -29860 80490 -29640 80540
rect -29860 80420 -29850 80490
rect -29650 80420 -29640 80490
rect -29860 80380 -29640 80420
rect -29860 80310 -29850 80380
rect -29650 80310 -29640 80380
rect -29860 80260 -29640 80310
rect -29360 80490 -29140 80540
rect -29360 80420 -29350 80490
rect -29150 80420 -29140 80490
rect -29360 80380 -29140 80420
rect -29360 80310 -29350 80380
rect -29150 80310 -29140 80380
rect -29360 80260 -29140 80310
rect -28860 80490 -28640 80540
rect -28860 80420 -28850 80490
rect -28650 80420 -28640 80490
rect -28860 80380 -28640 80420
rect -28860 80310 -28850 80380
rect -28650 80310 -28640 80380
rect -28860 80260 -28640 80310
rect -28360 80490 -28140 80540
rect -28360 80420 -28350 80490
rect -28150 80420 -28140 80490
rect -28360 80380 -28140 80420
rect -28360 80310 -28350 80380
rect -28150 80310 -28140 80380
rect -28360 80260 -28140 80310
rect -27860 80490 -27640 80540
rect -27860 80420 -27850 80490
rect -27650 80420 -27640 80490
rect -27860 80380 -27640 80420
rect -27860 80310 -27850 80380
rect -27650 80310 -27640 80380
rect -27860 80260 -27640 80310
rect -27360 80490 -27140 80540
rect -27360 80420 -27350 80490
rect -27150 80420 -27140 80490
rect -27360 80380 -27140 80420
rect -27360 80310 -27350 80380
rect -27150 80310 -27140 80380
rect -27360 80260 -27140 80310
rect -26860 80490 -26640 80540
rect -26860 80420 -26850 80490
rect -26650 80420 -26640 80490
rect -26860 80380 -26640 80420
rect -26860 80310 -26850 80380
rect -26650 80310 -26640 80380
rect -26860 80260 -26640 80310
rect -26360 80490 -26140 80540
rect -26360 80420 -26350 80490
rect -26150 80420 -26140 80490
rect -26360 80380 -26140 80420
rect -26360 80310 -26350 80380
rect -26150 80310 -26140 80380
rect -26360 80260 -26140 80310
rect -25860 80490 -25640 80540
rect -25860 80420 -25850 80490
rect -25650 80420 -25640 80490
rect -25860 80380 -25640 80420
rect -25860 80310 -25850 80380
rect -25650 80310 -25640 80380
rect -25860 80260 -25640 80310
rect -25360 80490 -25140 80540
rect -25360 80420 -25350 80490
rect -25150 80420 -25140 80490
rect -25360 80380 -25140 80420
rect -25360 80310 -25350 80380
rect -25150 80310 -25140 80380
rect -25360 80260 -25140 80310
rect -24860 80490 -24640 80540
rect -24860 80420 -24850 80490
rect -24650 80420 -24640 80490
rect -24860 80380 -24640 80420
rect -24860 80310 -24850 80380
rect -24650 80310 -24640 80380
rect -24860 80260 -24640 80310
rect -24360 80490 -24140 80540
rect -24360 80420 -24350 80490
rect -24150 80420 -24140 80490
rect -24360 80380 -24140 80420
rect -24360 80310 -24350 80380
rect -24150 80310 -24140 80380
rect -24360 80260 -24140 80310
rect -23860 80490 -23640 80540
rect -23860 80420 -23850 80490
rect -23650 80420 -23640 80490
rect -23860 80380 -23640 80420
rect -23860 80310 -23850 80380
rect -23650 80310 -23640 80380
rect -23860 80260 -23640 80310
rect -23360 80490 -23140 80540
rect -23360 80420 -23350 80490
rect -23150 80420 -23140 80490
rect -23360 80380 -23140 80420
rect -23360 80310 -23350 80380
rect -23150 80310 -23140 80380
rect -23360 80260 -23140 80310
rect -22860 80490 -22640 80540
rect -22860 80420 -22850 80490
rect -22650 80420 -22640 80490
rect -22860 80380 -22640 80420
rect -22860 80310 -22850 80380
rect -22650 80310 -22640 80380
rect -22860 80260 -22640 80310
rect -22360 80490 -22140 80540
rect -22360 80420 -22350 80490
rect -22150 80420 -22140 80490
rect -22360 80380 -22140 80420
rect -22360 80310 -22350 80380
rect -22150 80310 -22140 80380
rect -22360 80260 -22140 80310
rect -21860 80490 -21640 80540
rect -21860 80420 -21850 80490
rect -21650 80420 -21640 80490
rect -21860 80380 -21640 80420
rect -21860 80310 -21850 80380
rect -21650 80310 -21640 80380
rect -21860 80260 -21640 80310
rect -21360 80490 -21140 80540
rect -21360 80420 -21350 80490
rect -21150 80420 -21140 80490
rect -21360 80380 -21140 80420
rect -21360 80310 -21350 80380
rect -21150 80310 -21140 80380
rect -21360 80260 -21140 80310
rect -20860 80490 -20640 80540
rect -20860 80420 -20850 80490
rect -20650 80420 -20640 80490
rect -20860 80380 -20640 80420
rect -20860 80310 -20850 80380
rect -20650 80310 -20640 80380
rect -20860 80260 -20640 80310
rect -20360 80490 -20140 80540
rect -20360 80420 -20350 80490
rect -20150 80420 -20140 80490
rect -20360 80380 -20140 80420
rect -20360 80310 -20350 80380
rect -20150 80310 -20140 80380
rect -20360 80260 -20140 80310
rect -19860 80490 -19640 80540
rect -19860 80420 -19850 80490
rect -19650 80420 -19640 80490
rect -19860 80380 -19640 80420
rect -19860 80310 -19850 80380
rect -19650 80310 -19640 80380
rect -19860 80260 -19640 80310
rect -19360 80490 -19140 80540
rect -19360 80420 -19350 80490
rect -19150 80420 -19140 80490
rect -19360 80380 -19140 80420
rect -19360 80310 -19350 80380
rect -19150 80310 -19140 80380
rect -19360 80260 -19140 80310
rect -18860 80490 -18640 80540
rect -18860 80420 -18850 80490
rect -18650 80420 -18640 80490
rect -18860 80380 -18640 80420
rect -18860 80310 -18850 80380
rect -18650 80310 -18640 80380
rect -18860 80260 -18640 80310
rect -18360 80490 -18140 80540
rect -18360 80420 -18350 80490
rect -18150 80420 -18140 80490
rect -18360 80380 -18140 80420
rect -18360 80310 -18350 80380
rect -18150 80310 -18140 80380
rect -18360 80260 -18140 80310
rect -17860 80490 -17640 80540
rect -17860 80420 -17850 80490
rect -17650 80420 -17640 80490
rect -17860 80380 -17640 80420
rect -17860 80310 -17850 80380
rect -17650 80310 -17640 80380
rect -17860 80260 -17640 80310
rect -17360 80490 -17140 80540
rect -17360 80420 -17350 80490
rect -17150 80420 -17140 80490
rect -17360 80380 -17140 80420
rect -17360 80310 -17350 80380
rect -17150 80310 -17140 80380
rect -17360 80260 -17140 80310
rect -16860 80490 -16640 80540
rect -16860 80420 -16850 80490
rect -16650 80420 -16640 80490
rect -16860 80380 -16640 80420
rect -16860 80310 -16850 80380
rect -16650 80310 -16640 80380
rect -16860 80260 -16640 80310
rect -16360 80490 -16140 80540
rect -16360 80420 -16350 80490
rect -16150 80420 -16140 80490
rect -16360 80380 -16140 80420
rect -16360 80310 -16350 80380
rect -16150 80310 -16140 80380
rect -16360 80260 -16140 80310
rect -15860 80490 -15640 80540
rect -15860 80420 -15850 80490
rect -15650 80420 -15640 80490
rect -15860 80380 -15640 80420
rect -15860 80310 -15850 80380
rect -15650 80310 -15640 80380
rect -15860 80260 -15640 80310
rect -15360 80490 -15140 80540
rect -15360 80420 -15350 80490
rect -15150 80420 -15140 80490
rect -15360 80380 -15140 80420
rect -15360 80310 -15350 80380
rect -15150 80310 -15140 80380
rect -15360 80260 -15140 80310
rect -14860 80490 -14640 80540
rect -14860 80420 -14850 80490
rect -14650 80420 -14640 80490
rect -14860 80380 -14640 80420
rect -14860 80310 -14850 80380
rect -14650 80310 -14640 80380
rect -14860 80260 -14640 80310
rect -14360 80490 -14140 80540
rect -14360 80420 -14350 80490
rect -14150 80420 -14140 80490
rect -14360 80380 -14140 80420
rect -14360 80310 -14350 80380
rect -14150 80310 -14140 80380
rect -14360 80260 -14140 80310
rect -13860 80490 -13640 80540
rect -13860 80420 -13850 80490
rect -13650 80420 -13640 80490
rect -13860 80380 -13640 80420
rect -13860 80310 -13850 80380
rect -13650 80310 -13640 80380
rect -13860 80260 -13640 80310
rect -13360 80490 -13140 80540
rect -13360 80420 -13350 80490
rect -13150 80420 -13140 80490
rect -13360 80380 -13140 80420
rect -13360 80310 -13350 80380
rect -13150 80310 -13140 80380
rect -13360 80260 -13140 80310
rect -12860 80490 -12640 80540
rect -12860 80420 -12850 80490
rect -12650 80420 -12640 80490
rect -12860 80380 -12640 80420
rect -12860 80310 -12850 80380
rect -12650 80310 -12640 80380
rect -12860 80260 -12640 80310
rect -12360 80490 -12140 80540
rect -12360 80420 -12350 80490
rect -12150 80420 -12140 80490
rect -12360 80380 -12140 80420
rect -12360 80310 -12350 80380
rect -12150 80310 -12140 80380
rect -12360 80260 -12140 80310
rect -11860 80490 -11640 80540
rect -11860 80420 -11850 80490
rect -11650 80420 -11640 80490
rect -11860 80380 -11640 80420
rect -11860 80310 -11850 80380
rect -11650 80310 -11640 80380
rect -11860 80260 -11640 80310
rect -11360 80490 -11140 80540
rect -11360 80420 -11350 80490
rect -11150 80420 -11140 80490
rect -11360 80380 -11140 80420
rect -11360 80310 -11350 80380
rect -11150 80310 -11140 80380
rect -11360 80260 -11140 80310
rect -10860 80490 -10640 80540
rect -10860 80420 -10850 80490
rect -10650 80420 -10640 80490
rect -10860 80380 -10640 80420
rect -10860 80310 -10850 80380
rect -10650 80310 -10640 80380
rect -10860 80260 -10640 80310
rect -10360 80490 -10140 80540
rect -10360 80420 -10350 80490
rect -10150 80420 -10140 80490
rect -10360 80380 -10140 80420
rect -10360 80310 -10350 80380
rect -10150 80310 -10140 80380
rect -10360 80260 -10140 80310
rect -9860 80490 -9640 80540
rect -9860 80420 -9850 80490
rect -9650 80420 -9640 80490
rect -9860 80380 -9640 80420
rect -9860 80310 -9850 80380
rect -9650 80310 -9640 80380
rect -9860 80260 -9640 80310
rect -9360 80490 -9140 80540
rect -9360 80420 -9350 80490
rect -9150 80420 -9140 80490
rect -9360 80380 -9140 80420
rect -9360 80310 -9350 80380
rect -9150 80310 -9140 80380
rect -9360 80260 -9140 80310
rect -8860 80490 -8640 80540
rect -8860 80420 -8850 80490
rect -8650 80420 -8640 80490
rect -8860 80380 -8640 80420
rect -8860 80310 -8850 80380
rect -8650 80310 -8640 80380
rect -8860 80260 -8640 80310
rect -8360 80490 -8140 80540
rect -8360 80420 -8350 80490
rect -8150 80420 -8140 80490
rect -8360 80380 -8140 80420
rect -8360 80310 -8350 80380
rect -8150 80310 -8140 80380
rect -8360 80260 -8140 80310
rect -7860 80490 -7640 80540
rect -7860 80420 -7850 80490
rect -7650 80420 -7640 80490
rect -7860 80380 -7640 80420
rect -7860 80310 -7850 80380
rect -7650 80310 -7640 80380
rect -7860 80260 -7640 80310
rect -7360 80490 -7140 80540
rect -7360 80420 -7350 80490
rect -7150 80420 -7140 80490
rect -7360 80380 -7140 80420
rect -7360 80310 -7350 80380
rect -7150 80310 -7140 80380
rect -7360 80260 -7140 80310
rect -6860 80490 -6640 80540
rect -6860 80420 -6850 80490
rect -6650 80420 -6640 80490
rect -6860 80380 -6640 80420
rect -6860 80310 -6850 80380
rect -6650 80310 -6640 80380
rect -6860 80260 -6640 80310
rect -6360 80490 -6140 80540
rect -6360 80420 -6350 80490
rect -6150 80420 -6140 80490
rect -6360 80380 -6140 80420
rect -6360 80310 -6350 80380
rect -6150 80310 -6140 80380
rect -6360 80260 -6140 80310
rect -5860 80490 -5640 80540
rect -5860 80420 -5850 80490
rect -5650 80420 -5640 80490
rect -5860 80380 -5640 80420
rect -5860 80310 -5850 80380
rect -5650 80310 -5640 80380
rect -5860 80260 -5640 80310
rect -5360 80490 -5140 80540
rect -5360 80420 -5350 80490
rect -5150 80420 -5140 80490
rect -5360 80380 -5140 80420
rect -5360 80310 -5350 80380
rect -5150 80310 -5140 80380
rect -5360 80260 -5140 80310
rect -4860 80490 -4640 80540
rect -4860 80420 -4850 80490
rect -4650 80420 -4640 80490
rect -4860 80380 -4640 80420
rect -4860 80310 -4850 80380
rect -4650 80310 -4640 80380
rect -4860 80260 -4640 80310
rect -4360 80490 -4140 80540
rect -4360 80420 -4350 80490
rect -4150 80420 -4140 80490
rect -4360 80380 -4140 80420
rect -4360 80310 -4350 80380
rect -4150 80310 -4140 80380
rect -4360 80260 -4140 80310
rect -3860 80490 -3640 80540
rect -3860 80420 -3850 80490
rect -3650 80420 -3640 80490
rect -3860 80380 -3640 80420
rect -3860 80310 -3850 80380
rect -3650 80310 -3640 80380
rect -3860 80260 -3640 80310
rect -3360 80490 -3140 80540
rect -3360 80420 -3350 80490
rect -3150 80420 -3140 80490
rect -3360 80380 -3140 80420
rect -3360 80310 -3350 80380
rect -3150 80310 -3140 80380
rect -3360 80260 -3140 80310
rect -2860 80490 -2640 80540
rect -2860 80420 -2850 80490
rect -2650 80420 -2640 80490
rect -2860 80380 -2640 80420
rect -2860 80310 -2850 80380
rect -2650 80310 -2640 80380
rect -2860 80260 -2640 80310
rect -2360 80490 -2140 80540
rect -2360 80420 -2350 80490
rect -2150 80420 -2140 80490
rect -2360 80380 -2140 80420
rect -2360 80310 -2350 80380
rect -2150 80310 -2140 80380
rect -2360 80260 -2140 80310
rect -1860 80490 -1640 80540
rect -1860 80420 -1850 80490
rect -1650 80420 -1640 80490
rect -1860 80380 -1640 80420
rect -1860 80310 -1850 80380
rect -1650 80310 -1640 80380
rect -1860 80260 -1640 80310
rect -1360 80490 -1140 80540
rect -1360 80420 -1350 80490
rect -1150 80420 -1140 80490
rect -1360 80380 -1140 80420
rect -1360 80310 -1350 80380
rect -1150 80310 -1140 80380
rect -1360 80260 -1140 80310
rect -860 80490 -640 80540
rect -860 80420 -850 80490
rect -650 80420 -640 80490
rect -860 80380 -640 80420
rect -860 80310 -850 80380
rect -650 80310 -640 80380
rect -860 80260 -640 80310
rect -360 80490 -140 80540
rect -360 80420 -350 80490
rect -150 80420 -140 80490
rect -360 80380 -140 80420
rect -360 80310 -350 80380
rect -150 80310 -140 80380
rect -360 80260 -140 80310
rect 140 80490 360 80540
rect 140 80420 150 80490
rect 350 80420 360 80490
rect 140 80380 360 80420
rect 140 80310 150 80380
rect 350 80310 360 80380
rect 140 80260 360 80310
rect 640 80490 860 80540
rect 640 80420 650 80490
rect 850 80420 860 80490
rect 640 80380 860 80420
rect 640 80310 650 80380
rect 850 80310 860 80380
rect 640 80260 860 80310
rect 1140 80490 1360 80540
rect 1140 80420 1150 80490
rect 1350 80420 1360 80490
rect 1140 80380 1360 80420
rect 1140 80310 1150 80380
rect 1350 80310 1360 80380
rect 1140 80260 1360 80310
rect 1640 80490 1860 80540
rect 1640 80420 1650 80490
rect 1850 80420 1860 80490
rect 1640 80380 1860 80420
rect 1640 80310 1650 80380
rect 1850 80310 1860 80380
rect 1640 80260 1860 80310
rect 2140 80490 2360 80540
rect 2140 80420 2150 80490
rect 2350 80420 2360 80490
rect 2140 80380 2360 80420
rect 2140 80310 2150 80380
rect 2350 80310 2360 80380
rect 2140 80260 2360 80310
rect 2640 80490 2860 80540
rect 2640 80420 2650 80490
rect 2850 80420 2860 80490
rect 2640 80380 2860 80420
rect 2640 80310 2650 80380
rect 2850 80310 2860 80380
rect 2640 80260 2860 80310
rect 3140 80490 3360 80540
rect 3140 80420 3150 80490
rect 3350 80420 3360 80490
rect 3140 80380 3360 80420
rect 3140 80310 3150 80380
rect 3350 80310 3360 80380
rect 3140 80260 3360 80310
rect 3640 80490 3860 80540
rect 3640 80420 3650 80490
rect 3850 80420 3860 80490
rect 3640 80380 3860 80420
rect 3640 80310 3650 80380
rect 3850 80310 3860 80380
rect 3640 80260 3860 80310
rect 4140 80490 4360 80540
rect 4140 80420 4150 80490
rect 4350 80420 4360 80490
rect 4140 80380 4360 80420
rect 4140 80310 4150 80380
rect 4350 80310 4360 80380
rect 4140 80260 4360 80310
rect 4640 80490 4860 80540
rect 4640 80420 4650 80490
rect 4850 80420 4860 80490
rect 4640 80380 4860 80420
rect 4640 80310 4650 80380
rect 4850 80310 4860 80380
rect 4640 80260 4860 80310
rect 5140 80490 5360 80540
rect 5140 80420 5150 80490
rect 5350 80420 5360 80490
rect 5140 80380 5360 80420
rect 5140 80310 5150 80380
rect 5350 80310 5360 80380
rect 5140 80260 5360 80310
rect 5640 80490 5860 80540
rect 5640 80420 5650 80490
rect 5850 80420 5860 80490
rect 5640 80380 5860 80420
rect 5640 80310 5650 80380
rect 5850 80310 5860 80380
rect 5640 80260 5860 80310
rect 6140 80490 6360 80540
rect 6140 80420 6150 80490
rect 6350 80420 6360 80490
rect 6140 80380 6360 80420
rect 6140 80310 6150 80380
rect 6350 80310 6360 80380
rect 6140 80260 6360 80310
rect 6640 80490 6860 80540
rect 6640 80420 6650 80490
rect 6850 80420 6860 80490
rect 6640 80380 6860 80420
rect 6640 80310 6650 80380
rect 6850 80310 6860 80380
rect 6640 80260 6860 80310
rect 7140 80490 7360 80540
rect 7140 80420 7150 80490
rect 7350 80420 7360 80490
rect 7140 80380 7360 80420
rect 7140 80310 7150 80380
rect 7350 80310 7360 80380
rect 7140 80260 7360 80310
rect 7640 80490 7860 80540
rect 7640 80420 7650 80490
rect 7850 80420 7860 80490
rect 7640 80380 7860 80420
rect 7640 80310 7650 80380
rect 7850 80310 7860 80380
rect 7640 80260 7860 80310
rect 8140 80490 8360 80540
rect 8140 80420 8150 80490
rect 8350 80420 8360 80490
rect 8140 80380 8360 80420
rect 8140 80310 8150 80380
rect 8350 80310 8360 80380
rect 8140 80260 8360 80310
rect 8640 80490 8860 80540
rect 8640 80420 8650 80490
rect 8850 80420 8860 80490
rect 8640 80380 8860 80420
rect 8640 80310 8650 80380
rect 8850 80310 8860 80380
rect 8640 80260 8860 80310
rect 9140 80490 9360 80540
rect 9140 80420 9150 80490
rect 9350 80420 9360 80490
rect 9140 80380 9360 80420
rect 9140 80310 9150 80380
rect 9350 80310 9360 80380
rect 9140 80260 9360 80310
rect 9640 80490 9860 80540
rect 9640 80420 9650 80490
rect 9850 80420 9860 80490
rect 9640 80380 9860 80420
rect 9640 80310 9650 80380
rect 9850 80310 9860 80380
rect 9640 80260 9860 80310
rect 10140 80490 10360 80540
rect 10140 80420 10150 80490
rect 10350 80420 10360 80490
rect 10140 80380 10360 80420
rect 10140 80310 10150 80380
rect 10350 80310 10360 80380
rect 10140 80260 10360 80310
rect 10640 80490 10860 80540
rect 10640 80420 10650 80490
rect 10850 80420 10860 80490
rect 10640 80380 10860 80420
rect 10640 80310 10650 80380
rect 10850 80310 10860 80380
rect 10640 80260 10860 80310
rect 11140 80490 11360 80540
rect 11140 80420 11150 80490
rect 11350 80420 11360 80490
rect 11140 80380 11360 80420
rect 11140 80310 11150 80380
rect 11350 80310 11360 80380
rect 11140 80260 11360 80310
rect 11640 80490 11860 80540
rect 11640 80420 11650 80490
rect 11850 80420 11860 80490
rect 11640 80380 11860 80420
rect 11640 80310 11650 80380
rect 11850 80310 11860 80380
rect 11640 80260 11860 80310
rect 12140 80490 12360 80540
rect 12140 80420 12150 80490
rect 12350 80420 12360 80490
rect 12140 80380 12360 80420
rect 12140 80310 12150 80380
rect 12350 80310 12360 80380
rect 12140 80260 12360 80310
rect 12640 80490 12860 80540
rect 12640 80420 12650 80490
rect 12850 80420 12860 80490
rect 12640 80380 12860 80420
rect 12640 80310 12650 80380
rect 12850 80310 12860 80380
rect 12640 80260 12860 80310
rect 13140 80490 13360 80540
rect 13140 80420 13150 80490
rect 13350 80420 13360 80490
rect 13140 80380 13360 80420
rect 13140 80310 13150 80380
rect 13350 80310 13360 80380
rect 13140 80260 13360 80310
rect 13640 80490 13860 80540
rect 13640 80420 13650 80490
rect 13850 80420 13860 80490
rect 13640 80380 13860 80420
rect 13640 80310 13650 80380
rect 13850 80310 13860 80380
rect 13640 80260 13860 80310
rect 14140 80490 14360 80540
rect 14140 80420 14150 80490
rect 14350 80420 14360 80490
rect 14140 80380 14360 80420
rect 14140 80310 14150 80380
rect 14350 80310 14360 80380
rect 14140 80260 14360 80310
rect 14640 80490 14860 80540
rect 14640 80420 14650 80490
rect 14850 80420 14860 80490
rect 14640 80380 14860 80420
rect 14640 80310 14650 80380
rect 14850 80310 14860 80380
rect 14640 80260 14860 80310
rect 15140 80490 15360 80540
rect 15140 80420 15150 80490
rect 15350 80420 15360 80490
rect 15140 80380 15360 80420
rect 15140 80310 15150 80380
rect 15350 80310 15360 80380
rect 15140 80260 15360 80310
rect 15640 80490 15860 80540
rect 15640 80420 15650 80490
rect 15850 80420 15860 80490
rect 15640 80380 15860 80420
rect 15640 80310 15650 80380
rect 15850 80310 15860 80380
rect 15640 80260 15860 80310
rect 16140 80490 16360 80540
rect 16140 80420 16150 80490
rect 16350 80420 16360 80490
rect 16140 80380 16360 80420
rect 16140 80310 16150 80380
rect 16350 80310 16360 80380
rect 16140 80260 16360 80310
rect 16640 80490 16860 80540
rect 16640 80420 16650 80490
rect 16850 80420 16860 80490
rect 16640 80380 16860 80420
rect 16640 80310 16650 80380
rect 16850 80310 16860 80380
rect 16640 80260 16860 80310
rect 17140 80490 17360 80540
rect 17140 80420 17150 80490
rect 17350 80420 17360 80490
rect 17140 80380 17360 80420
rect 17140 80310 17150 80380
rect 17350 80310 17360 80380
rect 17140 80260 17360 80310
rect 17640 80490 17860 80540
rect 17640 80420 17650 80490
rect 17850 80420 17860 80490
rect 17640 80380 17860 80420
rect 17640 80310 17650 80380
rect 17850 80310 17860 80380
rect 17640 80260 17860 80310
rect 18140 80490 18360 80540
rect 18140 80420 18150 80490
rect 18350 80420 18360 80490
rect 18140 80380 18360 80420
rect 18140 80310 18150 80380
rect 18350 80310 18360 80380
rect 18140 80260 18360 80310
rect 18640 80490 18860 80540
rect 18640 80420 18650 80490
rect 18850 80420 18860 80490
rect 18640 80380 18860 80420
rect 18640 80310 18650 80380
rect 18850 80310 18860 80380
rect 18640 80260 18860 80310
rect 19140 80490 19360 80540
rect 19140 80420 19150 80490
rect 19350 80420 19360 80490
rect 19140 80380 19360 80420
rect 19140 80310 19150 80380
rect 19350 80310 19360 80380
rect 19140 80260 19360 80310
rect 19640 80490 19860 80540
rect 19640 80420 19650 80490
rect 19850 80420 19860 80490
rect 19640 80380 19860 80420
rect 19640 80310 19650 80380
rect 19850 80310 19860 80380
rect 19640 80260 19860 80310
rect 20140 80490 20360 80540
rect 20140 80420 20150 80490
rect 20350 80420 20360 80490
rect 20140 80380 20360 80420
rect 20140 80310 20150 80380
rect 20350 80310 20360 80380
rect 20140 80260 20360 80310
rect 20640 80490 20860 80540
rect 20640 80420 20650 80490
rect 20850 80420 20860 80490
rect 20640 80380 20860 80420
rect 20640 80310 20650 80380
rect 20850 80310 20860 80380
rect 20640 80260 20860 80310
rect 21140 80490 21360 80540
rect 21140 80420 21150 80490
rect 21350 80420 21360 80490
rect 21140 80380 21360 80420
rect 21140 80310 21150 80380
rect 21350 80310 21360 80380
rect 21140 80260 21360 80310
rect 21640 80490 21860 80540
rect 21640 80420 21650 80490
rect 21850 80420 21860 80490
rect 21640 80380 21860 80420
rect 21640 80310 21650 80380
rect 21850 80310 21860 80380
rect 21640 80260 21860 80310
rect 22140 80490 22360 80540
rect 22140 80420 22150 80490
rect 22350 80420 22360 80490
rect 22140 80380 22360 80420
rect 22140 80310 22150 80380
rect 22350 80310 22360 80380
rect 22140 80260 22360 80310
rect 22640 80490 22860 80540
rect 22640 80420 22650 80490
rect 22850 80420 22860 80490
rect 22640 80380 22860 80420
rect 22640 80310 22650 80380
rect 22850 80310 22860 80380
rect 22640 80260 22860 80310
rect 23140 80490 23360 80540
rect 23140 80420 23150 80490
rect 23350 80420 23360 80490
rect 23140 80380 23360 80420
rect 23140 80310 23150 80380
rect 23350 80310 23360 80380
rect 23140 80260 23360 80310
rect 23640 80490 23860 80540
rect 23640 80420 23650 80490
rect 23850 80420 23860 80490
rect 23640 80380 23860 80420
rect 23640 80310 23650 80380
rect 23850 80310 23860 80380
rect 23640 80260 23860 80310
rect 24140 80490 24360 80540
rect 24140 80420 24150 80490
rect 24350 80420 24360 80490
rect 24140 80380 24360 80420
rect 24140 80310 24150 80380
rect 24350 80310 24360 80380
rect 24140 80260 24360 80310
rect 24640 80490 24860 80540
rect 24640 80420 24650 80490
rect 24850 80420 24860 80490
rect 24640 80380 24860 80420
rect 24640 80310 24650 80380
rect 24850 80310 24860 80380
rect 24640 80260 24860 80310
rect 25140 80490 25360 80540
rect 25140 80420 25150 80490
rect 25350 80420 25360 80490
rect 25140 80380 25360 80420
rect 25140 80310 25150 80380
rect 25350 80310 25360 80380
rect 25140 80260 25360 80310
rect 25640 80490 25860 80540
rect 25640 80420 25650 80490
rect 25850 80420 25860 80490
rect 25640 80380 25860 80420
rect 25640 80310 25650 80380
rect 25850 80310 25860 80380
rect 25640 80260 25860 80310
rect 26140 80490 26360 80540
rect 26140 80420 26150 80490
rect 26350 80420 26360 80490
rect 26140 80380 26360 80420
rect 26140 80310 26150 80380
rect 26350 80310 26360 80380
rect 26140 80260 26360 80310
rect 26640 80490 26860 80540
rect 26640 80420 26650 80490
rect 26850 80420 26860 80490
rect 26640 80380 26860 80420
rect 26640 80310 26650 80380
rect 26850 80310 26860 80380
rect 26640 80260 26860 80310
rect 27140 80490 27360 80540
rect 27140 80420 27150 80490
rect 27350 80420 27360 80490
rect 27140 80380 27360 80420
rect 27140 80310 27150 80380
rect 27350 80310 27360 80380
rect 27140 80260 27360 80310
rect 27640 80490 27860 80540
rect 27640 80420 27650 80490
rect 27850 80420 27860 80490
rect 27640 80380 27860 80420
rect 27640 80310 27650 80380
rect 27850 80310 27860 80380
rect 27640 80260 27860 80310
rect 28140 80490 28360 80540
rect 28140 80420 28150 80490
rect 28350 80420 28360 80490
rect 28140 80380 28360 80420
rect 28140 80310 28150 80380
rect 28350 80310 28360 80380
rect 28140 80260 28360 80310
rect 28640 80490 28860 80540
rect 28640 80420 28650 80490
rect 28850 80420 28860 80490
rect 28640 80380 28860 80420
rect 28640 80310 28650 80380
rect 28850 80310 28860 80380
rect 28640 80260 28860 80310
rect 29140 80490 29360 80540
rect 29140 80420 29150 80490
rect 29350 80420 29360 80490
rect 29140 80380 29360 80420
rect 29140 80310 29150 80380
rect 29350 80310 29360 80380
rect 29140 80260 29360 80310
rect 29640 80490 29860 80540
rect 29640 80420 29650 80490
rect 29850 80420 29860 80490
rect 29640 80380 29860 80420
rect 29640 80310 29650 80380
rect 29850 80310 29860 80380
rect 29640 80260 29860 80310
rect 30140 80490 30360 80540
rect 30140 80420 30150 80490
rect 30350 80420 30360 80490
rect 30140 80380 30360 80420
rect 30140 80310 30150 80380
rect 30350 80310 30360 80380
rect 30140 80260 30360 80310
rect 30640 80490 30860 80540
rect 30640 80420 30650 80490
rect 30850 80420 30860 80490
rect 30640 80380 30860 80420
rect 30640 80310 30650 80380
rect 30850 80310 30860 80380
rect 30640 80260 30860 80310
rect 31140 80490 31360 80540
rect 31140 80420 31150 80490
rect 31350 80420 31360 80490
rect 31140 80380 31360 80420
rect 31140 80310 31150 80380
rect 31350 80310 31360 80380
rect 31140 80260 31360 80310
rect 31640 80490 31860 80540
rect 31640 80420 31650 80490
rect 31850 80420 31860 80490
rect 31640 80380 31860 80420
rect 31640 80310 31650 80380
rect 31850 80310 31860 80380
rect 31640 80260 31860 80310
rect 32140 80490 32360 80540
rect 32140 80420 32150 80490
rect 32350 80420 32360 80490
rect 32140 80380 32360 80420
rect 32140 80310 32150 80380
rect 32350 80310 32360 80380
rect 32140 80260 32360 80310
rect 32640 80490 32860 80540
rect 32640 80420 32650 80490
rect 32850 80420 32860 80490
rect 32640 80380 32860 80420
rect 32640 80310 32650 80380
rect 32850 80310 32860 80380
rect 32640 80260 32860 80310
rect 33140 80490 33360 80540
rect 33140 80420 33150 80490
rect 33350 80420 33360 80490
rect 33140 80380 33360 80420
rect 33140 80310 33150 80380
rect 33350 80310 33360 80380
rect 33140 80260 33360 80310
rect 33640 80490 33860 80540
rect 33640 80420 33650 80490
rect 33850 80420 33860 80490
rect 33640 80380 33860 80420
rect 33640 80310 33650 80380
rect 33850 80310 33860 80380
rect 33640 80260 33860 80310
rect 34140 80490 34360 80540
rect 34140 80420 34150 80490
rect 34350 80420 34360 80490
rect 34140 80380 34360 80420
rect 34140 80310 34150 80380
rect 34350 80310 34360 80380
rect 34140 80260 34360 80310
rect 34640 80490 34860 80540
rect 34640 80420 34650 80490
rect 34850 80420 34860 80490
rect 34640 80380 34860 80420
rect 34640 80310 34650 80380
rect 34850 80310 34860 80380
rect 34640 80260 34860 80310
rect 35140 80490 35360 80540
rect 35140 80420 35150 80490
rect 35350 80420 35360 80490
rect 35140 80380 35360 80420
rect 35140 80310 35150 80380
rect 35350 80310 35360 80380
rect 35140 80260 35360 80310
rect 35640 80490 35860 80540
rect 35640 80420 35650 80490
rect 35850 80420 35860 80490
rect 35640 80380 35860 80420
rect 35640 80310 35650 80380
rect 35850 80310 35860 80380
rect 35640 80260 35860 80310
rect 36140 80490 36360 80540
rect 36140 80420 36150 80490
rect 36350 80420 36360 80490
rect 36140 80380 36360 80420
rect 36140 80310 36150 80380
rect 36350 80310 36360 80380
rect 36140 80260 36360 80310
rect 36640 80490 36860 80540
rect 36640 80420 36650 80490
rect 36850 80420 36860 80490
rect 36640 80380 36860 80420
rect 36640 80310 36650 80380
rect 36850 80310 36860 80380
rect 36640 80260 36860 80310
rect 37140 80490 37360 80540
rect 37140 80420 37150 80490
rect 37350 80420 37360 80490
rect 37140 80380 37360 80420
rect 37140 80310 37150 80380
rect 37350 80310 37360 80380
rect 37140 80260 37360 80310
rect 37640 80490 37860 80540
rect 37640 80420 37650 80490
rect 37850 80420 37860 80490
rect 37640 80380 37860 80420
rect 37640 80310 37650 80380
rect 37850 80310 37860 80380
rect 37640 80260 37860 80310
rect 38140 80490 38360 80540
rect 38140 80420 38150 80490
rect 38350 80420 38360 80490
rect 38140 80380 38360 80420
rect 38140 80310 38150 80380
rect 38350 80310 38360 80380
rect 38140 80260 38360 80310
rect 38640 80490 38860 80540
rect 38640 80420 38650 80490
rect 38850 80420 38860 80490
rect 38640 80380 38860 80420
rect 38640 80310 38650 80380
rect 38850 80310 38860 80380
rect 38640 80260 38860 80310
rect 39140 80490 39360 80540
rect 39140 80420 39150 80490
rect 39350 80420 39360 80490
rect 39140 80380 39360 80420
rect 39140 80310 39150 80380
rect 39350 80310 39360 80380
rect 39140 80260 39360 80310
rect 39640 80490 39860 80540
rect 39640 80420 39650 80490
rect 39850 80420 39860 80490
rect 39640 80380 39860 80420
rect 39640 80310 39650 80380
rect 39850 80310 39860 80380
rect 39640 80260 39860 80310
rect 40140 80490 40360 80540
rect 40140 80420 40150 80490
rect 40350 80420 40360 80490
rect 40140 80380 40360 80420
rect 40140 80310 40150 80380
rect 40350 80310 40360 80380
rect 40140 80260 40360 80310
rect 40640 80490 40860 80540
rect 40640 80420 40650 80490
rect 40850 80420 40860 80490
rect 40640 80380 40860 80420
rect 40640 80310 40650 80380
rect 40850 80310 40860 80380
rect 40640 80260 40860 80310
rect 41140 80490 41360 80540
rect 41140 80420 41150 80490
rect 41350 80420 41360 80490
rect 41140 80380 41360 80420
rect 41140 80310 41150 80380
rect 41350 80310 41360 80380
rect 41140 80260 41360 80310
rect 41640 80490 41860 80540
rect 41640 80420 41650 80490
rect 41850 80420 41860 80490
rect 41640 80380 41860 80420
rect 41640 80310 41650 80380
rect 41850 80310 41860 80380
rect 41640 80260 41860 80310
rect 42140 80490 42360 80540
rect 42140 80420 42150 80490
rect 42350 80420 42360 80490
rect 42140 80380 42360 80420
rect 42140 80310 42150 80380
rect 42350 80310 42360 80380
rect 42140 80260 42360 80310
rect 42640 80490 42860 80540
rect 42640 80420 42650 80490
rect 42850 80420 42860 80490
rect 42640 80380 42860 80420
rect 42640 80310 42650 80380
rect 42850 80310 42860 80380
rect 42640 80260 42860 80310
rect 43140 80490 43360 80540
rect 43140 80420 43150 80490
rect 43350 80420 43360 80490
rect 43140 80380 43360 80420
rect 43140 80310 43150 80380
rect 43350 80310 43360 80380
rect 43140 80260 43360 80310
rect 43640 80490 43860 80540
rect 43640 80420 43650 80490
rect 43850 80420 43860 80490
rect 43640 80380 43860 80420
rect 43640 80310 43650 80380
rect 43850 80310 43860 80380
rect 43640 80260 43860 80310
rect 44140 80490 44360 80540
rect 44140 80420 44150 80490
rect 44350 80420 44360 80490
rect 44140 80380 44360 80420
rect 44140 80310 44150 80380
rect 44350 80310 44360 80380
rect 44140 80260 44360 80310
rect 44640 80490 44860 80540
rect 44640 80420 44650 80490
rect 44850 80420 44860 80490
rect 44640 80380 44860 80420
rect 44640 80310 44650 80380
rect 44850 80310 44860 80380
rect 44640 80260 44860 80310
rect 45140 80490 45360 80540
rect 45140 80420 45150 80490
rect 45350 80420 45360 80490
rect 45140 80380 45360 80420
rect 45140 80310 45150 80380
rect 45350 80310 45360 80380
rect 45140 80260 45360 80310
rect 45640 80490 45860 80540
rect 45640 80420 45650 80490
rect 45850 80420 45860 80490
rect 45640 80380 45860 80420
rect 45640 80310 45650 80380
rect 45850 80310 45860 80380
rect 45640 80260 45860 80310
rect 46140 80490 46360 80540
rect 46140 80420 46150 80490
rect 46350 80420 46360 80490
rect 46140 80380 46360 80420
rect 46140 80310 46150 80380
rect 46350 80310 46360 80380
rect 46140 80260 46360 80310
rect 46640 80490 46860 80540
rect 46640 80420 46650 80490
rect 46850 80420 46860 80490
rect 46640 80380 46860 80420
rect 46640 80310 46650 80380
rect 46850 80310 46860 80380
rect 46640 80260 46860 80310
rect 47140 80490 47360 80540
rect 47140 80420 47150 80490
rect 47350 80420 47360 80490
rect 47140 80380 47360 80420
rect 47140 80310 47150 80380
rect 47350 80310 47360 80380
rect 47140 80260 47360 80310
rect 47640 80490 47860 80540
rect 47640 80420 47650 80490
rect 47850 80420 47860 80490
rect 47640 80380 47860 80420
rect 47640 80310 47650 80380
rect 47850 80310 47860 80380
rect 47640 80260 47860 80310
rect 48140 80490 48360 80540
rect 48140 80420 48150 80490
rect 48350 80420 48360 80490
rect 48140 80380 48360 80420
rect 48140 80310 48150 80380
rect 48350 80310 48360 80380
rect 48140 80260 48360 80310
rect 48640 80490 48860 80540
rect 48640 80420 48650 80490
rect 48850 80420 48860 80490
rect 48640 80380 48860 80420
rect 48640 80310 48650 80380
rect 48850 80310 48860 80380
rect 48640 80260 48860 80310
rect 49140 80490 49360 80540
rect 49140 80420 49150 80490
rect 49350 80420 49360 80490
rect 49140 80380 49360 80420
rect 49140 80310 49150 80380
rect 49350 80310 49360 80380
rect 49140 80260 49360 80310
rect 49640 80490 49860 80540
rect 49640 80420 49650 80490
rect 49850 80420 49860 80490
rect 49640 80380 49860 80420
rect 49640 80310 49650 80380
rect 49850 80310 49860 80380
rect 49640 80260 49860 80310
rect 50140 80490 50360 80540
rect 50140 80420 50150 80490
rect 50350 80420 50360 80490
rect 50140 80380 50360 80420
rect 50140 80310 50150 80380
rect 50350 80310 50360 80380
rect 50140 80260 50360 80310
rect 50640 80490 50860 80540
rect 50640 80420 50650 80490
rect 50850 80420 50860 80490
rect 50640 80380 50860 80420
rect 50640 80310 50650 80380
rect 50850 80310 50860 80380
rect 50640 80260 50860 80310
rect 51140 80490 51360 80540
rect 51140 80420 51150 80490
rect 51350 80420 51360 80490
rect 51140 80380 51360 80420
rect 51140 80310 51150 80380
rect 51350 80310 51360 80380
rect 51140 80260 51360 80310
rect 51640 80490 51860 80540
rect 51640 80420 51650 80490
rect 51850 80420 51860 80490
rect 51640 80380 51860 80420
rect 51640 80310 51650 80380
rect 51850 80310 51860 80380
rect 51640 80260 51860 80310
rect 52140 80490 52360 80540
rect 52140 80420 52150 80490
rect 52350 80420 52360 80490
rect 52140 80380 52360 80420
rect 52140 80310 52150 80380
rect 52350 80310 52360 80380
rect 52140 80260 52360 80310
rect 52640 80490 52860 80540
rect 52640 80420 52650 80490
rect 52850 80420 52860 80490
rect 52640 80380 52860 80420
rect 52640 80310 52650 80380
rect 52850 80310 52860 80380
rect 52640 80260 52860 80310
rect 53140 80490 53360 80540
rect 53140 80420 53150 80490
rect 53350 80420 53360 80490
rect 53140 80380 53360 80420
rect 53140 80310 53150 80380
rect 53350 80310 53360 80380
rect 53140 80260 53360 80310
rect 53640 80490 53860 80540
rect 53640 80420 53650 80490
rect 53850 80420 53860 80490
rect 53640 80380 53860 80420
rect 53640 80310 53650 80380
rect 53850 80310 53860 80380
rect 53640 80260 53860 80310
rect 54140 80490 54360 80540
rect 54140 80420 54150 80490
rect 54350 80420 54360 80490
rect 54140 80380 54360 80420
rect 54140 80310 54150 80380
rect 54350 80310 54360 80380
rect 54140 80260 54360 80310
rect 54640 80490 54860 80540
rect 54640 80420 54650 80490
rect 54850 80420 54860 80490
rect 54640 80380 54860 80420
rect 54640 80310 54650 80380
rect 54850 80310 54860 80380
rect 54640 80260 54860 80310
rect 55140 80490 55360 80540
rect 55140 80420 55150 80490
rect 55350 80420 55360 80490
rect 55140 80380 55360 80420
rect 55140 80310 55150 80380
rect 55350 80310 55360 80380
rect 55140 80260 55360 80310
rect 55640 80490 55860 80540
rect 55640 80420 55650 80490
rect 55850 80420 55860 80490
rect 55640 80380 55860 80420
rect 55640 80310 55650 80380
rect 55850 80310 55860 80380
rect 55640 80260 55860 80310
rect 56140 80490 56360 80540
rect 56140 80420 56150 80490
rect 56350 80420 56360 80490
rect 56140 80380 56360 80420
rect 56140 80310 56150 80380
rect 56350 80310 56360 80380
rect 56140 80260 56360 80310
rect 56640 80490 56860 80540
rect 56640 80420 56650 80490
rect 56850 80420 56860 80490
rect 56640 80380 56860 80420
rect 56640 80310 56650 80380
rect 56850 80310 56860 80380
rect 56640 80260 56860 80310
rect 57140 80490 57360 80540
rect 57140 80420 57150 80490
rect 57350 80420 57360 80490
rect 57140 80380 57360 80420
rect 57140 80310 57150 80380
rect 57350 80310 57360 80380
rect 57140 80260 57360 80310
rect 57640 80490 57860 80540
rect 57640 80420 57650 80490
rect 57850 80420 57860 80490
rect 57640 80380 57860 80420
rect 57640 80310 57650 80380
rect 57850 80310 57860 80380
rect 57640 80260 57860 80310
rect 58140 80490 58360 80540
rect 58140 80420 58150 80490
rect 58350 80420 58360 80490
rect 58140 80380 58360 80420
rect 58140 80310 58150 80380
rect 58350 80310 58360 80380
rect 58140 80260 58360 80310
rect 58640 80490 58860 80540
rect 58640 80420 58650 80490
rect 58850 80420 58860 80490
rect 58640 80380 58860 80420
rect 58640 80310 58650 80380
rect 58850 80310 58860 80380
rect 58640 80260 58860 80310
rect 59140 80490 59360 80540
rect 59140 80420 59150 80490
rect 59350 80420 59360 80490
rect 59140 80380 59360 80420
rect 59140 80310 59150 80380
rect 59350 80310 59360 80380
rect 59140 80260 59360 80310
rect 59640 80490 59860 80540
rect 59640 80420 59650 80490
rect 59850 80420 59860 80490
rect 59640 80380 59860 80420
rect 59640 80310 59650 80380
rect 59850 80310 59860 80380
rect 59640 80260 59860 80310
rect 60140 80490 60360 80540
rect 60140 80420 60150 80490
rect 60350 80420 60360 80490
rect 60140 80380 60360 80420
rect 60140 80310 60150 80380
rect 60350 80310 60360 80380
rect 60140 80260 60360 80310
rect 60640 80490 60860 80540
rect 60640 80420 60650 80490
rect 60850 80420 60860 80490
rect 60640 80380 60860 80420
rect 60640 80310 60650 80380
rect 60850 80310 60860 80380
rect 60640 80260 60860 80310
rect 61140 80490 61360 80540
rect 61140 80420 61150 80490
rect 61350 80420 61360 80490
rect 61140 80380 61360 80420
rect 61140 80310 61150 80380
rect 61350 80310 61360 80380
rect 61140 80260 61360 80310
rect 61640 80490 61860 80540
rect 61640 80420 61650 80490
rect 61850 80420 61860 80490
rect 61640 80380 61860 80420
rect 61640 80310 61650 80380
rect 61850 80310 61860 80380
rect 61640 80260 61860 80310
rect 62140 80490 62360 80540
rect 62140 80420 62150 80490
rect 62350 80420 62360 80490
rect 62140 80380 62360 80420
rect 62140 80310 62150 80380
rect 62350 80310 62360 80380
rect 62140 80260 62360 80310
rect 62640 80490 62860 80540
rect 62640 80420 62650 80490
rect 62850 80420 62860 80490
rect 62640 80380 62860 80420
rect 62640 80310 62650 80380
rect 62850 80310 62860 80380
rect 62640 80260 62860 80310
rect 63140 80490 63360 80540
rect 63140 80420 63150 80490
rect 63350 80420 63360 80490
rect 63140 80380 63360 80420
rect 63140 80310 63150 80380
rect 63350 80310 63360 80380
rect 63140 80260 63360 80310
rect 63640 80490 63860 80540
rect 63640 80420 63650 80490
rect 63850 80420 63860 80490
rect 63640 80380 63860 80420
rect 63640 80310 63650 80380
rect 63850 80310 63860 80380
rect 63640 80260 63860 80310
rect 64140 80490 64360 80540
rect 64140 80420 64150 80490
rect 64350 80420 64360 80490
rect 64140 80380 64360 80420
rect 64140 80310 64150 80380
rect 64350 80310 64360 80380
rect 64140 80260 64360 80310
rect 64640 80490 64860 80540
rect 64640 80420 64650 80490
rect 64850 80420 64860 80490
rect 64640 80380 64860 80420
rect 64640 80310 64650 80380
rect 64850 80310 64860 80380
rect 64640 80260 64860 80310
rect 65140 80490 65360 80540
rect 65140 80420 65150 80490
rect 65350 80420 65360 80490
rect 65140 80380 65360 80420
rect 65140 80310 65150 80380
rect 65350 80310 65360 80380
rect 65140 80260 65360 80310
rect 65640 80490 65860 80540
rect 65640 80420 65650 80490
rect 65850 80420 65860 80490
rect 65640 80380 65860 80420
rect 65640 80310 65650 80380
rect 65850 80310 65860 80380
rect 65640 80260 65860 80310
rect 66140 80490 66360 80540
rect 66140 80420 66150 80490
rect 66350 80420 66360 80490
rect 66140 80380 66360 80420
rect 66140 80310 66150 80380
rect 66350 80310 66360 80380
rect 66140 80260 66360 80310
rect 66640 80490 66860 80540
rect 66640 80420 66650 80490
rect 66850 80420 66860 80490
rect 66640 80380 66860 80420
rect 66640 80310 66650 80380
rect 66850 80310 66860 80380
rect 66640 80260 66860 80310
rect 67140 80490 67360 80540
rect 67140 80420 67150 80490
rect 67350 80420 67360 80490
rect 67140 80380 67360 80420
rect 67140 80310 67150 80380
rect 67350 80310 67360 80380
rect 67140 80260 67360 80310
rect 67640 80490 67860 80540
rect 67640 80420 67650 80490
rect 67850 80420 67860 80490
rect 67640 80380 67860 80420
rect 67640 80310 67650 80380
rect 67850 80310 67860 80380
rect 67640 80260 67860 80310
rect 68140 80490 68360 80540
rect 68140 80420 68150 80490
rect 68350 80420 68360 80490
rect 68140 80380 68360 80420
rect 68140 80310 68150 80380
rect 68350 80310 68360 80380
rect 68140 80260 68360 80310
rect 68640 80490 68860 80540
rect 68640 80420 68650 80490
rect 68850 80420 68860 80490
rect 68640 80380 68860 80420
rect 68640 80310 68650 80380
rect 68850 80310 68860 80380
rect 68640 80260 68860 80310
rect 69140 80490 69360 80540
rect 69140 80420 69150 80490
rect 69350 80420 69360 80490
rect 69140 80380 69360 80420
rect 69140 80310 69150 80380
rect 69350 80310 69360 80380
rect 69140 80260 69360 80310
rect 69640 80490 69860 80540
rect 69640 80420 69650 80490
rect 69850 80420 69860 80490
rect 69640 80380 69860 80420
rect 69640 80310 69650 80380
rect 69850 80310 69860 80380
rect 69640 80260 69860 80310
rect 70140 80490 70360 80540
rect 70140 80420 70150 80490
rect 70350 80420 70360 80490
rect 70140 80380 70360 80420
rect 70140 80310 70150 80380
rect 70350 80310 70360 80380
rect 70140 80260 70360 80310
rect 70640 80490 70860 80540
rect 70640 80420 70650 80490
rect 70850 80420 70860 80490
rect 70640 80380 70860 80420
rect 70640 80310 70650 80380
rect 70850 80310 70860 80380
rect 70640 80260 70860 80310
rect 71140 80490 71360 80540
rect 71140 80420 71150 80490
rect 71350 80420 71360 80490
rect 71140 80380 71360 80420
rect 71140 80310 71150 80380
rect 71350 80310 71360 80380
rect 71140 80260 71360 80310
rect 71640 80490 71860 80540
rect 71640 80420 71650 80490
rect 71850 80420 71860 80490
rect 71640 80380 71860 80420
rect 71640 80310 71650 80380
rect 71850 80310 71860 80380
rect 71640 80260 71860 80310
rect 72140 80490 72360 80540
rect 72140 80420 72150 80490
rect 72350 80420 72360 80490
rect 72140 80380 72360 80420
rect 72140 80310 72150 80380
rect 72350 80310 72360 80380
rect 72140 80260 72360 80310
rect 72640 80490 72860 80540
rect 72640 80420 72650 80490
rect 72850 80420 72860 80490
rect 72640 80380 72860 80420
rect 72640 80310 72650 80380
rect 72850 80310 72860 80380
rect 72640 80260 72860 80310
rect 73140 80490 73360 80540
rect 73140 80420 73150 80490
rect 73350 80420 73360 80490
rect 73140 80380 73360 80420
rect 73140 80310 73150 80380
rect 73350 80310 73360 80380
rect 73140 80260 73360 80310
rect 73640 80490 73860 80540
rect 73640 80420 73650 80490
rect 73850 80420 73860 80490
rect 73640 80380 73860 80420
rect 73640 80310 73650 80380
rect 73850 80310 73860 80380
rect 73640 80260 73860 80310
rect 74140 80490 74360 80540
rect 74140 80420 74150 80490
rect 74350 80420 74360 80490
rect 74140 80380 74360 80420
rect 74140 80310 74150 80380
rect 74350 80310 74360 80380
rect 74140 80260 74360 80310
rect 74640 80490 74860 80540
rect 74640 80420 74650 80490
rect 74850 80420 74860 80490
rect 74640 80380 74860 80420
rect 74640 80310 74650 80380
rect 74850 80310 74860 80380
rect 74640 80260 74860 80310
rect 75140 80490 75360 80540
rect 75140 80420 75150 80490
rect 75350 80420 75360 80490
rect 75140 80380 75360 80420
rect 75140 80310 75150 80380
rect 75350 80310 75360 80380
rect 75140 80260 75360 80310
rect 75640 80490 75860 80540
rect 75640 80420 75650 80490
rect 75850 80420 75860 80490
rect 75640 80380 75860 80420
rect 75640 80310 75650 80380
rect 75850 80310 75860 80380
rect 75640 80260 75860 80310
rect 76140 80490 76360 80540
rect 76140 80420 76150 80490
rect 76350 80420 76360 80490
rect 76140 80380 76360 80420
rect 76140 80310 76150 80380
rect 76350 80310 76360 80380
rect 76140 80260 76360 80310
rect 76640 80490 76860 80540
rect 76640 80420 76650 80490
rect 76850 80420 76860 80490
rect 76640 80380 76860 80420
rect 76640 80310 76650 80380
rect 76850 80310 76860 80380
rect 76640 80260 76860 80310
rect 77140 80490 77360 80540
rect 77140 80420 77150 80490
rect 77350 80420 77360 80490
rect 77140 80380 77360 80420
rect 77140 80310 77150 80380
rect 77350 80310 77360 80380
rect 77140 80260 77360 80310
rect 77640 80490 77860 80540
rect 77640 80420 77650 80490
rect 77850 80420 77860 80490
rect 77640 80380 77860 80420
rect 77640 80310 77650 80380
rect 77850 80310 77860 80380
rect 77640 80260 77860 80310
rect 78140 80490 78360 80540
rect 78140 80420 78150 80490
rect 78350 80420 78360 80490
rect 78140 80380 78360 80420
rect 78140 80310 78150 80380
rect 78350 80310 78360 80380
rect 78140 80260 78360 80310
rect 78640 80490 78860 80540
rect 78640 80420 78650 80490
rect 78850 80420 78860 80490
rect 78640 80380 78860 80420
rect 78640 80310 78650 80380
rect 78850 80310 78860 80380
rect 78640 80260 78860 80310
rect 79140 80490 79360 80540
rect 79140 80420 79150 80490
rect 79350 80420 79360 80490
rect 79140 80380 79360 80420
rect 79140 80310 79150 80380
rect 79350 80310 79360 80380
rect 79140 80260 79360 80310
rect 79640 80490 79860 80540
rect 79640 80420 79650 80490
rect 79850 80420 79860 80490
rect 79640 80380 79860 80420
rect 79640 80310 79650 80380
rect 79850 80310 79860 80380
rect 79640 80260 79860 80310
rect 80140 80490 80360 80540
rect 80140 80420 80150 80490
rect 80350 80420 80360 80490
rect 80140 80380 80360 80420
rect 80140 80310 80150 80380
rect 80350 80310 80360 80380
rect 80140 80260 80360 80310
rect 80640 80490 80860 80540
rect 80640 80420 80650 80490
rect 80850 80420 80860 80490
rect 80640 80380 80860 80420
rect 80640 80310 80650 80380
rect 80850 80310 80860 80380
rect 80640 80260 80860 80310
rect 81140 80490 81360 80540
rect 81140 80420 81150 80490
rect 81350 80420 81360 80490
rect 81140 80380 81360 80420
rect 81140 80310 81150 80380
rect 81350 80310 81360 80380
rect 81140 80260 81360 80310
rect 81640 80490 81860 80540
rect 81640 80420 81650 80490
rect 81850 80420 81860 80490
rect 81640 80380 81860 80420
rect 81640 80310 81650 80380
rect 81850 80310 81860 80380
rect 81640 80260 81860 80310
rect 82140 80490 82360 80540
rect 82140 80420 82150 80490
rect 82350 80420 82360 80490
rect 82140 80380 82360 80420
rect 82140 80310 82150 80380
rect 82350 80310 82360 80380
rect 82140 80260 82360 80310
rect 82640 80490 82860 80540
rect 82640 80420 82650 80490
rect 82850 80420 82860 80490
rect 82640 80380 82860 80420
rect 82640 80310 82650 80380
rect 82850 80310 82860 80380
rect 82640 80260 82860 80310
rect 83140 80490 83360 80540
rect 83140 80420 83150 80490
rect 83350 80420 83360 80490
rect 83140 80380 83360 80420
rect 83140 80310 83150 80380
rect 83350 80310 83360 80380
rect 83140 80260 83360 80310
rect 83640 80490 83860 80540
rect 83640 80420 83650 80490
rect 83850 80420 83860 80490
rect 83640 80380 83860 80420
rect 83640 80310 83650 80380
rect 83850 80310 83860 80380
rect 83640 80260 83860 80310
rect 84140 80490 84360 80540
rect 84140 80420 84150 80490
rect 84350 80420 84360 80490
rect 84140 80380 84360 80420
rect 84140 80310 84150 80380
rect 84350 80310 84360 80380
rect 84140 80260 84360 80310
rect 84640 80490 84860 80540
rect 84640 80420 84650 80490
rect 84850 80420 84860 80490
rect 84640 80380 84860 80420
rect 84640 80310 84650 80380
rect 84850 80310 84860 80380
rect 84640 80260 84860 80310
rect 85140 80490 85360 80540
rect 85140 80420 85150 80490
rect 85350 80420 85360 80490
rect 85140 80380 85360 80420
rect 85140 80310 85150 80380
rect 85350 80310 85360 80380
rect 85140 80260 85360 80310
rect 85640 80490 85860 80540
rect 85640 80420 85650 80490
rect 85850 80420 85860 80490
rect 85640 80380 85860 80420
rect 85640 80310 85650 80380
rect 85850 80310 85860 80380
rect 85640 80260 85860 80310
rect 86140 80490 86360 80540
rect 86140 80420 86150 80490
rect 86350 80420 86360 80490
rect 86140 80380 86360 80420
rect 86140 80310 86150 80380
rect 86350 80310 86360 80380
rect 86140 80260 86360 80310
rect 86640 80490 86860 80540
rect 86640 80420 86650 80490
rect 86850 80420 86860 80490
rect 86640 80380 86860 80420
rect 86640 80310 86650 80380
rect 86850 80310 86860 80380
rect 86640 80260 86860 80310
rect 87140 80490 87360 80540
rect 87140 80420 87150 80490
rect 87350 80420 87360 80490
rect 87140 80380 87360 80420
rect 87140 80310 87150 80380
rect 87350 80310 87360 80380
rect 87140 80260 87360 80310
rect 87640 80490 87860 80540
rect 87640 80420 87650 80490
rect 87850 80420 87860 80490
rect 87640 80380 87860 80420
rect 87640 80310 87650 80380
rect 87850 80310 87860 80380
rect 87640 80260 87860 80310
rect 88140 80490 88360 80540
rect 88140 80420 88150 80490
rect 88350 80420 88360 80490
rect 88140 80380 88360 80420
rect 88140 80310 88150 80380
rect 88350 80310 88360 80380
rect 88140 80260 88360 80310
rect 88640 80490 88860 80540
rect 88640 80420 88650 80490
rect 88850 80420 88860 80490
rect 88640 80380 88860 80420
rect 88640 80310 88650 80380
rect 88850 80310 88860 80380
rect 88640 80260 88860 80310
rect 89140 80490 89360 80540
rect 89140 80420 89150 80490
rect 89350 80420 89360 80490
rect 89140 80380 89360 80420
rect 89140 80310 89150 80380
rect 89350 80310 89360 80380
rect 89140 80260 89360 80310
rect 89640 80490 89860 80540
rect 89640 80420 89650 80490
rect 89850 80420 89860 80490
rect 89640 80380 89860 80420
rect 89640 80310 89650 80380
rect 89850 80310 89860 80380
rect 89640 80260 89860 80310
rect 90140 80490 90360 80540
rect 90140 80420 90150 80490
rect 90350 80420 90360 80490
rect 90140 80380 90360 80420
rect 90140 80310 90150 80380
rect 90350 80310 90360 80380
rect 90140 80260 90360 80310
rect 90640 80490 90860 80540
rect 90640 80420 90650 80490
rect 90850 80420 90860 80490
rect 90640 80380 90860 80420
rect 90640 80310 90650 80380
rect 90850 80310 90860 80380
rect 90640 80260 90860 80310
rect 91140 80490 91360 80540
rect 91140 80420 91150 80490
rect 91350 80420 91360 80490
rect 91140 80380 91360 80420
rect 91140 80310 91150 80380
rect 91350 80310 91360 80380
rect 91140 80260 91360 80310
rect 91640 80490 91860 80540
rect 91640 80420 91650 80490
rect 91850 80420 91860 80490
rect 91640 80380 91860 80420
rect 91640 80310 91650 80380
rect 91850 80310 91860 80380
rect 91640 80260 91860 80310
rect 92140 80490 92360 80540
rect 92140 80420 92150 80490
rect 92350 80420 92360 80490
rect 92140 80380 92360 80420
rect 92140 80310 92150 80380
rect 92350 80310 92360 80380
rect 92140 80260 92360 80310
rect 92640 80490 92860 80540
rect 92640 80420 92650 80490
rect 92850 80420 92860 80490
rect 92640 80380 92860 80420
rect 92640 80310 92650 80380
rect 92850 80310 92860 80380
rect 92640 80260 92860 80310
rect 93140 80490 93360 80540
rect 93140 80420 93150 80490
rect 93350 80420 93360 80490
rect 93140 80380 93360 80420
rect 93140 80310 93150 80380
rect 93350 80310 93360 80380
rect 93140 80260 93360 80310
rect 93640 80490 93860 80540
rect 93640 80420 93650 80490
rect 93850 80420 93860 80490
rect 93640 80380 93860 80420
rect 93640 80310 93650 80380
rect 93850 80310 93860 80380
rect 93640 80260 93860 80310
rect 94140 80490 94360 80540
rect 94140 80420 94150 80490
rect 94350 80420 94360 80490
rect 94140 80380 94360 80420
rect 94140 80310 94150 80380
rect 94350 80310 94360 80380
rect 94140 80260 94360 80310
rect 94640 80490 94860 80540
rect 94640 80420 94650 80490
rect 94850 80420 94860 80490
rect 94640 80380 94860 80420
rect 94640 80310 94650 80380
rect 94850 80310 94860 80380
rect 94640 80260 94860 80310
rect 95140 80490 95360 80540
rect 95140 80420 95150 80490
rect 95350 80420 95360 80490
rect 95140 80380 95360 80420
rect 95140 80310 95150 80380
rect 95350 80310 95360 80380
rect 95140 80260 95360 80310
rect 95640 80490 95860 80540
rect 95640 80420 95650 80490
rect 95850 80420 95860 80490
rect 95640 80380 95860 80420
rect 95640 80310 95650 80380
rect 95850 80310 95860 80380
rect 95640 80260 95860 80310
rect 96140 80490 96360 80540
rect 96140 80420 96150 80490
rect 96350 80420 96360 80490
rect 96140 80380 96360 80420
rect 96140 80310 96150 80380
rect 96350 80310 96360 80380
rect 96140 80260 96360 80310
rect 96640 80490 96860 80540
rect 96640 80420 96650 80490
rect 96850 80420 96860 80490
rect 96640 80380 96860 80420
rect 96640 80310 96650 80380
rect 96850 80310 96860 80380
rect 96640 80260 96860 80310
rect 97140 80490 97360 80540
rect 97140 80420 97150 80490
rect 97350 80420 97360 80490
rect 97140 80380 97360 80420
rect 97140 80310 97150 80380
rect 97350 80310 97360 80380
rect 97140 80260 97360 80310
rect 97640 80490 97860 80540
rect 97640 80420 97650 80490
rect 97850 80420 97860 80490
rect 97640 80380 97860 80420
rect 97640 80310 97650 80380
rect 97850 80310 97860 80380
rect 97640 80260 97860 80310
rect 98140 80490 98360 80540
rect 98140 80420 98150 80490
rect 98350 80420 98360 80490
rect 98140 80380 98360 80420
rect 98140 80310 98150 80380
rect 98350 80310 98360 80380
rect 98140 80260 98360 80310
rect 98640 80490 98860 80540
rect 98640 80420 98650 80490
rect 98850 80420 98860 80490
rect 98640 80380 98860 80420
rect 98640 80310 98650 80380
rect 98850 80310 98860 80380
rect 98640 80260 98860 80310
rect 99140 80490 99360 80540
rect 99140 80420 99150 80490
rect 99350 80420 99360 80490
rect 99140 80380 99360 80420
rect 99140 80310 99150 80380
rect 99350 80310 99360 80380
rect 99140 80260 99360 80310
rect 99640 80490 99860 80540
rect 99640 80420 99650 80490
rect 99850 80420 99860 80490
rect 99640 80380 99860 80420
rect 99640 80310 99650 80380
rect 99850 80310 99860 80380
rect 99640 80260 99860 80310
rect 100140 80490 100360 80540
rect 100140 80420 100150 80490
rect 100350 80420 100360 80490
rect 100140 80380 100360 80420
rect 100140 80310 100150 80380
rect 100350 80310 100360 80380
rect 100140 80260 100360 80310
rect -83500 80250 100500 80260
rect -83500 80050 -83480 80250
rect -83410 80050 -83090 80250
rect -83020 80050 -82980 80250
rect -82910 80050 -82590 80250
rect -82520 80050 -82480 80250
rect -82410 80050 -82090 80250
rect -82020 80050 -81980 80250
rect -81910 80050 -81590 80250
rect -81520 80050 -81480 80250
rect -81410 80050 -81090 80250
rect -81020 80050 -80980 80250
rect -80910 80050 -80590 80250
rect -80520 80050 -80480 80250
rect -80410 80050 -80090 80250
rect -80020 80050 -79980 80250
rect -79910 80050 -79590 80250
rect -79520 80050 -79480 80250
rect -79410 80050 -79090 80250
rect -79020 80050 -78980 80250
rect -78910 80050 -78590 80250
rect -78520 80050 -78480 80250
rect -78410 80050 -78090 80250
rect -78020 80050 -77980 80250
rect -77910 80050 -77590 80250
rect -77520 80050 -77480 80250
rect -77410 80050 -77090 80250
rect -77020 80050 -76980 80250
rect -76910 80050 -76590 80250
rect -76520 80050 -76480 80250
rect -76410 80050 -76090 80250
rect -76020 80050 -75980 80250
rect -75910 80050 -75590 80250
rect -75520 80050 -75480 80250
rect -75410 80050 -75090 80250
rect -75020 80050 -74980 80250
rect -74910 80050 -74590 80250
rect -74520 80050 -74480 80250
rect -74410 80050 -74090 80250
rect -74020 80050 -73980 80250
rect -73910 80050 -73590 80250
rect -73520 80050 -73480 80250
rect -73410 80050 -73090 80250
rect -73020 80050 -72980 80250
rect -72910 80050 -72590 80250
rect -72520 80050 -72480 80250
rect -72410 80050 -72090 80250
rect -72020 80050 -71980 80250
rect -71910 80050 -71590 80250
rect -71520 80050 -71480 80250
rect -71410 80050 -71090 80250
rect -71020 80050 -70980 80250
rect -70910 80050 -70590 80250
rect -70520 80050 -70480 80250
rect -70410 80050 -70090 80250
rect -70020 80050 -69980 80250
rect -69910 80050 -69590 80250
rect -69520 80050 -69480 80250
rect -69410 80050 -69090 80250
rect -69020 80050 -68980 80250
rect -68910 80050 -68590 80250
rect -68520 80050 -68480 80250
rect -68410 80050 -68090 80250
rect -68020 80050 -67980 80250
rect -67910 80050 -67590 80250
rect -67520 80050 -67480 80250
rect -67410 80050 -67090 80250
rect -67020 80050 -66980 80250
rect -66910 80050 -66590 80250
rect -66520 80050 -66480 80250
rect -66410 80050 -66090 80250
rect -66020 80050 -65980 80250
rect -65910 80050 -65590 80250
rect -65520 80050 -65480 80250
rect -65410 80050 -65090 80250
rect -65020 80050 -64980 80250
rect -64910 80050 -64590 80250
rect -64520 80050 -64480 80250
rect -64410 80050 -64090 80250
rect -64020 80050 -63980 80250
rect -63910 80050 -63590 80250
rect -63520 80050 -63480 80250
rect -63410 80050 -63090 80250
rect -63020 80050 -62980 80250
rect -62910 80050 -62590 80250
rect -62520 80050 -62480 80250
rect -62410 80050 -62090 80250
rect -62020 80050 -61980 80250
rect -61910 80050 -61590 80250
rect -61520 80050 -61480 80250
rect -61410 80050 -61090 80250
rect -61020 80050 -60980 80250
rect -60910 80050 -60590 80250
rect -60520 80050 -60480 80250
rect -60410 80050 -60090 80250
rect -60020 80050 -59980 80250
rect -59910 80050 -59590 80250
rect -59520 80050 -59480 80250
rect -59410 80050 -59090 80250
rect -59020 80050 -58980 80250
rect -58910 80050 -58590 80250
rect -58520 80050 -58480 80250
rect -58410 80050 -58090 80250
rect -58020 80050 -57980 80250
rect -57910 80050 -57590 80250
rect -57520 80050 -57480 80250
rect -57410 80050 -57090 80250
rect -57020 80050 -56980 80250
rect -56910 80050 -56590 80250
rect -56520 80050 -56480 80250
rect -56410 80050 -56090 80250
rect -56020 80050 -55980 80250
rect -55910 80050 -55590 80250
rect -55520 80050 -55480 80250
rect -55410 80050 -55090 80250
rect -55020 80050 -54980 80250
rect -54910 80050 -54590 80250
rect -54520 80050 -54480 80250
rect -54410 80050 -54090 80250
rect -54020 80050 -53980 80250
rect -53910 80050 -53590 80250
rect -53520 80050 -53480 80250
rect -53410 80050 -53090 80250
rect -53020 80050 -52980 80250
rect -52910 80050 -52590 80250
rect -52520 80050 -52480 80250
rect -52410 80050 -52090 80250
rect -52020 80050 -51980 80250
rect -51910 80050 -51590 80250
rect -51520 80050 -51480 80250
rect -51410 80050 -51090 80250
rect -51020 80050 -50980 80250
rect -50910 80050 -50590 80250
rect -50520 80050 -50480 80250
rect -50410 80050 -50090 80250
rect -50020 80050 -49980 80250
rect -49910 80050 -49590 80250
rect -49520 80050 -49480 80250
rect -49410 80050 -49090 80250
rect -49020 80050 -48980 80250
rect -48910 80050 -48590 80250
rect -48520 80050 -48480 80250
rect -48410 80050 -48090 80250
rect -48020 80050 -47980 80250
rect -47910 80050 -47590 80250
rect -47520 80050 -47480 80250
rect -47410 80050 -47090 80250
rect -47020 80050 -46980 80250
rect -46910 80050 -46590 80250
rect -46520 80050 -46480 80250
rect -46410 80050 -46090 80250
rect -46020 80050 -45980 80250
rect -45910 80050 -45590 80250
rect -45520 80050 -45480 80250
rect -45410 80050 -45090 80250
rect -45020 80050 -44980 80250
rect -44910 80050 -44590 80250
rect -44520 80050 -44480 80250
rect -44410 80050 -44090 80250
rect -44020 80050 -43980 80250
rect -43910 80050 -43590 80250
rect -43520 80050 -43480 80250
rect -43410 80050 -43090 80250
rect -43020 80050 -42980 80250
rect -42910 80050 -42590 80250
rect -42520 80050 -42480 80250
rect -42410 80050 -42090 80250
rect -42020 80050 -41980 80250
rect -41910 80050 -41590 80250
rect -41520 80050 -41480 80250
rect -41410 80050 -41090 80250
rect -41020 80050 -40980 80250
rect -40910 80050 -40590 80250
rect -40520 80050 -40480 80250
rect -40410 80050 -40090 80250
rect -40020 80050 -39980 80250
rect -39910 80050 -39590 80250
rect -39520 80050 -39480 80250
rect -39410 80050 -39090 80250
rect -39020 80050 -38980 80250
rect -38910 80050 -38590 80250
rect -38520 80050 -38480 80250
rect -38410 80050 -38090 80250
rect -38020 80050 -37980 80250
rect -37910 80050 -37590 80250
rect -37520 80050 -37480 80250
rect -37410 80050 -37090 80250
rect -37020 80050 -36980 80250
rect -36910 80050 -36590 80250
rect -36520 80050 -36480 80250
rect -36410 80050 -36090 80250
rect -36020 80050 -35980 80250
rect -35910 80050 -35590 80250
rect -35520 80050 -35480 80250
rect -35410 80050 -35090 80250
rect -35020 80050 -34980 80250
rect -34910 80050 -34590 80250
rect -34520 80050 -34480 80250
rect -34410 80050 -34090 80250
rect -34020 80050 -33980 80250
rect -33910 80050 -33590 80250
rect -33520 80050 -33480 80250
rect -33410 80050 -33090 80250
rect -33020 80050 -32980 80250
rect -32910 80050 -32590 80250
rect -32520 80050 -32480 80250
rect -32410 80050 -32090 80250
rect -32020 80050 -31980 80250
rect -31910 80050 -31590 80250
rect -31520 80050 -31480 80250
rect -31410 80050 -31090 80250
rect -31020 80050 -30980 80250
rect -30910 80050 -30590 80250
rect -30520 80050 -30480 80250
rect -30410 80050 -30090 80250
rect -30020 80050 -29980 80250
rect -29910 80050 -29590 80250
rect -29520 80050 -29480 80250
rect -29410 80050 -29090 80250
rect -29020 80050 -28980 80250
rect -28910 80050 -28590 80250
rect -28520 80050 -28480 80250
rect -28410 80050 -28090 80250
rect -28020 80050 -27980 80250
rect -27910 80050 -27590 80250
rect -27520 80050 -27480 80250
rect -27410 80050 -27090 80250
rect -27020 80050 -26980 80250
rect -26910 80050 -26590 80250
rect -26520 80050 -26480 80250
rect -26410 80050 -26090 80250
rect -26020 80050 -25980 80250
rect -25910 80050 -25590 80250
rect -25520 80050 -25480 80250
rect -25410 80050 -25090 80250
rect -25020 80050 -24980 80250
rect -24910 80050 -24590 80250
rect -24520 80050 -24480 80250
rect -24410 80050 -24090 80250
rect -24020 80050 -23980 80250
rect -23910 80050 -23590 80250
rect -23520 80050 -23480 80250
rect -23410 80050 -23090 80250
rect -23020 80050 -22980 80250
rect -22910 80050 -22590 80250
rect -22520 80050 -22480 80250
rect -22410 80050 -22090 80250
rect -22020 80050 -21980 80250
rect -21910 80050 -21590 80250
rect -21520 80050 -21480 80250
rect -21410 80050 -21090 80250
rect -21020 80050 -20980 80250
rect -20910 80050 -20590 80250
rect -20520 80050 -20480 80250
rect -20410 80050 -20090 80250
rect -20020 80050 -19980 80250
rect -19910 80050 -19590 80250
rect -19520 80050 -19480 80250
rect -19410 80050 -19090 80250
rect -19020 80050 -18980 80250
rect -18910 80050 -18590 80250
rect -18520 80050 -18480 80250
rect -18410 80050 -18090 80250
rect -18020 80050 -17980 80250
rect -17910 80050 -17590 80250
rect -17520 80050 -17480 80250
rect -17410 80050 -17090 80250
rect -17020 80050 -16980 80250
rect -16910 80050 -16590 80250
rect -16520 80050 -16480 80250
rect -16410 80050 -16090 80250
rect -16020 80050 -15980 80250
rect -15910 80050 -15590 80250
rect -15520 80050 -15480 80250
rect -15410 80050 -15090 80250
rect -15020 80050 -14980 80250
rect -14910 80050 -14590 80250
rect -14520 80050 -14480 80250
rect -14410 80050 -14090 80250
rect -14020 80050 -13980 80250
rect -13910 80050 -13590 80250
rect -13520 80050 -13480 80250
rect -13410 80050 -13090 80250
rect -13020 80050 -12980 80250
rect -12910 80050 -12590 80250
rect -12520 80050 -12480 80250
rect -12410 80050 -12090 80250
rect -12020 80050 -11980 80250
rect -11910 80050 -11590 80250
rect -11520 80050 -11480 80250
rect -11410 80050 -11090 80250
rect -11020 80050 -10980 80250
rect -10910 80050 -10590 80250
rect -10520 80050 -10480 80250
rect -10410 80050 -10090 80250
rect -10020 80050 -9980 80250
rect -9910 80050 -9590 80250
rect -9520 80050 -9480 80250
rect -9410 80050 -9090 80250
rect -9020 80050 -8980 80250
rect -8910 80050 -8590 80250
rect -8520 80050 -8480 80250
rect -8410 80050 -8090 80250
rect -8020 80050 -7980 80250
rect -7910 80050 -7590 80250
rect -7520 80050 -7480 80250
rect -7410 80050 -7090 80250
rect -7020 80050 -6980 80250
rect -6910 80050 -6590 80250
rect -6520 80050 -6480 80250
rect -6410 80050 -6090 80250
rect -6020 80050 -5980 80250
rect -5910 80050 -5590 80250
rect -5520 80050 -5480 80250
rect -5410 80050 -5090 80250
rect -5020 80050 -4980 80250
rect -4910 80050 -4590 80250
rect -4520 80050 -4480 80250
rect -4410 80050 -4090 80250
rect -4020 80050 -3980 80250
rect -3910 80050 -3590 80250
rect -3520 80050 -3480 80250
rect -3410 80050 -3090 80250
rect -3020 80050 -2980 80250
rect -2910 80050 -2590 80250
rect -2520 80050 -2480 80250
rect -2410 80050 -2090 80250
rect -2020 80050 -1980 80250
rect -1910 80050 -1590 80250
rect -1520 80050 -1480 80250
rect -1410 80050 -1090 80250
rect -1020 80050 -980 80250
rect -910 80050 -590 80250
rect -520 80050 -480 80250
rect -410 80050 -90 80250
rect -20 80050 20 80250
rect 90 80050 410 80250
rect 480 80050 520 80250
rect 590 80050 910 80250
rect 980 80050 1020 80250
rect 1090 80050 1410 80250
rect 1480 80050 1520 80250
rect 1590 80050 1910 80250
rect 1980 80050 2020 80250
rect 2090 80050 2410 80250
rect 2480 80050 2520 80250
rect 2590 80050 2910 80250
rect 2980 80050 3020 80250
rect 3090 80050 3410 80250
rect 3480 80050 3520 80250
rect 3590 80050 3910 80250
rect 3980 80050 4020 80250
rect 4090 80050 4410 80250
rect 4480 80050 4520 80250
rect 4590 80050 4910 80250
rect 4980 80050 5020 80250
rect 5090 80050 5410 80250
rect 5480 80050 5520 80250
rect 5590 80050 5910 80250
rect 5980 80050 6020 80250
rect 6090 80050 6410 80250
rect 6480 80050 6520 80250
rect 6590 80050 6910 80250
rect 6980 80050 7020 80250
rect 7090 80050 7410 80250
rect 7480 80050 7520 80250
rect 7590 80050 7910 80250
rect 7980 80050 8020 80250
rect 8090 80050 8410 80250
rect 8480 80050 8520 80250
rect 8590 80050 8910 80250
rect 8980 80050 9020 80250
rect 9090 80050 9410 80250
rect 9480 80050 9520 80250
rect 9590 80050 9910 80250
rect 9980 80050 10020 80250
rect 10090 80050 10410 80250
rect 10480 80050 10520 80250
rect 10590 80050 10910 80250
rect 10980 80050 11020 80250
rect 11090 80050 11410 80250
rect 11480 80050 11520 80250
rect 11590 80050 11910 80250
rect 11980 80050 12020 80250
rect 12090 80050 12410 80250
rect 12480 80050 12520 80250
rect 12590 80050 12910 80250
rect 12980 80050 13020 80250
rect 13090 80050 13410 80250
rect 13480 80050 13520 80250
rect 13590 80050 13910 80250
rect 13980 80050 14020 80250
rect 14090 80050 14410 80250
rect 14480 80050 14520 80250
rect 14590 80050 14910 80250
rect 14980 80050 15020 80250
rect 15090 80050 15410 80250
rect 15480 80050 15520 80250
rect 15590 80050 15910 80250
rect 15980 80050 16020 80250
rect 16090 80050 16410 80250
rect 16480 80050 16520 80250
rect 16590 80050 16910 80250
rect 16980 80050 17020 80250
rect 17090 80050 17410 80250
rect 17480 80050 17520 80250
rect 17590 80050 17910 80250
rect 17980 80050 18020 80250
rect 18090 80050 18410 80250
rect 18480 80050 18520 80250
rect 18590 80050 18910 80250
rect 18980 80050 19020 80250
rect 19090 80050 19410 80250
rect 19480 80050 19520 80250
rect 19590 80050 19910 80250
rect 19980 80050 20020 80250
rect 20090 80050 20410 80250
rect 20480 80050 20520 80250
rect 20590 80050 20910 80250
rect 20980 80050 21020 80250
rect 21090 80050 21410 80250
rect 21480 80050 21520 80250
rect 21590 80050 21910 80250
rect 21980 80050 22020 80250
rect 22090 80050 22410 80250
rect 22480 80050 22520 80250
rect 22590 80050 22910 80250
rect 22980 80050 23020 80250
rect 23090 80050 23410 80250
rect 23480 80050 23520 80250
rect 23590 80050 23910 80250
rect 23980 80050 24020 80250
rect 24090 80050 24410 80250
rect 24480 80050 24520 80250
rect 24590 80050 24910 80250
rect 24980 80050 25020 80250
rect 25090 80050 25410 80250
rect 25480 80050 25520 80250
rect 25590 80050 25910 80250
rect 25980 80050 26020 80250
rect 26090 80050 26410 80250
rect 26480 80050 26520 80250
rect 26590 80050 26910 80250
rect 26980 80050 27020 80250
rect 27090 80050 27410 80250
rect 27480 80050 27520 80250
rect 27590 80050 27910 80250
rect 27980 80050 28020 80250
rect 28090 80050 28410 80250
rect 28480 80050 28520 80250
rect 28590 80050 28910 80250
rect 28980 80050 29020 80250
rect 29090 80050 29410 80250
rect 29480 80050 29520 80250
rect 29590 80050 29910 80250
rect 29980 80050 30020 80250
rect 30090 80050 30410 80250
rect 30480 80050 30520 80250
rect 30590 80050 30910 80250
rect 30980 80050 31020 80250
rect 31090 80050 31410 80250
rect 31480 80050 31520 80250
rect 31590 80050 31910 80250
rect 31980 80050 32020 80250
rect 32090 80050 32410 80250
rect 32480 80050 32520 80250
rect 32590 80050 32910 80250
rect 32980 80050 33020 80250
rect 33090 80050 33410 80250
rect 33480 80050 33520 80250
rect 33590 80050 33910 80250
rect 33980 80050 34020 80250
rect 34090 80050 34410 80250
rect 34480 80050 34520 80250
rect 34590 80050 34910 80250
rect 34980 80050 35020 80250
rect 35090 80050 35410 80250
rect 35480 80050 35520 80250
rect 35590 80050 35910 80250
rect 35980 80050 36020 80250
rect 36090 80050 36410 80250
rect 36480 80050 36520 80250
rect 36590 80050 36910 80250
rect 36980 80050 37020 80250
rect 37090 80050 37410 80250
rect 37480 80050 37520 80250
rect 37590 80050 37910 80250
rect 37980 80050 38020 80250
rect 38090 80050 38410 80250
rect 38480 80050 38520 80250
rect 38590 80050 38910 80250
rect 38980 80050 39020 80250
rect 39090 80050 39410 80250
rect 39480 80050 39520 80250
rect 39590 80050 39910 80250
rect 39980 80050 40020 80250
rect 40090 80050 40410 80250
rect 40480 80050 40520 80250
rect 40590 80050 40910 80250
rect 40980 80050 41020 80250
rect 41090 80050 41410 80250
rect 41480 80050 41520 80250
rect 41590 80050 41910 80250
rect 41980 80050 42020 80250
rect 42090 80050 42410 80250
rect 42480 80050 42520 80250
rect 42590 80050 42910 80250
rect 42980 80050 43020 80250
rect 43090 80050 43410 80250
rect 43480 80050 43520 80250
rect 43590 80050 43910 80250
rect 43980 80050 44020 80250
rect 44090 80050 44410 80250
rect 44480 80050 44520 80250
rect 44590 80050 44910 80250
rect 44980 80050 45020 80250
rect 45090 80050 45410 80250
rect 45480 80050 45520 80250
rect 45590 80050 45910 80250
rect 45980 80050 46020 80250
rect 46090 80050 46410 80250
rect 46480 80050 46520 80250
rect 46590 80050 46910 80250
rect 46980 80050 47020 80250
rect 47090 80050 47410 80250
rect 47480 80050 47520 80250
rect 47590 80050 47910 80250
rect 47980 80050 48020 80250
rect 48090 80050 48410 80250
rect 48480 80050 48520 80250
rect 48590 80050 48910 80250
rect 48980 80050 49020 80250
rect 49090 80050 49410 80250
rect 49480 80050 49520 80250
rect 49590 80050 49910 80250
rect 49980 80050 50020 80250
rect 50090 80050 50410 80250
rect 50480 80050 50520 80250
rect 50590 80050 50910 80250
rect 50980 80050 51020 80250
rect 51090 80050 51410 80250
rect 51480 80050 51520 80250
rect 51590 80050 51910 80250
rect 51980 80050 52020 80250
rect 52090 80050 52410 80250
rect 52480 80050 52520 80250
rect 52590 80050 52910 80250
rect 52980 80050 53020 80250
rect 53090 80050 53410 80250
rect 53480 80050 53520 80250
rect 53590 80050 53910 80250
rect 53980 80050 54020 80250
rect 54090 80050 54410 80250
rect 54480 80050 54520 80250
rect 54590 80050 54910 80250
rect 54980 80050 55020 80250
rect 55090 80050 55410 80250
rect 55480 80050 55520 80250
rect 55590 80050 55910 80250
rect 55980 80050 56020 80250
rect 56090 80050 56410 80250
rect 56480 80050 56520 80250
rect 56590 80050 56910 80250
rect 56980 80050 57020 80250
rect 57090 80050 57410 80250
rect 57480 80050 57520 80250
rect 57590 80050 57910 80250
rect 57980 80050 58020 80250
rect 58090 80050 58410 80250
rect 58480 80050 58520 80250
rect 58590 80050 58910 80250
rect 58980 80050 59020 80250
rect 59090 80050 59410 80250
rect 59480 80050 59520 80250
rect 59590 80050 59910 80250
rect 59980 80050 60020 80250
rect 60090 80050 60410 80250
rect 60480 80050 60520 80250
rect 60590 80050 60910 80250
rect 60980 80050 61020 80250
rect 61090 80050 61410 80250
rect 61480 80050 61520 80250
rect 61590 80050 61910 80250
rect 61980 80050 62020 80250
rect 62090 80050 62410 80250
rect 62480 80050 62520 80250
rect 62590 80050 62910 80250
rect 62980 80050 63020 80250
rect 63090 80050 63410 80250
rect 63480 80050 63520 80250
rect 63590 80050 63910 80250
rect 63980 80050 64020 80250
rect 64090 80050 64410 80250
rect 64480 80050 64520 80250
rect 64590 80050 64910 80250
rect 64980 80050 65020 80250
rect 65090 80050 65410 80250
rect 65480 80050 65520 80250
rect 65590 80050 65910 80250
rect 65980 80050 66020 80250
rect 66090 80050 66410 80250
rect 66480 80050 66520 80250
rect 66590 80050 66910 80250
rect 66980 80050 67020 80250
rect 67090 80050 67410 80250
rect 67480 80050 67520 80250
rect 67590 80050 67910 80250
rect 67980 80050 68020 80250
rect 68090 80050 68410 80250
rect 68480 80050 68520 80250
rect 68590 80050 68910 80250
rect 68980 80050 69020 80250
rect 69090 80050 69410 80250
rect 69480 80050 69520 80250
rect 69590 80050 69910 80250
rect 69980 80050 70020 80250
rect 70090 80050 70410 80250
rect 70480 80050 70520 80250
rect 70590 80050 70910 80250
rect 70980 80050 71020 80250
rect 71090 80050 71410 80250
rect 71480 80050 71520 80250
rect 71590 80050 71910 80250
rect 71980 80050 72020 80250
rect 72090 80050 72410 80250
rect 72480 80050 72520 80250
rect 72590 80050 72910 80250
rect 72980 80050 73020 80250
rect 73090 80050 73410 80250
rect 73480 80050 73520 80250
rect 73590 80050 73910 80250
rect 73980 80050 74020 80250
rect 74090 80050 74410 80250
rect 74480 80050 74520 80250
rect 74590 80050 74910 80250
rect 74980 80050 75020 80250
rect 75090 80050 75410 80250
rect 75480 80050 75520 80250
rect 75590 80050 75910 80250
rect 75980 80050 76020 80250
rect 76090 80050 76410 80250
rect 76480 80050 76520 80250
rect 76590 80050 76910 80250
rect 76980 80050 77020 80250
rect 77090 80050 77410 80250
rect 77480 80050 77520 80250
rect 77590 80050 77910 80250
rect 77980 80050 78020 80250
rect 78090 80050 78410 80250
rect 78480 80050 78520 80250
rect 78590 80050 78910 80250
rect 78980 80050 79020 80250
rect 79090 80050 79410 80250
rect 79480 80050 79520 80250
rect 79590 80050 79910 80250
rect 79980 80050 80020 80250
rect 80090 80050 80410 80250
rect 80480 80050 80520 80250
rect 80590 80050 80910 80250
rect 80980 80050 81020 80250
rect 81090 80050 81410 80250
rect 81480 80050 81520 80250
rect 81590 80050 81910 80250
rect 81980 80050 82020 80250
rect 82090 80050 82410 80250
rect 82480 80050 82520 80250
rect 82590 80050 82910 80250
rect 82980 80050 83020 80250
rect 83090 80050 83410 80250
rect 83480 80050 83520 80250
rect 83590 80050 83910 80250
rect 83980 80050 84020 80250
rect 84090 80050 84410 80250
rect 84480 80050 84520 80250
rect 84590 80050 84910 80250
rect 84980 80050 85020 80250
rect 85090 80050 85410 80250
rect 85480 80050 85520 80250
rect 85590 80050 85910 80250
rect 85980 80050 86020 80250
rect 86090 80050 86410 80250
rect 86480 80050 86520 80250
rect 86590 80050 86910 80250
rect 86980 80050 87020 80250
rect 87090 80050 87410 80250
rect 87480 80050 87520 80250
rect 87590 80050 87910 80250
rect 87980 80050 88020 80250
rect 88090 80050 88410 80250
rect 88480 80050 88520 80250
rect 88590 80050 88910 80250
rect 88980 80050 89020 80250
rect 89090 80050 89410 80250
rect 89480 80050 89520 80250
rect 89590 80050 89910 80250
rect 89980 80050 90020 80250
rect 90090 80050 90410 80250
rect 90480 80050 90520 80250
rect 90590 80050 90910 80250
rect 90980 80050 91020 80250
rect 91090 80050 91410 80250
rect 91480 80050 91520 80250
rect 91590 80050 91910 80250
rect 91980 80050 92020 80250
rect 92090 80050 92410 80250
rect 92480 80050 92520 80250
rect 92590 80050 92910 80250
rect 92980 80050 93020 80250
rect 93090 80050 93410 80250
rect 93480 80050 93520 80250
rect 93590 80050 93910 80250
rect 93980 80050 94020 80250
rect 94090 80050 94410 80250
rect 94480 80050 94520 80250
rect 94590 80050 94910 80250
rect 94980 80050 95020 80250
rect 95090 80050 95410 80250
rect 95480 80050 95520 80250
rect 95590 80050 95910 80250
rect 95980 80050 96020 80250
rect 96090 80050 96410 80250
rect 96480 80050 96520 80250
rect 96590 80050 96910 80250
rect 96980 80050 97020 80250
rect 97090 80050 97410 80250
rect 97480 80050 97520 80250
rect 97590 80050 97910 80250
rect 97980 80050 98020 80250
rect 98090 80050 98410 80250
rect 98480 80050 98520 80250
rect 98590 80050 98910 80250
rect 98980 80050 99020 80250
rect 99090 80050 99410 80250
rect 99480 80050 99520 80250
rect 99590 80050 99910 80250
rect 99980 80050 100020 80250
rect 100090 80050 100410 80250
rect 100480 80050 100500 80250
rect -83500 80040 100500 80050
rect -83360 79990 -83140 80040
rect -83360 79920 -83350 79990
rect -83150 79920 -83140 79990
rect -83360 79900 -83140 79920
rect -82860 79990 -82640 80040
rect -82860 79920 -82850 79990
rect -82650 79920 -82640 79990
rect -82860 79900 -82640 79920
rect -82360 79990 -82140 80040
rect -82360 79920 -82350 79990
rect -82150 79920 -82140 79990
rect -82360 79900 -82140 79920
rect -81860 79990 -81640 80040
rect -81860 79920 -81850 79990
rect -81650 79920 -81640 79990
rect -81860 79900 -81640 79920
rect -81360 79990 -81140 80040
rect -81360 79920 -81350 79990
rect -81150 79920 -81140 79990
rect -81360 79900 -81140 79920
rect -80860 79990 -80640 80040
rect -80860 79920 -80850 79990
rect -80650 79920 -80640 79990
rect -80860 79900 -80640 79920
rect -80360 79990 -80140 80040
rect -80360 79920 -80350 79990
rect -80150 79920 -80140 79990
rect -80360 79900 -80140 79920
rect -79860 79990 -79640 80040
rect -79860 79920 -79850 79990
rect -79650 79920 -79640 79990
rect -79860 79900 -79640 79920
rect -79360 79990 -79140 80040
rect -79360 79920 -79350 79990
rect -79150 79920 -79140 79990
rect -79360 79900 -79140 79920
rect -78860 79990 -78640 80040
rect -78860 79920 -78850 79990
rect -78650 79920 -78640 79990
rect -78860 79900 -78640 79920
rect -78360 79990 -78140 80040
rect -78360 79920 -78350 79990
rect -78150 79920 -78140 79990
rect -78360 79900 -78140 79920
rect -77860 79990 -77640 80040
rect -77860 79920 -77850 79990
rect -77650 79920 -77640 79990
rect -77860 79900 -77640 79920
rect -77360 79990 -77140 80040
rect -77360 79920 -77350 79990
rect -77150 79920 -77140 79990
rect -77360 79900 -77140 79920
rect -76860 79990 -76640 80040
rect -76860 79920 -76850 79990
rect -76650 79920 -76640 79990
rect -76860 79900 -76640 79920
rect -76360 79990 -76140 80040
rect -76360 79920 -76350 79990
rect -76150 79920 -76140 79990
rect -76360 79900 -76140 79920
rect -75860 79990 -75640 80040
rect -75860 79920 -75850 79990
rect -75650 79920 -75640 79990
rect -75860 79900 -75640 79920
rect -75360 79990 -75140 80040
rect -75360 79920 -75350 79990
rect -75150 79920 -75140 79990
rect -75360 79900 -75140 79920
rect -74860 79990 -74640 80040
rect -74860 79920 -74850 79990
rect -74650 79920 -74640 79990
rect -74860 79900 -74640 79920
rect -74360 79990 -74140 80040
rect -74360 79920 -74350 79990
rect -74150 79920 -74140 79990
rect -74360 79900 -74140 79920
rect -73860 79990 -73640 80040
rect -73860 79920 -73850 79990
rect -73650 79920 -73640 79990
rect -73860 79900 -73640 79920
rect -73360 79990 -73140 80040
rect -73360 79920 -73350 79990
rect -73150 79920 -73140 79990
rect -73360 79900 -73140 79920
rect -72860 79990 -72640 80040
rect -72860 79920 -72850 79990
rect -72650 79920 -72640 79990
rect -72860 79900 -72640 79920
rect -72360 79990 -72140 80040
rect -72360 79920 -72350 79990
rect -72150 79920 -72140 79990
rect -72360 79900 -72140 79920
rect -71860 79990 -71640 80040
rect -71860 79920 -71850 79990
rect -71650 79920 -71640 79990
rect -71860 79900 -71640 79920
rect -71360 79990 -71140 80040
rect -71360 79920 -71350 79990
rect -71150 79920 -71140 79990
rect -71360 79900 -71140 79920
rect -70860 79990 -70640 80040
rect -70860 79920 -70850 79990
rect -70650 79920 -70640 79990
rect -70860 79900 -70640 79920
rect -70360 79990 -70140 80040
rect -70360 79920 -70350 79990
rect -70150 79920 -70140 79990
rect -70360 79900 -70140 79920
rect -69860 79990 -69640 80040
rect -69860 79920 -69850 79990
rect -69650 79920 -69640 79990
rect -69860 79900 -69640 79920
rect -69360 79990 -69140 80040
rect -69360 79920 -69350 79990
rect -69150 79920 -69140 79990
rect -69360 79900 -69140 79920
rect -68860 79990 -68640 80040
rect -68860 79920 -68850 79990
rect -68650 79920 -68640 79990
rect -68860 79900 -68640 79920
rect -68360 79990 -68140 80040
rect -68360 79920 -68350 79990
rect -68150 79920 -68140 79990
rect -68360 79900 -68140 79920
rect -67860 79990 -67640 80040
rect -67860 79920 -67850 79990
rect -67650 79920 -67640 79990
rect -67860 79900 -67640 79920
rect -67360 79990 -67140 80040
rect -67360 79920 -67350 79990
rect -67150 79920 -67140 79990
rect -67360 79900 -67140 79920
rect -66860 79990 -66640 80040
rect -66860 79920 -66850 79990
rect -66650 79920 -66640 79990
rect -66860 79900 -66640 79920
rect -66360 79990 -66140 80040
rect -66360 79920 -66350 79990
rect -66150 79920 -66140 79990
rect -66360 79900 -66140 79920
rect -65860 79990 -65640 80040
rect -65860 79920 -65850 79990
rect -65650 79920 -65640 79990
rect -65860 79900 -65640 79920
rect -65360 79990 -65140 80040
rect -65360 79920 -65350 79990
rect -65150 79920 -65140 79990
rect -65360 79900 -65140 79920
rect -64860 79990 -64640 80040
rect -64860 79920 -64850 79990
rect -64650 79920 -64640 79990
rect -64860 79900 -64640 79920
rect -64360 79990 -64140 80040
rect -64360 79920 -64350 79990
rect -64150 79920 -64140 79990
rect -64360 79900 -64140 79920
rect -63860 79990 -63640 80040
rect -63860 79920 -63850 79990
rect -63650 79920 -63640 79990
rect -63860 79900 -63640 79920
rect -63360 79990 -63140 80040
rect -63360 79920 -63350 79990
rect -63150 79920 -63140 79990
rect -63360 79900 -63140 79920
rect -62860 79990 -62640 80040
rect -62860 79920 -62850 79990
rect -62650 79920 -62640 79990
rect -62860 79900 -62640 79920
rect -62360 79990 -62140 80040
rect -62360 79920 -62350 79990
rect -62150 79920 -62140 79990
rect -62360 79900 -62140 79920
rect -61860 79990 -61640 80040
rect -61860 79920 -61850 79990
rect -61650 79920 -61640 79990
rect -61860 79900 -61640 79920
rect -61360 79990 -61140 80040
rect -61360 79920 -61350 79990
rect -61150 79920 -61140 79990
rect -61360 79900 -61140 79920
rect -60860 79990 -60640 80040
rect -60860 79920 -60850 79990
rect -60650 79920 -60640 79990
rect -60860 79900 -60640 79920
rect -60360 79990 -60140 80040
rect -60360 79920 -60350 79990
rect -60150 79920 -60140 79990
rect -60360 79900 -60140 79920
rect -59860 79990 -59640 80040
rect -59860 79920 -59850 79990
rect -59650 79920 -59640 79990
rect -59860 79900 -59640 79920
rect -59360 79990 -59140 80040
rect -59360 79920 -59350 79990
rect -59150 79920 -59140 79990
rect -59360 79900 -59140 79920
rect -58860 79990 -58640 80040
rect -58860 79920 -58850 79990
rect -58650 79920 -58640 79990
rect -58860 79900 -58640 79920
rect -58360 79990 -58140 80040
rect -58360 79920 -58350 79990
rect -58150 79920 -58140 79990
rect -58360 79900 -58140 79920
rect -57860 79990 -57640 80040
rect -57860 79920 -57850 79990
rect -57650 79920 -57640 79990
rect -57860 79900 -57640 79920
rect -57360 79990 -57140 80040
rect -57360 79920 -57350 79990
rect -57150 79920 -57140 79990
rect -57360 79900 -57140 79920
rect -56860 79990 -56640 80040
rect -56860 79920 -56850 79990
rect -56650 79920 -56640 79990
rect -56860 79900 -56640 79920
rect -56360 79990 -56140 80040
rect -56360 79920 -56350 79990
rect -56150 79920 -56140 79990
rect -56360 79900 -56140 79920
rect -55860 79990 -55640 80040
rect -55860 79920 -55850 79990
rect -55650 79920 -55640 79990
rect -55860 79900 -55640 79920
rect -55360 79990 -55140 80040
rect -55360 79920 -55350 79990
rect -55150 79920 -55140 79990
rect -55360 79900 -55140 79920
rect -54860 79990 -54640 80040
rect -54860 79920 -54850 79990
rect -54650 79920 -54640 79990
rect -54860 79900 -54640 79920
rect -54360 79990 -54140 80040
rect -54360 79920 -54350 79990
rect -54150 79920 -54140 79990
rect -54360 79900 -54140 79920
rect -53860 79990 -53640 80040
rect -53860 79920 -53850 79990
rect -53650 79920 -53640 79990
rect -53860 79900 -53640 79920
rect -53360 79990 -53140 80040
rect -53360 79920 -53350 79990
rect -53150 79920 -53140 79990
rect -53360 79900 -53140 79920
rect -52860 79990 -52640 80040
rect -52860 79920 -52850 79990
rect -52650 79920 -52640 79990
rect -52860 79900 -52640 79920
rect -52360 79990 -52140 80040
rect -52360 79920 -52350 79990
rect -52150 79920 -52140 79990
rect -52360 79900 -52140 79920
rect -51860 79990 -51640 80040
rect -51860 79920 -51850 79990
rect -51650 79920 -51640 79990
rect -51860 79900 -51640 79920
rect -51360 79990 -51140 80040
rect -51360 79920 -51350 79990
rect -51150 79920 -51140 79990
rect -51360 79900 -51140 79920
rect -50860 79990 -50640 80040
rect -50860 79920 -50850 79990
rect -50650 79920 -50640 79990
rect -50860 79900 -50640 79920
rect -50360 79990 -50140 80040
rect -50360 79920 -50350 79990
rect -50150 79920 -50140 79990
rect -50360 79900 -50140 79920
rect -49860 79990 -49640 80040
rect -49860 79920 -49850 79990
rect -49650 79920 -49640 79990
rect -49860 79900 -49640 79920
rect -49360 79990 -49140 80040
rect -49360 79920 -49350 79990
rect -49150 79920 -49140 79990
rect -49360 79900 -49140 79920
rect -48860 79990 -48640 80040
rect -48860 79920 -48850 79990
rect -48650 79920 -48640 79990
rect -48860 79900 -48640 79920
rect -48360 79990 -48140 80040
rect -48360 79920 -48350 79990
rect -48150 79920 -48140 79990
rect -48360 79900 -48140 79920
rect -47860 79990 -47640 80040
rect -47860 79920 -47850 79990
rect -47650 79920 -47640 79990
rect -47860 79900 -47640 79920
rect -47360 79990 -47140 80040
rect -47360 79920 -47350 79990
rect -47150 79920 -47140 79990
rect -47360 79900 -47140 79920
rect -46860 79990 -46640 80040
rect -46860 79920 -46850 79990
rect -46650 79920 -46640 79990
rect -46860 79900 -46640 79920
rect -46360 79990 -46140 80040
rect -46360 79920 -46350 79990
rect -46150 79920 -46140 79990
rect -46360 79900 -46140 79920
rect -45860 79990 -45640 80040
rect -45860 79920 -45850 79990
rect -45650 79920 -45640 79990
rect -45860 79900 -45640 79920
rect -45360 79990 -45140 80040
rect -45360 79920 -45350 79990
rect -45150 79920 -45140 79990
rect -45360 79900 -45140 79920
rect -44860 79990 -44640 80040
rect -44860 79920 -44850 79990
rect -44650 79920 -44640 79990
rect -44860 79900 -44640 79920
rect -44360 79990 -44140 80040
rect -44360 79920 -44350 79990
rect -44150 79920 -44140 79990
rect -44360 79900 -44140 79920
rect -43860 79990 -43640 80040
rect -43860 79920 -43850 79990
rect -43650 79920 -43640 79990
rect -43860 79900 -43640 79920
rect -43360 79990 -43140 80040
rect -43360 79920 -43350 79990
rect -43150 79920 -43140 79990
rect -43360 79900 -43140 79920
rect -42860 79990 -42640 80040
rect -42860 79920 -42850 79990
rect -42650 79920 -42640 79990
rect -42860 79900 -42640 79920
rect -42360 79990 -42140 80040
rect -42360 79920 -42350 79990
rect -42150 79920 -42140 79990
rect -42360 79900 -42140 79920
rect -41860 79990 -41640 80040
rect -41860 79920 -41850 79990
rect -41650 79920 -41640 79990
rect -41860 79900 -41640 79920
rect -41360 79990 -41140 80040
rect -41360 79920 -41350 79990
rect -41150 79920 -41140 79990
rect -41360 79900 -41140 79920
rect -40860 79990 -40640 80040
rect -40860 79920 -40850 79990
rect -40650 79920 -40640 79990
rect -40860 79900 -40640 79920
rect -40360 79990 -40140 80040
rect -40360 79920 -40350 79990
rect -40150 79920 -40140 79990
rect -40360 79900 -40140 79920
rect -39860 79990 -39640 80040
rect -39860 79920 -39850 79990
rect -39650 79920 -39640 79990
rect -39860 79900 -39640 79920
rect -39360 79990 -39140 80040
rect -39360 79920 -39350 79990
rect -39150 79920 -39140 79990
rect -39360 79900 -39140 79920
rect -38860 79990 -38640 80040
rect -38860 79920 -38850 79990
rect -38650 79920 -38640 79990
rect -38860 79900 -38640 79920
rect -38360 79990 -38140 80040
rect -38360 79920 -38350 79990
rect -38150 79920 -38140 79990
rect -38360 79900 -38140 79920
rect -37860 79990 -37640 80040
rect -37860 79920 -37850 79990
rect -37650 79920 -37640 79990
rect -37860 79900 -37640 79920
rect -37360 79990 -37140 80040
rect -37360 79920 -37350 79990
rect -37150 79920 -37140 79990
rect -37360 79900 -37140 79920
rect -36860 79990 -36640 80040
rect -36860 79920 -36850 79990
rect -36650 79920 -36640 79990
rect -36860 79900 -36640 79920
rect -36360 79990 -36140 80040
rect -36360 79920 -36350 79990
rect -36150 79920 -36140 79990
rect -36360 79900 -36140 79920
rect -35860 79990 -35640 80040
rect -35860 79920 -35850 79990
rect -35650 79920 -35640 79990
rect -35860 79900 -35640 79920
rect -35360 79990 -35140 80040
rect -35360 79920 -35350 79990
rect -35150 79920 -35140 79990
rect -35360 79900 -35140 79920
rect -34860 79990 -34640 80040
rect -34860 79920 -34850 79990
rect -34650 79920 -34640 79990
rect -34860 79900 -34640 79920
rect -34360 79990 -34140 80040
rect -34360 79920 -34350 79990
rect -34150 79920 -34140 79990
rect -34360 79900 -34140 79920
rect -33860 79990 -33640 80040
rect -33860 79920 -33850 79990
rect -33650 79920 -33640 79990
rect -33860 79900 -33640 79920
rect -33360 79990 -33140 80040
rect -33360 79920 -33350 79990
rect -33150 79920 -33140 79990
rect -33360 79900 -33140 79920
rect -32860 79990 -32640 80040
rect -32860 79920 -32850 79990
rect -32650 79920 -32640 79990
rect -32860 79900 -32640 79920
rect -32360 79990 -32140 80040
rect -32360 79920 -32350 79990
rect -32150 79920 -32140 79990
rect -32360 79900 -32140 79920
rect -31860 79990 -31640 80040
rect -31860 79920 -31850 79990
rect -31650 79920 -31640 79990
rect -31860 79900 -31640 79920
rect -31360 79990 -31140 80040
rect -31360 79920 -31350 79990
rect -31150 79920 -31140 79990
rect -31360 79900 -31140 79920
rect -30860 79990 -30640 80040
rect -30860 79920 -30850 79990
rect -30650 79920 -30640 79990
rect -30860 79900 -30640 79920
rect -30360 79990 -30140 80040
rect -30360 79920 -30350 79990
rect -30150 79920 -30140 79990
rect -30360 79900 -30140 79920
rect -29860 79990 -29640 80040
rect -29860 79920 -29850 79990
rect -29650 79920 -29640 79990
rect -29860 79900 -29640 79920
rect -29360 79990 -29140 80040
rect -29360 79920 -29350 79990
rect -29150 79920 -29140 79990
rect -29360 79900 -29140 79920
rect -28860 79990 -28640 80040
rect -28860 79920 -28850 79990
rect -28650 79920 -28640 79990
rect -28860 79900 -28640 79920
rect -28360 79990 -28140 80040
rect -28360 79920 -28350 79990
rect -28150 79920 -28140 79990
rect -28360 79900 -28140 79920
rect -27860 79990 -27640 80040
rect -27860 79920 -27850 79990
rect -27650 79920 -27640 79990
rect -27860 79900 -27640 79920
rect -27360 79990 -27140 80040
rect -27360 79920 -27350 79990
rect -27150 79920 -27140 79990
rect -27360 79900 -27140 79920
rect -26860 79990 -26640 80040
rect -26860 79920 -26850 79990
rect -26650 79920 -26640 79990
rect -26860 79900 -26640 79920
rect -26360 79990 -26140 80040
rect -26360 79920 -26350 79990
rect -26150 79920 -26140 79990
rect -26360 79900 -26140 79920
rect -25860 79990 -25640 80040
rect -25860 79920 -25850 79990
rect -25650 79920 -25640 79990
rect -25860 79900 -25640 79920
rect -25360 79990 -25140 80040
rect -25360 79920 -25350 79990
rect -25150 79920 -25140 79990
rect -25360 79900 -25140 79920
rect -24860 79990 -24640 80040
rect -24860 79920 -24850 79990
rect -24650 79920 -24640 79990
rect -24860 79900 -24640 79920
rect -24360 79990 -24140 80040
rect -24360 79920 -24350 79990
rect -24150 79920 -24140 79990
rect -24360 79900 -24140 79920
rect -23860 79990 -23640 80040
rect -23860 79920 -23850 79990
rect -23650 79920 -23640 79990
rect -23860 79900 -23640 79920
rect -23360 79990 -23140 80040
rect -23360 79920 -23350 79990
rect -23150 79920 -23140 79990
rect -23360 79900 -23140 79920
rect -22860 79990 -22640 80040
rect -22860 79920 -22850 79990
rect -22650 79920 -22640 79990
rect -22860 79900 -22640 79920
rect -22360 79990 -22140 80040
rect -22360 79920 -22350 79990
rect -22150 79920 -22140 79990
rect -22360 79900 -22140 79920
rect -21860 79990 -21640 80040
rect -21860 79920 -21850 79990
rect -21650 79920 -21640 79990
rect -21860 79900 -21640 79920
rect -21360 79990 -21140 80040
rect -21360 79920 -21350 79990
rect -21150 79920 -21140 79990
rect -21360 79900 -21140 79920
rect -20860 79990 -20640 80040
rect -20860 79920 -20850 79990
rect -20650 79920 -20640 79990
rect -20860 79900 -20640 79920
rect -20360 79990 -20140 80040
rect -20360 79920 -20350 79990
rect -20150 79920 -20140 79990
rect -20360 79900 -20140 79920
rect -19860 79990 -19640 80040
rect -19860 79920 -19850 79990
rect -19650 79920 -19640 79990
rect -19860 79900 -19640 79920
rect -19360 79990 -19140 80040
rect -19360 79920 -19350 79990
rect -19150 79920 -19140 79990
rect -19360 79900 -19140 79920
rect -18860 79990 -18640 80040
rect -18860 79920 -18850 79990
rect -18650 79920 -18640 79990
rect -18860 79900 -18640 79920
rect -18360 79990 -18140 80040
rect -18360 79920 -18350 79990
rect -18150 79920 -18140 79990
rect -18360 79900 -18140 79920
rect -17860 79990 -17640 80040
rect -17860 79920 -17850 79990
rect -17650 79920 -17640 79990
rect -17860 79900 -17640 79920
rect -17360 79990 -17140 80040
rect -17360 79920 -17350 79990
rect -17150 79920 -17140 79990
rect -17360 79900 -17140 79920
rect -16860 79990 -16640 80040
rect -16860 79920 -16850 79990
rect -16650 79920 -16640 79990
rect -16860 79900 -16640 79920
rect -16360 79990 -16140 80040
rect -16360 79920 -16350 79990
rect -16150 79920 -16140 79990
rect -16360 79900 -16140 79920
rect -15860 79990 -15640 80040
rect -15860 79920 -15850 79990
rect -15650 79920 -15640 79990
rect -15860 79900 -15640 79920
rect -15360 79990 -15140 80040
rect -15360 79920 -15350 79990
rect -15150 79920 -15140 79990
rect -15360 79900 -15140 79920
rect -14860 79990 -14640 80040
rect -14860 79920 -14850 79990
rect -14650 79920 -14640 79990
rect -14860 79900 -14640 79920
rect -14360 79990 -14140 80040
rect -14360 79920 -14350 79990
rect -14150 79920 -14140 79990
rect -14360 79900 -14140 79920
rect -13860 79990 -13640 80040
rect -13860 79920 -13850 79990
rect -13650 79920 -13640 79990
rect -13860 79900 -13640 79920
rect -13360 79990 -13140 80040
rect -13360 79920 -13350 79990
rect -13150 79920 -13140 79990
rect -13360 79900 -13140 79920
rect -12860 79990 -12640 80040
rect -12860 79920 -12850 79990
rect -12650 79920 -12640 79990
rect -12860 79900 -12640 79920
rect -12360 79990 -12140 80040
rect -12360 79920 -12350 79990
rect -12150 79920 -12140 79990
rect -12360 79900 -12140 79920
rect -11860 79990 -11640 80040
rect -11860 79920 -11850 79990
rect -11650 79920 -11640 79990
rect -11860 79900 -11640 79920
rect -11360 79990 -11140 80040
rect -11360 79920 -11350 79990
rect -11150 79920 -11140 79990
rect -11360 79900 -11140 79920
rect -10860 79990 -10640 80040
rect -10860 79920 -10850 79990
rect -10650 79920 -10640 79990
rect -10860 79900 -10640 79920
rect -10360 79990 -10140 80040
rect -10360 79920 -10350 79990
rect -10150 79920 -10140 79990
rect -10360 79900 -10140 79920
rect -9860 79990 -9640 80040
rect -9860 79920 -9850 79990
rect -9650 79920 -9640 79990
rect -9860 79900 -9640 79920
rect -9360 79990 -9140 80040
rect -9360 79920 -9350 79990
rect -9150 79920 -9140 79990
rect -9360 79900 -9140 79920
rect -8860 79990 -8640 80040
rect -8860 79920 -8850 79990
rect -8650 79920 -8640 79990
rect -8860 79900 -8640 79920
rect -8360 79990 -8140 80040
rect -8360 79920 -8350 79990
rect -8150 79920 -8140 79990
rect -8360 79900 -8140 79920
rect -7860 79990 -7640 80040
rect -7860 79920 -7850 79990
rect -7650 79920 -7640 79990
rect -7860 79900 -7640 79920
rect -7360 79990 -7140 80040
rect -7360 79920 -7350 79990
rect -7150 79920 -7140 79990
rect -7360 79900 -7140 79920
rect -6860 79990 -6640 80040
rect -6860 79920 -6850 79990
rect -6650 79920 -6640 79990
rect -6860 79900 -6640 79920
rect -6360 79990 -6140 80040
rect -6360 79920 -6350 79990
rect -6150 79920 -6140 79990
rect -6360 79900 -6140 79920
rect -5860 79990 -5640 80040
rect -5860 79920 -5850 79990
rect -5650 79920 -5640 79990
rect -5860 79900 -5640 79920
rect -5360 79990 -5140 80040
rect -5360 79920 -5350 79990
rect -5150 79920 -5140 79990
rect -5360 79900 -5140 79920
rect -4860 79990 -4640 80040
rect -4860 79920 -4850 79990
rect -4650 79920 -4640 79990
rect -4860 79900 -4640 79920
rect -4360 79990 -4140 80040
rect -4360 79920 -4350 79990
rect -4150 79920 -4140 79990
rect -4360 79900 -4140 79920
rect -3860 79990 -3640 80040
rect -3860 79920 -3850 79990
rect -3650 79920 -3640 79990
rect -3860 79900 -3640 79920
rect -3360 79990 -3140 80040
rect -3360 79920 -3350 79990
rect -3150 79920 -3140 79990
rect -3360 79900 -3140 79920
rect -2860 79990 -2640 80040
rect -2860 79920 -2850 79990
rect -2650 79920 -2640 79990
rect -2860 79900 -2640 79920
rect -2360 79990 -2140 80040
rect -2360 79920 -2350 79990
rect -2150 79920 -2140 79990
rect -2360 79900 -2140 79920
rect -1860 79990 -1640 80040
rect -1860 79920 -1850 79990
rect -1650 79920 -1640 79990
rect -1860 79900 -1640 79920
rect -1360 79990 -1140 80040
rect -1360 79920 -1350 79990
rect -1150 79920 -1140 79990
rect -1360 79900 -1140 79920
rect -860 79990 -640 80040
rect -860 79920 -850 79990
rect -650 79920 -640 79990
rect -860 79900 -640 79920
rect -360 79990 -140 80040
rect -360 79920 -350 79990
rect -150 79920 -140 79990
rect -360 79900 -140 79920
rect 140 79990 360 80040
rect 140 79920 150 79990
rect 350 79920 360 79990
rect 140 79900 360 79920
rect 640 79990 860 80040
rect 640 79920 650 79990
rect 850 79920 860 79990
rect 640 79900 860 79920
rect 1140 79990 1360 80040
rect 1140 79920 1150 79990
rect 1350 79920 1360 79990
rect 1140 79900 1360 79920
rect 1640 79990 1860 80040
rect 1640 79920 1650 79990
rect 1850 79920 1860 79990
rect 1640 79900 1860 79920
rect 2140 79990 2360 80040
rect 2140 79920 2150 79990
rect 2350 79920 2360 79990
rect 2140 79900 2360 79920
rect 2640 79990 2860 80040
rect 2640 79920 2650 79990
rect 2850 79920 2860 79990
rect 2640 79900 2860 79920
rect 3140 79990 3360 80040
rect 3140 79920 3150 79990
rect 3350 79920 3360 79990
rect 3140 79900 3360 79920
rect 3640 79990 3860 80040
rect 3640 79920 3650 79990
rect 3850 79920 3860 79990
rect 3640 79900 3860 79920
rect 4140 79990 4360 80040
rect 4140 79920 4150 79990
rect 4350 79920 4360 79990
rect 4140 79900 4360 79920
rect 4640 79990 4860 80040
rect 4640 79920 4650 79990
rect 4850 79920 4860 79990
rect 4640 79900 4860 79920
rect 5140 79990 5360 80040
rect 5140 79920 5150 79990
rect 5350 79920 5360 79990
rect 5140 79900 5360 79920
rect 5640 79990 5860 80040
rect 5640 79920 5650 79990
rect 5850 79920 5860 79990
rect 5640 79900 5860 79920
rect 6140 79990 6360 80040
rect 6140 79920 6150 79990
rect 6350 79920 6360 79990
rect 6140 79900 6360 79920
rect 6640 79990 6860 80040
rect 6640 79920 6650 79990
rect 6850 79920 6860 79990
rect 6640 79900 6860 79920
rect 7140 79990 7360 80040
rect 7140 79920 7150 79990
rect 7350 79920 7360 79990
rect 7140 79900 7360 79920
rect 7640 79990 7860 80040
rect 7640 79920 7650 79990
rect 7850 79920 7860 79990
rect 7640 79900 7860 79920
rect 8140 79990 8360 80040
rect 8140 79920 8150 79990
rect 8350 79920 8360 79990
rect 8140 79900 8360 79920
rect 8640 79990 8860 80040
rect 8640 79920 8650 79990
rect 8850 79920 8860 79990
rect 8640 79900 8860 79920
rect 9140 79990 9360 80040
rect 9140 79920 9150 79990
rect 9350 79920 9360 79990
rect 9140 79900 9360 79920
rect 9640 79990 9860 80040
rect 9640 79920 9650 79990
rect 9850 79920 9860 79990
rect 9640 79900 9860 79920
rect 10140 79990 10360 80040
rect 10140 79920 10150 79990
rect 10350 79920 10360 79990
rect 10140 79900 10360 79920
rect 10640 79990 10860 80040
rect 10640 79920 10650 79990
rect 10850 79920 10860 79990
rect 10640 79900 10860 79920
rect 11140 79990 11360 80040
rect 11140 79920 11150 79990
rect 11350 79920 11360 79990
rect 11140 79900 11360 79920
rect 11640 79990 11860 80040
rect 11640 79920 11650 79990
rect 11850 79920 11860 79990
rect 11640 79900 11860 79920
rect 12140 79990 12360 80040
rect 12140 79920 12150 79990
rect 12350 79920 12360 79990
rect 12140 79900 12360 79920
rect 12640 79990 12860 80040
rect 12640 79920 12650 79990
rect 12850 79920 12860 79990
rect 12640 79900 12860 79920
rect 13140 79990 13360 80040
rect 13140 79920 13150 79990
rect 13350 79920 13360 79990
rect 13140 79900 13360 79920
rect 13640 79990 13860 80040
rect 13640 79920 13650 79990
rect 13850 79920 13860 79990
rect 13640 79900 13860 79920
rect 14140 79990 14360 80040
rect 14140 79920 14150 79990
rect 14350 79920 14360 79990
rect 14140 79900 14360 79920
rect 14640 79990 14860 80040
rect 14640 79920 14650 79990
rect 14850 79920 14860 79990
rect 14640 79900 14860 79920
rect 15140 79990 15360 80040
rect 15140 79920 15150 79990
rect 15350 79920 15360 79990
rect 15140 79900 15360 79920
rect 15640 79990 15860 80040
rect 15640 79920 15650 79990
rect 15850 79920 15860 79990
rect 15640 79900 15860 79920
rect 16140 79990 16360 80040
rect 16140 79920 16150 79990
rect 16350 79920 16360 79990
rect 16140 79900 16360 79920
rect 16640 79990 16860 80040
rect 16640 79920 16650 79990
rect 16850 79920 16860 79990
rect 16640 79900 16860 79920
rect 17140 79990 17360 80040
rect 17140 79920 17150 79990
rect 17350 79920 17360 79990
rect 17140 79900 17360 79920
rect 17640 79990 17860 80040
rect 17640 79920 17650 79990
rect 17850 79920 17860 79990
rect 17640 79900 17860 79920
rect 18140 79990 18360 80040
rect 18140 79920 18150 79990
rect 18350 79920 18360 79990
rect 18140 79900 18360 79920
rect 18640 79990 18860 80040
rect 18640 79920 18650 79990
rect 18850 79920 18860 79990
rect 18640 79900 18860 79920
rect 19140 79990 19360 80040
rect 19140 79920 19150 79990
rect 19350 79920 19360 79990
rect 19140 79900 19360 79920
rect 19640 79990 19860 80040
rect 19640 79920 19650 79990
rect 19850 79920 19860 79990
rect 19640 79900 19860 79920
rect 20140 79990 20360 80040
rect 20140 79920 20150 79990
rect 20350 79920 20360 79990
rect 20140 79900 20360 79920
rect 20640 79990 20860 80040
rect 20640 79920 20650 79990
rect 20850 79920 20860 79990
rect 20640 79900 20860 79920
rect 21140 79990 21360 80040
rect 21140 79920 21150 79990
rect 21350 79920 21360 79990
rect 21140 79900 21360 79920
rect 21640 79990 21860 80040
rect 21640 79920 21650 79990
rect 21850 79920 21860 79990
rect 21640 79900 21860 79920
rect 22140 79990 22360 80040
rect 22140 79920 22150 79990
rect 22350 79920 22360 79990
rect 22140 79900 22360 79920
rect 22640 79990 22860 80040
rect 22640 79920 22650 79990
rect 22850 79920 22860 79990
rect 22640 79900 22860 79920
rect 23140 79990 23360 80040
rect 23140 79920 23150 79990
rect 23350 79920 23360 79990
rect 23140 79900 23360 79920
rect 23640 79990 23860 80040
rect 23640 79920 23650 79990
rect 23850 79920 23860 79990
rect 23640 79900 23860 79920
rect 24140 79990 24360 80040
rect 24140 79920 24150 79990
rect 24350 79920 24360 79990
rect 24140 79900 24360 79920
rect 24640 79990 24860 80040
rect 24640 79920 24650 79990
rect 24850 79920 24860 79990
rect 24640 79900 24860 79920
rect 25140 79990 25360 80040
rect 25140 79920 25150 79990
rect 25350 79920 25360 79990
rect 25140 79900 25360 79920
rect 25640 79990 25860 80040
rect 25640 79920 25650 79990
rect 25850 79920 25860 79990
rect 25640 79900 25860 79920
rect 26140 79990 26360 80040
rect 26140 79920 26150 79990
rect 26350 79920 26360 79990
rect 26140 79900 26360 79920
rect 26640 79990 26860 80040
rect 26640 79920 26650 79990
rect 26850 79920 26860 79990
rect 26640 79900 26860 79920
rect 27140 79990 27360 80040
rect 27140 79920 27150 79990
rect 27350 79920 27360 79990
rect 27140 79900 27360 79920
rect 27640 79990 27860 80040
rect 27640 79920 27650 79990
rect 27850 79920 27860 79990
rect 27640 79900 27860 79920
rect 28140 79990 28360 80040
rect 28140 79920 28150 79990
rect 28350 79920 28360 79990
rect 28140 79900 28360 79920
rect 28640 79990 28860 80040
rect 28640 79920 28650 79990
rect 28850 79920 28860 79990
rect 28640 79900 28860 79920
rect 29140 79990 29360 80040
rect 29140 79920 29150 79990
rect 29350 79920 29360 79990
rect 29140 79900 29360 79920
rect 29640 79990 29860 80040
rect 29640 79920 29650 79990
rect 29850 79920 29860 79990
rect 29640 79900 29860 79920
rect 30140 79990 30360 80040
rect 30140 79920 30150 79990
rect 30350 79920 30360 79990
rect 30140 79900 30360 79920
rect 30640 79990 30860 80040
rect 30640 79920 30650 79990
rect 30850 79920 30860 79990
rect 30640 79900 30860 79920
rect 31140 79990 31360 80040
rect 31140 79920 31150 79990
rect 31350 79920 31360 79990
rect 31140 79900 31360 79920
rect 31640 79990 31860 80040
rect 31640 79920 31650 79990
rect 31850 79920 31860 79990
rect 31640 79900 31860 79920
rect 32140 79990 32360 80040
rect 32140 79920 32150 79990
rect 32350 79920 32360 79990
rect 32140 79900 32360 79920
rect 32640 79990 32860 80040
rect 32640 79920 32650 79990
rect 32850 79920 32860 79990
rect 32640 79900 32860 79920
rect 33140 79990 33360 80040
rect 33140 79920 33150 79990
rect 33350 79920 33360 79990
rect 33140 79900 33360 79920
rect 33640 79990 33860 80040
rect 33640 79920 33650 79990
rect 33850 79920 33860 79990
rect 33640 79900 33860 79920
rect 34140 79990 34360 80040
rect 34140 79920 34150 79990
rect 34350 79920 34360 79990
rect 34140 79900 34360 79920
rect 34640 79990 34860 80040
rect 34640 79920 34650 79990
rect 34850 79920 34860 79990
rect 34640 79900 34860 79920
rect 35140 79990 35360 80040
rect 35140 79920 35150 79990
rect 35350 79920 35360 79990
rect 35140 79900 35360 79920
rect 35640 79990 35860 80040
rect 35640 79920 35650 79990
rect 35850 79920 35860 79990
rect 35640 79900 35860 79920
rect 36140 79990 36360 80040
rect 36140 79920 36150 79990
rect 36350 79920 36360 79990
rect 36140 79900 36360 79920
rect 36640 79990 36860 80040
rect 36640 79920 36650 79990
rect 36850 79920 36860 79990
rect 36640 79900 36860 79920
rect 37140 79990 37360 80040
rect 37140 79920 37150 79990
rect 37350 79920 37360 79990
rect 37140 79900 37360 79920
rect 37640 79990 37860 80040
rect 37640 79920 37650 79990
rect 37850 79920 37860 79990
rect 37640 79900 37860 79920
rect 38140 79990 38360 80040
rect 38140 79920 38150 79990
rect 38350 79920 38360 79990
rect 38140 79900 38360 79920
rect 38640 79990 38860 80040
rect 38640 79920 38650 79990
rect 38850 79920 38860 79990
rect 38640 79900 38860 79920
rect 39140 79990 39360 80040
rect 39140 79920 39150 79990
rect 39350 79920 39360 79990
rect 39140 79900 39360 79920
rect 39640 79990 39860 80040
rect 39640 79920 39650 79990
rect 39850 79920 39860 79990
rect 39640 79900 39860 79920
rect 40140 79990 40360 80040
rect 40140 79920 40150 79990
rect 40350 79920 40360 79990
rect 40140 79900 40360 79920
rect 40640 79990 40860 80040
rect 40640 79920 40650 79990
rect 40850 79920 40860 79990
rect 40640 79900 40860 79920
rect 41140 79990 41360 80040
rect 41140 79920 41150 79990
rect 41350 79920 41360 79990
rect 41140 79900 41360 79920
rect 41640 79990 41860 80040
rect 41640 79920 41650 79990
rect 41850 79920 41860 79990
rect 41640 79900 41860 79920
rect 42140 79990 42360 80040
rect 42140 79920 42150 79990
rect 42350 79920 42360 79990
rect 42140 79900 42360 79920
rect 42640 79990 42860 80040
rect 42640 79920 42650 79990
rect 42850 79920 42860 79990
rect 42640 79900 42860 79920
rect 43140 79990 43360 80040
rect 43140 79920 43150 79990
rect 43350 79920 43360 79990
rect 43140 79900 43360 79920
rect 43640 79990 43860 80040
rect 43640 79920 43650 79990
rect 43850 79920 43860 79990
rect 43640 79900 43860 79920
rect 44140 79990 44360 80040
rect 44140 79920 44150 79990
rect 44350 79920 44360 79990
rect 44140 79900 44360 79920
rect 44640 79990 44860 80040
rect 44640 79920 44650 79990
rect 44850 79920 44860 79990
rect 44640 79900 44860 79920
rect 45140 79990 45360 80040
rect 45140 79920 45150 79990
rect 45350 79920 45360 79990
rect 45140 79900 45360 79920
rect 45640 79990 45860 80040
rect 45640 79920 45650 79990
rect 45850 79920 45860 79990
rect 45640 79900 45860 79920
rect 46140 79990 46360 80040
rect 46140 79920 46150 79990
rect 46350 79920 46360 79990
rect 46140 79900 46360 79920
rect 46640 79990 46860 80040
rect 46640 79920 46650 79990
rect 46850 79920 46860 79990
rect 46640 79900 46860 79920
rect 47140 79990 47360 80040
rect 47140 79920 47150 79990
rect 47350 79920 47360 79990
rect 47140 79900 47360 79920
rect 47640 79990 47860 80040
rect 47640 79920 47650 79990
rect 47850 79920 47860 79990
rect 47640 79900 47860 79920
rect 48140 79990 48360 80040
rect 48140 79920 48150 79990
rect 48350 79920 48360 79990
rect 48140 79900 48360 79920
rect 48640 79990 48860 80040
rect 48640 79920 48650 79990
rect 48850 79920 48860 79990
rect 48640 79900 48860 79920
rect 49140 79990 49360 80040
rect 49140 79920 49150 79990
rect 49350 79920 49360 79990
rect 49140 79900 49360 79920
rect 49640 79990 49860 80040
rect 49640 79920 49650 79990
rect 49850 79920 49860 79990
rect 49640 79900 49860 79920
rect 50140 79990 50360 80040
rect 50140 79920 50150 79990
rect 50350 79920 50360 79990
rect 50140 79900 50360 79920
rect 50640 79990 50860 80040
rect 50640 79920 50650 79990
rect 50850 79920 50860 79990
rect 50640 79900 50860 79920
rect 51140 79990 51360 80040
rect 51140 79920 51150 79990
rect 51350 79920 51360 79990
rect 51140 79900 51360 79920
rect 51640 79990 51860 80040
rect 51640 79920 51650 79990
rect 51850 79920 51860 79990
rect 51640 79900 51860 79920
rect 52140 79990 52360 80040
rect 52140 79920 52150 79990
rect 52350 79920 52360 79990
rect 52140 79900 52360 79920
rect 52640 79990 52860 80040
rect 52640 79920 52650 79990
rect 52850 79920 52860 79990
rect 52640 79900 52860 79920
rect 53140 79990 53360 80040
rect 53140 79920 53150 79990
rect 53350 79920 53360 79990
rect 53140 79900 53360 79920
rect 53640 79990 53860 80040
rect 53640 79920 53650 79990
rect 53850 79920 53860 79990
rect 53640 79900 53860 79920
rect 54140 79990 54360 80040
rect 54140 79920 54150 79990
rect 54350 79920 54360 79990
rect 54140 79900 54360 79920
rect 54640 79990 54860 80040
rect 54640 79920 54650 79990
rect 54850 79920 54860 79990
rect 54640 79900 54860 79920
rect 55140 79990 55360 80040
rect 55140 79920 55150 79990
rect 55350 79920 55360 79990
rect 55140 79900 55360 79920
rect 55640 79990 55860 80040
rect 55640 79920 55650 79990
rect 55850 79920 55860 79990
rect 55640 79900 55860 79920
rect 56140 79990 56360 80040
rect 56140 79920 56150 79990
rect 56350 79920 56360 79990
rect 56140 79900 56360 79920
rect 56640 79990 56860 80040
rect 56640 79920 56650 79990
rect 56850 79920 56860 79990
rect 56640 79900 56860 79920
rect 57140 79990 57360 80040
rect 57140 79920 57150 79990
rect 57350 79920 57360 79990
rect 57140 79900 57360 79920
rect 57640 79990 57860 80040
rect 57640 79920 57650 79990
rect 57850 79920 57860 79990
rect 57640 79900 57860 79920
rect 58140 79990 58360 80040
rect 58140 79920 58150 79990
rect 58350 79920 58360 79990
rect 58140 79900 58360 79920
rect 58640 79990 58860 80040
rect 58640 79920 58650 79990
rect 58850 79920 58860 79990
rect 58640 79900 58860 79920
rect 59140 79990 59360 80040
rect 59140 79920 59150 79990
rect 59350 79920 59360 79990
rect 59140 79900 59360 79920
rect 59640 79990 59860 80040
rect 59640 79920 59650 79990
rect 59850 79920 59860 79990
rect 59640 79900 59860 79920
rect 60140 79990 60360 80040
rect 60140 79920 60150 79990
rect 60350 79920 60360 79990
rect 60140 79900 60360 79920
rect 60640 79990 60860 80040
rect 60640 79920 60650 79990
rect 60850 79920 60860 79990
rect 60640 79900 60860 79920
rect 61140 79990 61360 80040
rect 61140 79920 61150 79990
rect 61350 79920 61360 79990
rect 61140 79900 61360 79920
rect 61640 79990 61860 80040
rect 61640 79920 61650 79990
rect 61850 79920 61860 79990
rect 61640 79900 61860 79920
rect 62140 79990 62360 80040
rect 62140 79920 62150 79990
rect 62350 79920 62360 79990
rect 62140 79900 62360 79920
rect 62640 79990 62860 80040
rect 62640 79920 62650 79990
rect 62850 79920 62860 79990
rect 62640 79900 62860 79920
rect 63140 79990 63360 80040
rect 63140 79920 63150 79990
rect 63350 79920 63360 79990
rect 63140 79900 63360 79920
rect 63640 79990 63860 80040
rect 63640 79920 63650 79990
rect 63850 79920 63860 79990
rect 63640 79900 63860 79920
rect 64140 79990 64360 80040
rect 64140 79920 64150 79990
rect 64350 79920 64360 79990
rect 64140 79900 64360 79920
rect 64640 79990 64860 80040
rect 64640 79920 64650 79990
rect 64850 79920 64860 79990
rect 64640 79900 64860 79920
rect 65140 79990 65360 80040
rect 65140 79920 65150 79990
rect 65350 79920 65360 79990
rect 65140 79900 65360 79920
rect 65640 79990 65860 80040
rect 65640 79920 65650 79990
rect 65850 79920 65860 79990
rect 65640 79900 65860 79920
rect 66140 79990 66360 80040
rect 66140 79920 66150 79990
rect 66350 79920 66360 79990
rect 66140 79900 66360 79920
rect 66640 79990 66860 80040
rect 66640 79920 66650 79990
rect 66850 79920 66860 79990
rect 66640 79900 66860 79920
rect 67140 79990 67360 80040
rect 67140 79920 67150 79990
rect 67350 79920 67360 79990
rect 67140 79900 67360 79920
rect 67640 79990 67860 80040
rect 67640 79920 67650 79990
rect 67850 79920 67860 79990
rect 67640 79900 67860 79920
rect 68140 79990 68360 80040
rect 68140 79920 68150 79990
rect 68350 79920 68360 79990
rect 68140 79900 68360 79920
rect 68640 79990 68860 80040
rect 68640 79920 68650 79990
rect 68850 79920 68860 79990
rect 68640 79900 68860 79920
rect 69140 79990 69360 80040
rect 69140 79920 69150 79990
rect 69350 79920 69360 79990
rect 69140 79900 69360 79920
rect 69640 79990 69860 80040
rect 69640 79920 69650 79990
rect 69850 79920 69860 79990
rect 69640 79900 69860 79920
rect 70140 79990 70360 80040
rect 70140 79920 70150 79990
rect 70350 79920 70360 79990
rect 70140 79900 70360 79920
rect 70640 79990 70860 80040
rect 70640 79920 70650 79990
rect 70850 79920 70860 79990
rect 70640 79900 70860 79920
rect 71140 79990 71360 80040
rect 71140 79920 71150 79990
rect 71350 79920 71360 79990
rect 71140 79900 71360 79920
rect 71640 79990 71860 80040
rect 71640 79920 71650 79990
rect 71850 79920 71860 79990
rect 71640 79900 71860 79920
rect 72140 79990 72360 80040
rect 72140 79920 72150 79990
rect 72350 79920 72360 79990
rect 72140 79900 72360 79920
rect 72640 79990 72860 80040
rect 72640 79920 72650 79990
rect 72850 79920 72860 79990
rect 72640 79900 72860 79920
rect 73140 79990 73360 80040
rect 73140 79920 73150 79990
rect 73350 79920 73360 79990
rect 73140 79900 73360 79920
rect 73640 79990 73860 80040
rect 73640 79920 73650 79990
rect 73850 79920 73860 79990
rect 73640 79900 73860 79920
rect 74140 79990 74360 80040
rect 74140 79920 74150 79990
rect 74350 79920 74360 79990
rect 74140 79900 74360 79920
rect 74640 79990 74860 80040
rect 74640 79920 74650 79990
rect 74850 79920 74860 79990
rect 74640 79900 74860 79920
rect 75140 79990 75360 80040
rect 75140 79920 75150 79990
rect 75350 79920 75360 79990
rect 75140 79900 75360 79920
rect 75640 79990 75860 80040
rect 75640 79920 75650 79990
rect 75850 79920 75860 79990
rect 75640 79900 75860 79920
rect 76140 79990 76360 80040
rect 76140 79920 76150 79990
rect 76350 79920 76360 79990
rect 76140 79900 76360 79920
rect 76640 79990 76860 80040
rect 76640 79920 76650 79990
rect 76850 79920 76860 79990
rect 76640 79900 76860 79920
rect 77140 79990 77360 80040
rect 77140 79920 77150 79990
rect 77350 79920 77360 79990
rect 77140 79900 77360 79920
rect 77640 79990 77860 80040
rect 77640 79920 77650 79990
rect 77850 79920 77860 79990
rect 77640 79900 77860 79920
rect 78140 79990 78360 80040
rect 78140 79920 78150 79990
rect 78350 79920 78360 79990
rect 78140 79900 78360 79920
rect 78640 79990 78860 80040
rect 78640 79920 78650 79990
rect 78850 79920 78860 79990
rect 78640 79900 78860 79920
rect 79140 79990 79360 80040
rect 79140 79920 79150 79990
rect 79350 79920 79360 79990
rect 79140 79900 79360 79920
rect 79640 79990 79860 80040
rect 79640 79920 79650 79990
rect 79850 79920 79860 79990
rect 79640 79900 79860 79920
rect 80140 79990 80360 80040
rect 80140 79920 80150 79990
rect 80350 79920 80360 79990
rect 80140 79900 80360 79920
rect 80640 79990 80860 80040
rect 80640 79920 80650 79990
rect 80850 79920 80860 79990
rect 80640 79900 80860 79920
rect 81140 79990 81360 80040
rect 81140 79920 81150 79990
rect 81350 79920 81360 79990
rect 81140 79900 81360 79920
rect 81640 79990 81860 80040
rect 81640 79920 81650 79990
rect 81850 79920 81860 79990
rect 81640 79900 81860 79920
rect 82140 79990 82360 80040
rect 82140 79920 82150 79990
rect 82350 79920 82360 79990
rect 82140 79900 82360 79920
rect 82640 79990 82860 80040
rect 82640 79920 82650 79990
rect 82850 79920 82860 79990
rect 82640 79900 82860 79920
rect 83140 79990 83360 80040
rect 83140 79920 83150 79990
rect 83350 79920 83360 79990
rect 83140 79900 83360 79920
rect 83640 79990 83860 80040
rect 83640 79920 83650 79990
rect 83850 79920 83860 79990
rect 83640 79900 83860 79920
rect 84140 79990 84360 80040
rect 84140 79920 84150 79990
rect 84350 79920 84360 79990
rect 84140 79900 84360 79920
rect 84640 79990 84860 80040
rect 84640 79920 84650 79990
rect 84850 79920 84860 79990
rect 84640 79900 84860 79920
rect 85140 79990 85360 80040
rect 85140 79920 85150 79990
rect 85350 79920 85360 79990
rect 85140 79900 85360 79920
rect 85640 79990 85860 80040
rect 85640 79920 85650 79990
rect 85850 79920 85860 79990
rect 85640 79900 85860 79920
rect 86140 79990 86360 80040
rect 86140 79920 86150 79990
rect 86350 79920 86360 79990
rect 86140 79900 86360 79920
rect 86640 79990 86860 80040
rect 86640 79920 86650 79990
rect 86850 79920 86860 79990
rect 86640 79900 86860 79920
rect 87140 79990 87360 80040
rect 87140 79920 87150 79990
rect 87350 79920 87360 79990
rect 87140 79900 87360 79920
rect 87640 79990 87860 80040
rect 87640 79920 87650 79990
rect 87850 79920 87860 79990
rect 87640 79900 87860 79920
rect 88140 79990 88360 80040
rect 88140 79920 88150 79990
rect 88350 79920 88360 79990
rect 88140 79900 88360 79920
rect 88640 79990 88860 80040
rect 88640 79920 88650 79990
rect 88850 79920 88860 79990
rect 88640 79900 88860 79920
rect 89140 79990 89360 80040
rect 89140 79920 89150 79990
rect 89350 79920 89360 79990
rect 89140 79900 89360 79920
rect 89640 79990 89860 80040
rect 89640 79920 89650 79990
rect 89850 79920 89860 79990
rect 89640 79900 89860 79920
rect 90140 79990 90360 80040
rect 90140 79920 90150 79990
rect 90350 79920 90360 79990
rect 90140 79900 90360 79920
rect 90640 79990 90860 80040
rect 90640 79920 90650 79990
rect 90850 79920 90860 79990
rect 90640 79900 90860 79920
rect 91140 79990 91360 80040
rect 91140 79920 91150 79990
rect 91350 79920 91360 79990
rect 91140 79900 91360 79920
rect 91640 79990 91860 80040
rect 91640 79920 91650 79990
rect 91850 79920 91860 79990
rect 91640 79900 91860 79920
rect 92140 79990 92360 80040
rect 92140 79920 92150 79990
rect 92350 79920 92360 79990
rect 92140 79900 92360 79920
rect 92640 79990 92860 80040
rect 92640 79920 92650 79990
rect 92850 79920 92860 79990
rect 92640 79900 92860 79920
rect 93140 79990 93360 80040
rect 93140 79920 93150 79990
rect 93350 79920 93360 79990
rect 93140 79900 93360 79920
rect 93640 79990 93860 80040
rect 93640 79920 93650 79990
rect 93850 79920 93860 79990
rect 93640 79900 93860 79920
rect 94140 79990 94360 80040
rect 94140 79920 94150 79990
rect 94350 79920 94360 79990
rect 94140 79900 94360 79920
rect 94640 79990 94860 80040
rect 94640 79920 94650 79990
rect 94850 79920 94860 79990
rect 94640 79900 94860 79920
rect 95140 79990 95360 80040
rect 95140 79920 95150 79990
rect 95350 79920 95360 79990
rect 95140 79900 95360 79920
rect 95640 79990 95860 80040
rect 95640 79920 95650 79990
rect 95850 79920 95860 79990
rect 95640 79900 95860 79920
rect 96140 79990 96360 80040
rect 96140 79920 96150 79990
rect 96350 79920 96360 79990
rect 96140 79900 96360 79920
rect 96640 79990 96860 80040
rect 96640 79920 96650 79990
rect 96850 79920 96860 79990
rect 96640 79900 96860 79920
rect 97140 79990 97360 80040
rect 97140 79920 97150 79990
rect 97350 79920 97360 79990
rect 97140 79900 97360 79920
rect 97640 79990 97860 80040
rect 97640 79920 97650 79990
rect 97850 79920 97860 79990
rect 97640 79900 97860 79920
rect 98140 79990 98360 80040
rect 98140 79920 98150 79990
rect 98350 79920 98360 79990
rect 98140 79900 98360 79920
rect 98640 79990 98860 80040
rect 98640 79920 98650 79990
rect 98850 79920 98860 79990
rect 98640 79900 98860 79920
rect 99140 79990 99360 80040
rect 99140 79920 99150 79990
rect 99350 79920 99360 79990
rect 99140 79900 99360 79920
rect 99640 79990 99860 80040
rect 99640 79920 99650 79990
rect 99850 79920 99860 79990
rect 99640 79900 99860 79920
rect 100140 79990 100360 80040
rect 100140 79920 100150 79990
rect 100350 79920 100360 79990
rect 100140 79900 100360 79920
rect 16000 13700 20000 13900
rect 13400 10200 14200 10220
rect 13400 9900 13560 10200
rect 14180 9900 14200 10200
rect 13400 9160 14200 9900
rect 13400 1800 13700 9160
rect 13400 1400 15300 1800
rect -23500 -12000 -22700 -11950
rect -23700 -16300 -23450 -12000
rect -22750 -16300 -22700 -12000
rect 14700 -12300 15300 1400
rect 14700 -12900 18300 -12300
rect -23700 -16350 -22700 -16300
rect -23700 -17000 -23000 -16350
rect -23700 -17200 -22700 -17000
rect -23700 -17400 -23000 -17200
rect -23700 -17600 -22700 -17400
rect -23700 -17800 -23000 -17600
rect -23700 -18000 -22700 -17800
rect -23700 -18200 -23000 -18000
rect -23700 -18400 -22700 -18200
rect -23700 -18600 -23000 -18400
rect -23700 -18800 -22700 -18600
rect -23700 -19000 -23000 -18800
rect -23700 -19200 -22700 -19000
rect -23700 -19400 -23000 -19200
rect -23700 -19600 -22700 -19400
rect -23700 -19800 -23000 -19600
rect -23700 -20000 -22700 -19800
rect -23700 -20200 -23000 -20000
rect -23700 -20400 -22700 -20200
rect 17700 -20300 18300 -12900
rect -23700 -20600 -23000 -20400
rect -23700 -20800 -22700 -20600
rect 17700 -20900 20300 -20300
rect 19700 -28300 20300 -20900
rect 23500 -28200 24000 -5600
rect 32800 -28200 34000 -20100
rect 19700 -28700 22300 -28300
rect 23500 -28500 26000 -28200
rect 30800 -28500 34000 -28200
rect 34900 -28400 36300 -28300
rect 34900 -28700 35000 -28400
rect 19700 -28800 35000 -28700
rect 36200 -28800 36300 -28400
rect 19700 -28900 36300 -28800
rect 22640 -29120 22860 -29100
rect 22640 -29190 22650 -29120
rect 22850 -29190 22860 -29120
rect 22640 -29240 22860 -29190
rect 23140 -29120 23360 -29100
rect 23140 -29190 23150 -29120
rect 23350 -29190 23360 -29120
rect 23140 -29240 23360 -29190
rect 23500 -29240 24000 -29100
rect 22500 -29250 24000 -29240
rect 22500 -29450 22520 -29250
rect 22590 -29450 22910 -29250
rect 22980 -29450 23020 -29250
rect 23090 -29450 23410 -29250
rect 23480 -29450 24000 -29250
rect 22500 -29460 24000 -29450
rect 22640 -29510 22860 -29460
rect 22640 -29580 22650 -29510
rect 22850 -29580 22860 -29510
rect 22640 -29600 22860 -29580
rect 23140 -29510 23360 -29460
rect 23140 -29580 23150 -29510
rect 23350 -29580 23360 -29510
rect 23140 -29600 23360 -29580
rect 23500 -30500 24000 -29460
rect 32800 -30500 34000 -29100
rect 23500 -30700 26000 -30500
rect 23500 -33200 24200 -30700
rect 25800 -31000 26000 -30700
rect 30800 -30700 34000 -30500
rect 30800 -31000 31000 -30700
rect 25800 -33200 31000 -31000
rect 32600 -32100 34000 -30700
rect 32600 -33200 32800 -32100
rect 23500 -33600 32800 -33200
rect -19600 -38100 -19500 -35700
<< via2 >>
rect 13560 9900 14180 10200
rect -23450 -16300 -22750 -12000
rect 35000 -28800 36200 -28400
rect 22650 -29190 22850 -29120
rect 23150 -29190 23350 -29120
rect 22520 -29450 22590 -29250
rect 22910 -29450 22980 -29250
rect 23020 -29450 23090 -29250
rect 23410 -29450 23480 -29250
rect 22650 -29580 22850 -29510
rect 23150 -29580 23350 -29510
rect 24200 -33200 25800 -30700
rect 31000 -33200 32600 -30700
<< metal3 >>
rect -30500 62700 -6500 74900
rect -30500 61100 -30300 62700
rect -20300 61100 -16700 62700
rect -6700 61100 -6500 62700
rect -30500 60100 -6500 61100
rect -30500 49100 -19300 60100
rect -17700 49100 -6500 60100
rect 9500 64700 35500 64900
rect 9500 54700 21700 64700
rect 23300 54700 35500 64700
rect 9500 53700 35500 54700
rect 9500 52100 9700 53700
rect 20700 52100 35500 53700
rect 9500 51900 35500 52100
rect 37500 64700 63500 64900
rect 37500 54700 49700 64700
rect 51300 54700 63500 64700
rect 37500 53700 63500 54700
rect 37500 52100 37700 53700
rect 48700 52100 63500 53700
rect -30500 48900 -6500 49100
rect 37500 51100 63500 52100
rect 37500 41100 49700 51100
rect 51300 41100 63500 51100
rect 37500 40900 63500 41100
rect 65500 64700 91500 64900
rect 65500 54700 77700 64700
rect 79300 54700 91500 64700
rect 65500 53700 91500 54700
rect 65500 52100 65700 53700
rect 76700 52100 91500 53700
rect 65500 51100 91500 52100
rect 65500 41100 77700 51100
rect 79300 41100 91500 51100
rect 65500 40900 91500 41100
rect -22500 26700 -12500 37900
rect 136700 36700 141500 36900
rect 136700 27100 136900 36700
rect 141300 34300 141500 36700
rect 141300 29300 143500 34300
rect 141300 27100 141500 29300
rect 136700 26900 141500 27100
rect -22500 25100 -22300 26700
rect -12700 25100 -12500 26700
rect -22500 24900 -12500 25100
rect -14700 13850 -14300 13900
rect -14700 12650 -14650 13850
rect -14350 13000 -14300 13850
rect 16000 13700 20000 13900
rect -14350 12650 -12000 13000
rect -14700 12600 -12000 12650
rect -13200 11850 -12800 12000
rect -14850 11550 -12800 11850
rect -13200 9600 -12800 11550
rect -12400 10400 -12000 12600
rect -12400 10000 -3800 10400
rect -13200 9200 -4600 9600
rect -18300 8200 -18100 8800
rect -22600 8000 -18100 8200
rect -22600 -1300 -22400 8000
rect -17600 7900 -17400 8800
rect -23400 -1400 -22400 -1300
rect -22300 7700 -17400 7900
rect -28000 -8100 -27500 -7600
rect -23400 -8300 -23200 -1400
rect -22300 -1500 -22100 7700
rect -17200 7600 -17000 8800
rect -27200 -8400 -23200 -8300
rect -23100 -1600 -22100 -1500
rect -22000 7400 -17000 7600
rect -27200 -16400 -27000 -8400
rect -23100 -8500 -22900 -1600
rect -22000 -1700 -21800 7400
rect -16400 7300 -16200 8800
rect -31300 -16500 -27000 -16400
rect -26900 -8600 -22900 -8500
rect -22800 -1800 -21800 -1700
rect -21700 7100 -16200 7300
rect -31300 -28500 -31100 -16500
rect -26900 -16600 -26700 -8600
rect -22800 -8700 -22600 -1800
rect -21700 -1900 -21500 7100
rect -16000 7000 -15800 8800
rect -31000 -16700 -26700 -16600
rect -26600 -8800 -22600 -8700
rect -22500 -2000 -21500 -1900
rect -21400 6800 -15800 7000
rect -31000 -28900 -30800 -16700
rect -26600 -16800 -26400 -8800
rect -22500 -8900 -22300 -2000
rect -21400 -2100 -21200 6800
rect -21000 5900 -15800 6500
rect -5000 6000 -4600 9200
rect -4200 6000 -3800 10000
rect 10700 4500 12500 8600
rect 10700 700 12400 4500
rect -13100 -1300 -13000 400
rect -30700 -16900 -26400 -16800
rect -26300 -9000 -22300 -8900
rect -22200 -2200 -21200 -2100
rect -21000 -1400 -13000 -1300
rect -30700 -29300 -30500 -16900
rect -26300 -17000 -26100 -9000
rect -22200 -9100 -22000 -2200
rect -21000 -2400 -20800 -1400
rect -12900 -1500 -12800 400
rect -30400 -17100 -26100 -17000
rect -26000 -9200 -22000 -9100
rect -21900 -2500 -20800 -2400
rect -20700 -1600 -12800 -1500
rect -30400 -29700 -30200 -17100
rect -26000 -17200 -25800 -9200
rect -21900 -9400 -21700 -2500
rect -20700 -2600 -20500 -1600
rect -12700 -1700 -12600 400
rect -30100 -17300 -25800 -17200
rect -25300 -9500 -21700 -9400
rect -21600 -2700 -20500 -2600
rect -20400 -1800 -12600 -1700
rect -30100 -30100 -29900 -17300
rect -25300 -30000 -25100 -9500
rect -21600 -9600 -21400 -2700
rect -20400 -2800 -20200 -1800
rect -12500 -1900 -12400 400
rect -25000 -9700 -21400 -9600
rect -21300 -2900 -20200 -2800
rect -20100 -2000 -12400 -1900
rect -25000 -30000 -24800 -9700
rect -21300 -9800 -21100 -2900
rect -20100 -3000 -19900 -2000
rect -12300 -2100 -12200 400
rect -24700 -9900 -21100 -9800
rect -21000 -3100 -19900 -3000
rect -19800 -2200 -12200 -2100
rect -24700 -30000 -24500 -9900
rect -21000 -10000 -20800 -3100
rect -19800 -3200 -19600 -2200
rect -24400 -10100 -20800 -10000
rect -20700 -3300 -19600 -3200
rect -24400 -30000 -24200 -10100
rect -20700 -10200 -20500 -3300
rect -24100 -10300 -20500 -10200
rect -24100 -30000 -23900 -10300
rect -23500 -12000 -22700 -11950
rect -23500 -16300 -23450 -12000
rect -22750 -16300 -22700 -12000
rect -23500 -16350 -22700 -16300
rect -22500 -16400 -18000 -11900
rect -23600 -19600 -22400 -19400
rect -23600 -21400 -23500 -19600
rect -23800 -21600 -23500 -21400
rect -23400 -19900 -22400 -19700
rect -23800 -30000 -23600 -21600
rect -23400 -21700 -23300 -19900
rect -23500 -30000 -23300 -21700
rect -23200 -20200 -22400 -20000
rect -23200 -21900 -23100 -20200
rect -23000 -20500 -22400 -20300
rect -23000 -21700 -22900 -20500
rect -22800 -20800 -22400 -20600
rect -22800 -21400 -22700 -20800
rect -22800 -21600 -22400 -21400
rect -23000 -21800 -22700 -21700
rect -23200 -30000 -23000 -21900
rect -22900 -30000 -22700 -21800
rect -22600 -30000 -22400 -21600
rect 23500 -28200 24000 -5600
rect 32800 -28200 34000 -20100
rect 23500 -28600 26000 -28200
rect 23500 -29100 24200 -28600
rect 22500 -29120 24200 -29100
rect 22500 -29190 22650 -29120
rect 22850 -29190 23150 -29120
rect 23350 -29190 24200 -29120
rect 22500 -29200 24200 -29190
rect 22500 -29220 22620 -29200
rect 22880 -29220 23120 -29200
rect 23380 -29220 24200 -29200
rect 22500 -29250 22600 -29220
rect 22500 -29450 22520 -29250
rect 22590 -29450 22600 -29250
rect 22500 -29480 22600 -29450
rect 22900 -29250 23100 -29220
rect 22900 -29450 22910 -29250
rect 22980 -29450 23020 -29250
rect 23090 -29450 23100 -29250
rect 22900 -29480 23100 -29450
rect 23400 -29250 24200 -29220
rect 23400 -29450 23410 -29250
rect 23480 -29450 24200 -29250
rect 23400 -29480 24200 -29450
rect 22500 -29500 22620 -29480
rect 22880 -29500 23120 -29480
rect 23380 -29500 24200 -29480
rect 22500 -29510 24200 -29500
rect 22500 -29580 22650 -29510
rect 22850 -29580 23150 -29510
rect 23350 -29580 24200 -29510
rect 22500 -29600 24200 -29580
rect 23500 -33200 24200 -29600
rect 25800 -31000 26000 -28600
rect 30800 -28600 34000 -28200
rect 30800 -31000 31000 -28600
rect 25800 -33200 31000 -31000
rect 32600 -32100 34000 -28600
rect 34900 -28400 36300 -28300
rect 34900 -28800 35000 -28400
rect 36200 -28800 36300 -28400
rect 34900 -28900 36300 -28800
rect 32600 -33200 32800 -32100
rect 23500 -33600 32800 -33200
rect 124700 -32600 134300 -32500
rect 26600 -34100 30200 -34000
rect -22500 -35000 -21900 -34900
rect -22500 -35400 -22400 -35000
rect -22000 -35400 -21900 -35000
rect 26600 -35300 26700 -34100
rect 30100 -35300 30200 -34100
rect 26600 -35400 30200 -35300
rect 124700 -35400 124800 -32600
rect 125100 -35400 134300 -32600
rect -22500 -35500 -21900 -35400
rect 124700 -35500 134300 -35400
rect -27300 -36030 -25140 -35840
rect -27300 -36100 -25500 -36030
rect -27300 -37700 -27100 -36100
rect -25900 -36220 -25500 -36100
rect -25900 -36460 -25140 -36220
rect -25900 -36740 -25500 -36460
rect -22500 -36700 -22100 -35500
rect -25900 -37000 -25140 -36740
rect -25900 -37280 -25500 -37000
rect -25900 -37540 -25150 -37280
rect -25900 -37700 -25500 -37540
rect -27300 -37730 -25500 -37700
rect -27300 -37920 -25290 -37730
rect -22530 -40060 -22020 -37560
rect -19600 -38100 -19500 -35700
rect 127200 -36300 127700 -35500
<< via3 >>
rect -30300 61100 -20300 62700
rect -16700 61100 -6700 62700
rect -19300 49100 -17700 60100
rect 21700 54700 23300 64700
rect 9700 52100 20700 53700
rect 49700 54700 51300 64700
rect 37700 52100 48700 53700
rect 49700 41100 51300 51100
rect 77700 54700 79300 64700
rect 65700 52100 76700 53700
rect 77700 41100 79300 51100
rect 136900 27100 141300 36700
rect -22300 25100 -12700 26700
rect -14650 12650 -14350 13850
rect -23450 -16300 -22750 -12000
rect 24200 -30700 25800 -28600
rect 24200 -33200 25800 -30700
rect 31000 -30700 32600 -28600
rect 31000 -33200 32600 -30700
rect 35000 -28800 36200 -28400
rect -22400 -35400 -22000 -35000
rect 26700 -35300 30100 -34100
rect 124800 -35400 125100 -32600
rect -27100 -37700 -25900 -36100
<< mimcap >>
rect -30300 74500 -20300 74700
rect -30300 63900 -30100 74500
rect -20500 63900 -20300 74500
rect -30300 63700 -20300 63900
rect -16700 74500 -6700 74700
rect -16700 63900 -16500 74500
rect -6900 63900 -6700 74500
rect -16700 63700 -6700 63900
rect 9700 64500 20700 64700
rect -30300 59900 -20300 60100
rect -30300 49300 -30100 59900
rect -20500 49300 -20300 59900
rect -30300 49100 -20300 49300
rect -16700 59900 -6700 60100
rect -16700 49300 -16500 59900
rect -6900 49300 -6700 59900
rect 9700 54900 9900 64500
rect 20500 54900 20700 64500
rect 9700 54700 20700 54900
rect 24300 64500 35300 64700
rect 24300 54900 24500 64500
rect 35100 54900 35300 64500
rect 24300 54700 35300 54900
rect 37700 64500 48700 64700
rect 37700 54900 37900 64500
rect 48500 54900 48700 64500
rect 37700 54700 48700 54900
rect 52300 64500 63300 64700
rect 52300 54900 52500 64500
rect 63100 54900 63300 64500
rect 52300 54700 63300 54900
rect 65700 64500 76700 64700
rect 65700 54900 65900 64500
rect 76500 54900 76700 64500
rect 65700 54700 76700 54900
rect 80300 64500 91300 64700
rect 80300 54900 80500 64500
rect 91100 54900 91300 64500
rect 80300 54700 91300 54900
rect -16700 49100 -6700 49300
rect 37700 50900 48700 51100
rect 37700 41300 37900 50900
rect 48500 41300 48700 50900
rect 37700 41100 48700 41300
rect 52300 50900 63300 51100
rect 52300 41300 52500 50900
rect 63100 41300 63300 50900
rect 52300 41100 63300 41300
rect 65700 50900 76700 51100
rect 65700 41300 65900 50900
rect 76500 41300 76700 50900
rect 65700 41100 76700 41300
rect 80300 50900 91300 51100
rect 80300 41300 80500 50900
rect 91100 41300 91300 50900
rect 80300 41100 91300 41300
rect -22300 37500 -12700 37700
rect -22300 27900 -22100 37500
rect -12900 27900 -12700 37500
rect -22300 27700 -12700 27900
rect -22400 -12100 -18300 -12000
rect -22400 -16200 -22300 -12100
rect -18400 -16200 -18300 -12100
rect -22400 -16300 -18300 -16200
rect 125700 -32700 134200 -32600
rect 125700 -35300 125800 -32700
rect 134100 -35300 134200 -32700
rect 125700 -35400 134200 -35300
<< mimcapcontact >>
rect -30100 63900 -20500 74500
rect -16500 63900 -6900 74500
rect -30100 49300 -20500 59900
rect -16500 49300 -6900 59900
rect 9900 54900 20500 64500
rect 24500 54900 35100 64500
rect 37900 54900 48500 64500
rect 52500 54900 63100 64500
rect 65900 54900 76500 64500
rect 80500 54900 91100 64500
rect 37900 41300 48500 50900
rect 52500 41300 63100 50900
rect 65900 41300 76500 50900
rect 80500 41300 91100 50900
rect -22100 27900 -12900 37500
rect -22300 -16200 -18400 -12100
rect 125800 -35300 134100 -32700
<< metal4 >>
rect 113500 82700 113900 82900
rect 114500 82700 115500 82900
rect 115900 82700 116900 82900
rect 113300 82500 114100 82700
rect 114500 82500 115700 82700
rect 113100 82300 114300 82500
rect 113100 81300 113500 82300
rect 113900 81300 114300 82300
rect 114500 81700 114900 82500
rect 115300 81700 115700 82500
rect 114500 81500 115700 81700
rect 115900 82500 117100 82700
rect 115900 81700 116300 82500
rect 116700 81700 117100 82500
rect 115900 81500 117100 81700
rect 117300 82500 117700 82900
rect 118700 82500 119100 82900
rect 119500 82500 119900 82900
rect 117300 82300 118300 82500
rect 117300 82100 118500 82300
rect 117300 81700 117700 82100
rect 118100 81700 118500 82100
rect 117300 81500 118500 81700
rect 118700 82100 119900 82500
rect 118700 81700 119100 82100
rect 119500 81700 119900 82100
rect 118700 81500 119900 81700
rect 120100 82700 121100 82900
rect 120100 82500 121300 82700
rect 120100 81700 120500 82500
rect 120900 81700 121300 82500
rect 120100 81500 121300 81700
rect 121500 82500 121900 82900
rect 122300 82700 122700 82900
rect 123300 82700 123700 82900
rect 122100 82500 122700 82700
rect 123100 82500 123900 82700
rect 121500 82100 122500 82500
rect 122900 82300 124100 82500
rect 121500 81700 121900 82100
rect 122300 81700 122700 82100
rect 121500 81500 122700 81700
rect 114500 81300 115500 81500
rect 115900 81300 116900 81500
rect 117300 81300 118300 81500
rect 118900 81300 119700 81500
rect 120100 81300 121100 81500
rect 121500 81300 122500 81500
rect 122900 81300 123300 82300
rect 123700 81300 124100 82300
rect 124900 81900 132300 83800
rect 124900 80300 133500 81900
rect 116500 77900 133500 80300
rect -29500 74900 -21500 75900
rect -15500 74900 -7500 75900
rect -30500 74500 -20100 74900
rect -30500 73900 -30100 74500
rect -31500 64900 -30100 73900
rect -30500 63900 -30100 64900
rect -20500 63900 -20100 74500
rect -30500 63500 -20100 63900
rect -19500 74700 -17500 74900
rect -19500 63700 -19300 74700
rect -17700 63700 -17500 74700
rect -19500 63500 -17500 63700
rect -16900 74500 -6500 74900
rect -16900 63900 -16500 74500
rect -6900 73900 -6500 74500
rect -6900 64900 -5500 73900
rect 10500 64900 19500 65900
rect 25500 64900 34500 65900
rect 38500 64900 47500 65900
rect 53500 64900 62500 65900
rect 66500 64900 75500 65900
rect 81500 64900 90500 65900
rect -6900 63900 -6500 64900
rect 9500 64500 20900 64900
rect 9500 63900 9900 64500
rect -16900 63500 -6500 63900
rect -30500 62700 -20100 62900
rect -30500 61100 -30300 62700
rect -20300 62500 -20100 62700
rect -19100 62500 -17900 63500
rect -16900 62700 -6500 62900
rect -16900 62500 -16700 62700
rect -20300 61300 -16700 62500
rect -20300 61100 -20100 61300
rect -30500 60900 -20100 61100
rect -19100 60300 -17900 61300
rect -16900 61100 -16700 61300
rect -6700 61100 -6500 62700
rect -16900 60900 -6500 61100
rect -30500 59900 -20100 60300
rect -30500 58900 -30100 59900
rect -31500 49900 -30100 58900
rect -30500 49300 -30100 49900
rect -20500 49300 -20100 59900
rect -30500 48900 -20100 49300
rect -19500 60100 -17500 60300
rect -19500 49100 -19300 60100
rect -17700 49100 -17500 60100
rect -19500 48900 -17500 49100
rect -16900 59900 -6500 60300
rect -16900 49300 -16500 59900
rect -6900 58900 -6500 59900
rect -6900 49900 -5500 58900
rect 8500 55900 9900 63900
rect 9500 54900 9900 55900
rect 20500 54900 20900 64500
rect 9500 54500 20900 54900
rect 21500 64700 23500 64900
rect 21500 54700 21700 64700
rect 23300 54700 23500 64700
rect 21500 54500 23500 54700
rect 24100 64500 35500 64900
rect 24100 54900 24500 64500
rect 35100 63900 35500 64500
rect 37500 64500 48900 64900
rect 37500 63900 37900 64500
rect 35100 55900 37900 63900
rect 35100 54900 35500 55900
rect 24100 54500 35500 54900
rect 37500 54900 37900 55900
rect 48500 54900 48900 64500
rect 37500 54500 48900 54900
rect 49500 64700 51500 64900
rect 49500 54700 49700 64700
rect 51300 54700 51500 64700
rect 49500 54500 51500 54700
rect 52100 64500 63500 64900
rect 52100 54900 52500 64500
rect 63100 63900 63500 64500
rect 65500 64500 76900 64900
rect 65500 63900 65900 64500
rect 63100 55900 65900 63900
rect 63100 54900 63500 55900
rect 52100 54500 63500 54900
rect 65500 54900 65900 55900
rect 76500 54900 76900 64500
rect 65500 54500 76900 54900
rect 77500 64700 79500 64900
rect 77500 54700 77700 64700
rect 79300 54700 79500 64700
rect 77500 54500 79500 54700
rect 80100 64500 91500 64900
rect 80100 54900 80500 64500
rect 91100 63900 91500 64500
rect 91100 55900 92500 63900
rect 116500 59900 121500 77900
rect 122500 59900 127500 77900
rect 128500 59900 133500 77900
rect 116500 59700 133500 59900
rect 91100 54900 91500 55900
rect 80100 54500 91500 54900
rect 9500 53700 20900 53900
rect 9500 52100 9700 53700
rect 20700 53500 20900 53700
rect 21900 53500 23100 54500
rect 24100 53700 35500 53900
rect 24100 53500 24300 53700
rect 20700 52300 24300 53500
rect 20700 52100 20900 52300
rect 9500 51900 20900 52100
rect 21900 51900 23100 52300
rect 24100 52100 24300 52300
rect 35300 52100 35500 53700
rect 24100 51900 35500 52100
rect 37500 53700 48900 53900
rect 37500 52100 37700 53700
rect 48700 53500 48900 53700
rect 49900 53500 51100 54500
rect 52100 53700 63500 53900
rect 52100 53500 52300 53700
rect 48700 52300 52300 53500
rect 48700 52100 48900 52300
rect 37500 51900 48900 52100
rect 49900 51300 51100 52300
rect 52100 52100 52300 52300
rect 63300 52100 63500 53700
rect 52100 51900 63500 52100
rect 65500 53700 76900 53900
rect 65500 52100 65700 53700
rect 76700 53500 76900 53700
rect 77900 53500 79100 54500
rect 116500 54100 116700 59700
rect 127300 54100 133500 59700
rect 116500 53900 133500 54100
rect 80100 53700 91500 53900
rect 80100 53500 80300 53700
rect 76700 52300 80300 53500
rect 76700 52100 76900 52300
rect 65500 51900 76900 52100
rect 77900 51300 79100 52300
rect 80100 52100 80300 52300
rect 91300 52100 91500 53700
rect 80100 51900 91500 52100
rect 116500 51900 121500 53900
rect 122500 51900 127500 53900
rect 128500 51900 133500 53900
rect 116500 51700 133500 51900
rect 37500 50900 48900 51300
rect 37500 49900 37900 50900
rect -6900 49300 -6500 49900
rect -16900 48900 -6500 49300
rect -29500 47900 -23500 48900
rect -15500 47900 -7500 48900
rect 36500 41900 37900 49900
rect 37500 41300 37900 41900
rect 48500 41300 48900 50900
rect 37500 40900 48900 41300
rect 49500 51100 51500 51300
rect 49500 41100 49700 51100
rect 51300 41100 51500 51100
rect 49500 40900 51500 41100
rect 52100 50900 63500 51300
rect 52100 41300 52500 50900
rect 63100 49900 63500 50900
rect 65500 50900 76900 51300
rect 65500 49900 65900 50900
rect 63100 41900 65900 49900
rect 63100 41300 63500 41900
rect 52100 40900 63500 41300
rect 65500 41300 65900 41900
rect 76500 41300 76900 50900
rect 65500 40900 76900 41300
rect 77500 51100 79500 51300
rect 77500 41100 77700 51100
rect 79300 41100 79500 51100
rect 77500 40900 79500 41100
rect 80100 50900 91500 51300
rect 80100 41300 80500 50900
rect 91100 49900 91500 50900
rect 91100 41900 92500 49900
rect 116500 46100 116700 51700
rect 127300 46100 133500 51700
rect 116500 45900 133500 46100
rect 91100 41300 91500 41900
rect 80100 40900 91500 41300
rect 38500 39900 47500 40900
rect 53500 39900 62500 40900
rect 66500 39900 75500 40900
rect 81500 39900 90500 40900
rect -22500 37500 -12500 37900
rect -22500 36900 -22100 37500
rect -23500 28900 -22100 36900
rect -22500 27900 -22100 28900
rect -12900 36900 -12500 37500
rect -12900 28900 -11500 36900
rect 129500 36700 141500 36900
rect -12900 27900 -12500 28900
rect -22500 27500 -12500 27900
rect 129500 27100 129700 36700
rect 135300 33900 136700 36700
rect 135300 29900 135500 33900
rect 136500 29900 136700 33900
rect 135300 27100 136700 29900
rect 141300 27100 141500 36700
rect 129500 26900 141500 27100
rect -22500 26700 -12500 26900
rect -22500 25100 -22300 26700
rect -12700 25100 -12500 26700
rect 133900 26100 134300 26300
rect 134900 26100 135900 26300
rect 136300 26100 137300 26300
rect 133700 25900 134500 26100
rect 134900 25900 136100 26100
rect -22500 24900 -12500 25100
rect 24600 21300 26100 25900
rect 133500 25700 134700 25900
rect 133500 24700 133900 25700
rect 134300 24700 134700 25700
rect 134900 25100 135300 25900
rect 135700 25100 136100 25900
rect 134900 24900 136100 25100
rect 136300 25900 137500 26100
rect 136300 25100 136700 25900
rect 137100 25100 137500 25900
rect 136300 24900 137500 25100
rect 137700 25900 138100 26300
rect 139100 25900 139500 26300
rect 139900 25900 140300 26300
rect 137700 25700 138700 25900
rect 137700 25500 138900 25700
rect 137700 25100 138100 25500
rect 138500 25100 138900 25500
rect 137700 24900 138900 25100
rect 139100 25500 140300 25900
rect 139100 25100 139500 25500
rect 139900 25100 140300 25500
rect 139100 24900 140300 25100
rect 134900 24700 135900 24900
rect 136300 24700 137300 24900
rect 137700 24700 138700 24900
rect 139300 24700 140100 24900
rect 24600 19900 26400 21300
rect 24500 13900 26300 19900
rect -14700 13850 -14300 13900
rect -14700 12650 -14650 13850
rect -14350 12650 -14300 13850
rect 16000 13700 20000 13900
rect -14700 12600 -14300 12650
rect 25900 8000 30500 8100
rect -21800 7700 -18800 7800
rect -21800 4700 -21700 7700
rect -18900 4700 -18800 7700
rect -21800 4600 -18800 4700
rect 1600 300 3600 700
rect 17500 -1300 17900 2400
rect 25900 -1800 26000 8000
rect 30400 -1800 30500 8000
rect 25900 -1900 30500 -1800
rect -22700 -11950 -18100 -11900
rect -23600 -12000 -18100 -11950
rect -23600 -16300 -23450 -12000
rect -22750 -12100 -18100 -12000
rect -22750 -16200 -22300 -12100
rect -18400 -16200 -18100 -12100
rect -22750 -16300 -18100 -16200
rect -23600 -16400 -18100 -16300
rect -20500 -21400 -19900 -21300
rect -20500 -21500 -20400 -21400
rect -22100 -21800 -20400 -21500
rect -20000 -21800 -19900 -21400
rect -22100 -21900 -19900 -21800
rect -25100 -28100 -22900 -27900
rect -25100 -29900 -24900 -28100
rect -23100 -29900 -22900 -28100
rect -25100 -30300 -22900 -29900
rect -27300 -31500 -22900 -30300
rect -27300 -31900 -25700 -31500
rect -24500 -31900 -22900 -31500
rect -27300 -33100 -22900 -31900
rect -27300 -36100 -25700 -33100
rect -22100 -34900 -21700 -21900
rect 23500 -28200 24000 -5600
rect 32800 -28200 34000 -20100
rect 23500 -28600 26000 -28200
rect 23500 -33200 24200 -28600
rect 25800 -33200 26000 -28600
rect 23500 -33600 26000 -33200
rect 30800 -28600 34000 -28200
rect 30800 -33200 31000 -28600
rect 32600 -32100 34000 -28600
rect 34900 -28400 36300 -28300
rect 34900 -28800 35000 -28400
rect 36200 -28800 36300 -28400
rect 34900 -28900 36300 -28800
rect 32600 -33200 32800 -32100
rect 30800 -33600 32800 -33200
rect 124700 -32600 125200 -32500
rect -22500 -35000 -21700 -34900
rect -22500 -35400 -22400 -35000
rect -22000 -35400 -21700 -35000
rect 26600 -34100 30200 -34000
rect 26600 -35300 26700 -34100
rect 30100 -35300 30200 -34100
rect 26600 -35400 30200 -35300
rect 124700 -35400 124800 -32600
rect 125100 -35400 125200 -32600
rect -22500 -35500 -21700 -35400
rect 124700 -35500 125200 -35400
rect 125600 -32700 134300 -32500
rect 125600 -35300 125800 -32700
rect 134100 -35300 134300 -32700
rect 125600 -35500 134300 -35300
rect -27300 -37700 -27100 -36100
rect -25900 -37700 -25700 -36100
rect 130800 -36500 132400 -35500
rect -27300 -37920 -25700 -37700
<< via4 >>
rect -19300 63700 -17700 74700
rect -30300 61100 -20300 62700
rect -16700 61100 -6700 62700
rect -19300 49100 -17700 60100
rect 21700 54700 23300 64700
rect 49700 54700 51300 64700
rect 77700 54700 79300 64700
rect 9700 52100 20700 53700
rect 24300 52100 35300 53700
rect 37700 52100 48700 53700
rect 52300 52100 63300 53700
rect 65700 52100 76700 53700
rect 116700 54100 127300 59700
rect 80300 52100 91300 53700
rect 49700 41100 51300 51100
rect 77700 41100 79300 51100
rect 116700 46100 127300 51700
rect 129700 27100 135300 36700
rect 136700 27100 136900 36700
rect 136900 27100 141300 36700
rect -22300 25100 -12700 26700
rect -21700 4700 -18900 7700
rect 26000 -1800 30400 8000
rect -20400 -21800 -20000 -21400
rect -24900 -29900 -23100 -28100
rect 24200 -33200 25800 -28600
rect 31000 -33200 32600 -28600
rect 26700 -35300 30100 -34100
rect 124800 -35400 125100 -32600
<< mimcap2 >>
rect -30300 74500 -20300 74700
rect -30300 63900 -30100 74500
rect -20500 63900 -20300 74500
rect -30300 63700 -20300 63900
rect -16700 74500 -6700 74700
rect -16700 63900 -16500 74500
rect -6900 63900 -6700 74500
rect -16700 63700 -6700 63900
rect 9700 64500 20700 64700
rect -30300 59900 -20300 60100
rect -30300 49300 -30100 59900
rect -20500 49300 -20300 59900
rect -30300 49100 -20300 49300
rect -16700 59900 -6700 60100
rect -16700 49300 -16500 59900
rect -6900 49300 -6700 59900
rect 9700 54900 9900 64500
rect 20500 54900 20700 64500
rect 9700 54700 20700 54900
rect 24300 64500 35300 64700
rect 24300 54900 24500 64500
rect 35100 54900 35300 64500
rect 24300 54700 35300 54900
rect 37700 64500 48700 64700
rect 37700 54900 37900 64500
rect 48500 54900 48700 64500
rect 37700 54700 48700 54900
rect 52300 64500 63300 64700
rect 52300 54900 52500 64500
rect 63100 54900 63300 64500
rect 52300 54700 63300 54900
rect 65700 64500 76700 64700
rect 65700 54900 65900 64500
rect 76500 54900 76700 64500
rect 65700 54700 76700 54900
rect 80300 64500 91300 64700
rect 80300 54900 80500 64500
rect 91100 54900 91300 64500
rect 80300 54700 91300 54900
rect -16700 49100 -6700 49300
rect 37700 50900 48700 51100
rect 37700 41300 37900 50900
rect 48500 41300 48700 50900
rect 37700 41100 48700 41300
rect 52300 50900 63300 51100
rect 52300 41300 52500 50900
rect 63100 41300 63300 50900
rect 52300 41100 63300 41300
rect 65700 50900 76700 51100
rect 65700 41300 65900 50900
rect 76500 41300 76700 50900
rect 65700 41100 76700 41300
rect 80300 50900 91300 51100
rect 80300 41300 80500 50900
rect 91100 41300 91300 50900
rect 80300 41100 91300 41300
rect -22300 37500 -12700 37700
rect -22300 27900 -22100 37500
rect -12900 27900 -12700 37500
rect -22300 27700 -12700 27900
rect -22400 -12100 -18300 -12000
rect -22400 -16200 -22300 -12100
rect -18400 -16200 -18300 -12100
rect -22400 -16300 -18300 -16200
rect 125700 -32700 134200 -32600
rect 125700 -35300 125800 -32700
rect 134100 -35300 134200 -32700
rect 125700 -35400 134200 -35300
<< mimcap2contact >>
rect -30100 63900 -20500 74500
rect -16500 63900 -6900 74500
rect -30100 49300 -20500 59900
rect -16500 49300 -6900 59900
rect 9900 54900 20500 64500
rect 24500 54900 35100 64500
rect 37900 54900 48500 64500
rect 52500 54900 63100 64500
rect 65900 54900 76500 64500
rect 80500 54900 91100 64500
rect 37900 41300 48500 50900
rect 52500 41300 63100 50900
rect 65900 41300 76500 50900
rect 80500 41300 91100 50900
rect -22100 27900 -12900 37500
rect -22300 -16200 -18400 -12100
rect 125800 -35300 134100 -32700
<< metal5 >>
rect -30500 80300 112500 81900
rect -30500 76900 142500 80300
rect -30500 74900 -26500 76900
rect -20500 74900 -16500 76900
rect -10500 75900 -2500 76900
rect 10500 75900 14500 76900
rect 26500 75900 30500 76900
rect 42500 75900 46500 76900
rect 58500 75900 62500 76900
rect 74500 75900 78500 76900
rect 90500 75900 94500 76900
rect 106500 75900 110500 76900
rect 122500 75900 126500 76900
rect 129500 75900 135500 76900
rect -10500 74900 135500 75900
rect -30500 74700 135500 74900
rect -30500 74500 -19300 74700
rect -30500 63900 -30100 74500
rect -20500 63900 -19300 74500
rect -30500 63700 -19300 63900
rect -17700 74500 135500 74700
rect -17700 63900 -16500 74500
rect -6900 70900 135500 74500
rect -6900 63900 -6500 70900
rect 10500 66900 84500 68900
rect 10500 64900 14500 66900
rect 24500 64900 28500 66900
rect 38500 64900 42500 66900
rect 52500 64900 56500 66900
rect 66500 64900 70500 66900
rect 80500 64900 84500 66900
rect 129500 64900 135500 70900
rect 136500 64900 142500 76900
rect -17700 63700 -6500 63900
rect -30500 62700 -6500 63700
rect -30500 61100 -30300 62700
rect -20300 61100 -16700 62700
rect -6700 61100 -6500 62700
rect -30500 60100 -6500 61100
rect -30500 59900 -19300 60100
rect -30500 49300 -30100 59900
rect -20500 49300 -19300 59900
rect -30500 49100 -19300 49300
rect -17700 59900 -6500 60100
rect -17700 49300 -16500 59900
rect -6900 49300 -6500 59900
rect 9500 64700 98500 64900
rect 9500 64500 21700 64700
rect 9500 54900 9900 64500
rect 20500 54900 21700 64500
rect 9500 54700 21700 54900
rect 23300 64500 49700 64700
rect 23300 54900 24500 64500
rect 35100 60900 37900 64500
rect 35100 55900 35500 60900
rect 37500 55900 37900 60900
rect 35100 54900 37900 55900
rect 48500 54900 49700 64500
rect 23300 54700 49700 54900
rect 51300 64500 77700 64700
rect 51300 54900 52500 64500
rect 63100 60900 65900 64500
rect 63100 55900 63500 60900
rect 65500 55900 65900 60900
rect 63100 54900 65900 55900
rect 76500 54900 77700 64500
rect 51300 54700 77700 54900
rect 79300 64500 98500 64700
rect 79300 54900 80500 64500
rect 91100 60900 98500 64500
rect 91100 54900 91500 60900
rect 92500 59900 98500 60900
rect 129500 60900 142500 64900
rect 92500 59700 127500 59900
rect 92500 54900 116700 59700
rect 79300 54700 116700 54900
rect 9500 54100 116700 54700
rect 127300 54100 127500 59700
rect 9500 53900 127500 54100
rect 9500 53700 98500 53900
rect 9500 52100 9700 53700
rect 20700 52100 24300 53700
rect 35300 52100 37700 53700
rect 48700 52100 52300 53700
rect 63300 52100 65700 53700
rect 76700 52100 80300 53700
rect 91300 52100 98500 53700
rect 9500 51900 98500 52100
rect 105500 51900 110500 53900
rect 116500 51900 121500 53900
rect 122500 51900 127500 53900
rect -17700 49100 -6500 49300
rect -30500 48900 -6500 49100
rect -22500 46900 -15500 48900
rect -22500 39900 -19500 46900
rect -18500 39900 -15500 46900
rect -22500 37900 -15500 39900
rect 28500 45900 31500 51900
rect 32500 45900 35500 51900
rect 28500 43900 35500 45900
rect 28500 37900 31500 43900
rect 32500 38900 35500 43900
rect 37500 51700 127500 51900
rect 37500 51100 116700 51700
rect 37500 50900 49700 51100
rect 37500 41300 37900 50900
rect 48500 41300 49700 50900
rect 37500 41100 49700 41300
rect 51300 50900 77700 51100
rect 51300 41300 52500 50900
rect 63100 49900 65900 50900
rect 63100 44900 63500 49900
rect 65500 44900 65900 49900
rect 63100 41300 65900 44900
rect 76500 41300 77700 50900
rect 51300 41100 77700 41300
rect 79300 50900 116700 51100
rect 79300 41300 80500 50900
rect 91100 45900 91500 50900
rect 92500 46100 116700 50900
rect 127300 46100 127500 51700
rect 92500 45900 127500 46100
rect 129500 48900 135500 60900
rect 136500 48900 142500 60900
rect 91100 41300 98500 45900
rect 79300 41100 98500 41300
rect 37500 40900 98500 41100
rect 129500 44900 142500 48900
rect 38500 38900 46500 40900
rect 59500 38900 63500 40900
rect 72500 38900 76500 40900
rect 87500 38900 91500 40900
rect 32500 37900 91500 38900
rect -22500 37500 -12500 37900
rect -22500 27900 -22100 37500
rect -12900 28900 -12500 37500
rect 28500 36900 91500 37900
rect 129500 36900 135500 44900
rect 136500 36900 142500 44900
rect 28500 35900 47500 36900
rect 129500 36700 141500 36900
rect 28500 29900 31500 35900
rect 32500 29900 39500 35900
rect 40500 34900 46500 35900
rect 40500 33900 45500 34900
rect 40500 29900 44500 33900
rect -12900 27900 -10500 28900
rect 28500 27900 44500 29900
rect -22500 26700 -10500 27900
rect 33500 26900 39500 27900
rect -22500 25100 -22300 26700
rect -12700 25100 -10500 26700
rect -22500 24900 -10500 25100
rect -18500 15900 -16500 24900
rect -15500 15900 -13500 24900
rect -15500 7900 -13500 9900
rect -12500 7900 -10500 24900
rect 34500 21900 39500 26900
rect 40500 21900 44500 27900
rect 129500 27100 129700 36700
rect 135300 33900 136700 36700
rect 135300 29900 135500 33900
rect 136500 29900 136700 33900
rect 135300 27100 136700 29900
rect 141300 27100 141500 36700
rect 129500 26900 141500 27100
rect -19500 7800 -10500 7900
rect -21800 7700 -10500 7800
rect -21800 4700 -21700 7700
rect -18900 5900 -10500 7700
rect 25900 8000 30500 8100
rect -18900 4700 -18800 5900
rect -21800 4600 -18800 4700
rect -21800 800 -19800 4600
rect -13100 1500 -10700 1900
rect -25100 -2300 -23100 -2200
rect -21800 -2300 -18800 800
rect -13100 -300 -12700 1500
rect -25100 -4100 -18800 -2300
rect -25100 -7100 -23100 -4100
rect -21800 -7100 -18800 -4100
rect -25100 -8900 -18800 -7100
rect -25100 -11900 -23100 -8900
rect -21800 -11900 -18800 -8900
rect -17500 -1100 -12700 -300
rect -25100 -12100 -18100 -11900
rect -25100 -16200 -22300 -12100
rect -18400 -16200 -18100 -12100
rect -25100 -16400 -18100 -16200
rect -25100 -28100 -22900 -16400
rect -17500 -19500 -16700 -1100
rect 25900 -1600 26000 8000
rect 25800 -1800 26000 -1600
rect 30400 -1600 30500 8000
rect 30400 -1800 30600 -1600
rect 25800 -2000 30600 -1800
rect 26600 -4200 30200 -2000
rect -20300 -19900 -16700 -19500
rect -20300 -21300 -19900 -19900
rect -20500 -21400 -19900 -21300
rect -20500 -21800 -20400 -21400
rect -20000 -21800 -19900 -21400
rect -20500 -21900 -19900 -21800
rect -25100 -29900 -24900 -28100
rect -23100 -29900 -22900 -28100
rect -25100 -30100 -22900 -29900
rect 24000 -28600 26000 -28200
rect 24000 -33200 24200 -28600
rect 25800 -33200 26000 -28600
rect 24000 -33600 26000 -33200
rect 26600 -34100 30200 -28200
rect 30800 -28600 32800 -28200
rect 30800 -33200 31000 -28600
rect 32600 -33200 32800 -28600
rect 130500 -30100 132500 26900
rect 130500 -31600 136300 -30100
rect 30800 -33600 32800 -33200
rect 124700 -32600 134300 -32500
rect 26600 -35300 26700 -34100
rect 30100 -35300 30200 -34100
rect 26600 -35400 30200 -35300
rect 124700 -35400 124800 -32600
rect 125100 -32700 134300 -32600
rect 125100 -35300 125800 -32700
rect 134100 -35300 134300 -32700
rect 125100 -35400 134300 -35300
rect 124700 -35500 134300 -35400
rect 134900 -36200 136300 -31600
rect 132500 -38000 136300 -36200
use CPW_chunk_1_W20  CPW_chunk_1_W20_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660959839
transform 1 0 26000 0 1 -11600
box -2000 -600 6800 7400
use CPW_chunk_1_W20  CPW_chunk_1_W20_1
timestamp 1660959839
transform 1 0 26000 0 1 -19600
box -2000 -600 6800 7400
use CPW_chunk_1_W20  CPW_chunk_1_W20_2
timestamp 1660959839
transform 1 0 26000 0 1 -27600
box -2000 -600 6800 7400
use ESD_diode_DNW  ESD_diode_DNW_0
timestamp 1662581340
transform 1 0 -25090 0 -1 -34100
box -210 1600 5580 3948
use OSC_5GHz_1  OSC_5GHz_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/OSC
timestamp 1662654558
transform -1 0 -3300 0 1 5900
box 10000 -21000 68022 34000
use PA_complete  PA_complete_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/PA
timestamp 1662263286
transform 1 0 14099 0 1 2080
box -18800 -26000 70600 43800
use VGA_complete_1  VGA_complete_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/PA
timestamp 1662654558
transform 1 0 500 0 1 -15300
box -21500 -7100 11600 21400
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660275339
transform 1 0 -24600 0 1 4500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_1
timestamp 1660275339
transform 1 0 -24100 0 1 4500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_2
timestamp 1660275339
transform 1 0 -23600 0 1 4500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_3
timestamp 1660275339
transform 1 0 -24600 0 1 4000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_4
timestamp 1660275339
transform 1 0 -24100 0 1 4000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_5
timestamp 1660275339
transform 1 0 -23600 0 1 4000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_6
timestamp 1660275339
transform 1 0 -24600 0 1 3500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_7
timestamp 1660275339
transform 1 0 -24100 0 1 3500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_8
timestamp 1660275339
transform 1 0 -23600 0 1 3500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_9
timestamp 1660275339
transform 1 0 -24600 0 1 3000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_10
timestamp 1660275339
transform 1 0 -24100 0 1 3000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_11
timestamp 1660275339
transform 1 0 -23600 0 1 3000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_12
timestamp 1660275339
transform 1 0 -24600 0 1 2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_13
timestamp 1660275339
transform 1 0 -24100 0 1 2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_14
timestamp 1660275339
transform 1 0 -23600 0 1 2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_15
timestamp 1660275339
transform 1 0 -24600 0 1 2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_16
timestamp 1660275339
transform 1 0 -24100 0 1 2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_17
timestamp 1660275339
transform 1 0 -23600 0 1 2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_18
timestamp 1660275339
transform 1 0 -24600 0 1 1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_19
timestamp 1660275339
transform 1 0 -24100 0 1 1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_20
timestamp 1660275339
transform 1 0 -23600 0 1 1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_21
timestamp 1660275339
transform 1 0 -24600 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_22
timestamp 1660275339
transform 1 0 -24100 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_23
timestamp 1660275339
transform 1 0 -23600 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_24
timestamp 1660275339
transform 1 0 -24600 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_25
timestamp 1660275339
transform 1 0 -24100 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_26
timestamp 1660275339
transform 1 0 -23600 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_27
timestamp 1660275339
transform 1 0 -24600 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_28
timestamp 1660275339
transform 1 0 -24100 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_29
timestamp 1660275339
transform 1 0 -23600 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_30
timestamp 1660275339
transform 1 0 -12100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_31
timestamp 1660275339
transform 1 0 -10600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_32
timestamp 1660275339
transform 1 0 -10100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_33
timestamp 1660275339
transform 1 0 -10600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_34
timestamp 1660275339
transform 1 0 -10100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_35
timestamp 1660275339
transform 1 0 -11600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_36
timestamp 1660275339
transform 1 0 -11100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_37
timestamp 1660275339
transform 1 0 -11600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_38
timestamp 1660275339
transform 1 0 -15600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_39
timestamp 1660275339
transform 1 0 -15100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_40
timestamp 1660275339
transform 1 0 -15600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_41
timestamp 1660275339
transform 1 0 -15100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_42
timestamp 1660275339
transform 1 0 -14600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_43
timestamp 1660275339
transform 1 0 -14600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_44
timestamp 1660275339
transform 1 0 -14100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_45
timestamp 1660275339
transform 1 0 -14100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_46
timestamp 1660275339
transform 1 0 -11100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_47
timestamp 1660275339
transform 1 0 -12600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_48
timestamp 1660275339
transform 1 0 -13100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_49
timestamp 1660275339
transform 1 0 -13600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_50
timestamp 1660275339
transform 1 0 -8600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_51
timestamp 1660275339
transform 1 0 -8100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_52
timestamp 1660275339
transform 1 0 -9600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_53
timestamp 1660275339
transform 1 0 -9100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_54
timestamp 1660275339
transform 1 0 -8600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_55
timestamp 1660275339
transform 1 0 -13600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_56
timestamp 1660275339
transform 1 0 -8100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_57
timestamp 1660275339
transform 1 0 -9600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_58
timestamp 1660275339
transform 1 0 -9100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_59
timestamp 1660275339
transform 1 0 -6100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_60
timestamp 1660275339
transform 1 0 -6600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_61
timestamp 1660275339
transform 1 0 -7600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_62
timestamp 1660275339
transform 1 0 -7100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_63
timestamp 1660275339
transform 1 0 -6100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_64
timestamp 1660275339
transform 1 0 -6600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_65
timestamp 1660275339
transform 1 0 -7600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_66
timestamp 1660275339
transform 1 0 -7100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_67
timestamp 1660275339
transform 1 0 -8600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_68
timestamp 1660275339
transform 1 0 -8100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_69
timestamp 1660275339
transform 1 0 -12100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_70
timestamp 1660275339
transform 1 0 -8600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_71
timestamp 1660275339
transform 1 0 -12600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_72
timestamp 1660275339
transform 1 0 -13100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_73
timestamp 1660275339
transform 1 0 -8100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_74
timestamp 1660275339
transform 1 0 -9100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_75
timestamp 1660275339
transform 1 0 -9600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_76
timestamp 1660275339
transform 1 0 -9600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_77
timestamp 1660275339
transform 1 0 -9100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_78
timestamp 1660275339
transform 1 0 -6100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_79
timestamp 1660275339
transform 1 0 -6100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_80
timestamp 1660275339
transform 1 0 -6600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_81
timestamp 1660275339
transform 1 0 -6600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_82
timestamp 1660275339
transform 1 0 -7100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_83
timestamp 1660275339
transform 1 0 -7600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_84
timestamp 1660275339
transform 1 0 -7600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_85
timestamp 1660275339
transform 1 0 -7100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_86
timestamp 1660275339
transform 1 0 -10100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_87
timestamp 1660275339
transform 1 0 -10100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_88
timestamp 1660275339
transform 1 0 -10600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_89
timestamp 1660275339
transform 1 0 -10600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_90
timestamp 1660275339
transform 1 0 -11100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_91
timestamp 1660275339
transform 1 0 -11600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_92
timestamp 1660275339
transform 1 0 -11600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_93
timestamp 1660275339
transform 1 0 -11100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_94
timestamp 1660275339
transform 1 0 -10100 0 1 13500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_95
timestamp 1660275339
transform 1 0 -10100 0 1 13000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_96
timestamp 1660275339
transform 1 0 -10600 0 1 13500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_97
timestamp 1660275339
transform 1 0 -10600 0 1 13000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_98
timestamp 1660275339
transform 1 0 -11100 0 1 13500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_99
timestamp 1660275339
transform 1 0 -11600 0 1 13500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_100
timestamp 1660275339
transform 1 0 -11600 0 1 13000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_101
timestamp 1660275339
transform 1 0 -11100 0 1 13000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_102
timestamp 1660275339
transform 1 0 -10100 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_103
timestamp 1660275339
transform 1 0 -10100 0 1 14000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_104
timestamp 1660275339
transform 1 0 -10600 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_105
timestamp 1660275339
transform 1 0 -10600 0 1 14000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_106
timestamp 1660275339
transform 1 0 -11100 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_107
timestamp 1660275339
transform 1 0 -11600 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_108
timestamp 1660275339
transform 1 0 -11600 0 1 14000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_109
timestamp 1660275339
transform 1 0 -11100 0 1 14000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_110
timestamp 1660275339
transform 1 0 -11600 0 1 15000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_111
timestamp 1660275339
transform 1 0 -12100 0 1 15000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_112
timestamp 1660275339
transform 1 0 -12100 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_113
timestamp 1660275339
transform 1 0 -12600 0 1 15000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_114
timestamp 1660275339
transform 1 0 -13100 0 1 15000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_115
timestamp 1660275339
transform 1 0 -13100 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_116
timestamp 1660275339
transform 1 0 -12600 0 1 14500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_117
timestamp 1660275339
transform 1 0 -5600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_118
timestamp 1660275339
transform 1 0 -5100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_119
timestamp 1660275339
transform 1 0 -4600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_120
timestamp 1660275339
transform 1 0 -4100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_121
timestamp 1660275339
transform 1 0 -3600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_122
timestamp 1660275339
transform 1 0 -3100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_123
timestamp 1660275339
transform 1 0 -5600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_124
timestamp 1660275339
transform 1 0 -5100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_125
timestamp 1660275339
transform 1 0 -4600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_126
timestamp 1660275339
transform 1 0 -4100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_127
timestamp 1660275339
transform 1 0 -3600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_128
timestamp 1660275339
transform 1 0 -3100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_129
timestamp 1660275339
transform 1 0 -2600 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_130
timestamp 1660275339
transform 1 0 -2100 0 1 12000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_131
timestamp 1660275339
transform 1 0 -2600 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_132
timestamp 1660275339
transform 1 0 -2100 0 1 12500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_133
timestamp 1660275339
transform 1 0 -2600 0 1 11500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_134
timestamp 1660275339
transform 1 0 -2100 0 1 11500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_135
timestamp 1660275339
transform 1 0 -2600 0 1 11000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_136
timestamp 1660275339
transform 1 0 -2100 0 1 11000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_137
timestamp 1660275339
transform 1 0 -2600 0 1 10500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_138
timestamp 1660275339
transform 1 0 -2100 0 1 10500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_139
timestamp 1660275339
transform 1 0 -2600 0 1 10000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_140
timestamp 1660275339
transform 1 0 -2100 0 1 10000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_141
timestamp 1660275339
transform 1 0 -2600 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_142
timestamp 1660275339
transform 1 0 -2100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_143
timestamp 1660275339
transform 1 0 -2600 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_144
timestamp 1660275339
transform 1 0 -2100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_145
timestamp 1660275339
transform 1 0 -2600 0 1 8500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_146
timestamp 1660275339
transform 1 0 -2100 0 1 8500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_147
timestamp 1660275339
transform 1 0 -2600 0 1 8000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_148
timestamp 1660275339
transform 1 0 -2100 0 1 8000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_149
timestamp 1660275339
transform 1 0 -2600 0 1 7500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_150
timestamp 1660275339
transform 1 0 -2100 0 1 7500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_151
timestamp 1660275339
transform 1 0 -2600 0 1 7000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_152
timestamp 1660275339
transform 1 0 -2100 0 1 7000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_153
timestamp 1660275339
transform 1 0 -3100 0 1 11500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_154
timestamp 1660275339
transform 1 0 -3100 0 1 11000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_155
timestamp 1660275339
transform 1 0 -3100 0 1 10500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_156
timestamp 1660275339
transform 1 0 -24100 0 1 5000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_157
timestamp 1660275339
transform 1 0 -24600 0 1 5000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_158
timestamp 1660275339
transform 1 0 -24600 0 1 5500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_159
timestamp 1660275339
transform 1 0 -24100 0 1 5500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_160
timestamp 1660275339
transform 1 0 -3100 0 1 10000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_161
timestamp 1660275339
transform 1 0 -23600 0 1 5000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_162
timestamp 1660275339
transform 1 0 -23600 0 1 5500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_163
timestamp 1660275339
transform 1 0 -3100 0 1 9500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_164
timestamp 1660275339
transform 1 0 -3100 0 1 9000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_165
timestamp 1660275339
transform 1 0 -3100 0 1 8500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_166
timestamp 1660275339
transform 1 0 -3100 0 1 8000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_167
timestamp 1660275339
transform 1 0 -3100 0 1 7000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_168
timestamp 1660275339
transform 1 0 -3100 0 1 7500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_169
timestamp 1660275339
transform 1 0 13400 0 1 -1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_170
timestamp 1660275339
transform 1 0 13400 0 1 -1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_171
timestamp 1660275339
transform 1 0 13400 0 1 -2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_172
timestamp 1660275339
transform 1 0 13400 0 1 -2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_173
timestamp 1660275339
transform 1 0 13400 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_174
timestamp 1660275339
transform 1 0 13400 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_175
timestamp 1660275339
transform 1 0 13400 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_176
timestamp 1660275339
transform 1 0 13400 0 1 -500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_177
timestamp 1660275339
transform 1 0 13900 0 1 500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_178
timestamp 1660275339
transform 1 0 13900 0 1 1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_179
timestamp 1660275339
transform 1 0 13900 0 1 0
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_180
timestamp 1660275339
transform 1 0 13900 0 1 -500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_181
timestamp 1660275339
transform 1 0 13900 0 1 -1500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_182
timestamp 1660275339
transform 1 0 13900 0 1 -1000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_183
timestamp 1660275339
transform 1 0 13900 0 1 -2000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_184
timestamp 1660275339
transform 1 0 13900 0 1 -2500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_185
timestamp 1660275339
transform 1 0 15400 0 1 -3500
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_186
timestamp 1660275339
transform 1 0 15400 0 1 -3000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_187
timestamp 1660275339
transform 1 0 15400 0 1 -4000
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_188
timestamp 1660275339
transform 1 0 15400 0 1 -4500
box 100 -1100 600 -600
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660789662
transform 1 0 22500 0 1 -11900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_1
timestamp 1660789662
transform 1 0 14500 0 1 -12400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_2
timestamp 1660789662
transform 1 0 15500 0 1 -12400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_3
timestamp 1660789662
transform 1 0 16500 0 1 -12400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_4
timestamp 1660789662
transform 1 0 16500 0 1 -13400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_5
timestamp 1660789662
transform 1 0 16500 0 1 -14400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_6
timestamp 1660789662
transform 1 0 16500 0 1 -15400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_7
timestamp 1660789662
transform 1 0 16500 0 1 -16400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_8
timestamp 1660789662
transform 1 0 16500 0 1 -17400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_9
timestamp 1660789662
transform 1 0 16500 0 1 -18400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_10
timestamp 1660789662
transform 1 0 16500 0 1 -19400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_11
timestamp 1660789662
transform 1 0 16500 0 1 -20400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_12
timestamp 1660789662
transform 1 0 17500 0 1 -20400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_13
timestamp 1660789662
transform 1 0 18500 0 1 -20400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_14
timestamp 1660789662
transform 1 0 18500 0 1 -21400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_15
timestamp 1660789662
transform 1 0 18500 0 1 -22400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_16
timestamp 1660789662
transform 1 0 18500 0 1 -23400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_17
timestamp 1660789662
transform 1 0 18500 0 1 -24400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_18
timestamp 1660789662
transform 1 0 18500 0 1 -25400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_19
timestamp 1660789662
transform 1 0 18500 0 1 -26400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_20
timestamp 1660789662
transform 1 0 18500 0 1 -27400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_21
timestamp 1660789662
transform 1 0 18500 0 1 -28400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_22
timestamp 1660789662
transform 1 0 19500 0 1 -28400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_23
timestamp 1660789662
transform 1 0 20500 0 1 -28400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_24
timestamp 1660789662
transform 1 0 21500 0 1 -28400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_25
timestamp 1660789662
transform 1 0 34500 0 1 -28400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_26
timestamp 1660789662
transform 1 0 35500 0 1 -28400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_0
timestamp 1660789662
transform 1 0 22500 0 1 -8900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_1
timestamp 1660789662
transform 1 0 22500 0 1 -9900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_2
timestamp 1660789662
transform 1 0 22500 0 1 -10900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_4
timestamp 1660789662
transform 1 0 22500 0 1 -14900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_5
timestamp 1660789662
transform 1 0 22500 0 1 -13900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_6
timestamp 1660789662
transform 1 0 22500 0 1 -12900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_7
timestamp 1660789662
transform 1 0 22500 0 1 -17900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_8
timestamp 1660789662
transform 1 0 22500 0 1 -16900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_9
timestamp 1660789662
transform 1 0 22500 0 1 -15900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_10
timestamp 1660789662
transform 1 0 22500 0 1 -20900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_11
timestamp 1660789662
transform 1 0 22500 0 1 -19900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_12
timestamp 1660789662
transform 1 0 22500 0 1 -18900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_13
timestamp 1660789662
transform 1 0 22500 0 1 -23900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_14
timestamp 1660789662
transform 1 0 22500 0 1 -22900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_15
timestamp 1660789662
transform 1 0 22500 0 1 -21900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_16
timestamp 1660789662
transform 1 0 22500 0 1 -26900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_17
timestamp 1660789662
transform 1 0 22500 0 1 -25900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_18
timestamp 1660789662
transform 1 0 22500 0 1 -24900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_19
timestamp 1660789662
transform 1 0 22500 0 1 -29900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_20
timestamp 1660789662
transform 1 0 22500 0 1 -28900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_22
timestamp 1660789662
transform 1 0 -17000 0 1 -2400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_23
timestamp 1660789662
transform 1 0 22500 0 1 -31900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_24
timestamp 1660789662
transform 1 0 22500 0 1 -30900
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_25
timestamp 1660789662
transform 1 0 -16000 0 1 -2400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_26
timestamp 1660789662
transform 1 0 -16500 0 1 -18400
box 0 -1700 1000 -700
use hash_m1m2m3_W5L5  hash_m1m2m3_W5L5_27
timestamp 1660789662
transform 1 0 -16500 0 1 -17400
box 0 -1700 1000 -700
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660789662
transform 1 0 -11500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_1
timestamp 1660789662
transform 1 0 -15500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_2
timestamp 1660789662
transform 1 0 -13500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_3
timestamp 1660789662
transform 1 0 -9500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_4
timestamp 1660789662
transform 1 0 -7500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_5
timestamp 1660789662
transform 1 0 -7500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_6
timestamp 1660789662
transform 1 0 -9500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_7
timestamp 1660789662
transform 1 0 500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_8
timestamp 1660789662
transform 1 0 500 0 1 9600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_9
timestamp 1660789662
transform 1 0 -3500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_10
timestamp 1660789662
transform 1 0 -5500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_11
timestamp 1660789662
transform 1 0 500 0 1 11600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_12
timestamp 1660789662
transform 1 0 -1500 0 1 13600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_13
timestamp 1660789662
transform 1 0 2500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_14
timestamp 1660789662
transform 1 0 -1500 0 1 11600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_15
timestamp 1660789662
transform 1 0 2500 0 1 9600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_16
timestamp 1660789662
transform 1 0 -1500 0 1 9600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_17
timestamp 1660789662
transform 1 0 2500 0 1 11600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_18
timestamp 1660789662
transform 1 0 -1500 0 1 7600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_19
timestamp 1660789662
transform 1 0 16000 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_20
timestamp 1660789662
transform 1 0 -3500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_21
timestamp 1660789662
transform 1 0 -5500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_22
timestamp 1660789662
transform 1 0 -7500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_23
timestamp 1660789662
transform 1 0 -9500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_24
timestamp 1660789662
transform 1 0 -11500 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_25
timestamp 1660789662
transform 1 0 -11500 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_26
timestamp 1660789662
transform 1 0 -9500 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_27
timestamp 1660789662
transform 1 0 -7500 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_28
timestamp 1660789662
transform 1 0 -5500 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_29
timestamp 1660789662
transform 1 0 18000 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_30
timestamp 1660789662
transform 1 0 -11500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_31
timestamp 1660789662
transform 1 0 -9500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_32
timestamp 1660789662
transform 1 0 -7500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_33
timestamp 1660789662
transform 1 0 20000 0 1 15600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_34
timestamp 1660789662
transform 1 0 26500 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_35
timestamp 1660789662
transform 1 0 9500 0 1 100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_36
timestamp 1660789662
transform 1 0 11500 0 1 100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_37
timestamp 1660789662
transform 1 0 11500 0 1 -1900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_38
timestamp 1660789662
transform 1 0 19500 0 1 -3900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_39
timestamp 1660789662
transform 1 0 15500 0 1 100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_40
timestamp 1660789662
transform 1 0 15500 0 1 -1900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_41
timestamp 1660789662
transform 1 0 15500 0 1 2100
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_42
timestamp 1660789662
transform 1 0 21500 0 1 -3900
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_43
timestamp 1660789662
transform 1 0 28500 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_44
timestamp 1660789662
transform 1 0 24000 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_45
timestamp 1660789662
transform 1 0 22000 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_46
timestamp 1660789662
transform 1 0 20000 0 1 17600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_47
timestamp 1660789662
transform 1 0 30500 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_48
timestamp 1660789662
transform 1 0 32500 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_49
timestamp 1660789662
transform 1 0 26500 0 1 29600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_50
timestamp 1660789662
transform 1 0 26500 0 1 31600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_51
timestamp 1660789662
transform 1 0 26500 0 1 33600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_52
timestamp 1660789662
transform 1 0 26500 0 1 35600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_53
timestamp 1660789662
transform 1 0 26500 0 1 37600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_54
timestamp 1660789662
transform 1 0 26500 0 1 39600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_55
timestamp 1660789662
transform 1 0 34500 0 1 -24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_56
timestamp 1660789662
transform 1 0 34500 0 1 -26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_57
timestamp 1660789662
transform 1 0 34500 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_59
timestamp 1660789662
transform 1 0 26500 0 1 41600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_60
timestamp 1660789662
transform 1 0 26500 0 1 43600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_61
timestamp 1660789662
transform 1 0 34000 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_62
timestamp 1660789662
transform 1 0 34000 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_63
timestamp 1660789662
transform 1 0 34000 0 1 -24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_64
timestamp 1660789662
transform 1 0 34000 0 1 -26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_66
timestamp 1660789662
transform 1 0 34000 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_67
timestamp 1660789662
transform 1 0 34500 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_68
timestamp 1660789662
transform 1 0 -15500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_69
timestamp 1660789662
transform 1 0 -13500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_70
timestamp 1660789662
transform 1 0 -19500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_71
timestamp 1660789662
transform 1 0 -17500 0 1 19600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_72
timestamp 1660789662
transform 1 0 22500 0 1 47600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_73
timestamp 1660789662
transform 1 0 -3500 0 1 47600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_74
timestamp 1660789662
transform 1 0 -7500 0 1 43600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_75
timestamp 1660789662
transform 1 0 22500 0 1 45600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_76
timestamp 1660789662
transform 1 0 24500 0 1 43600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_77
timestamp 1660789662
transform 1 0 20500 0 1 47600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_78
timestamp 1660789662
transform 1 0 36500 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_79
timestamp 1660789662
transform 1 0 38500 0 1 27600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_80
timestamp 1660789662
transform 1 0 -17500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_81
timestamp 1660789662
transform 1 0 -17500 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_82
timestamp 1660789662
transform 1 0 -19500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_83
timestamp 1660789662
transform 1 0 -21500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_84
timestamp 1660789662
transform 1 0 -21500 0 1 -24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_85
timestamp 1660789662
transform 1 0 -21500 0 1 -26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_86
timestamp 1660789662
transform 1 0 -21500 0 1 -28400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_87
timestamp 1660789662
transform 1 0 -21500 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_88
timestamp 1660789662
transform 1 0 36500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_89
timestamp 1660789662
transform 1 0 38500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_90
timestamp 1660789662
transform 1 0 40500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_91
timestamp 1660789662
transform 1 0 42500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_92
timestamp 1660789662
transform 1 0 44500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_93
timestamp 1660789662
transform 1 0 46500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_94
timestamp 1660789662
transform 1 0 58500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_95
timestamp 1660789662
transform 1 0 56500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_96
timestamp 1660789662
transform 1 0 54500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_97
timestamp 1660789662
transform 1 0 52500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_98
timestamp 1660789662
transform 1 0 50500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_99
timestamp 1660789662
transform 1 0 48500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_100
timestamp 1660789662
transform 1 0 70500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_101
timestamp 1660789662
transform 1 0 68500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_102
timestamp 1660789662
transform 1 0 66500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_103
timestamp 1660789662
transform 1 0 64500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_104
timestamp 1660789662
transform 1 0 62500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_105
timestamp 1660789662
transform 1 0 60500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_106
timestamp 1660789662
transform 1 0 82500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_107
timestamp 1660789662
transform 1 0 80500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_108
timestamp 1660789662
transform 1 0 78500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_109
timestamp 1660789662
transform 1 0 76500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_110
timestamp 1660789662
transform 1 0 74500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_111
timestamp 1660789662
transform 1 0 72500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_112
timestamp 1660789662
transform 1 0 90500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_113
timestamp 1660789662
transform 1 0 86500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_114
timestamp 1660789662
transform 1 0 88500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_115
timestamp 1660789662
transform 1 0 84500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_116
timestamp 1660789662
transform 1 0 -5500 0 1 75600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_117
timestamp 1660789662
transform 1 0 -5500 0 1 73600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_118
timestamp 1660789662
transform 1 0 -5500 0 1 71600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_119
timestamp 1660789662
transform 1 0 -5500 0 1 69600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_120
timestamp 1660789662
transform 1 0 -5500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_121
timestamp 1660789662
transform 1 0 -5500 0 1 65600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_122
timestamp 1660789662
transform 1 0 -5500 0 1 63600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_123
timestamp 1660789662
transform 1 0 -5500 0 1 61600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_124
timestamp 1660789662
transform 1 0 -5500 0 1 59600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_125
timestamp 1660789662
transform 1 0 -5500 0 1 57600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_126
timestamp 1660789662
transform 1 0 -5500 0 1 55600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_127
timestamp 1660789662
transform 1 0 -5500 0 1 53600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_128
timestamp 1660789662
transform 1 0 -5500 0 1 51600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_129
timestamp 1660789662
transform 1 0 -5500 0 1 49600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_130
timestamp 1660789662
transform 1 0 8500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_131
timestamp 1660789662
transform 1 0 10500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_132
timestamp 1660789662
transform 1 0 12500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_133
timestamp 1660789662
transform 1 0 14500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_134
timestamp 1660789662
transform 1 0 22500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_135
timestamp 1660789662
transform 1 0 16500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_136
timestamp 1660789662
transform 1 0 18500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_137
timestamp 1660789662
transform 1 0 20500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_138
timestamp 1660789662
transform 1 0 30500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_139
timestamp 1660789662
transform 1 0 24500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_140
timestamp 1660789662
transform 1 0 26500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_141
timestamp 1660789662
transform 1 0 28500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_142
timestamp 1660789662
transform 1 0 34500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_143
timestamp 1660789662
transform 1 0 32500 0 1 67600
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_144
timestamp 1660789662
transform 1 0 14500 0 1 -14400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_145
timestamp 1660789662
transform 1 0 14500 0 1 -16400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_146
timestamp 1660789662
transform 1 0 14500 0 1 -18400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_147
timestamp 1660789662
transform 1 0 14500 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_148
timestamp 1660789662
transform 1 0 14500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_149
timestamp 1660789662
transform 1 0 16500 0 1 -24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_150
timestamp 1660789662
transform 1 0 16500 0 1 -26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_151
timestamp 1660789662
transform 1 0 20500 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_152
timestamp 1660789662
transform 1 0 20500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_153
timestamp 1660789662
transform 1 0 20500 0 1 -24400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_154
timestamp 1660789662
transform 1 0 20500 0 1 -26400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_155
timestamp 1660789662
transform 1 0 16500 0 1 -28400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_156
timestamp 1660789662
transform 1 0 16500 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_157
timestamp 1660789662
transform 1 0 18500 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_158
timestamp 1660789662
transform 1 0 20500 0 1 -30400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_159
timestamp 1660789662
transform 1 0 16500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_160
timestamp 1660789662
transform 1 0 34500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_168
timestamp 1660789662
transform 1 0 34500 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_183
timestamp 1660789662
transform 1 0 12500 0 1 -20400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_185
timestamp 1660789662
transform 1 0 12500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_186
timestamp 1660789662
transform 1 0 10500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_255
timestamp 1660789662
transform 1 0 -11500 0 1 -22400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_256
timestamp 1660789662
transform 1 0 -15500 0 1 -18400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_258
timestamp 1660789662
transform 1 0 -17000 0 1 -16400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_259
timestamp 1660789662
transform 1 0 -17000 0 1 -14400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_260
timestamp 1660789662
transform 1 0 -17000 0 1 -12400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_261
timestamp 1660789662
transform 1 0 -17000 0 1 -4400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_262
timestamp 1660789662
transform 1 0 -17000 0 1 -8400
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10  hash_m1m2m3m4_W10L10_263
timestamp 1660789662
transform 1 0 -17000 0 1 -6400
box 0 -1700 2000 300
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1662263286
transform 1 0 -11500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_1
timestamp 1662263286
transform 1 0 -7500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_2
timestamp 1662263286
transform 1 0 24500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_3
timestamp 1662263286
transform 1 0 -27500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_4
timestamp 1662263286
transform 1 0 -83500 0 1 31900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_5
timestamp 1662263286
transform 1 0 -15500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_6
timestamp 1662263286
transform 1 0 -19500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_7
timestamp 1662263286
transform 1 0 -27500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_8
timestamp 1662263286
transform 1 0 -23500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_9
timestamp 1662263286
transform 1 0 28500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_10
timestamp 1662263286
transform 1 0 22000 0 1 13900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_11
timestamp 1662263286
transform 1 0 32500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_12
timestamp 1662263286
transform 1 0 36500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_13
timestamp 1662263286
transform 1 0 -31500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_14
timestamp 1662263286
transform 1 0 -19500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_15
timestamp 1662263286
transform 1 0 -29500 0 1 -21600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_16
timestamp 1662263286
transform 1 0 -19500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_17
timestamp 1662263286
transform 1 0 -29500 0 1 -25600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_18
timestamp 1662263286
transform 1 0 15500 0 1 -5600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_19
timestamp 1662263286
transform 1 0 15500 0 1 -9600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_20
timestamp 1662263286
transform 1 0 19500 0 1 -9600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_21
timestamp 1662263286
transform 1 0 -83500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_22
timestamp 1662263286
transform 1 0 -71500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_23
timestamp 1662263286
transform 1 0 -83500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_24
timestamp 1662263286
transform 1 0 -83500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_25
timestamp 1662263286
transform 1 0 -83500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_26
timestamp 1662263286
transform 1 0 4500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_27
timestamp 1662263286
transform 1 0 -29500 0 1 -29600
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_28
timestamp 1662263286
transform 1 0 8500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_29
timestamp 1662263286
transform 1 0 -83500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_30
timestamp 1662263286
transform 1 0 -83500 0 1 -20100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_31
timestamp 1662263286
transform 1 0 -83500 0 1 -24100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_32
timestamp 1662263286
transform 1 0 -35500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_33
timestamp 1662263286
transform 1 0 -83500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_34
timestamp 1662263286
transform 1 0 -27500 0 1 23900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_35
timestamp 1662263286
transform 1 0 -31500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_36
timestamp 1662263286
transform 1 0 -63500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_37
timestamp 1662263286
transform 1 0 -27500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_38
timestamp 1662263286
transform 1 0 -27500 0 1 -8100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_39
timestamp 1662263286
transform 1 0 -59500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_40
timestamp 1662263286
transform 1 0 -27500 0 1 -4100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_41
timestamp 1662263286
transform 1 0 -55500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_42
timestamp 1662263286
transform 1 0 -51500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_43
timestamp 1662263286
transform 1 0 -47500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_44
timestamp 1662263286
transform 1 0 -43500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_45
timestamp 1662263286
transform 1 0 -71500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_46
timestamp 1662263286
transform 1 0 -31500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_47
timestamp 1662263286
transform 1 0 -39500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_48
timestamp 1662263286
transform 1 0 -27500 0 1 -100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_49
timestamp 1662263286
transform 1 0 76500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_50
timestamp 1662263286
transform 1 0 -19500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_51
timestamp 1662263286
transform 1 0 84500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_52
timestamp 1662263286
transform 1 0 -19500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_53
timestamp 1662263286
transform 1 0 -27500 0 1 31900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_54
timestamp 1662263286
transform 1 0 88500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_55
timestamp 1662263286
transform 1 0 76500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_56
timestamp 1662263286
transform 1 0 -15500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_57
timestamp 1662263286
transform 1 0 -3500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_58
timestamp 1662263286
transform 1 0 -7500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_59
timestamp 1662263286
transform 1 0 12500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_60
timestamp 1662263286
transform 1 0 8500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_61
timestamp 1662263286
transform 1 0 88500 0 1 23900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_62
timestamp 1662263286
transform 1 0 4500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_63
timestamp 1662263286
transform 1 0 500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_64
timestamp 1662263286
transform 1 0 88500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_65
timestamp 1662263286
transform 1 0 -11500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_66
timestamp 1662263286
transform 1 0 18500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_67
timestamp 1662263286
transform 1 0 84500 0 1 -20100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_71
timestamp 1662263286
transform 1 0 36500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_72
timestamp 1662263286
transform 1 0 92500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_74
timestamp 1662263286
transform 1 0 18500 0 1 -20100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_75
timestamp 1662263286
transform 1 0 84500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_76
timestamp 1662263286
transform 1 0 88500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_77
timestamp 1662263286
transform 1 0 92500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_78
timestamp 1662263286
transform 1 0 80500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_79
timestamp 1662263286
transform 1 0 76500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_80
timestamp 1662263286
transform 1 0 72500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_81
timestamp 1662263286
transform 1 0 68500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_82
timestamp 1662263286
transform 1 0 64500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_83
timestamp 1662263286
transform 1 0 60500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_84
timestamp 1662263286
transform 1 0 56500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_85
timestamp 1662263286
transform 1 0 52500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_86
timestamp 1662263286
transform 1 0 36500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_87
timestamp 1662263286
transform 1 0 36500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_88
timestamp 1662263286
transform 1 0 40500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_89
timestamp 1662263286
transform 1 0 44500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_90
timestamp 1662263286
transform 1 0 48500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_95
timestamp 1662263286
transform 1 0 8500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_96
timestamp 1662263286
transform 1 0 12500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_97
timestamp 1662263286
transform 1 0 12500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_98
timestamp 1662263286
transform 1 0 16500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_99
timestamp 1662263286
transform 1 0 18500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_100
timestamp 1662263286
transform 1 0 16500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_101
timestamp 1662263286
transform 1 0 96500 0 1 19900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_102
timestamp 1662263286
transform 1 0 -39500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_103
timestamp 1662263286
transform 1 0 -35500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_104
timestamp 1662263286
transform 1 0 96500 0 1 15900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_105
timestamp 1662263286
transform 1 0 96500 0 1 11900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_106
timestamp 1662263286
transform 1 0 96500 0 1 7900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_107
timestamp 1662263286
transform 1 0 96500 0 1 3900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_108
timestamp 1662263286
transform 1 0 96500 0 1 -100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_109
timestamp 1662263286
transform 1 0 96500 0 1 -4100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_110
timestamp 1662263286
transform 1 0 -71500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_111
timestamp 1662263286
transform 1 0 -67500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_112
timestamp 1662263286
transform 1 0 -79500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_113
timestamp 1662263286
transform 1 0 -75500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_114
timestamp 1662263286
transform 1 0 96500 0 1 -8100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_115
timestamp 1662263286
transform 1 0 96500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_116
timestamp 1662263286
transform 1 0 -11500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_117
timestamp 1662263286
transform 1 0 -15500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_118
timestamp 1662263286
transform 1 0 -15500 0 1 -24100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_119
timestamp 1662263286
transform 1 0 -7500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_120
timestamp 1662263286
transform 1 0 -3500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_121
timestamp 1662263286
transform 1 0 500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_122
timestamp 1662263286
transform 1 0 4500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_123
timestamp 1662263286
transform 1 0 96500 0 1 -16100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_124
timestamp 1662263286
transform 1 0 96500 0 1 -20100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_125
timestamp 1662263286
transform 1 0 96500 0 1 -24100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_126
timestamp 1662263286
transform 1 0 96500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_127
timestamp 1662263286
transform 1 0 96500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_128
timestamp 1662263286
transform 1 0 40500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_129
timestamp 1662263286
transform 1 0 44500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_130
timestamp 1662263286
transform 1 0 48500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_131
timestamp 1662263286
transform 1 0 52500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_132
timestamp 1662263286
transform 1 0 56500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_133
timestamp 1662263286
transform 1 0 60500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_134
timestamp 1662263286
transform 1 0 76500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_135
timestamp 1662263286
transform 1 0 72500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_136
timestamp 1662263286
transform 1 0 68500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_137
timestamp 1662263286
transform 1 0 64500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_138
timestamp 1662263286
transform 1 0 84500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_139
timestamp 1662263286
transform 1 0 80500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_140
timestamp 1662263286
transform 1 0 88500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_141
timestamp 1662263286
transform 1 0 -11500 0 1 23900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_142
timestamp 1662263286
transform 1 0 -11500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_143
timestamp 1662263286
transform 1 0 -11500 0 1 31900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_144
timestamp 1662263286
transform 1 0 -11500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_145
timestamp 1662263286
transform 1 0 -35500 0 1 71900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_146
timestamp 1662263286
transform 1 0 -35500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_147
timestamp 1662263286
transform 1 0 -35500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_148
timestamp 1662263286
transform 1 0 -31500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_149
timestamp 1662263286
transform 1 0 -27500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_150
timestamp 1662263286
transform 1 0 -23500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_151
timestamp 1662263286
transform 1 0 -19500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_152
timestamp 1662263286
transform 1 0 -15500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_153
timestamp 1662263286
transform 1 0 -11500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_154
timestamp 1662263286
transform 1 0 -7500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_155
timestamp 1662263286
transform 1 0 20500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_156
timestamp 1662263286
transform 1 0 24500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_157
timestamp 1662263286
transform 1 0 -35500 0 1 63900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_158
timestamp 1662263286
transform 1 0 -35500 0 1 59900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_159
timestamp 1662263286
transform 1 0 -35500 0 1 55900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_160
timestamp 1662263286
transform 1 0 28500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_161
timestamp 1662263286
transform 1 0 32500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_162
timestamp 1662263286
transform 1 0 -35500 0 1 51900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_163
timestamp 1662263286
transform 1 0 -35500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_164
timestamp 1662263286
transform 1 0 4500 0 1 51900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_165
timestamp 1662263286
transform 1 0 4500 0 1 55900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_166
timestamp 1662263286
transform 1 0 4500 0 1 59900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_167
timestamp 1662263286
transform 1 0 8500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_168
timestamp 1662263286
transform 1 0 4500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_169
timestamp 1662263286
transform 1 0 16500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_170
timestamp 1662263286
transform 1 0 12500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_171
timestamp 1662263286
transform 1 0 24500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_172
timestamp 1662263286
transform 1 0 20500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_173
timestamp 1662263286
transform 1 0 32500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_174
timestamp 1662263286
transform 1 0 28500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_175
timestamp 1662263286
transform 1 0 4500 0 1 63900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_176
timestamp 1662263286
transform 1 0 108500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_177
timestamp 1662263286
transform 1 0 112500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_178
timestamp 1662263286
transform 1 0 116500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_179
timestamp 1662263286
transform 1 0 120500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_180
timestamp 1662263286
transform 1 0 124500 0 1 39900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_181
timestamp 1662263286
transform 1 0 124500 0 1 35900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_182
timestamp 1662263286
transform 1 0 124500 0 1 31900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_183
timestamp 1662263286
transform 1 0 124500 0 1 27900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_184
timestamp 1662263286
transform 1 0 124500 0 1 23900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_188
timestamp 1662263286
transform 1 0 136500 0 1 -36100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_189
timestamp 1662263286
transform 1 0 136500 0 1 -40100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_190
timestamp 1662263286
transform 1 0 140500 0 1 -40100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_191
timestamp 1662263286
transform 1 0 140500 0 1 -36100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_192
timestamp 1662263286
transform 1 0 140500 0 1 -32100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_193
timestamp 1662263286
transform 1 0 140500 0 1 -28100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_194
timestamp 1662263286
transform 1 0 140500 0 1 -24100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_195
timestamp 1662263286
transform 1 0 140500 0 1 -12100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_196
timestamp 1662263286
transform 1 0 140500 0 1 -8100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_197
timestamp 1662263286
transform 1 0 140500 0 1 -4100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_198
timestamp 1662263286
transform 1 0 140500 0 1 -100
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_199
timestamp 1662263286
transform 1 0 140500 0 1 3900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_200
timestamp 1662263286
transform 1 0 140500 0 1 7900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_201
timestamp 1662263286
transform 1 0 140500 0 1 11900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_202
timestamp 1662263286
transform 1 0 108500 0 1 59900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_203
timestamp 1662263286
transform 1 0 108500 0 1 63900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_204
timestamp 1662263286
transform 1 0 108500 0 1 67900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_205
timestamp 1662263286
transform 1 0 108500 0 1 71900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_206
timestamp 1662263286
transform 1 0 108500 0 1 75900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_207
timestamp 1662263286
transform 1 0 108500 0 1 55900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_208
timestamp 1662263286
transform 1 0 108500 0 1 51900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_209
timestamp 1662263286
transform 1 0 108500 0 1 47900
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_210
timestamp 1662263286
transform 1 0 108500 0 1 43900
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660792292
transform 1 0 -43500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_1
timestamp 1660792292
transform 1 0 -43500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_2
timestamp 1660792292
transform 1 0 -43500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_3
timestamp 1660792292
transform 1 0 -43500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_4
timestamp 1660792292
transform 1 0 -35500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_5
timestamp 1660792292
transform 1 0 -27500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_6
timestamp 1660792292
transform 1 0 -15500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_7
timestamp 1660792292
transform 1 0 -83500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_8
timestamp 1660792292
transform 1 0 -75500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_9
timestamp 1660792292
transform 1 0 -67500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_10
timestamp 1660792292
transform 1 0 -59500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_11
timestamp 1660792292
transform 1 0 -3500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_12
timestamp 1660792292
transform 1 0 100500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_13
timestamp 1660792292
transform 1 0 100500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_14
timestamp 1660792292
transform 1 0 100500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_15
timestamp 1660792292
transform 1 0 -63500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_16
timestamp 1660792292
transform 1 0 -51500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_17
timestamp 1660792292
transform 1 0 -55500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_18
timestamp 1660792292
transform 1 0 100500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_19
timestamp 1660792292
transform 1 0 -47500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_20
timestamp 1660792292
transform 1 0 100500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_21
timestamp 1660792292
transform 1 0 100500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_22
timestamp 1660792292
transform 1 0 108500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_23
timestamp 1660792292
transform 1 0 -71500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_24
timestamp 1660792292
transform 1 0 116500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_25
timestamp 1660792292
transform 1 0 -79500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_26
timestamp 1660792292
transform 1 0 44500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_27
timestamp 1660792292
transform 1 0 -83500 0 1 -8100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_28
timestamp 1660792292
transform 1 0 -83500 0 1 -100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_29
timestamp 1660792292
transform 1 0 -83500 0 1 7900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_30
timestamp 1660792292
transform 1 0 -83500 0 1 15900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_31
timestamp 1660792292
transform 1 0 -83500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_32
timestamp 1660792292
transform 1 0 -79500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_33
timestamp 1660792292
transform 1 0 52500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_34
timestamp 1660792292
transform 1 0 60500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_35
timestamp 1660792292
transform 1 0 68500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_36
timestamp 1660792292
transform 1 0 -79500 0 1 -16100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_37
timestamp 1660792292
transform 1 0 -79500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_38
timestamp 1660792292
transform 1 0 -71500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_39
timestamp 1660792292
transform 1 0 76500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_40
timestamp 1660792292
transform 1 0 -67500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_41
timestamp 1660792292
transform 1 0 -83500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_42
timestamp 1660792292
transform 1 0 -39500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_43
timestamp 1660792292
transform 1 0 -75500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_44
timestamp 1660792292
transform 1 0 -59500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_45
timestamp 1660792292
transform 1 0 100500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_46
timestamp 1660792292
transform 1 0 -51500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_47
timestamp 1660792292
transform 1 0 108500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_48
timestamp 1660792292
transform 1 0 116500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_49
timestamp 1660792292
transform 1 0 108500 0 1 7900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_50
timestamp 1660792292
transform 1 0 100500 0 1 7900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_51
timestamp 1660792292
transform 1 0 92500 0 1 47900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_52
timestamp 1660792292
transform 1 0 28500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_53
timestamp 1660792292
transform 1 0 100500 0 1 15900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_54
timestamp 1660792292
transform 1 0 -3500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_55
timestamp 1660792292
transform 1 0 -83500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_56
timestamp 1660792292
transform 1 0 100500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_57
timestamp 1660792292
transform 1 0 108500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_58
timestamp 1660792292
transform 1 0 108500 0 1 15900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_59
timestamp 1660792292
transform 1 0 92500 0 1 39900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_60
timestamp 1660792292
transform 1 0 92500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_61
timestamp 1660792292
transform 1 0 92500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_62
timestamp 1660792292
transform 1 0 88500 0 1 11900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_63
timestamp 1660792292
transform 1 0 88500 0 1 3900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_64
timestamp 1660792292
transform 1 0 88500 0 1 -4100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_65
timestamp 1660792292
transform 1 0 88500 0 1 -12100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_66
timestamp 1660792292
transform 1 0 88500 0 1 -20100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_67
timestamp 1660792292
transform 1 0 -75500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_68
timestamp 1660792292
transform 1 0 88500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_69
timestamp 1660792292
transform 1 0 -83500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_70
timestamp 1660792292
transform 1 0 -75500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_71
timestamp 1660792292
transform 1 0 -59500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_72
timestamp 1660792292
transform 1 0 84500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_73
timestamp 1660792292
transform 1 0 -59500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_74
timestamp 1660792292
transform 1 0 -67500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_75
timestamp 1660792292
transform 1 0 36500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_76
timestamp 1660792292
transform 1 0 28500 0 1 31900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_77
timestamp 1660792292
transform 1 0 80500 0 1 -28100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_78
timestamp 1660792292
transform 1 0 80500 0 1 23900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_79
timestamp 1660792292
transform 1 0 92500 0 1 55900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_80
timestamp 1660792292
transform 1 0 -67500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_81
timestamp 1660792292
transform 1 0 116500 0 1 15900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_82
timestamp 1660792292
transform 1 0 124500 0 1 15900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_83
timestamp 1660792292
transform 1 0 -51500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_84
timestamp 1660792292
transform 1 0 -51500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_85
timestamp 1660792292
transform 1 0 124500 0 1 7900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_86
timestamp 1660792292
transform 1 0 116500 0 1 7900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_87
timestamp 1660792292
transform 1 0 132500 0 1 15900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_88
timestamp 1660792292
transform 1 0 132500 0 1 7900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_89
timestamp 1660792292
transform 1 0 100500 0 1 -100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_90
timestamp 1660792292
transform 1 0 108500 0 1 -100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_91
timestamp 1660792292
transform 1 0 116500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_92
timestamp 1660792292
transform 1 0 108500 0 1 -8100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_93
timestamp 1660792292
transform 1 0 4500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_94
timestamp 1660792292
transform 1 0 100500 0 1 -8100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_95
timestamp 1660792292
transform 1 0 -3500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_96
timestamp 1660792292
transform 1 0 -3500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_97
timestamp 1660792292
transform 1 0 20500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_98
timestamp 1660792292
transform 1 0 124500 0 1 -8100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_99
timestamp 1660792292
transform 1 0 12500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_100
timestamp 1660792292
transform 1 0 116500 0 1 -8100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_101
timestamp 1660792292
transform 1 0 116500 0 1 -100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_102
timestamp 1660792292
transform 1 0 28500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_103
timestamp 1660792292
transform 1 0 36500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_104
timestamp 1660792292
transform 1 0 44500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_105
timestamp 1660792292
transform 1 0 60500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_106
timestamp 1660792292
transform 1 0 52500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_107
timestamp 1660792292
transform 1 0 76500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_108
timestamp 1660792292
transform 1 0 68500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_109
timestamp 1660792292
transform 1 0 92500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_110
timestamp 1660792292
transform 1 0 84500 0 1 71900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_111
timestamp 1660792292
transform 1 0 92500 0 1 63900
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_112
timestamp 1660792292
transform 1 0 34500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_113
timestamp 1660792292
transform 1 0 42500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_114
timestamp 1660792292
transform 1 0 50500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_115
timestamp 1660792292
transform 1 0 58500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_116
timestamp 1660792292
transform 1 0 62500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_117
timestamp 1660792292
transform 1 0 88500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_118
timestamp 1660792292
transform 1 0 92500 0 1 -40100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_119
timestamp 1660792292
transform 1 0 124500 0 1 -100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_120
timestamp 1660792292
transform 1 0 132500 0 1 -8100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_121
timestamp 1660792292
transform 1 0 132500 0 1 -100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_122
timestamp 1660792292
transform 1 0 108500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_123
timestamp 1660792292
transform 1 0 100500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_124
timestamp 1660792292
transform 1 0 108500 0 1 -16100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_125
timestamp 1660792292
transform 1 0 100500 0 1 -16100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_126
timestamp 1660792292
transform 1 0 116500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_127
timestamp 1660792292
transform 1 0 116500 0 1 -16100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_128
timestamp 1660792292
transform 1 0 132500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_129
timestamp 1660792292
transform 1 0 124500 0 1 -24100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_130
timestamp 1660792292
transform 1 0 132500 0 1 -16100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_131
timestamp 1660792292
transform 1 0 124500 0 1 -16100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_132
timestamp 1660792292
transform 1 0 108500 0 1 -32100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_133
timestamp 1660792292
transform 1 0 100500 0 1 -32100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_134
timestamp 1660792292
transform 1 0 116500 0 1 -32100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_135
timestamp 1660792292
transform 1 0 132500 0 1 -32100
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_136
timestamp 1660792292
transform 1 0 124500 0 1 -32100
box 0 0 8000 8000
<< labels >>
rlabel metal4 -23600 -16400 -22500 -16300 1 VHI
rlabel metal3 -23600 -21300 -23500 -21100 1 G32
rlabel metal3 -23400 -21300 -23300 -21100 1 G16
rlabel metal3 -23200 -21300 -23100 -21100 1 G2
rlabel metal3 -23000 -21300 -22900 -21100 1 G4
rlabel metal3 -22800 -21300 -22700 -21100 1 G8
rlabel metal5 -21700 -20050 -20900 -19450 3 IREF
<< end >>
