* SPICE3 file created from PA_core_1.ext - technology: sky130B

X0 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X1 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X2 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X3 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X4 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X5 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X6 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X7 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X8 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X9 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X10 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X11 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X12 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X13 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X14 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X15 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X16 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X17 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X18 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X19 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X20 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X21 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X22 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X23 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X24 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X25 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X26 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X27 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X28 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X29 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X30 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X31 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X32 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X33 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X34 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X35 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X36 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X37 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X38 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X39 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X40 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X41 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X42 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X43 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X44 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X45 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X46 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X47 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X48 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X49 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X50 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X51 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X52 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X53 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X54 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X55 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X56 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X57 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X58 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X59 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X60 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X61 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X62 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X63 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X64 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X65 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X66 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X67 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X68 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X69 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X70 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X71 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X72 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X73 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X74 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X75 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X76 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X77 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X78 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X79 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X80 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X81 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X82 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X83 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X84 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X85 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X86 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X87 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X88 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X89 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X90 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X91 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X92 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X93 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X94 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X95 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X96 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X97 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X98 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X99 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X100 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X101 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X102 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X103 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X104 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X105 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X106 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X107 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X108 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X109 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X110 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X111 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X112 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X113 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X114 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X115 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X116 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X117 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X118 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X119 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X120 MID RF_nfet_3v_dnwell_cascode_0/G2 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X121 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X122 MID RF_nfet_3v_dnwell_cascode_0/G1 DRAIN MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X123 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X124 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X125 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X126 DRAIN RF_nfet_3v_dnwell_cascode_0/G1 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X127 DRAIN RF_nfet_3v_dnwell_cascode_0/G2 MID MID sky130_fd_pr__nfet_03v3_nvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=500000u
X128 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X129 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X130 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X131 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X132 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X133 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X134 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X135 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X136 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X137 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X138 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X139 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X140 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X141 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X142 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X143 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X144 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X145 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X146 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X147 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X148 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X149 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X150 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X151 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X152 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X153 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X154 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X155 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X156 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X157 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X158 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X159 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X160 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X161 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X162 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X163 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X164 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X165 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X166 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X167 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X168 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X169 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X170 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X171 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X172 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X173 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X174 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X175 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X176 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X177 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X178 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X179 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X180 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X181 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X182 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X183 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X184 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X185 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X186 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X187 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X188 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X189 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X190 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X191 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X192 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X193 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X194 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X195 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X196 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X197 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X198 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X199 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X200 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X201 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X202 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X203 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X204 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X205 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X206 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X207 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X208 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X209 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X210 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X211 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X212 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X213 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X214 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X215 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X216 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X217 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X218 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X219 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X220 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X221 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X222 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X223 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X224 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X225 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X226 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X227 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X228 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X229 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X230 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X231 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X232 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X233 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X234 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X235 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X236 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X237 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X238 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X239 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X240 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X241 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X242 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X243 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X244 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X245 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X246 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X247 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X248 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X249 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X250 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X251 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X252 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X253 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X254 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X255 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X256 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X257 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X258 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X259 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X260 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X261 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X262 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X263 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X264 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X265 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X266 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X267 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X268 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X269 VSUB GATE MID VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X270 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X271 MID GATE VSUB VSUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X272 TOPBIAS_L RF_nfet_3v_dnwell_cascode_0/G2 VSUB sky130_fd_pr__res_high_po_0p35 l=3e+06u
X273 RF_nfet_3v_dnwell_cascode_0/G1 TOPBIAS_R VSUB sky130_fd_pr__res_high_po_0p35 l=3e+06u
C0 RF_nfet_3v_dnwell_cascode_0/G1 DRAIN 22.62fF
C1 RF_nfet_3v_dnwell_cascode_0/G1 VSUB 4.64fF
C2 RF_nfet_3v_dnwell_cascode_0/G1 MID 27.80fF
C3 GATE VSUB 27.73fF
C4 GATE MID 34.68fF
C5 VSUB DRAIN 3.98fF
C6 MID DRAIN 194.17fF
C7 VSUB MID 355.73fF
C8 RF_nfet_3v_dnwell_cascode_0/G2 DRAIN 22.66fF
C9 RF_nfet_3v_dnwell_cascode_0/G2 VSUB 4.80fF
C10 RF_nfet_3v_dnwell_cascode_0/G2 MID 29.29fF
C11 GATE 0 17.76fF **FLOATING
C12 VSUB 0 85.58fF **FLOATING
C13 RF_nfet_3v_dnwell_cascode_0/G1 0 4.12fF **FLOATING
C14 RF_nfet_3v_dnwell_cascode_0/G2 0 4.07fF **FLOATING
