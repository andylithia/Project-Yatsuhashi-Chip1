magic
tech sky130A
magscale 1 2
timestamp 1665275542
<< pwell >>
rect 29802 38680 30200 40458
rect 30802 25480 31200 27258
rect 30798 12500 31200 14016
<< psubdiff >>
rect 29838 40388 29934 40422
rect 30068 40388 30164 40422
rect 29838 40326 29872 40388
rect 30130 40326 30164 40388
rect 29838 38750 29872 38812
rect 30130 38750 30164 38812
rect 29838 38716 29934 38750
rect 30068 38716 30164 38750
rect 30838 27188 30934 27222
rect 31068 27188 31164 27222
rect 30838 27126 30872 27188
rect 31130 27126 31164 27188
rect 30838 25550 30872 25612
rect 31130 25550 31164 25612
rect 30838 25516 30934 25550
rect 31068 25516 31164 25550
rect 30834 13946 30930 13980
rect 31068 13946 31164 13980
rect 30834 13884 30868 13946
rect 31130 13884 31164 13946
rect 30834 12570 30868 12632
rect 31130 12570 31164 12632
rect 30834 12536 30930 12570
rect 31068 12536 31164 12570
<< psubdiffcont >>
rect 29934 40388 30068 40422
rect 29838 38812 29872 40326
rect 30130 38812 30164 40326
rect 29934 38716 30068 38750
rect 30934 27188 31068 27222
rect 30838 25612 30872 27126
rect 31130 25612 31164 27126
rect 30934 25516 31068 25550
rect 30930 13946 31068 13980
rect 30834 12632 30868 13884
rect 31130 12632 31164 13884
rect 30930 12536 31068 12570
<< poly >>
rect 29968 40276 30034 40292
rect 29968 40242 29984 40276
rect 30018 40242 30034 40276
rect 29968 40219 30034 40242
rect 29968 38896 30034 38919
rect 29968 38862 29984 38896
rect 30018 38862 30034 38896
rect 29968 38846 30034 38862
rect 30968 27076 31034 27092
rect 30968 27042 30984 27076
rect 31018 27042 31034 27076
rect 30968 27019 31034 27042
rect 30968 25696 31034 25719
rect 30968 25662 30984 25696
rect 31018 25662 31034 25696
rect 30968 25646 31034 25662
<< polycont >>
rect 29984 40242 30018 40276
rect 29984 38862 30018 38896
rect 30984 27042 31018 27076
rect 30984 25662 31018 25696
<< xpolycontact >>
rect 30964 13418 31034 13850
rect 30964 12666 31034 13098
<< npolyres >>
rect 29968 38919 30034 40219
rect 30968 25719 31034 27019
<< ppolyres >>
rect 30964 13098 31034 13418
<< locali >>
rect 29838 40420 29934 40422
rect -3060 40400 -2980 40420
rect -3060 38740 -3040 40400
rect -3000 38740 -2980 40400
rect -3060 38720 -2980 38740
rect 29780 40400 29934 40420
rect 29780 38720 29800 40400
rect 29840 40388 29934 40400
rect 30068 40388 30164 40422
rect 29840 40326 29872 40388
rect 30130 40326 30164 40388
rect 29968 40242 29984 40276
rect 30018 40242 30034 40276
rect 29968 38862 29984 38896
rect 30018 38862 30034 38896
rect 29840 38750 29872 38812
rect 30130 38750 30164 38812
rect 29840 38720 29934 38750
rect 29780 38716 29934 38720
rect 30068 38716 30164 38750
rect 29780 38700 29860 38716
rect -4060 27200 -3980 27220
rect -4060 25540 -4040 27200
rect -4000 25540 -3980 27200
rect 30838 27188 30934 27222
rect 31068 27188 31164 27222
rect 30838 27126 30872 27188
rect 30780 26980 30838 27000
rect 31130 27126 31164 27188
rect 30968 27042 30984 27076
rect 31018 27042 31034 27076
rect 30780 26020 30800 26980
rect 30780 26000 30838 26020
rect -4060 25520 -3980 25540
rect 30968 25662 30984 25696
rect 31018 25662 31034 25696
rect 30838 25550 30872 25612
rect 31130 25550 31164 25612
rect 30838 25516 30934 25550
rect 31068 25516 31164 25550
rect 30780 13980 30860 14000
rect -4060 13940 -3980 13960
rect -4060 12560 -4040 13940
rect -4000 12560 -3980 13940
rect -4060 12540 -3980 12560
rect 30780 12520 30800 13980
rect 30840 13946 30930 13980
rect 31068 13946 31164 13980
rect 30840 13884 30868 13946
rect 31130 13884 31164 13946
rect 30840 12570 30868 12632
rect 31130 12570 31164 12632
rect 30840 12536 30930 12570
rect 31068 12536 31164 12570
rect 30840 12520 30860 12536
rect 30780 12500 30860 12520
<< viali >>
rect -3040 38740 -3000 40400
rect 29800 40326 29840 40400
rect 29800 38812 29838 40326
rect 29838 38812 29840 40326
rect 29984 40242 30018 40276
rect 29984 40236 30018 40242
rect 29984 38896 30018 38902
rect 29984 38862 30018 38896
rect 29800 38720 29840 38812
rect -4040 25540 -4000 27200
rect 30984 27042 31018 27076
rect 30984 27036 31018 27042
rect 30800 26020 30838 26980
rect 30838 26020 30840 26980
rect 30984 25696 31018 25702
rect 30984 25662 31018 25696
rect -4040 12560 -4000 13940
rect 30800 13884 30840 13980
rect 30800 12632 30834 13884
rect 30834 12632 30840 13884
rect 30980 13435 31018 13832
rect 30980 12684 31018 13081
rect 30800 12520 30840 12632
<< metal1 >>
rect -3300 40450 -3100 40460
rect -3300 40190 -3290 40450
rect -3110 40190 -3100 40450
rect -3300 40180 -3100 40190
rect -3060 40400 -2980 40420
rect -3300 38910 -3100 38920
rect -3300 38690 -3290 38910
rect -3110 38690 -3100 38910
rect -3060 38740 -3040 40400
rect -3000 38740 -2980 40400
rect -3060 38720 -2980 38740
rect -3300 38680 -3100 38690
rect 1000 32500 1340 46500
rect 25260 32500 25500 46500
rect 29900 40450 30100 40460
rect 29780 40400 29860 40420
rect 29780 40000 29800 40400
rect 29500 39000 29800 40000
rect 29780 38720 29800 39000
rect 29840 38720 29860 40400
rect 29900 40190 29910 40450
rect 30090 40190 30100 40450
rect 29900 40180 30100 40190
rect 29780 38700 29860 38720
rect 29900 38910 30100 38920
rect 29900 38690 29910 38910
rect 30090 38690 30100 38910
rect 29900 38680 30100 38690
rect -4300 27250 -4100 27260
rect -4300 27030 -4290 27250
rect -4110 27030 -4100 27250
rect -4300 27020 -4100 27030
rect -4060 27200 -3980 27220
rect -4300 25710 -4100 25720
rect -4300 25490 -4290 25710
rect -4110 25490 -4100 25710
rect -4060 25540 -4040 27200
rect -4000 25540 -3980 27200
rect -4060 25520 -3980 25540
rect -4300 25480 -4100 25490
rect 1000 17000 1340 31500
rect 25260 17000 25500 31500
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect 30500 26980 30860 27000
rect 30500 26020 30800 26980
rect 30840 26020 30860 26980
rect 30500 26000 30860 26020
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect -4060 13940 -3980 13960
rect -4300 13900 -4100 13910
rect -4300 13420 -4290 13900
rect -4110 13420 -4100 13900
rect -4300 13410 -4100 13420
rect -4300 13090 -4100 13100
rect -4300 12610 -4290 13090
rect -4110 12610 -4100 13090
rect -4300 12600 -4100 12610
rect -4060 12560 -4040 13940
rect -4000 12560 -3980 13940
rect -3920 13900 -3540 14000
rect -4060 12540 -3980 12560
rect 1000 2180 1340 16000
rect 6360 2180 6500 2500
rect 1000 2000 6500 2180
rect 7500 2180 7640 2500
rect 12700 2180 13000 2500
rect 7500 2000 13000 2180
rect 13500 2180 14000 2500
rect 18980 2180 19500 2500
rect 13500 2000 19500 2180
rect 20000 2160 20260 2500
rect 25260 2160 25500 16000
rect 30500 13980 30860 14000
rect 30500 13000 30800 13980
rect 30780 12520 30800 13000
rect 30840 12520 30860 13980
rect 30900 13900 31100 13910
rect 30900 13420 30910 13900
rect 31090 13420 31100 13900
rect 30900 13410 31100 13420
rect 30900 13090 31100 13100
rect 30900 12610 30910 13090
rect 31090 12610 31100 13090
rect 30900 12600 31100 12610
rect 30780 12500 30860 12520
rect 20000 2000 25500 2160
<< via1 >>
rect -3290 40190 -3110 40450
rect -3290 38690 -3110 38910
rect 29910 40276 30090 40450
rect 29910 40236 29984 40276
rect 29984 40236 30018 40276
rect 30018 40236 30090 40276
rect 29910 40190 30090 40236
rect 29910 38902 30090 38910
rect 29910 38862 29984 38902
rect 29984 38862 30018 38902
rect 30018 38862 30090 38902
rect 29910 38690 30090 38862
rect -4290 27030 -4110 27250
rect -4290 25490 -4110 25710
rect 30910 27076 31090 27250
rect 30910 27036 30984 27076
rect 30984 27036 31018 27076
rect 31018 27036 31090 27076
rect 30910 27030 31090 27036
rect 30910 25702 31090 25710
rect 30910 25662 30984 25702
rect 30984 25662 31018 25702
rect 31018 25662 31090 25702
rect 30910 25490 31090 25662
rect -4290 13420 -4110 13900
rect -4290 12610 -4110 13090
rect 30910 13832 31090 13900
rect 30910 13435 30980 13832
rect 30980 13435 31018 13832
rect 31018 13435 31090 13832
rect 30910 13420 31090 13435
rect 30910 13081 31090 13090
rect 30910 12684 30980 13081
rect 30980 12684 31018 13081
rect 31018 12684 31090 13081
rect 30910 12610 31090 12684
<< metal2 >>
rect -3300 40450 -3100 40460
rect -3300 40190 -3290 40450
rect -3110 40190 -3100 40450
rect -3300 40180 -3100 40190
rect 29900 40450 30100 40460
rect 29900 40190 29910 40450
rect 30090 40190 30100 40450
rect 29900 40180 30100 40190
rect -3300 38910 -3100 38920
rect -3300 38690 -3290 38910
rect -3110 38690 -3100 38910
rect -3300 38680 -3100 38690
rect 29900 38910 30100 38920
rect 29900 38690 29910 38910
rect 30090 38690 30100 38910
rect 29900 38680 30100 38690
rect -4300 27250 -4100 27260
rect -4300 27030 -4290 27250
rect -4110 27030 -4100 27250
rect -4300 27020 -4100 27030
rect 30900 27250 31100 27260
rect 30900 27030 30910 27250
rect 31090 27030 31100 27250
rect 30900 27020 31100 27030
rect -4300 25710 -4100 25720
rect -4300 25490 -4290 25710
rect -4110 25490 -4100 25710
rect -4300 25480 -4100 25490
rect 30900 25710 31100 25720
rect 30900 25490 30910 25710
rect 31090 25490 31100 25710
rect 30900 25480 31100 25490
rect -4300 13900 -4100 13910
rect -4300 13420 -4290 13900
rect -4110 13420 -4100 13900
rect -4300 13410 -4100 13420
rect 30900 13900 31100 13910
rect 30900 13420 30910 13900
rect 31090 13420 31100 13900
rect 30900 13410 31100 13420
rect -4300 13090 -4100 13100
rect -4300 12610 -4290 13090
rect -4110 12610 -4100 13090
rect -4300 12600 -4100 12610
rect 30900 13090 31100 13100
rect 30900 12610 30910 13090
rect 31090 12610 31100 13090
rect 30900 12600 31100 12610
<< via2 >>
rect -3290 40190 -3110 40450
rect 29910 40190 30090 40450
rect -3290 38690 -3110 38910
rect 29910 38690 30090 38910
rect -4290 27030 -4110 27250
rect 30910 27030 31090 27250
rect -4290 25490 -4110 25710
rect 30910 25490 31090 25710
rect -4290 13420 -4110 13900
rect 30910 13420 31090 13900
rect -4290 12610 -4110 13090
rect 30910 12610 31090 13090
<< metal3 >>
rect -3400 40480 -3000 40500
rect -3400 40410 -3380 40480
rect -3400 40190 -3390 40410
rect -3020 40410 -3000 40480
rect -3010 40190 -3000 40410
rect -3400 40180 -3000 40190
rect 29800 40480 30200 40500
rect 29800 40410 29820 40480
rect 29800 40190 29810 40410
rect 30180 40410 30200 40480
rect 30190 40190 30200 40410
rect 29800 40180 30200 40190
rect -3400 38910 -3000 38920
rect -3400 38690 -3390 38910
rect -3010 38690 -3000 38910
rect -3400 38680 -3000 38690
rect 29800 38910 30200 38920
rect 29800 38690 29810 38910
rect 30190 38690 30200 38910
rect 29800 38680 30200 38690
rect -4400 31700 2800 31800
rect -4400 31100 1400 31700
rect 2700 31100 2800 31700
rect -4400 31000 2800 31100
rect 24000 31700 31200 31800
rect 24000 31100 24100 31700
rect 25400 31100 31200 31700
rect 24000 31000 31200 31100
rect -4400 27250 -3900 31000
rect -4400 27030 -4290 27250
rect -4110 27030 -3900 27250
rect -4400 27000 -3900 27030
rect 30700 27250 31200 31000
rect 30700 27030 30910 27250
rect 31090 27030 31200 27250
rect 30700 27000 31200 27030
rect -4400 25710 -4000 25720
rect -4400 25490 -4390 25710
rect -4010 25490 -4000 25710
rect -4400 25480 -4000 25490
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25480 31200 25490
rect -4400 14000 -4000 14010
rect -4400 13420 -4390 14000
rect -4010 13420 -4000 14000
rect -4400 13410 -4000 13420
rect 30800 14000 31200 14010
rect 30800 13420 30810 14000
rect 31190 13420 31200 14000
rect 30800 13410 31200 13420
rect -4400 13090 -4000 13100
rect -4400 12510 -4390 13090
rect -4010 12510 -4000 13090
rect -4400 12500 -4000 12510
rect 30800 13090 31200 13100
rect 30800 12510 30810 13090
rect 31190 12510 31200 13090
rect 30800 12500 31200 12510
<< via3 >>
rect -3380 40450 -3020 40480
rect -3380 40410 -3290 40450
rect -3390 40190 -3290 40410
rect -3290 40190 -3110 40450
rect -3110 40410 -3020 40450
rect -3110 40190 -3010 40410
rect 29820 40450 30180 40480
rect 29820 40410 29910 40450
rect 29810 40190 29910 40410
rect 29910 40190 30090 40450
rect 30090 40410 30180 40450
rect 30090 40190 30190 40410
rect -3390 38690 -3290 38910
rect -3290 38690 -3110 38910
rect -3110 38690 -3010 38910
rect 29810 38690 29910 38910
rect 29910 38690 30090 38910
rect 30090 38690 30190 38910
rect 1400 31100 2700 31700
rect 24100 31100 25400 31700
rect -4390 25490 -4290 25710
rect -4290 25490 -4110 25710
rect -4110 25490 -4010 25710
rect 30810 25490 30910 25710
rect 30910 25490 31090 25710
rect 31090 25490 31190 25710
rect -4390 13900 -4010 14000
rect -4390 13420 -4290 13900
rect -4290 13420 -4110 13900
rect -4110 13420 -4010 13900
rect 30810 13900 31190 14000
rect 30810 13420 30910 13900
rect 30910 13420 31090 13900
rect 31090 13420 31190 13900
rect -4390 12610 -4290 13090
rect -4290 12610 -4110 13090
rect -4110 12610 -4010 13090
rect -4390 12510 -4010 12610
rect 30810 12610 30910 13090
rect 30910 12610 31090 13090
rect 31090 12610 31190 13090
rect 30810 12510 31190 12610
<< metal4 >>
rect -3400 40800 800 46000
rect -3400 40480 -3000 40500
rect -3400 40410 -3380 40480
rect -3400 40190 -3390 40410
rect -3020 40410 -3000 40480
rect -3010 40190 -3000 40410
rect -3400 40100 -3000 40190
rect -1000 39100 800 40800
rect -3440 38960 -3000 39000
rect -3440 38700 -3400 38960
rect -3020 38910 -3000 38960
rect -3010 38700 -3000 38910
rect -3440 38690 -3390 38700
rect -3010 38690 -1600 38700
rect -3440 38660 -1600 38690
rect -3400 38600 -1600 38660
rect -3400 37600 -3300 38600
rect -1700 37600 -1600 38600
rect -3400 37500 -1600 37600
rect -4400 25710 -4000 25720
rect -4400 25490 -4390 25710
rect -4010 25490 -4000 25710
rect -4400 25450 -4370 25490
rect -4030 25450 -4000 25490
rect -4400 25430 -4000 25450
rect -3400 24900 -1600 37100
rect -6400 14300 -1600 24900
rect -1000 25500 -600 39100
rect 700 25500 800 39100
rect 26000 40800 30200 46000
rect 26000 38100 27800 40800
rect 29800 40480 30200 40500
rect 29800 40410 29820 40480
rect 29800 40190 29810 40410
rect 30180 40410 30200 40480
rect 30190 40190 30200 40410
rect 29800 40100 30200 40190
rect 29700 38960 30200 39000
rect 29700 38910 29820 38960
rect 30180 38910 30200 38960
rect 29700 38700 29810 38910
rect -1000 23200 800 25500
rect -1000 18500 -600 23200
rect 700 18500 800 23200
rect -1000 17800 800 18500
rect -1000 16600 -900 17800
rect 700 16600 800 17800
rect -1000 16500 800 16600
rect 26000 25500 26100 38100
rect 27400 25500 27800 38100
rect 28400 38690 29810 38700
rect 30190 38690 30200 38910
rect 28400 38600 30200 38690
rect 28400 37600 28500 38600
rect 30100 37600 30200 38600
rect 28400 37500 30200 37600
rect 26000 23200 27800 25500
rect 26000 16300 26100 23200
rect 27400 16300 27800 23200
rect 26000 15600 27800 16300
rect 26000 14400 26100 15600
rect 27700 14400 27800 15600
rect 26000 14300 27800 14400
rect 28400 24900 30200 37100
rect 30800 25710 31200 25720
rect 30800 25490 30810 25710
rect 31190 25490 31200 25710
rect 30800 25450 30830 25490
rect 31170 25450 31200 25490
rect 30800 25430 31200 25450
rect 28400 14300 33200 24900
rect -4400 14000 -4000 14010
rect -4400 13420 -4390 14000
rect -4010 13420 -4000 14000
rect -4400 13410 -4000 13420
rect -3400 13900 -1600 14300
rect -3400 13100 800 13900
rect 28400 13400 30200 14300
rect 30800 14000 31200 14010
rect 30800 13420 30810 14000
rect 31190 13420 31200 14000
rect 30800 13410 31200 13420
rect -4400 13090 800 13100
rect -4400 12510 -4390 13090
rect -4010 12510 800 13090
rect -4400 12500 800 12510
rect -3400 12100 800 12500
rect -3400 11100 -600 12100
rect -1000 8000 -600 11100
rect 700 10100 800 12100
rect 200 10000 800 10100
rect 26000 13100 30200 13400
rect 26000 13090 31200 13100
rect 26000 12510 30810 13090
rect 31190 12510 31200 13090
rect 26000 12500 31200 12510
rect 26000 12100 30200 12500
rect 26000 10100 26100 12100
rect 27400 11100 30200 12100
rect 26000 10000 26600 10100
rect 200 8000 300 10000
rect -1000 7900 300 8000
rect 26500 8000 26600 10000
rect 27400 8000 27800 11100
rect 26500 7900 27800 8000
rect -1000 7400 800 7900
rect -7200 3600 800 7400
rect 26000 7400 27800 7900
rect 26000 3600 34000 7400
rect -7200 1200 2800 3600
rect -7200 400 -7100 1200
rect 2600 400 2800 1200
rect 24000 1200 34000 3600
rect 24000 400 25600 1200
rect 33900 400 34000 1200
rect -7200 200 2800 400
rect 25500 200 34000 400
<< via4 >>
rect -3370 40210 -3030 40450
rect -3400 38910 -3020 38960
rect -3400 38700 -3390 38910
rect -3390 38700 -3020 38910
rect -3300 37600 -1700 38600
rect -4370 25490 -4030 25690
rect -4370 25450 -4030 25490
rect -600 25500 700 39100
rect 29830 40210 30170 40450
rect 29820 38910 30180 38960
rect 29820 38720 30180 38910
rect -600 18500 700 23200
rect -900 16600 700 17800
rect 26100 25500 27400 38100
rect 28500 37600 30100 38600
rect 26100 16300 27400 23200
rect 26100 14400 27700 15600
rect 30830 25490 31170 25690
rect 30830 25450 31170 25490
rect -4370 13440 -4030 13980
rect 30830 13440 31170 13980
rect -600 10100 700 12100
rect -600 8000 200 10100
rect 26100 10100 27400 12100
rect 26600 8000 27400 10100
rect -7100 400 2600 1200
rect 25600 400 33900 1200
<< mimcap2 >>
rect -3300 45800 700 45900
rect -3300 41000 -3200 45800
rect 600 41000 700 45800
rect -3300 40900 700 41000
rect 26100 45800 30100 45900
rect 26100 41000 26200 45800
rect 30000 41000 30100 45800
rect 26100 40900 30100 41000
rect -3300 36900 -1700 37000
rect -3300 26700 -3200 36900
rect -1800 26700 -1700 36900
rect -3300 26600 -1700 26700
rect 28500 36900 30100 37000
rect 28500 26700 28600 36900
rect 30000 26700 30100 36900
rect 28500 26600 30100 26700
rect -6300 24700 -1700 24800
rect -6300 14500 -6200 24700
rect -1800 14500 -1700 24700
rect -6300 14400 -1700 14500
rect 28500 24700 33100 24800
rect 28500 14500 28600 24700
rect 33000 14500 33100 24700
rect 28500 14400 33100 14500
rect -7100 7200 700 7300
rect -7100 2400 -7000 7200
rect 600 2400 700 7200
rect -7100 2300 700 2400
rect 26100 7200 33900 7300
rect 26100 2400 26200 7200
rect 33800 2400 33900 7200
rect 26100 2300 33900 2400
<< mimcap2contact >>
rect -3200 41000 600 45800
rect 26200 41000 30000 45800
rect -3200 26700 -1800 36900
rect 28600 26700 30000 36900
rect -6200 14500 -1800 24700
rect 28600 14500 33000 24700
rect -7000 2400 600 7200
rect 26200 2400 33800 7200
<< metal5 >>
rect 1300 47600 2800 48500
rect -600 46700 2800 47600
rect 24000 47600 25500 48500
rect 24000 46700 27400 47600
rect -600 46000 800 46700
rect -3400 45800 800 46000
rect -3400 41000 -3200 45800
rect 600 41000 800 45800
rect -3400 40800 800 41000
rect 26000 46000 27400 46700
rect 26000 45800 30200 46000
rect 26000 41000 26200 45800
rect 30000 41000 30200 45800
rect 26000 40800 30200 41000
rect -3400 40450 -3000 40800
rect -3400 40210 -3370 40450
rect -3030 40210 -3000 40450
rect -3400 40100 -3000 40210
rect 29800 40450 30200 40800
rect 29800 40210 29830 40450
rect 30170 40210 30200 40450
rect -2400 40100 1200 40200
rect 29800 40100 30200 40210
rect -2500 40000 1200 40100
rect -2600 39900 1200 40000
rect -2700 39800 1200 39900
rect -2800 39700 1200 39800
rect -2900 39600 -1400 39700
rect -3000 39500 -1500 39600
rect -3000 39000 -1600 39500
rect 25400 39200 29200 39300
rect -3440 38960 -1600 39000
rect -3440 38700 -3400 38960
rect -3020 38700 -1600 38960
rect -3440 38660 -1600 38700
rect -3400 38600 -1600 38660
rect -3400 37600 -3300 38600
rect -1700 37600 -1600 38600
rect -3400 36900 -1600 37600
rect -3400 26700 -3200 36900
rect -1800 26700 -1600 36900
rect -3400 26500 -1600 26700
rect -700 39100 800 39200
rect -4400 25690 -4000 25720
rect -4400 25450 -4370 25690
rect -4030 25450 -4000 25690
rect -4400 24900 -4000 25450
rect -700 25500 -600 39100
rect 700 25500 800 39100
rect 25400 39100 29300 39200
rect 25400 39000 29400 39100
rect 25400 38960 30220 39000
rect 25400 38800 29820 38960
rect 28200 38720 29820 38800
rect 30180 38720 30220 38960
rect 28200 38700 30220 38720
rect 28300 38660 30220 38700
rect 28300 38600 30200 38660
rect -700 25400 800 25500
rect 26000 38100 27500 38200
rect 26000 25500 26100 38100
rect 27400 25500 27500 38100
rect 28400 37600 28500 38600
rect 30100 37600 30200 38600
rect 28400 36900 30200 37600
rect 28400 26700 28600 36900
rect 30000 26700 30200 36900
rect 28400 26500 30200 26700
rect 26000 25400 27500 25500
rect 30800 25690 31200 25720
rect 30800 25450 30830 25690
rect 31170 25450 31200 25690
rect 30800 24900 31200 25450
rect -6400 24700 1200 24900
rect 25280 24700 33200 24900
rect -6400 14500 -6200 24700
rect -1800 24000 2100 24700
rect 24700 24000 28600 24700
rect -1800 23800 1200 24000
rect 25320 23800 28600 24000
rect -1800 14500 -1600 23800
rect -700 23200 800 23300
rect -700 18500 -600 23200
rect 700 18500 800 23200
rect -700 18400 800 18500
rect 26000 23200 27500 23300
rect -6400 14300 -1600 14500
rect -1200 17800 1300 17900
rect -1200 16600 -900 17800
rect 700 16600 1300 17800
rect -1200 16500 1300 16600
rect -4400 13980 -4000 14300
rect -4400 13440 -4370 13980
rect -4030 13440 -4000 13980
rect -1200 13900 0 16500
rect 26000 16300 26100 23200
rect 27400 16300 27500 23200
rect 26000 16200 27500 16300
rect 25500 15600 28000 15700
rect 25500 14400 26100 15600
rect 27700 14400 28000 15600
rect 25500 14300 28000 14400
rect 28400 14500 28600 23800
rect 33000 14500 33200 24700
rect 28400 14300 33200 14500
rect -4400 13410 -4000 13440
rect -3400 12600 0 13900
rect 26800 13900 28000 14300
rect 30800 13980 31200 14300
rect 26800 12600 30200 13900
rect 30800 13440 30830 13980
rect 31170 13440 31200 13980
rect 30800 13410 31200 13440
rect -3400 7400 -1600 12600
rect -700 12100 800 12200
rect -700 8000 -600 12100
rect 700 10100 800 12100
rect 200 10000 800 10100
rect 26000 12100 27500 12200
rect 26000 10100 26100 12100
rect 26000 10000 26600 10100
rect 200 8000 300 10000
rect 700 9100 1200 9600
rect 25400 8200 25900 8700
rect -700 7900 300 8000
rect 26500 8000 26600 10000
rect 27400 8000 27500 12100
rect 26500 7900 27500 8000
rect 28400 7400 30200 12600
rect -7200 7200 800 7400
rect -7200 2400 -7000 7200
rect 600 2400 800 7200
rect -7200 2200 800 2400
rect 26000 7200 34000 7400
rect 26000 2400 26200 7200
rect 33800 2400 34000 7200
rect 26000 2200 34000 2400
rect -7200 1200 1400 1400
rect 25400 1200 34000 1400
rect -7200 400 -7100 1200
rect 24200 400 25600 1200
rect 33900 400 34000 1200
rect -7200 200 2800 400
rect 1300 0 2800 200
rect 24000 200 34000 400
rect 24000 0 25500 200
use cascode_1  cascode_1_0
timestamp 1664506494
transform 1 0 14700 0 1 -3700
box -14700 3700 10800 52200
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660275339
transform 1 0 12900 0 1 33600
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_1
timestamp 1660275339
transform 1 0 6900 0 1 33600
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_2
timestamp 1660275339
transform 1 0 6400 0 1 33600
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_3
timestamp 1660275339
transform 1 0 6400 0 1 32100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_4
timestamp 1660275339
transform 1 0 6900 0 1 32100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_5
timestamp 1660275339
transform 1 0 6400 0 1 31600
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_6
timestamp 1660275339
transform 1 0 6900 0 1 31600
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_7
timestamp 1660275339
transform 1 0 19400 0 1 33600
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_8
timestamp 1660275339
transform 1 0 19400 0 1 32100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_9
timestamp 1660275339
transform 1 0 19400 0 1 31600
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_10
timestamp 1660275339
transform 1 0 12900 0 1 32100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_11
timestamp 1660275339
transform 1 0 12900 0 1 3100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_12
timestamp 1660275339
transform 1 0 19400 0 1 3100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_13
timestamp 1660275339
transform 1 0 6400 0 1 47100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_14
timestamp 1660275339
transform 1 0 6900 0 1 47100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_15
timestamp 1660275339
transform 1 0 12900 0 1 47100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_16
timestamp 1660275339
transform 1 0 13400 0 1 47100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_17
timestamp 1660275339
transform 1 0 18900 0 1 47100
box 100 -1100 600 -600
use hash_m1m2_W2p5L2p5#0  hash_m1m2_W2p5L2p5_18
timestamp 1660275339
transform 1 0 19400 0 1 47100
box 100 -1100 600 -600
use hash_m1m2_W5L5  hash_m1m2_W5L5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660789662
transform 1 0 1500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_1
timestamp 1660789662
transform 1 0 2500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_2
timestamp 1660789662
transform 1 0 3500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_3
timestamp 1660789662
transform 1 0 4500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_4
timestamp 1660789662
transform 1 0 5500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_5
timestamp 1660789662
transform 1 0 6500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_6
timestamp 1660789662
transform 1 0 7500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_7
timestamp 1660789662
transform 1 0 8500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_8
timestamp 1660789662
transform 1 0 9500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_9
timestamp 1660789662
transform 1 0 10500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_10
timestamp 1660789662
transform 1 0 11500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_11
timestamp 1660789662
transform 1 0 12500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_12
timestamp 1660789662
transform 1 0 13500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_13
timestamp 1660789662
transform 1 0 14500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_14
timestamp 1660789662
transform 1 0 15500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_15
timestamp 1660789662
transform 1 0 16500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_16
timestamp 1660789662
transform 1 0 17500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_17
timestamp 1660789662
transform 1 0 18500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_18
timestamp 1660789662
transform 1 0 19500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_19
timestamp 1660789662
transform 1 0 20500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_20
timestamp 1660789662
transform 1 0 21500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_21
timestamp 1660789662
transform 1 0 22500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_22
timestamp 1660789662
transform 1 0 23500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_23
timestamp 1660789662
transform 1 0 24500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_24
timestamp 1660789662
transform 1 0 500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_25
timestamp 1660789662
transform 1 0 0 0 1 4700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_26
timestamp 1660789662
transform 1 0 0 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_27
timestamp 1660789662
transform 1 0 0 0 1 3700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_28
timestamp 1660789662
transform 1 0 0 0 1 5700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_29
timestamp 1660789662
transform 1 0 0 0 1 6700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_30
timestamp 1660789662
transform 1 0 0 0 1 7700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_31
timestamp 1660789662
transform 1 0 0 0 1 8700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_32
timestamp 1660789662
transform 1 0 0 0 1 9700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_33
timestamp 1660789662
transform 1 0 0 0 1 10700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_34
timestamp 1660789662
transform 1 0 0 0 1 11700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_35
timestamp 1660789662
transform 1 0 0 0 1 12700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_36
timestamp 1660789662
transform 1 0 0 0 1 13700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_37
timestamp 1660789662
transform 1 0 0 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_38
timestamp 1660789662
transform 1 0 0 0 1 15700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_39
timestamp 1660789662
transform 1 0 0 0 1 16700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_40
timestamp 1660789662
transform 1 0 0 0 1 20700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_41
timestamp 1660789662
transform 1 0 0 0 1 19700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_42
timestamp 1660789662
transform 1 0 0 0 1 18700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_43
timestamp 1660789662
transform 1 0 0 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_44
timestamp 1660789662
transform 1 0 0 0 1 24700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_45
timestamp 1660789662
transform 1 0 0 0 1 23700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_46
timestamp 1660789662
transform 1 0 0 0 1 22700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_47
timestamp 1660789662
transform 1 0 0 0 1 21700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_48
timestamp 1660789662
transform 1 0 0 0 1 28700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_49
timestamp 1660789662
transform 1 0 0 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_50
timestamp 1660789662
transform 1 0 0 0 1 26700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_51
timestamp 1660789662
transform 1 0 0 0 1 25700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_52
timestamp 1660789662
transform 1 0 0 0 1 32700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_53
timestamp 1660789662
transform 1 0 0 0 1 31700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_54
timestamp 1660789662
transform 1 0 0 0 1 30700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_55
timestamp 1660789662
transform 1 0 0 0 1 29700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_56
timestamp 1660789662
transform 1 0 0 0 1 36700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_57
timestamp 1660789662
transform 1 0 0 0 1 35700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_58
timestamp 1660789662
transform 1 0 0 0 1 34700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_59
timestamp 1660789662
transform 1 0 0 0 1 33700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_60
timestamp 1660789662
transform 1 0 0 0 1 40700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_61
timestamp 1660789662
transform 1 0 0 0 1 39700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_62
timestamp 1660789662
transform 1 0 0 0 1 38700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_63
timestamp 1660789662
transform 1 0 0 0 1 37700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_64
timestamp 1660789662
transform 1 0 0 0 1 44700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_65
timestamp 1660789662
transform 1 0 0 0 1 43700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_66
timestamp 1660789662
transform 1 0 0 0 1 42700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_67
timestamp 1660789662
transform 1 0 0 0 1 41700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_68
timestamp 1660789662
transform 1 0 0 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_69
timestamp 1660789662
transform 1 0 0 0 1 47700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_70
timestamp 1660789662
transform 1 0 0 0 1 46700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_71
timestamp 1660789662
transform 1 0 0 0 1 45700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_72
timestamp 1660789662
transform 1 0 25500 0 1 5700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_73
timestamp 1660789662
transform 1 0 25500 0 1 4700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_74
timestamp 1660789662
transform 1 0 25500 0 1 3700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_75
timestamp 1660789662
transform 1 0 25500 0 1 2700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_76
timestamp 1660789662
transform 1 0 25500 0 1 9700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_77
timestamp 1660789662
transform 1 0 25500 0 1 8700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_78
timestamp 1660789662
transform 1 0 25500 0 1 7700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_79
timestamp 1660789662
transform 1 0 25500 0 1 6700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_80
timestamp 1660789662
transform 1 0 25500 0 1 13700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_81
timestamp 1660789662
transform 1 0 25500 0 1 12700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_82
timestamp 1660789662
transform 1 0 25500 0 1 11700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_83
timestamp 1660789662
transform 1 0 25500 0 1 10700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_84
timestamp 1660789662
transform 1 0 25500 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_85
timestamp 1660789662
transform 1 0 25500 0 1 16700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_86
timestamp 1660789662
transform 1 0 25500 0 1 15700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_87
timestamp 1660789662
transform 1 0 25500 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_88
timestamp 1660789662
transform 1 0 25500 0 1 21700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_89
timestamp 1660789662
transform 1 0 25500 0 1 20700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_90
timestamp 1660789662
transform 1 0 25500 0 1 19700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_91
timestamp 1660789662
transform 1 0 25500 0 1 18700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_92
timestamp 1660789662
transform 1 0 25500 0 1 25700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_93
timestamp 1660789662
transform 1 0 25500 0 1 24700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_94
timestamp 1660789662
transform 1 0 25500 0 1 23700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_95
timestamp 1660789662
transform 1 0 25500 0 1 22700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_96
timestamp 1660789662
transform 1 0 25500 0 1 29700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_97
timestamp 1660789662
transform 1 0 25500 0 1 28700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_98
timestamp 1660789662
transform 1 0 25500 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_99
timestamp 1660789662
transform 1 0 25500 0 1 26700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_100
timestamp 1660789662
transform 1 0 25500 0 1 33700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_101
timestamp 1660789662
transform 1 0 25500 0 1 32700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_102
timestamp 1660789662
transform 1 0 25500 0 1 31700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_103
timestamp 1660789662
transform 1 0 25500 0 1 30700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_104
timestamp 1660789662
transform 1 0 25500 0 1 37700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_105
timestamp 1660789662
transform 1 0 25500 0 1 36700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_106
timestamp 1660789662
transform 1 0 25500 0 1 35700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_107
timestamp 1660789662
transform 1 0 25500 0 1 34700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_108
timestamp 1660789662
transform 1 0 25500 0 1 41700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_109
timestamp 1660789662
transform 1 0 25500 0 1 40700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_110
timestamp 1660789662
transform 1 0 25500 0 1 39700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_111
timestamp 1660789662
transform 1 0 25500 0 1 38700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_112
timestamp 1660789662
transform 1 0 25500 0 1 45700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_113
timestamp 1660789662
transform 1 0 25500 0 1 44700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_114
timestamp 1660789662
transform 1 0 25500 0 1 43700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_115
timestamp 1660789662
transform 1 0 25500 0 1 42700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_116
timestamp 1660789662
transform 1 0 25500 0 1 46700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_117
timestamp 1660789662
transform 1 0 25500 0 1 47700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_118
timestamp 1660789662
transform 1 0 1000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_119
timestamp 1660789662
transform 1 0 500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_120
timestamp 1660789662
transform 1 0 1500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_121
timestamp 1660789662
transform 1 0 2500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_122
timestamp 1660789662
transform 1 0 3500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_123
timestamp 1660789662
transform 1 0 4500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_124
timestamp 1660789662
transform 1 0 5500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_125
timestamp 1660789662
transform 1 0 6500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_126
timestamp 1660789662
transform 1 0 10500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_127
timestamp 1660789662
transform 1 0 8500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_128
timestamp 1660789662
transform 1 0 9500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_129
timestamp 1660789662
transform 1 0 7500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_130
timestamp 1660789662
transform 1 0 14500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_131
timestamp 1660789662
transform 1 0 12500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_132
timestamp 1660789662
transform 1 0 13500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_133
timestamp 1660789662
transform 1 0 11500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_134
timestamp 1660789662
transform 1 0 18500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_135
timestamp 1660789662
transform 1 0 16500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_136
timestamp 1660789662
transform 1 0 17500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_137
timestamp 1660789662
transform 1 0 15500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_138
timestamp 1660789662
transform 1 0 22500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_139
timestamp 1660789662
transform 1 0 20500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_140
timestamp 1660789662
transform 1 0 21500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_141
timestamp 1660789662
transform 1 0 19500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_142
timestamp 1660789662
transform 1 0 2000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_143
timestamp 1660789662
transform 1 0 24500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_144
timestamp 1660789662
transform 1 0 25500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_145
timestamp 1660789662
transform 1 0 23500 0 1 48200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_146
timestamp 1660789662
transform 1 0 3000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_147
timestamp 1660789662
transform 1 0 6000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_148
timestamp 1660789662
transform 1 0 5000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_149
timestamp 1660789662
transform 1 0 4000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_150
timestamp 1660789662
transform 1 0 9000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_151
timestamp 1660789662
transform 1 0 8000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_152
timestamp 1660789662
transform 1 0 7000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_153
timestamp 1660789662
transform 1 0 12000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_154
timestamp 1660789662
transform 1 0 11000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_155
timestamp 1660789662
transform 1 0 10000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_156
timestamp 1660789662
transform 1 0 15000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_157
timestamp 1660789662
transform 1 0 14000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_158
timestamp 1660789662
transform 1 0 13000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_159
timestamp 1660789662
transform 1 0 18000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_160
timestamp 1660789662
transform 1 0 17000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_161
timestamp 1660789662
transform 1 0 16000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_162
timestamp 1660789662
transform 1 0 21000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_163
timestamp 1660789662
transform 1 0 20000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_164
timestamp 1660789662
transform 1 0 19000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_165
timestamp 1660789662
transform 1 0 24000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_166
timestamp 1660789662
transform 1 0 23000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_167
timestamp 1660789662
transform 1 0 22000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_168
timestamp 1660789662
transform 1 0 25000 0 1 33200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_169
timestamp 1660789662
transform 1 0 3000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_170
timestamp 1660789662
transform 1 0 2000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_171
timestamp 1660789662
transform 1 0 1000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_172
timestamp 1660789662
transform 1 0 6000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_173
timestamp 1660789662
transform 1 0 5000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_174
timestamp 1660789662
transform 1 0 4000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_175
timestamp 1660789662
transform 1 0 9000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_176
timestamp 1660789662
transform 1 0 8000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_177
timestamp 1660789662
transform 1 0 7000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_178
timestamp 1660789662
transform 1 0 12000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_179
timestamp 1660789662
transform 1 0 11000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_180
timestamp 1660789662
transform 1 0 10000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_181
timestamp 1660789662
transform 1 0 15000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_182
timestamp 1660789662
transform 1 0 14000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_183
timestamp 1660789662
transform 1 0 13000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_184
timestamp 1660789662
transform 1 0 18000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_185
timestamp 1660789662
transform 1 0 17000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_186
timestamp 1660789662
transform 1 0 16000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_187
timestamp 1660789662
transform 1 0 21000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_188
timestamp 1660789662
transform 1 0 20000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_189
timestamp 1660789662
transform 1 0 19000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_190
timestamp 1660789662
transform 1 0 24000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_191
timestamp 1660789662
transform 1 0 23000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_192
timestamp 1660789662
transform 1 0 22000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_193
timestamp 1660789662
transform 1 0 25000 0 1 17700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_194
timestamp 1660789662
transform 1 0 19000 0 1 18200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_195
timestamp 1660789662
transform 1 0 13000 0 1 18200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_196
timestamp 1660789662
transform 1 0 6500 0 1 18200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_197
timestamp 1660789662
transform 1 0 6500 0 1 17200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_198
timestamp 1660789662
transform 1 0 13000 0 1 17200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_199
timestamp 1660789662
transform 1 0 19000 0 1 17200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_200
timestamp 1660789662
transform 1 0 6500 0 1 3200
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_201
timestamp 1660789662
transform 1 0 -1000 0 1 40700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_202
timestamp 1660789662
transform 1 0 -2000 0 1 40700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_203
timestamp 1660789662
transform 1 0 -3000 0 1 40700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_204
timestamp 1660789662
transform 1 0 -1000 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_205
timestamp 1660789662
transform 1 0 -2000 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_206
timestamp 1660789662
transform 1 0 -3000 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_207
timestamp 1660789662
transform 1 0 -4000 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_208
timestamp 1660789662
transform 1 0 -1000 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_209
timestamp 1660789662
transform 1 0 -2000 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_210
timestamp 1660789662
transform 1 0 -3000 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_211
timestamp 1660789662
transform 1 0 -4000 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_212
timestamp 1660789662
transform 1 0 26500 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_213
timestamp 1660789662
transform 1 0 27500 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_214
timestamp 1660789662
transform 1 0 28500 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_215
timestamp 1660789662
transform 1 0 29500 0 1 14700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_216
timestamp 1660789662
transform 1 0 26500 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_217
timestamp 1660789662
transform 1 0 27500 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_218
timestamp 1660789662
transform 1 0 28500 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_219
timestamp 1660789662
transform 1 0 29500 0 1 27700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_220
timestamp 1660789662
transform 1 0 26500 0 1 40700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_221
timestamp 1660789662
transform 1 0 27500 0 1 40700
box 0 -1700 1000 -700
use hash_m1m2_W5L5  hash_m1m2_W5L5_222
timestamp 1660789662
transform 1 0 28500 0 1 40700
box 0 -1700 1000 -700
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_1
timestamp 1664814488
transform 1 0 -4201 0 1 26369
box -199 -889 199 889
use sky130_fd_pr__res_generic_po_63AFTY  sky130_fd_pr__res_generic_po_63AFTY_3
timestamp 1664814488
transform 1 0 -3201 0 1 39569
box -199 -889 199 889
use sky130_fd_pr__res_high_po_0p35_FFWWQH  sky130_fd_pr__res_high_po_0p35_FFWWQH_0
timestamp 1664805031
transform 1 0 -4199 0 1 13258
box -201 -758 201 758
<< labels >>
rlabel metal5 1300 48100 2800 48500 1 VDN
rlabel metal5 900 39700 1200 40200 1 VGN
rlabel metal3 800 31000 1000 31800 1 N2
rlabel metal5 700 9100 1000 9600 1 VINN
rlabel metal5 1300 0 2800 400 1 VSS
rlabel metal5 800 23800 1000 24800 1 MIDGATE
rlabel metal5 24000 48300 25500 48500 1 VDP
rlabel metal3 25600 31100 25900 31700 1 P2
rlabel metal5 24000 0 25500 200 1 VSSH
rlabel metal5 25700 38800 25900 39300 1 VGP
rlabel metal5 25700 8200 25900 8700 1 VINP
rlabel metal1 -3920 13900 -3540 14000 1 SUB
rlabel metal5 900 16500 1200 17900 1 N
rlabel metal5 25600 14300 25900 15700 1 P
<< end >>
