magic
tech sky130A
timestamp 1664716557
<< metal4 >>
rect -300 7850 400 7900
rect -300 7350 -250 7850
rect 350 7350 400 7850
rect -300 7300 400 7350
rect -1700 7100 -800 7300
rect -500 1800 400 7300
rect 13000 7800 13900 7850
rect 13000 7350 13050 7800
rect 13850 7350 13900 7800
rect 13000 1800 13900 7350
<< via4 >>
rect -250 7350 350 7850
rect 13050 7350 13850 7800
<< mimcap2 >>
rect -450 7000 350 7050
rect -450 1900 -400 7000
rect 300 1900 350 7000
rect -450 1850 350 1900
rect 13050 7000 13850 7050
rect 13050 1900 13100 7000
rect 13800 1900 13850 7000
rect 13050 1850 13850 1900
<< mimcap2contact >>
rect -400 1900 300 7000
rect 13100 1900 13800 7000
<< metal5 >>
rect -200 9450 150 12450
rect -1700 9200 150 9450
rect -1700 7300 -800 9200
rect -300 8250 650 8950
rect -300 7850 400 8250
rect -300 7350 -250 7850
rect 350 7350 400 7850
rect -300 7300 400 7350
rect 12750 7800 13900 7850
rect 12750 7350 13050 7800
rect 13850 7350 13900 7800
rect 12750 7300 13900 7350
rect -3050 1800 -800 7100
rect -500 7000 400 7100
rect -500 1900 -400 7000
rect 300 1900 400 7000
rect -500 1800 400 1900
rect 13000 7000 13900 7100
rect 13000 1900 13100 7000
rect 13800 1900 13900 7000
rect 13000 1800 13900 1900
rect 14200 1800 15100 7100
rect -1700 1100 700 1800
rect 12000 1100 15100 1800
rect 12000 850 12750 1100
use cascode_1  cascode_1_0
timestamp 1664506494
transform 1 0 7350 0 1 -1850
box -7350 1850 5400 26100
<< end >>
