magic
tech sky130A
timestamp 1664247701
<< metal2 >>
rect 3250 3050 3900 3250
rect 6400 3100 7050 3300
rect 9550 3050 10200 3250
rect 3250 2750 3900 2950
rect 6400 2800 7050 3000
rect 9550 2750 10200 2950
rect 3250 2450 3900 2650
rect 6400 2500 7050 2700
rect 9550 2450 10200 2650
rect 3250 2150 3900 2350
rect 6400 2200 7050 2400
rect 9550 2150 10200 2350
rect 3250 1850 3900 2050
rect 6400 1900 7050 2100
rect 9550 1850 10200 2050
rect 3250 1550 3900 1750
rect 6400 1600 7050 1800
rect 9550 1550 10200 1750
rect 3250 1250 3900 1450
rect 6400 1300 7050 1500
rect 9550 1250 10200 1450
rect 3250 950 3900 1150
rect 6400 1000 7050 1200
rect 9550 950 10200 1150
rect 3250 650 3900 850
rect 6400 700 7050 900
rect 9550 650 10200 850
rect 3250 350 3900 550
rect 6400 400 7050 600
rect 9550 350 10200 550
rect 3250 50 3900 250
rect 6400 100 7050 300
rect 3450 -250 3700 50
rect 6600 -250 6850 100
rect 9550 50 10200 250
rect 9750 -250 10000 50
rect 3250 -450 3900 -250
rect 6400 -450 7050 -250
rect 9550 -450 10200 -250
rect 3250 -750 3900 -550
rect 6400 -750 7050 -550
rect 9550 -750 10200 -550
rect 3250 -1050 3900 -850
rect 6400 -1050 7050 -850
rect 9550 -1050 10200 -850
rect 3250 -1350 3900 -1150
rect 6400 -1350 7050 -1150
rect 9550 -1350 10200 -1150
rect 3250 -1650 3900 -1450
rect 6400 -1650 7050 -1450
rect 9550 -1650 10200 -1450
rect 3250 -1950 3900 -1750
rect 6400 -1950 7050 -1750
rect 9550 -1950 10200 -1750
rect 3250 -2250 3900 -2050
rect 6400 -2250 7050 -2050
rect 9550 -2250 10200 -2050
rect 3250 -2550 3900 -2350
rect 6400 -2550 7050 -2350
rect 9550 -2550 10200 -2350
rect 3250 -2850 3900 -2650
rect 6400 -2850 7050 -2650
rect 9550 -2850 10200 -2650
rect 3250 -3150 3900 -2950
rect 6400 -3150 7050 -2950
rect 9550 -3150 10200 -2950
rect 3250 -3450 3900 -3250
rect 6400 -3450 7050 -3250
rect 9550 -3450 10200 -3250
<< metal3 >>
rect 700 2850 2550 2900
rect 700 1950 750 2850
rect 1400 1950 2550 2850
rect 700 1900 2550 1950
rect 3850 2850 4600 2900
rect 3850 1950 3900 2850
rect 4500 1950 4600 2850
rect 3850 1900 4600 1950
rect 7000 2850 7750 2900
rect 7000 1950 7050 2850
rect 7700 1950 7750 2850
rect 7000 1900 7750 1950
rect 10150 2850 10900 2900
rect 10150 1950 10200 2850
rect 10800 1950 10900 2850
rect 10150 1900 10900 1950
rect 700 1350 2550 1400
rect 700 450 750 1350
rect 1400 450 2550 1350
rect 700 400 2550 450
rect 5750 1350 6500 1400
rect 5750 450 5800 1350
rect 6450 450 6500 1350
rect 5750 400 6500 450
rect 7000 1350 7750 1400
rect 7000 450 7050 1350
rect 7700 450 7750 1350
rect 7000 400 7750 450
rect 12050 1350 12800 1400
rect 12050 450 12100 1350
rect 12750 450 12800 1350
rect 12050 400 12800 450
rect 1550 200 2500 250
rect 1550 150 1650 200
rect 700 50 1650 150
rect 2400 150 2500 200
rect 7850 200 8800 250
rect 7850 150 7950 200
rect 2400 90 3700 150
rect 2400 50 3510 90
rect 700 10 3510 50
rect 3690 10 3700 90
rect 700 0 3700 10
rect 3800 90 6850 150
rect 3800 10 6660 90
rect 6840 10 6850 90
rect 3800 0 6850 10
rect 6950 50 7950 150
rect 8700 150 8800 200
rect 8700 90 10000 150
rect 8700 50 9810 90
rect 6950 10 9810 50
rect 9990 10 10000 90
rect 6950 0 10000 10
rect 10100 0 12700 150
rect 3800 -100 3950 0
rect 4700 -50 6000 0
rect 6950 -50 7050 0
rect 10100 -50 10250 0
rect 11000 -50 12300 0
rect 3250 -200 3950 -100
rect 6400 -150 7050 -50
rect 9550 -150 10250 -50
rect 1550 -250 2500 -200
rect 3250 -250 3400 -200
rect 4700 -250 6000 -200
rect 6400 -250 6550 -150
rect 7850 -250 8800 -200
rect 9550 -250 9700 -150
rect 11000 -250 12300 -200
rect 700 -400 1650 -250
rect 2400 -400 3400 -250
rect 3500 -260 6550 -250
rect 3500 -340 3510 -260
rect 3690 -340 6550 -260
rect 3500 -400 6550 -340
rect 6650 -260 7950 -250
rect 6650 -340 6660 -260
rect 6840 -340 7950 -260
rect 6650 -400 7950 -340
rect 8700 -400 9700 -250
rect 9800 -260 12700 -250
rect 9800 -340 9810 -260
rect 9990 -340 12700 -260
rect 9800 -400 12700 -340
rect 1550 -450 2500 -400
rect 7850 -450 8800 -400
rect 1650 -650 2400 -600
rect 1650 -1550 1700 -650
rect 2350 -1550 2400 -650
rect 1650 -1600 2400 -1550
rect 3850 -650 4600 -600
rect 3850 -1550 3900 -650
rect 4550 -1550 4600 -650
rect 3850 -1600 4600 -1550
rect 7950 -650 8700 -600
rect 7950 -1550 8000 -650
rect 8650 -1550 8700 -650
rect 7950 -1600 8700 -1550
rect 10150 -650 10900 -600
rect 10150 -1550 10200 -650
rect 10850 -1550 10900 -650
rect 10150 -1600 10900 -1550
rect 800 -2150 3350 -2100
rect 800 -3050 2650 -2150
rect 3300 -3050 3350 -2150
rect 800 -3100 3350 -3050
rect 3950 -2150 6400 -2100
rect 3950 -3050 4850 -2150
rect 5500 -3050 6400 -2150
rect 3950 -3100 6400 -3050
rect 8900 -2150 9650 -2100
rect 8900 -3050 8950 -2150
rect 9600 -3050 9650 -2150
rect 8900 -3100 9650 -3050
rect 10150 -2150 12800 -2100
rect 10150 -3050 11150 -2150
rect 11800 -3050 12800 -2150
rect 10150 -3100 12800 -3050
<< via3 >>
rect 750 1950 1400 2850
rect 3900 1950 4500 2850
rect 7050 1950 7700 2850
rect 10200 1950 10800 2850
rect 750 450 1400 1350
rect 5800 450 6450 1350
rect 7050 450 7700 1350
rect 12100 450 12750 1350
rect 1650 50 2400 200
rect 3510 10 3690 90
rect 6660 10 6840 90
rect 7950 50 8700 200
rect 9810 10 9990 90
rect 1650 -400 2400 -250
rect 3510 -340 3690 -260
rect 6660 -340 6840 -260
rect 7950 -400 8700 -250
rect 9810 -340 9990 -260
rect 1700 -1550 2350 -650
rect 3900 -1550 4550 -650
rect 8000 -1550 8650 -650
rect 10200 -1550 10850 -650
rect 2650 -3050 3300 -2150
rect 4850 -3050 5500 -2150
rect 8950 -3050 9600 -2150
rect 11150 -3050 11800 -2150
<< metal4 >>
rect 2600 5550 3350 5600
rect 2600 4750 2650 5550
rect 3300 4750 3350 5550
rect 700 4000 1450 4100
rect 700 3300 800 4000
rect 1400 3300 1450 4000
rect 700 2850 1450 3300
rect 700 1950 750 2850
rect 1400 1950 1450 2850
rect 700 1900 1450 1950
rect 700 1350 1450 1400
rect 700 450 750 1350
rect 1400 450 1450 1350
rect 700 -4950 1450 450
rect 1600 200 2450 250
rect 1600 50 1650 200
rect 2400 50 2450 200
rect 1600 0 2450 50
rect 1600 -250 2450 -200
rect 1600 -400 1650 -250
rect 2400 -400 2450 -250
rect 1600 -450 2450 -400
rect 1650 -650 2400 -600
rect 1650 -1550 1700 -650
rect 2350 -1550 2400 -650
rect 1650 -3450 2400 -1550
rect 2600 -2150 3350 4750
rect 3850 5550 4600 5600
rect 3850 4750 3900 5550
rect 4550 4750 4600 5550
rect 3850 2850 4600 4750
rect 8900 5550 9650 5600
rect 8900 4750 8950 5550
rect 9600 4750 9650 5550
rect 3850 1950 3900 2850
rect 4500 1950 4600 2850
rect 3850 1900 4600 1950
rect 4800 4050 5550 4100
rect 4800 3250 4900 4050
rect 5500 3250 5550 4050
rect 3500 90 3700 100
rect 3500 10 3510 90
rect 3690 10 3700 90
rect 3500 -260 3700 10
rect 3500 -340 3510 -260
rect 3690 -340 3700 -260
rect 3500 -350 3700 -340
rect 2600 -3050 2650 -2150
rect 3300 -3050 3350 -2150
rect 2600 -3100 3350 -3050
rect 3850 -650 4600 -600
rect 3850 -1550 3900 -650
rect 4550 -1550 4600 -650
rect 1650 -4250 1700 -3450
rect 2350 -4250 2400 -3450
rect 1650 -4300 2400 -4250
rect 700 -5750 750 -4950
rect 1400 -5750 1450 -4950
rect 700 -5800 1450 -5750
rect 3850 -4950 4600 -1550
rect 4800 -2150 5550 3250
rect 7000 4000 7750 4100
rect 7000 3300 7100 4000
rect 7700 3300 7750 4000
rect 7000 2850 7750 3300
rect 7000 1950 7050 2850
rect 7700 1950 7750 2850
rect 7000 1900 7750 1950
rect 4800 -3050 4850 -2150
rect 5500 -3050 5550 -2150
rect 4800 -3100 5550 -3050
rect 5750 1350 6500 1400
rect 5750 450 5800 1350
rect 6450 450 6500 1350
rect 5750 -3450 6500 450
rect 7000 1350 7750 1400
rect 7000 450 7050 1350
rect 7700 450 7750 1350
rect 6650 90 6850 100
rect 6650 10 6660 90
rect 6840 10 6850 90
rect 6650 -260 6850 10
rect 6650 -340 6660 -260
rect 6840 -340 6850 -260
rect 6650 -350 6850 -340
rect 5750 -4250 5800 -3450
rect 6450 -4250 6500 -3450
rect 5750 -4300 6500 -4250
rect 7000 -4950 7750 450
rect 7900 200 8750 250
rect 7900 50 7950 200
rect 8700 50 8750 200
rect 7900 0 8750 50
rect 7900 -250 8750 -200
rect 7900 -400 7950 -250
rect 8700 -400 8750 -250
rect 7900 -450 8750 -400
rect 7950 -650 8700 -600
rect 7950 -1550 8000 -650
rect 8650 -1550 8700 -650
rect 7950 -3450 8700 -1550
rect 8900 -2150 9650 4750
rect 10150 5550 10900 5600
rect 10150 4750 10200 5550
rect 10850 4750 10900 5550
rect 10150 4100 10900 4750
rect 10150 3300 10950 4100
rect 11100 4050 11850 4100
rect 10150 2850 10900 3300
rect 10150 1950 10200 2850
rect 10800 1950 10900 2850
rect 10150 1900 10900 1950
rect 11100 3250 11200 4050
rect 11800 3250 11850 4050
rect 9800 90 10000 100
rect 9800 10 9810 90
rect 9990 10 10000 90
rect 9800 -260 10000 10
rect 9800 -340 9810 -260
rect 9990 -340 10000 -260
rect 9800 -350 10000 -340
rect 8900 -3050 8950 -2150
rect 9600 -3050 9650 -2150
rect 8900 -3100 9650 -3050
rect 10150 -650 10900 -600
rect 10150 -1550 10200 -650
rect 10850 -1550 10900 -650
rect 7950 -4250 8000 -3450
rect 8650 -4250 8700 -3450
rect 7950 -4300 8700 -4250
rect 3850 -5750 3900 -4950
rect 4550 -5750 4600 -4950
rect 3850 -5800 4600 -5750
rect 5750 -5750 5800 -4950
rect 6400 -5750 6500 -4950
rect 5750 -5800 6500 -5750
rect 7000 -5750 7050 -4950
rect 7700 -5750 7750 -4950
rect 7000 -5800 7750 -5750
rect 10150 -4950 10900 -1550
rect 11100 -2150 11850 3250
rect 11100 -3050 11150 -2150
rect 11800 -3050 11850 -2150
rect 11100 -3100 11850 -3050
rect 12050 1350 12800 1400
rect 12050 450 12100 1350
rect 12750 450 12800 1350
rect 12050 -3450 12800 450
rect 12050 -4250 12100 -3450
rect 12750 -4250 12800 -3450
rect 12050 -4300 12800 -4250
rect 10150 -5750 10200 -4950
rect 10850 -5750 10900 -4950
rect 10150 -5800 10900 -5750
<< via4 >>
rect 2650 4750 3300 5550
rect 800 3300 1400 4000
rect 1650 50 2400 200
rect 1650 -400 2400 -250
rect 3900 4750 4550 5550
rect 8950 4750 9600 5550
rect 4900 3250 5500 4050
rect 1700 -4250 2350 -3450
rect 750 -5750 1400 -4950
rect 7100 3300 7700 4000
rect 5800 -4250 6450 -3450
rect 7950 50 8700 200
rect 7950 -400 8700 -250
rect 10200 4750 10850 5550
rect 11200 3250 11800 4050
rect 8000 -4250 8650 -3450
rect 3900 -5750 4550 -4950
rect 7050 -5750 7700 -4950
rect 12100 -4250 12750 -3450
rect 10200 -5750 10850 -4950
<< metal5 >>
rect 700 4100 2100 5700
rect 11400 5600 12800 5700
rect 2600 5550 12800 5600
rect 2600 4750 2650 5550
rect 3300 4750 3900 5550
rect 4550 4750 8950 5550
rect 9600 4750 10200 5550
rect 10850 4750 12800 5550
rect 2600 4700 12800 4750
rect 700 4050 11850 4100
rect 700 4000 4900 4050
rect 700 3300 800 4000
rect 1400 3300 4900 4000
rect 700 3250 4900 3300
rect 5500 4000 11200 4050
rect 5500 3300 7100 4000
rect 7700 3300 11200 4000
rect 5500 3250 11200 3300
rect 11800 3250 11850 4050
rect 700 3200 11850 3250
rect 650 200 12750 250
rect 650 50 1650 200
rect 2400 50 7950 200
rect 8700 50 12750 200
rect 650 0 12750 50
rect 650 -250 12750 -200
rect 650 -400 1650 -250
rect 2400 -400 7950 -250
rect 8700 -400 12750 -250
rect 650 -450 12750 -400
rect 1650 -3450 12800 -3400
rect 1650 -4250 1700 -3450
rect 2350 -4250 5800 -3450
rect 6450 -4250 8000 -3450
rect 8650 -4250 12100 -3450
rect 12750 -4250 12800 -3450
rect 1650 -4300 12800 -4250
rect 700 -4950 10900 -4900
rect 700 -5750 750 -4950
rect 1400 -5750 3900 -4950
rect 4550 -5750 7050 -4950
rect 7700 -5750 10200 -4950
rect 10850 -5750 10900 -4950
rect 700 -5800 10900 -5750
rect 700 -5900 2100 -5800
rect 11400 -5900 12800 -4300
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_0
timestamp 1663721312
transform 1 0 700 0 1 0
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_1
timestamp 1663721312
transform 1 0 3850 0 1 0
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_2
timestamp 1663721312
transform 1 0 7000 0 1 0
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_3
timestamp 1663721312
transform 1 0 10150 0 1 0
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_4
timestamp 1663721312
transform 1 0 10150 0 1 -3500
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_5
timestamp 1663721312
transform 1 0 7000 0 1 -3500
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_6
timestamp 1663721312
transform 1 0 3850 0 1 -3500
box 0 0 2569 3258
use NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_7
timestamp 1663721312
transform 1 0 700 0 1 -3500
box 0 0 2569 3258
<< labels >>
rlabel metal5 650 0 700 250 1 GL
rlabel metal5 650 -450 700 -200 1 GR
rlabel metal5 700 -5900 2100 -5800 1 SD2L
rlabel metal5 11400 -5900 12800 -5800 1 SD2R
rlabel metal5 11400 5600 12800 5700 1 SD1R
rlabel metal5 700 5600 2100 5700 1 SD1L
rlabel metal2 7015 -290 7050 -260 1 SUB
<< end >>
