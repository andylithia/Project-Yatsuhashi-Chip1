magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< locali >>
rect 7212 25454 7452 25488
rect 8854 25383 11071 25417
rect 6844 25143 7045 25177
rect 11043 25143 11077 25177
rect 7011 24998 7045 25143
rect 7011 24964 7436 24998
rect 7011 24772 7436 24806
rect 7011 24627 7045 24772
rect 6844 24593 7045 24627
rect 11043 24593 11077 24627
rect 6844 24353 7045 24387
rect 11043 24353 11077 24387
rect 7011 24208 7045 24353
rect 7011 24174 7436 24208
rect 7011 23982 7436 24016
rect 7011 23837 7045 23982
rect 6844 23803 7045 23837
rect 11043 23803 11077 23837
rect 6844 23563 7045 23597
rect 11043 23563 11077 23597
rect 7011 23418 7045 23563
rect 7011 23384 7436 23418
rect 7011 23192 7436 23226
rect 7011 23047 7045 23192
rect 6844 23013 7045 23047
rect 11043 23013 11077 23047
rect 6844 22773 7045 22807
rect 11043 22773 11077 22807
rect 7011 22628 7045 22773
rect 7011 22594 7436 22628
rect 7011 22402 7436 22436
rect 7011 22257 7045 22402
rect 6844 22223 7045 22257
rect 11043 22223 11077 22257
rect 6844 21983 7045 22017
rect 11043 21983 11077 22017
rect 7011 21838 7045 21983
rect 7011 21804 7436 21838
rect 7011 21612 7436 21646
rect 7011 21467 7045 21612
rect 6844 21433 7045 21467
rect 11043 21433 11077 21467
rect 6844 21193 7045 21227
rect 11043 21193 11077 21227
rect 7011 21048 7045 21193
rect 7011 21014 7436 21048
rect 7011 20822 7436 20856
rect 7011 20677 7045 20822
rect 6844 20643 7045 20677
rect 11043 20643 11077 20677
rect 6844 20403 7045 20437
rect 11043 20403 11077 20437
rect 7011 20258 7045 20403
rect 7011 20224 7436 20258
rect 7011 20032 7436 20066
rect 7011 19887 7045 20032
rect 6844 19853 7045 19887
rect 11043 19853 11077 19887
rect 6844 19613 7045 19647
rect 11043 19613 11077 19647
rect 7011 19468 7045 19613
rect 7011 19434 7436 19468
rect 7011 19242 7436 19276
rect 7011 19097 7045 19242
rect 6844 19063 7045 19097
rect 11043 19063 11077 19097
rect 6844 18823 7045 18857
rect 11043 18823 11077 18857
rect 7011 18678 7045 18823
rect 7011 18644 7436 18678
rect 7011 18452 7436 18486
rect 7011 18307 7045 18452
rect 6844 18273 7045 18307
rect 11043 18273 11077 18307
rect 6844 18033 7045 18067
rect 11043 18033 11077 18067
rect 7011 17888 7045 18033
rect 7011 17854 7436 17888
rect 7011 17662 7436 17696
rect 7011 17517 7045 17662
rect 6844 17483 7045 17517
rect 11043 17483 11077 17517
rect 6844 17243 7045 17277
rect 11043 17243 11077 17277
rect 7011 17098 7045 17243
rect 7011 17064 7436 17098
rect 7011 16872 7436 16906
rect 7011 16727 7045 16872
rect 6844 16693 7045 16727
rect 11043 16693 11077 16727
rect 6844 16453 7045 16487
rect 11043 16453 11077 16487
rect 7011 16308 7045 16453
rect 7011 16274 7436 16308
rect 7011 16082 7436 16116
rect 7011 15937 7045 16082
rect 6844 15903 7045 15937
rect 11043 15903 11077 15937
rect 6844 15663 7045 15697
rect 11043 15663 11077 15697
rect 7011 15518 7045 15663
rect 7011 15484 7436 15518
rect 7011 15292 7436 15326
rect 7011 15147 7045 15292
rect 6844 15113 7045 15147
rect 11043 15113 11077 15147
rect 6844 14873 7045 14907
rect 11043 14873 11077 14907
rect 7011 14728 7045 14873
rect 7011 14694 7436 14728
rect 7011 14502 7436 14536
rect 7011 14357 7045 14502
rect 6844 14323 7045 14357
rect 11043 14323 11077 14357
rect 6844 14083 7045 14117
rect 11043 14083 11077 14117
rect 7011 13938 7045 14083
rect 7011 13904 7436 13938
rect 7011 13712 7436 13746
rect 7011 13567 7045 13712
rect 6844 13533 7045 13567
rect 11043 13533 11077 13567
rect 6844 13293 7045 13327
rect 11043 13293 11077 13327
rect 7011 13148 7045 13293
rect 7011 13114 7436 13148
rect 7011 12922 7436 12956
rect 7011 12777 7045 12922
rect 6844 12743 7045 12777
rect 11043 12743 11077 12777
rect 6844 12503 7045 12537
rect 11043 12503 11077 12537
rect 7011 12358 7045 12503
rect 7011 12324 7436 12358
rect 7011 12132 7436 12166
rect 7011 11987 7045 12132
rect 6844 11953 7045 11987
rect 11043 11953 11077 11987
rect 6844 11713 7045 11747
rect 11043 11713 11077 11747
rect 7011 11568 7045 11713
rect 7011 11534 7436 11568
rect 7011 11342 7436 11376
rect 7011 11197 7045 11342
rect 6844 11163 7045 11197
rect 11043 11163 11077 11197
rect 6844 10923 7045 10957
rect 11043 10923 11077 10957
rect 7011 10778 7045 10923
rect 7011 10744 7436 10778
rect 7011 10552 7436 10586
rect 7011 10407 7045 10552
rect 6844 10373 7045 10407
rect 11043 10373 11077 10407
rect 6844 10133 7045 10167
rect 11043 10133 11077 10167
rect 7011 9988 7045 10133
rect 7011 9954 7436 9988
rect 7011 9762 7436 9796
rect 7011 9617 7045 9762
rect 6844 9583 7045 9617
rect 11043 9583 11077 9617
rect 6844 9343 7045 9377
rect 11043 9343 11077 9377
rect 7011 9198 7045 9343
rect 7011 9164 7436 9198
rect 7011 8972 7436 9006
rect 7011 8827 7045 8972
rect 6844 8793 7045 8827
rect 11043 8793 11077 8827
rect 6844 8553 7045 8587
rect 11043 8553 11077 8587
rect 7011 8408 7045 8553
rect 7011 8374 7436 8408
rect 7011 8182 7436 8216
rect 7011 8037 7045 8182
rect 6844 8003 7045 8037
rect 11043 8003 11077 8037
rect 6844 7763 7045 7797
rect 11043 7763 11077 7797
rect 7011 7618 7045 7763
rect 7011 7584 7436 7618
rect 7011 7392 7436 7426
rect 7011 7247 7045 7392
rect 6844 7213 7045 7247
rect 11043 7213 11077 7247
rect 6844 6973 7045 7007
rect 11043 6973 11077 7007
rect 7011 6828 7045 6973
rect 7011 6794 7436 6828
rect 7011 6602 7436 6636
rect 7011 6457 7045 6602
rect 6844 6423 7045 6457
rect 11043 6423 11077 6457
rect 6844 6183 7045 6217
rect 11043 6183 11077 6217
rect 7011 6038 7045 6183
rect 7011 6004 7436 6038
rect 7011 5812 7436 5846
rect 7011 5667 7045 5812
rect 6844 5633 7045 5667
rect 11043 5633 11077 5667
rect 6844 5393 7045 5427
rect 11043 5393 11077 5427
rect 7011 5248 7045 5393
rect 7011 5214 7436 5248
rect 7011 5022 7436 5056
rect 7011 4877 7045 5022
rect 6844 4843 7045 4877
rect 11043 4843 11077 4877
rect 6844 4603 7045 4637
rect 11043 4603 11077 4637
rect 7011 4458 7045 4603
rect 7011 4424 7436 4458
rect 7011 4232 7436 4266
rect 7011 4087 7045 4232
rect 6844 4053 7045 4087
rect 11043 4053 11077 4087
rect 6844 3813 7045 3847
rect 11043 3813 11077 3847
rect 7011 3668 7045 3813
rect 7011 3634 7436 3668
rect 7011 3442 7436 3476
rect 7011 3297 7045 3442
rect 6844 3263 7045 3297
rect 11043 3263 11077 3297
rect 6844 3023 7045 3057
rect 11043 3023 11077 3057
rect 7011 2878 7045 3023
rect 7011 2844 7436 2878
rect 7011 2652 7436 2686
rect 7011 2507 7045 2652
rect 6844 2473 7045 2507
rect 11043 2473 11077 2507
rect 6844 2233 7045 2267
rect 11043 2233 11077 2267
rect 7011 2088 7045 2233
rect 7011 2054 7436 2088
rect 7011 1862 7436 1896
rect 7011 1717 7045 1862
rect 6844 1683 7045 1717
rect 11043 1683 11077 1717
rect 6844 1443 7045 1477
rect 11043 1443 11077 1477
rect 7011 1298 7045 1443
rect 7011 1264 7436 1298
rect 7011 1072 7436 1106
rect 7011 927 7045 1072
rect 6844 893 7045 927
rect 11043 893 11077 927
rect 6844 653 7045 687
rect 11043 653 11077 687
rect 7011 508 7045 653
rect 7011 474 7436 508
rect 7011 282 7436 316
rect 7011 137 7045 282
rect 6844 103 7045 137
rect 11043 103 11077 137
<< metal1 >>
rect 7420 25553 7484 25605
rect 7180 25445 7244 25497
rect 8019 25248 8069 25682
rect 10321 25280 10349 25675
rect 19 0 47 6320
rect 99 0 127 6320
rect 179 0 207 6320
rect 259 0 287 6320
rect 339 0 367 6320
rect 419 0 447 6320
<< metal2 >>
rect 7184 25447 7240 25495
rect 7438 25280 7466 25593
<< metal3 >>
rect 7163 25422 7261 25520
rect 2290 5883 2388 5981
rect 2715 5883 2813 5981
rect 3094 5876 3192 5974
rect 3490 5876 3588 5974
rect 996 5086 1094 5184
rect 1392 5086 1490 5184
rect 2290 5093 2388 5191
rect 2715 5093 2813 5191
rect 3094 5086 3192 5184
rect 3490 5086 3588 5184
rect 2290 3513 2388 3611
rect 2715 3513 2813 3611
rect 3094 3506 3192 3604
rect 3490 3506 3588 3604
rect 996 2716 1094 2814
rect 1392 2716 1490 2814
rect 2290 2723 2388 2821
rect 2715 2723 2813 2821
rect 3094 2716 3192 2814
rect 3490 2716 3588 2814
rect 2290 1143 2388 1241
rect 2715 1143 2813 1241
rect 3094 1136 3192 1234
rect 3490 1136 3588 1234
rect 996 346 1094 444
rect 1392 346 1490 444
rect 2290 353 2388 451
rect 2715 353 2813 451
rect 3094 346 3192 444
rect 3490 346 3588 444
<< metal4 >>
rect 5022 -33 5088 25341
rect 5494 -33 5560 25341
rect 5926 -33 5992 25341
rect 6270 -33 6336 25341
rect 6694 -33 6760 25341
rect 7586 -63 7652 25343
rect 8011 -65 8077 25345
rect 8854 -33 8920 25313
rect 10302 -33 10368 25313
use sky130_sram_1r1w_24x128_8_and2_dec_0  sky130_sram_1r1w_24x128_8_and2_dec_0_0
timestamp 1661296025
transform 1 0 7349 0 1 25280
box 70 -56 3740 490
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_0
timestamp 1661296025
transform 1 0 7183 0 1 25438
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_13  sky130_sram_1r1w_24x128_8_contact_13_1
timestamp 1661296025
transform 1 0 7423 0 1 25546
box 0 0 58 66
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_0
timestamp 1661296025
transform 1 0 7180 0 1 25439
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_18  sky130_sram_1r1w_24x128_8_contact_18_1
timestamp 1661296025
transform 1 0 7420 0 1 25547
box 0 0 64 64
use sky130_sram_1r1w_24x128_8_contact_21  sky130_sram_1r1w_24x128_8_contact_21_0
timestamp 1661296025
transform 1 0 7179 0 1 25434
box 0 0 66 74
use sky130_sram_1r1w_24x128_8_hierarchical_decoder  sky130_sram_1r1w_24x128_8_hierarchical_decoder_0
timestamp 1661296025
transform 1 0 0 0 1 0
box 0 -60 6879 25341
use sky130_sram_1r1w_24x128_8_wordline_driver_array  sky130_sram_1r1w_24x128_8_wordline_driver_array_0
timestamp 1661296025
transform 1 0 6861 0 1 0
box 558 -65 4228 25345
<< labels >>
rlabel metal1 s 19 0 47 6320 4 addr_0
port 1 nsew
rlabel metal1 s 99 0 127 6320 4 addr_1
port 2 nsew
rlabel metal1 s 179 0 207 6320 4 addr_2
port 3 nsew
rlabel metal1 s 259 0 287 6320 4 addr_3
port 4 nsew
rlabel metal1 s 339 0 367 6320 4 addr_4
port 5 nsew
rlabel metal1 s 419 0 447 6320 4 addr_5
port 6 nsew
rlabel locali s 11060 120 11060 120 4 wl_0
port 7 nsew
rlabel locali s 11060 670 11060 670 4 wl_1
port 8 nsew
rlabel locali s 11060 910 11060 910 4 wl_2
port 9 nsew
rlabel locali s 11060 1460 11060 1460 4 wl_3
port 10 nsew
rlabel locali s 11060 1700 11060 1700 4 wl_4
port 11 nsew
rlabel locali s 11060 2250 11060 2250 4 wl_5
port 12 nsew
rlabel locali s 11060 2490 11060 2490 4 wl_6
port 13 nsew
rlabel locali s 11060 3040 11060 3040 4 wl_7
port 14 nsew
rlabel locali s 11060 3280 11060 3280 4 wl_8
port 15 nsew
rlabel locali s 11060 3830 11060 3830 4 wl_9
port 16 nsew
rlabel locali s 11060 4070 11060 4070 4 wl_10
port 17 nsew
rlabel locali s 11060 4620 11060 4620 4 wl_11
port 18 nsew
rlabel locali s 11060 4860 11060 4860 4 wl_12
port 19 nsew
rlabel locali s 11060 5410 11060 5410 4 wl_13
port 20 nsew
rlabel locali s 11060 5650 11060 5650 4 wl_14
port 21 nsew
rlabel locali s 11060 6200 11060 6200 4 wl_15
port 22 nsew
rlabel locali s 11060 6440 11060 6440 4 wl_16
port 23 nsew
rlabel locali s 11060 6990 11060 6990 4 wl_17
port 24 nsew
rlabel locali s 11060 7230 11060 7230 4 wl_18
port 25 nsew
rlabel locali s 11060 7780 11060 7780 4 wl_19
port 26 nsew
rlabel locali s 11060 8020 11060 8020 4 wl_20
port 27 nsew
rlabel locali s 11060 8570 11060 8570 4 wl_21
port 28 nsew
rlabel locali s 11060 8810 11060 8810 4 wl_22
port 29 nsew
rlabel locali s 11060 9360 11060 9360 4 wl_23
port 30 nsew
rlabel locali s 11060 9600 11060 9600 4 wl_24
port 31 nsew
rlabel locali s 11060 10150 11060 10150 4 wl_25
port 32 nsew
rlabel locali s 11060 10390 11060 10390 4 wl_26
port 33 nsew
rlabel locali s 11060 10940 11060 10940 4 wl_27
port 34 nsew
rlabel locali s 11060 11180 11060 11180 4 wl_28
port 35 nsew
rlabel locali s 11060 11730 11060 11730 4 wl_29
port 36 nsew
rlabel locali s 11060 11970 11060 11970 4 wl_30
port 37 nsew
rlabel locali s 11060 12520 11060 12520 4 wl_31
port 38 nsew
rlabel locali s 11060 12760 11060 12760 4 wl_32
port 39 nsew
rlabel locali s 11060 13310 11060 13310 4 wl_33
port 40 nsew
rlabel locali s 11060 13550 11060 13550 4 wl_34
port 41 nsew
rlabel locali s 11060 14100 11060 14100 4 wl_35
port 42 nsew
rlabel locali s 11060 14340 11060 14340 4 wl_36
port 43 nsew
rlabel locali s 11060 14890 11060 14890 4 wl_37
port 44 nsew
rlabel locali s 11060 15130 11060 15130 4 wl_38
port 45 nsew
rlabel locali s 11060 15680 11060 15680 4 wl_39
port 46 nsew
rlabel locali s 11060 15920 11060 15920 4 wl_40
port 47 nsew
rlabel locali s 11060 16470 11060 16470 4 wl_41
port 48 nsew
rlabel locali s 11060 16710 11060 16710 4 wl_42
port 49 nsew
rlabel locali s 11060 17260 11060 17260 4 wl_43
port 50 nsew
rlabel locali s 11060 17500 11060 17500 4 wl_44
port 51 nsew
rlabel locali s 11060 18050 11060 18050 4 wl_45
port 52 nsew
rlabel locali s 11060 18290 11060 18290 4 wl_46
port 53 nsew
rlabel locali s 11060 18840 11060 18840 4 wl_47
port 54 nsew
rlabel locali s 11060 19080 11060 19080 4 wl_48
port 55 nsew
rlabel locali s 11060 19630 11060 19630 4 wl_49
port 56 nsew
rlabel locali s 11060 19870 11060 19870 4 wl_50
port 57 nsew
rlabel locali s 11060 20420 11060 20420 4 wl_51
port 58 nsew
rlabel locali s 11060 20660 11060 20660 4 wl_52
port 59 nsew
rlabel locali s 11060 21210 11060 21210 4 wl_53
port 60 nsew
rlabel locali s 11060 21450 11060 21450 4 wl_54
port 61 nsew
rlabel locali s 11060 22000 11060 22000 4 wl_55
port 62 nsew
rlabel locali s 11060 22240 11060 22240 4 wl_56
port 63 nsew
rlabel locali s 11060 22790 11060 22790 4 wl_57
port 64 nsew
rlabel locali s 11060 23030 11060 23030 4 wl_58
port 65 nsew
rlabel locali s 11060 23580 11060 23580 4 wl_59
port 66 nsew
rlabel locali s 11060 23820 11060 23820 4 wl_60
port 67 nsew
rlabel locali s 11060 24370 11060 24370 4 wl_61
port 68 nsew
rlabel locali s 11060 24610 11060 24610 4 wl_62
port 69 nsew
rlabel locali s 11060 25160 11060 25160 4 wl_63
port 70 nsew
rlabel locali s 9962 25400 9962 25400 4 rbl_wl
port 71 nsew
rlabel metal2 s 7438 25565 7466 25593 4 wl_en
port 72 nsew
rlabel metal3 s 1392 346 1490 444 4 vdd
port 73 nsew
rlabel metal3 s 2715 3513 2813 3611 4 vdd
port 73 nsew
rlabel metal3 s 2715 1143 2813 1241 4 vdd
port 73 nsew
rlabel metal3 s 3490 346 3588 444 4 vdd
port 73 nsew
rlabel metal4 s 8011 -65 8077 25345 4 vdd
port 73 nsew
rlabel metal3 s 1392 5086 1490 5184 4 vdd
port 73 nsew
rlabel metal3 s 2715 2723 2813 2821 4 vdd
port 73 nsew
rlabel metal3 s 3490 1136 3588 1234 4 vdd
port 73 nsew
rlabel metal4 s 5494 -33 5560 25341 4 vdd
port 73 nsew
rlabel metal3 s 3490 3506 3588 3604 4 vdd
port 73 nsew
rlabel metal3 s 3490 5086 3588 5184 4 vdd
port 73 nsew
rlabel metal3 s 2715 353 2813 451 4 vdd
port 73 nsew
rlabel metal3 s 7163 25422 7261 25520 4 vdd
port 73 nsew
rlabel metal3 s 2715 5093 2813 5191 4 vdd
port 73 nsew
rlabel metal4 s 6694 -33 6760 25341 4 vdd
port 73 nsew
rlabel metal3 s 3490 5876 3588 5974 4 vdd
port 73 nsew
rlabel metal1 s 8019 25248 8069 25682 4 vdd
port 73 nsew
rlabel metal3 s 1392 2716 1490 2814 4 vdd
port 73 nsew
rlabel metal1 s 10321 25280 10349 25675 4 vdd
port 73 nsew
rlabel metal4 s 5926 -33 5992 25341 4 vdd
port 73 nsew
rlabel metal4 s 10302 -33 10368 25313 4 vdd
port 73 nsew
rlabel metal3 s 3490 2716 3588 2814 4 vdd
port 73 nsew
rlabel metal3 s 2715 5883 2813 5981 4 vdd
port 73 nsew
rlabel metal3 s 3094 3506 3192 3604 4 gnd
port 74 nsew
rlabel metal3 s 3094 346 3192 444 4 gnd
port 74 nsew
rlabel metal3 s 3094 5086 3192 5184 4 gnd
port 74 nsew
rlabel metal3 s 996 5086 1094 5184 4 gnd
port 74 nsew
rlabel metal3 s 3094 1136 3192 1234 4 gnd
port 74 nsew
rlabel metal4 s 7586 -63 7652 25343 4 gnd
port 74 nsew
rlabel metal4 s 5022 -33 5088 25341 4 gnd
port 74 nsew
rlabel metal3 s 3094 5876 3192 5974 4 gnd
port 74 nsew
rlabel metal4 s 8854 -33 8920 25313 4 gnd
port 74 nsew
rlabel metal3 s 2290 1143 2388 1241 4 gnd
port 74 nsew
rlabel metal3 s 996 346 1094 444 4 gnd
port 74 nsew
rlabel metal3 s 996 2716 1094 2814 4 gnd
port 74 nsew
rlabel metal4 s 6270 -33 6336 25341 4 gnd
port 74 nsew
rlabel metal3 s 2290 2723 2388 2821 4 gnd
port 74 nsew
rlabel metal3 s 2290 353 2388 451 4 gnd
port 74 nsew
rlabel metal3 s 3094 2716 3192 2814 4 gnd
port 74 nsew
rlabel metal3 s 2290 3513 2388 3611 4 gnd
port 74 nsew
rlabel metal3 s 2290 5883 2388 5981 4 gnd
port 74 nsew
rlabel metal3 s 2290 5093 2388 5191 4 gnd
port 74 nsew
<< properties >>
string FIXED_BBOX 0 0 11107 25308
<< end >>
