** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/untitled-6.sch
**.subckt untitled-6
XM3 net2 net4 vmid GND sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext w=5.05u l=0.15u m=12
V2 net3 GND DC 0.9 AC 0 portnum 2 z0 50
V1 net1 GND DC 1.8 AC 0 portnum 1 z0 50
L1 vmid net5 5n m=1
V3 net2 GND DC 1.8
C1 net3 vmid 1p m=1
L2 net4 net6 1n m=1
R1 net5 GND 500 m=1
C2 net6 net1 1p m=1
R2 net2 net6 2k m=1
**** begin user architecture code


.subckt sky130_fd_pr__rf_nfet_01v8_bM04W5p00L0p15_ext DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=4.242e+12p
+ ps=3.198e+07u w=5.05e+06u l=150000u
X1 SOURCE SUBSTRATE SUBSTRATE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.03e+12p
+ ps=2.14e+07u w=5.05e+06u l=150000u
X2 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 SUBSTRATE SUBSTRATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X5 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends
* .options savecurrents
.sp dec 1000 1e9 10e9 1
.control
run
display
*let vo = v(von)-v(vop)
*plot v(von) v(vop)
*plot vo
*fft vo
*plot db(vo)

.endc


.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
* .include
*+ /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
