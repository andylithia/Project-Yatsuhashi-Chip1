magic
tech sky130B
magscale 1 2
timestamp 1663980778
<< metal4 >>
rect -57000 -28112 -38500 -28000
rect -57000 -35888 -46388 -28112
rect -38612 -35888 -38500 -28112
rect -57000 -36000 -38500 -35888
<< via4 >>
rect -46388 -35888 -38612 -28112
<< metal5 >>
tri -49069 12000 -41069 20000 se
rect -41069 12000 -7931 20000
tri -7931 12000 69 20000 sw
tri -56655 4414 -49069 12000 se
rect -49069 11000 -38755 12000
tri -38755 11000 -37755 12000 nw
tri -11245 11000 -10245 12000 ne
rect -10245 11000 69 12000
rect -49069 9586 -40169 11000
tri -40169 9586 -38755 11000 nw
tri -38755 9586 -37341 11000 se
rect -37341 9586 -11659 11000
tri -11659 9586 -10245 11000 sw
tri -10245 9586 -8831 11000 ne
rect -8831 9586 69 11000
rect -49069 8172 -41583 9586
tri -41583 8172 -40169 9586 nw
tri -40169 8172 -38755 9586 se
rect -38755 8172 -10245 9586
tri -10245 8172 -8831 9586 sw
tri -8831 8172 -7417 9586 ne
rect -7417 8172 69 9586
rect -49069 7242 -42513 8172
tri -42513 7242 -41583 8172 nw
tri -41099 7242 -40169 8172 se
rect -40169 7242 -8831 8172
rect -49069 5828 -43927 7242
tri -43927 5828 -42513 7242 nw
tri -42513 5828 -41099 7242 se
rect -41099 6758 -8831 7242
tri -8831 6758 -7417 8172 sw
tri -7417 6758 -6003 8172 ne
rect -6003 6758 69 8172
rect -41099 5828 -7417 6758
tri -7417 5828 -6487 6758 sw
tri -6003 5828 -5073 6758 ne
rect -5073 5828 69 6758
rect -49069 4414 -45341 5828
tri -45341 4414 -43927 5828 nw
tri -43927 4414 -42513 5828 se
rect -42513 4414 -6487 5828
tri -6487 4414 -5073 5828 sw
tri -5073 4414 -3659 5828 ne
rect -3659 4414 69 5828
tri -64500 -3431 -56655 4414 se
rect -56655 3000 -46755 4414
tri -46755 3000 -45341 4414 nw
tri -45341 3000 -43927 4414 se
rect -43927 3000 -5073 4414
tri -5073 3000 -3659 4414 sw
tri -3659 3000 -2245 4414 ne
rect -2245 3000 69 4414
rect -56655 1586 -48169 3000
tri -48169 1586 -46755 3000 nw
tri -46755 1586 -45341 3000 se
rect -56655 172 -49583 1586
tri -49583 172 -48169 1586 nw
tri -48169 172 -46755 1586 se
rect -46755 172 -45341 1586
rect -56655 -1172 -50927 172
tri -50927 -1172 -49583 172 nw
tri -49513 -1172 -48169 172 se
rect -48169 -1172 -45341 172
rect -56655 -2586 -52341 -1172
tri -52341 -2586 -50927 -1172 nw
tri -50927 -2586 -49513 -1172 se
rect -49513 -2586 -45341 -1172
rect -56655 -3431 -53755 -2586
rect -64500 -4000 -53755 -3431
tri -53755 -4000 -52341 -2586 nw
tri -52341 -4000 -50927 -2586 se
rect -50927 -4000 -45341 -2586
rect -66000 -5414 -55169 -4000
tri -55169 -5414 -53755 -4000 nw
tri -53755 -5414 -52341 -4000 se
rect -52341 -5414 -45341 -4000
rect -66000 -12000 -56500 -5414
tri -56500 -6745 -55169 -5414 nw
tri -55086 -6745 -53755 -5414 se
rect -53755 -6745 -45341 -5414
tri -55500 -7159 -55086 -6745 se
rect -55086 -7159 -45341 -6745
rect -55500 -8314 -45341 -7159
tri -45341 -8314 -34027 3000 nw
tri -14973 -8314 -3659 3000 ne
tri -3659 2255 -2914 3000 sw
tri -2245 2255 -1500 3000 ne
rect -1500 2255 69 3000
rect -3659 841 -2914 2255
tri -2914 841 -1500 2255 sw
tri -1500 841 -86 2255 ne
rect -86 841 69 2255
tri 69 841 11228 12000 sw
rect -3659 -573 -1500 841
tri -1500 -573 -86 841 sw
tri -86 -573 1328 841 ne
rect 1328 -573 11228 841
rect -3659 -1987 -86 -573
tri -86 -1987 1328 -573 sw
tri 1328 -1987 2742 -573 ne
rect 2742 -1987 11228 -573
rect -3659 -2917 1328 -1987
tri 1328 -2917 2258 -1987 sw
tri 2742 -2917 3672 -1987 ne
rect 3672 -2917 11228 -1987
rect -3659 -4331 2258 -2917
tri 2258 -4331 3672 -2917 sw
tri 3672 -4331 5086 -2917 ne
rect 5086 -3431 11228 -2917
tri 11228 -3431 15500 841 sw
rect 5086 -4331 15500 -3431
rect -3659 -5745 3672 -4331
tri 3672 -5745 5086 -4331 sw
tri 5086 -5745 6500 -4331 ne
rect 6500 -5745 15500 -4331
rect -3659 -7159 5086 -5745
tri 5086 -7159 6500 -5745 sw
tri 6500 -6745 7500 -5745 ne
rect -3659 -8314 6500 -7159
rect -55500 -36891 -47500 -8314
tri -47500 -10473 -45341 -8314 nw
tri -3659 -10473 -1500 -8314 ne
rect -46500 -28112 -38500 -28000
rect -46500 -35888 -46388 -28112
rect -38612 -35888 -38500 -28112
tri -47500 -36891 -46500 -35891 sw
rect -46500 -36000 -38500 -35888
tri -45977 -36891 -45086 -36000 ne
rect -45086 -36891 -38500 -36000
rect -55500 -38305 -46500 -36891
tri -46500 -38305 -45086 -36891 sw
tri -45086 -38305 -43672 -36891 ne
rect -43672 -38305 -38500 -36891
rect -55500 -39205 -45086 -38305
tri -55500 -43000 -51705 -39205 ne
rect -51705 -39719 -45086 -39205
tri -45086 -39719 -43672 -38305 sw
tri -43672 -39719 -42258 -38305 ne
rect -42258 -39719 -38500 -38305
rect -51705 -40172 -43672 -39719
tri -43672 -40172 -43219 -39719 sw
tri -42258 -40172 -41805 -39719 ne
rect -41805 -40172 -38500 -39719
rect -51705 -41586 -43219 -40172
tri -43219 -41586 -41805 -40172 sw
tri -41805 -41586 -40391 -40172 ne
rect -40391 -41586 -38500 -40172
rect -51705 -43000 -41805 -41586
tri -41805 -43000 -40391 -41586 sw
tri -40391 -43000 -38977 -41586 ne
rect -38977 -43000 -38500 -41586
tri -38500 -43000 -27663 -32163 sw
tri -12337 -43000 -1500 -32163 se
rect -1500 -35477 6500 -8314
rect -1500 -36891 5086 -35477
tri 5086 -36891 6500 -35477 nw
tri 6500 -36891 7500 -35891 se
rect 7500 -36891 15500 -5745
rect -1500 -38305 3672 -36891
tri 3672 -38305 5086 -36891 nw
tri 5086 -38305 6500 -36891 se
rect 6500 -38305 15500 -36891
rect -1500 -39719 2258 -38305
tri 2258 -39719 3672 -38305 nw
tri 3672 -39719 5086 -38305 se
rect 5086 -39205 15500 -38305
rect 5086 -39719 7500 -39205
rect -1500 -40172 1805 -39719
tri 1805 -40172 2258 -39719 nw
tri 3219 -40172 3672 -39719 se
rect 3672 -40172 7500 -39719
rect -1500 -41586 391 -40172
tri 391 -41586 1805 -40172 nw
tri 1805 -41586 3219 -40172 se
rect 3219 -41586 7500 -40172
rect -1500 -43000 -1023 -41586
tri -1023 -43000 391 -41586 nw
tri 391 -43000 1805 -41586 se
rect 1805 -43000 7500 -41586
tri -51705 -52000 -42705 -43000 ne
rect -42705 -44414 -40391 -43000
tri -40391 -44414 -38977 -43000 sw
tri -38977 -44414 -37563 -43000 ne
rect -37563 -43477 -1500 -43000
tri -1500 -43477 -1023 -43000 nw
tri -86 -43477 391 -43000 se
rect 391 -43477 7500 -43000
rect -37563 -44414 -2914 -43477
rect -42705 -45828 -38977 -44414
tri -38977 -45828 -37563 -44414 sw
tri -37563 -45828 -36149 -44414 ne
rect -36149 -44891 -2914 -44414
tri -2914 -44891 -1500 -43477 nw
tri -1500 -44891 -86 -43477 se
rect -86 -44891 7500 -43477
rect -36149 -45828 -4328 -44891
rect -42705 -47242 -37563 -45828
tri -37563 -47242 -36149 -45828 sw
tri -36149 -47242 -34735 -45828 ne
rect -34735 -46305 -4328 -45828
tri -4328 -46305 -2914 -44891 nw
tri -2914 -46305 -1500 -44891 se
rect -1500 -46305 7500 -44891
rect -34735 -47242 -5742 -46305
rect -42705 -48172 -36149 -47242
tri -36149 -48172 -35219 -47242 sw
tri -34735 -48172 -33805 -47242 ne
rect -33805 -47719 -5742 -47242
tri -5742 -47719 -4328 -46305 nw
tri -4328 -47719 -2914 -46305 se
rect -2914 -47205 7500 -46305
tri 7500 -47205 15500 -39205 nw
rect -2914 -47719 -1500 -47205
rect -33805 -48172 -6195 -47719
tri -6195 -48172 -5742 -47719 nw
tri -4781 -48172 -4328 -47719 se
rect -4328 -48172 -1500 -47719
rect -42705 -49586 -35219 -48172
tri -35219 -49586 -33805 -48172 sw
tri -33805 -49586 -32391 -48172 ne
rect -32391 -49586 -7609 -48172
tri -7609 -49586 -6195 -48172 nw
tri -6195 -49586 -4781 -48172 se
rect -4781 -49586 -1500 -48172
rect -42705 -51000 -33805 -49586
tri -33805 -51000 -32391 -49586 sw
tri -32391 -51000 -30977 -49586 ne
rect -30977 -51000 -9023 -49586
tri -9023 -51000 -7609 -49586 nw
tri -7609 -51000 -6195 -49586 se
rect -6195 -51000 -1500 -49586
rect -42705 -52000 -32391 -51000
tri -32391 -52000 -31391 -51000 sw
tri -8609 -52000 -7609 -51000 se
rect -7609 -52000 -1500 -51000
tri -42705 -60000 -34705 -52000 ne
rect -34705 -56205 -1500 -52000
tri -1500 -56205 7500 -47205 nw
rect -34705 -60000 -5295 -56205
tri -5295 -60000 -1500 -56205 nw
<< end >>
