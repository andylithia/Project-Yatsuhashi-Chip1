magic
tech sky130B
timestamp 1658693857
<< metal4 >>
rect 900 150 1400 2200
rect 900 0 950 150
rect 1100 0 1150 150
rect 1300 0 1400 150
rect 900 -50 1400 0
rect 900 -200 1000 -50
rect 1150 -200 1200 -50
rect 1350 -200 1400 -50
rect 900 -250 1400 -200
<< via4 >>
rect 950 0 1100 150
rect 1150 0 1300 150
rect 1000 -200 1150 -50
rect 1200 -200 1350 -50
<< metal5 >>
rect 100 1300 8100 1800
rect 100 500 7300 1000
rect 100 -5700 600 500
rect 900 150 1400 200
rect 900 0 950 150
rect 1100 0 1150 150
rect 1300 0 1400 150
rect 900 -50 1400 0
rect 900 -200 1000 -50
rect 1150 -200 1200 -50
rect 1350 -200 1400 -50
rect 900 -4900 1400 -200
rect 6800 -4900 7300 500
rect 900 -5400 7300 -4900
rect 7600 -5700 8100 1300
rect 100 -6200 8100 -5700
<< labels >>
rlabel metal5 100 1300 600 1800 1 A
rlabel metal4 900 1850 1400 2100 1 B
<< end >>
