magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< error_s >>
rect 182 26465 224 26491
rect 544 26482 586 26491
rect 186 26457 220 26465
rect 186 26450 190 26457
rect 216 26450 220 26457
rect 170 26449 236 26450
rect 120 26435 170 26437
rect 76 26431 130 26435
rect 110 26426 130 26431
rect 60 26401 67 26411
rect 76 26401 77 26421
rect 96 26392 99 26426
rect 109 26401 110 26421
rect 119 26401 126 26411
rect 76 26385 92 26391
rect 94 26385 110 26391
rect 170 26385 172 26435
rect 213 26337 224 26375
rect 251 26337 287 26365
rect 12 26332 62 26334
rect 28 26323 59 26325
rect 62 26323 64 26332
rect 251 26331 263 26337
rect 28 26315 64 26323
rect 127 26323 161 26325
rect 127 26316 182 26323
rect 127 26315 161 26316
rect 59 26299 64 26315
rect 253 26303 263 26331
rect 273 26303 287 26337
rect 28 26291 64 26299
rect 127 26298 161 26299
rect 127 26291 182 26298
rect 62 26282 64 26291
rect 120 26229 170 26231
rect 76 26223 92 26229
rect 94 26223 110 26229
rect 76 26213 99 26222
rect 60 26203 67 26213
rect 76 26193 77 26213
rect 96 26188 99 26213
rect 109 26193 110 26213
rect 119 26203 126 26213
rect 76 26179 110 26183
rect 170 26179 172 26229
rect 182 26173 224 26174
rect 186 26132 220 26166
rect 223 26132 257 26166
rect 160 26125 182 26131
rect 224 26125 246 26131
rect 288 26125 292 26465
rect 439 26448 444 26482
rect 468 26448 473 26482
rect 511 26465 586 26482
rect 476 26411 480 26465
rect 511 26448 582 26465
rect 544 26441 548 26448
rect 476 26331 480 26399
rect 544 26361 548 26411
rect 544 26321 553 26349
rect 599 26332 649 26334
rect 607 26323 624 26325
rect 476 26253 480 26321
rect 485 26277 495 26311
rect 505 26277 519 26311
rect 544 26277 555 26321
rect 586 26316 641 26323
rect 607 26315 641 26316
rect 616 26299 641 26315
rect 607 26298 641 26299
rect 586 26291 641 26298
rect 649 26282 651 26332
rect 485 26253 492 26277
rect 476 26173 480 26241
rect 544 26203 548 26253
rect 544 26168 548 26173
rect 295 26132 300 26166
rect 324 26132 329 26166
rect 544 26164 582 26168
rect 544 26134 552 26164
rect 578 26134 582 26164
rect 544 26131 548 26134
rect 522 26125 548 26131
rect 586 26125 608 26131
rect 182 26109 224 26125
rect 544 26109 586 26125
rect 17 26095 67 26097
rect 119 26095 169 26097
rect 599 26095 649 26097
rect 42 26053 59 26087
rect 67 26045 69 26095
rect 160 26087 246 26095
rect 522 26087 608 26095
rect 76 26053 110 26087
rect 127 26053 144 26087
rect 152 26053 161 26087
rect 162 26085 195 26087
rect 224 26085 244 26087
rect 162 26053 244 26085
rect 524 26085 548 26087
rect 573 26085 582 26087
rect 586 26085 606 26087
rect 160 26045 246 26053
rect 186 26029 220 26031
rect 182 26015 224 26016
rect 160 26009 182 26015
rect 224 26009 246 26015
rect 186 25974 220 26008
rect 223 25974 257 26008
rect 120 25961 170 25963
rect 76 25957 130 25961
rect 110 25952 130 25957
rect 60 25927 67 25937
rect 76 25927 77 25947
rect 96 25918 99 25952
rect 109 25927 110 25947
rect 119 25927 126 25937
rect 76 25911 92 25917
rect 94 25911 110 25917
rect 170 25911 172 25961
rect 186 25895 190 25929
rect 216 25895 220 25929
rect 288 25895 292 26083
rect 476 26015 480 26083
rect 524 26053 606 26085
rect 607 26053 616 26087
rect 522 26045 608 26053
rect 649 26045 651 26095
rect 548 26029 582 26031
rect 522 26010 548 26015
rect 522 26009 582 26010
rect 586 26009 608 26015
rect 295 25974 300 26008
rect 324 25974 329 26008
rect 544 26006 582 26009
rect 378 25969 450 25977
rect 428 25939 430 25955
rect 400 25931 430 25939
rect 476 25937 480 26005
rect 544 25976 552 26006
rect 578 25976 582 26006
rect 544 25967 548 25976
rect 400 25927 434 25931
rect 400 25897 408 25927
rect 420 25897 434 25927
rect 544 25929 548 25937
rect 12 25858 62 25860
rect 28 25849 59 25851
rect 62 25849 64 25858
rect 28 25841 64 25849
rect 127 25849 158 25851
rect 127 25842 182 25849
rect 215 25847 224 25875
rect 127 25841 161 25842
rect 59 25825 64 25841
rect 158 25825 161 25841
rect 28 25817 64 25825
rect 127 25824 161 25825
rect 127 25817 182 25824
rect 62 25808 64 25817
rect 213 25809 224 25847
rect 282 25837 292 25895
rect 296 25889 368 25897
rect 319 25860 335 25862
rect 251 25803 263 25837
rect 273 25803 292 25837
rect 303 25830 316 25846
rect 303 25812 316 25828
rect 120 25755 170 25757
rect 76 25749 92 25755
rect 94 25749 110 25755
rect 76 25739 99 25748
rect 60 25729 67 25739
rect 76 25719 77 25739
rect 96 25714 99 25739
rect 109 25719 110 25739
rect 119 25729 126 25739
rect 76 25705 110 25709
rect 170 25705 172 25755
rect 186 25737 190 25771
rect 216 25737 220 25771
rect 186 25660 220 25694
rect 282 25691 292 25803
rect 318 25806 324 25859
rect 346 25846 348 25859
rect 428 25850 430 25897
rect 443 25887 450 25889
rect 476 25857 480 25925
rect 544 25895 552 25929
rect 578 25895 582 25929
rect 481 25863 517 25891
rect 481 25857 495 25863
rect 333 25812 353 25846
rect 367 25816 380 25850
rect 396 25816 408 25850
rect 420 25816 434 25850
rect 318 25796 335 25806
rect 318 25727 324 25796
rect 346 25727 348 25812
rect 428 25769 430 25816
rect 476 25779 480 25847
rect 485 25829 495 25857
rect 505 25829 519 25863
rect 544 25857 555 25895
rect 544 25829 553 25857
rect 544 25809 548 25829
rect 579 25788 582 25878
rect 599 25858 649 25860
rect 610 25850 624 25851
rect 607 25849 624 25850
rect 586 25842 644 25849
rect 607 25841 644 25842
rect 607 25825 610 25841
rect 616 25825 644 25841
rect 607 25824 644 25825
rect 586 25817 644 25824
rect 607 25816 610 25817
rect 649 25808 651 25858
rect 544 25771 548 25779
rect 400 25739 408 25769
rect 420 25739 434 25769
rect 400 25735 434 25739
rect 400 25727 430 25735
rect 428 25711 430 25727
rect 476 25699 480 25767
rect 544 25737 552 25771
rect 578 25737 582 25771
rect 544 25729 548 25737
rect 544 25699 586 25700
rect 288 25659 292 25691
rect 296 25689 368 25697
rect 378 25689 450 25697
rect 544 25692 548 25699
rect 439 25661 444 25689
rect 120 25645 170 25647
rect 76 25641 130 25645
rect 110 25636 130 25641
rect 60 25611 67 25621
rect 76 25611 77 25631
rect 96 25602 99 25636
rect 109 25611 110 25631
rect 119 25611 126 25621
rect 76 25595 92 25601
rect 94 25595 110 25601
rect 170 25595 172 25645
rect 186 25579 190 25613
rect 216 25579 220 25613
rect 213 25547 224 25579
rect 282 25575 292 25659
rect 296 25653 368 25661
rect 378 25653 450 25661
rect 468 25658 473 25692
rect 428 25623 430 25639
rect 251 25547 292 25575
rect 12 25542 62 25544
rect 28 25533 59 25535
rect 62 25533 64 25542
rect 251 25541 263 25547
rect 28 25525 64 25533
rect 127 25533 158 25535
rect 127 25526 182 25533
rect 127 25525 161 25526
rect 59 25509 64 25525
rect 158 25509 161 25525
rect 253 25513 263 25541
rect 273 25513 292 25547
rect 318 25554 324 25623
rect 318 25544 335 25554
rect 303 25522 316 25538
rect 28 25501 64 25509
rect 127 25508 161 25509
rect 127 25501 182 25508
rect 62 25492 64 25501
rect 282 25455 292 25513
rect 303 25504 316 25520
rect 318 25491 324 25544
rect 346 25538 348 25623
rect 400 25615 430 25623
rect 476 25621 480 25689
rect 511 25658 582 25692
rect 544 25651 548 25658
rect 400 25611 434 25615
rect 400 25581 408 25611
rect 420 25581 434 25611
rect 544 25613 548 25621
rect 333 25504 353 25538
rect 428 25534 430 25581
rect 476 25541 480 25609
rect 544 25579 552 25613
rect 578 25579 582 25613
rect 544 25571 548 25579
rect 346 25491 348 25504
rect 367 25500 380 25534
rect 396 25500 408 25534
rect 420 25500 434 25534
rect 544 25531 553 25559
rect 319 25488 335 25490
rect 120 25439 170 25441
rect 76 25433 92 25439
rect 94 25433 110 25439
rect 76 25423 99 25432
rect 60 25413 67 25423
rect 76 25403 77 25423
rect 96 25398 99 25423
rect 109 25403 110 25423
rect 119 25413 126 25423
rect 76 25389 110 25393
rect 170 25389 172 25439
rect 186 25421 190 25455
rect 216 25421 220 25455
rect 182 25383 224 25384
rect 186 25342 220 25376
rect 223 25342 257 25376
rect 160 25335 182 25341
rect 224 25335 246 25341
rect 288 25335 292 25455
rect 296 25453 368 25461
rect 428 25453 430 25500
rect 476 25463 480 25531
rect 485 25487 495 25521
rect 505 25487 519 25521
rect 544 25487 555 25531
rect 485 25463 492 25487
rect 579 25472 582 25562
rect 599 25542 649 25544
rect 610 25534 624 25535
rect 607 25533 624 25534
rect 586 25526 644 25533
rect 607 25525 644 25526
rect 607 25509 610 25525
rect 616 25509 644 25525
rect 607 25508 644 25509
rect 586 25501 644 25508
rect 607 25500 610 25501
rect 649 25492 651 25542
rect 544 25455 548 25463
rect 400 25423 408 25453
rect 420 25423 434 25453
rect 400 25419 434 25423
rect 400 25411 430 25419
rect 428 25395 430 25411
rect 476 25383 480 25451
rect 544 25421 552 25455
rect 578 25421 582 25455
rect 544 25413 548 25421
rect 295 25342 300 25376
rect 324 25342 329 25376
rect 378 25373 450 25381
rect 544 25378 548 25383
rect 544 25374 582 25378
rect 544 25344 552 25374
rect 578 25344 582 25374
rect 544 25341 548 25344
rect 522 25335 548 25341
rect 586 25335 608 25341
rect 182 25319 224 25335
rect 544 25319 586 25335
rect 17 25305 67 25307
rect 119 25305 169 25307
rect 599 25305 649 25307
rect 42 25263 59 25297
rect 67 25255 69 25305
rect 160 25297 246 25305
rect 522 25297 608 25305
rect 76 25263 110 25297
rect 127 25263 144 25297
rect 152 25263 161 25297
rect 162 25295 195 25297
rect 224 25295 244 25297
rect 162 25263 244 25295
rect 524 25295 548 25297
rect 573 25295 582 25297
rect 586 25295 606 25297
rect 160 25255 246 25263
rect 186 25239 220 25241
rect 182 25225 224 25226
rect 160 25219 182 25225
rect 224 25219 246 25225
rect 186 25184 220 25218
rect 223 25184 257 25218
rect 120 25171 170 25173
rect 76 25167 130 25171
rect 110 25162 130 25167
rect 60 25137 67 25147
rect 76 25137 77 25157
rect 96 25128 99 25162
rect 109 25137 110 25157
rect 119 25137 126 25147
rect 76 25121 92 25127
rect 94 25121 110 25127
rect 170 25121 172 25171
rect 186 25105 190 25139
rect 216 25105 220 25139
rect 288 25105 292 25293
rect 476 25225 480 25293
rect 524 25263 606 25295
rect 607 25263 616 25297
rect 522 25255 608 25263
rect 649 25255 651 25305
rect 548 25239 582 25241
rect 522 25220 548 25225
rect 522 25219 582 25220
rect 586 25219 608 25225
rect 295 25184 300 25218
rect 324 25184 329 25218
rect 544 25216 582 25219
rect 378 25179 450 25187
rect 428 25149 430 25165
rect 400 25141 430 25149
rect 476 25147 480 25215
rect 544 25186 552 25216
rect 578 25186 582 25216
rect 544 25177 548 25186
rect 400 25137 434 25141
rect 400 25107 408 25137
rect 420 25107 434 25137
rect 544 25139 548 25147
rect 12 25068 62 25070
rect 28 25059 59 25061
rect 62 25059 64 25068
rect 28 25051 64 25059
rect 127 25059 158 25061
rect 127 25052 182 25059
rect 215 25057 224 25085
rect 127 25051 161 25052
rect 59 25035 64 25051
rect 158 25035 161 25051
rect 28 25027 64 25035
rect 127 25034 161 25035
rect 127 25027 182 25034
rect 62 25018 64 25027
rect 213 25019 224 25057
rect 282 25047 292 25105
rect 296 25099 368 25107
rect 319 25070 335 25072
rect 251 25013 263 25047
rect 273 25013 292 25047
rect 303 25040 316 25056
rect 303 25022 316 25038
rect 120 24965 170 24967
rect 76 24959 92 24965
rect 94 24959 110 24965
rect 76 24949 99 24958
rect 60 24939 67 24949
rect 76 24929 77 24949
rect 96 24924 99 24949
rect 109 24929 110 24949
rect 119 24939 126 24949
rect 76 24915 110 24919
rect 170 24915 172 24965
rect 186 24947 190 24981
rect 216 24947 220 24981
rect 186 24870 220 24904
rect 282 24901 292 25013
rect 318 25016 324 25069
rect 346 25056 348 25069
rect 428 25060 430 25107
rect 443 25097 450 25099
rect 476 25067 480 25135
rect 544 25105 552 25139
rect 578 25105 582 25139
rect 481 25073 517 25101
rect 481 25067 495 25073
rect 333 25022 353 25056
rect 367 25026 380 25060
rect 396 25026 408 25060
rect 420 25026 434 25060
rect 318 25006 335 25016
rect 318 24937 324 25006
rect 346 24937 348 25022
rect 428 24979 430 25026
rect 476 24989 480 25057
rect 485 25039 495 25067
rect 505 25039 519 25073
rect 544 25067 555 25105
rect 544 25039 553 25067
rect 544 25019 548 25039
rect 579 24998 582 25088
rect 599 25068 649 25070
rect 610 25060 624 25061
rect 607 25059 624 25060
rect 586 25052 644 25059
rect 607 25051 644 25052
rect 607 25035 610 25051
rect 616 25035 644 25051
rect 607 25034 644 25035
rect 586 25027 644 25034
rect 607 25026 610 25027
rect 649 25018 651 25068
rect 544 24981 548 24989
rect 400 24949 408 24979
rect 420 24949 434 24979
rect 400 24945 434 24949
rect 400 24937 430 24945
rect 428 24921 430 24937
rect 476 24909 480 24977
rect 544 24947 552 24981
rect 578 24947 582 24981
rect 544 24939 548 24947
rect 544 24909 586 24910
rect 288 24869 292 24901
rect 296 24899 368 24907
rect 378 24899 450 24907
rect 544 24902 548 24909
rect 439 24871 444 24899
rect 120 24855 170 24857
rect 76 24851 130 24855
rect 110 24846 130 24851
rect 60 24821 67 24831
rect 76 24821 77 24841
rect 96 24812 99 24846
rect 109 24821 110 24841
rect 119 24821 126 24831
rect 76 24805 92 24811
rect 94 24805 110 24811
rect 170 24805 172 24855
rect 186 24789 190 24823
rect 216 24789 220 24823
rect 213 24757 224 24789
rect 282 24785 292 24869
rect 296 24863 368 24871
rect 378 24863 450 24871
rect 468 24868 473 24902
rect 428 24833 430 24849
rect 251 24757 292 24785
rect 12 24752 62 24754
rect 28 24743 59 24745
rect 62 24743 64 24752
rect 251 24751 263 24757
rect 28 24735 64 24743
rect 127 24743 158 24745
rect 127 24736 182 24743
rect 127 24735 161 24736
rect 59 24719 64 24735
rect 158 24719 161 24735
rect 253 24723 263 24751
rect 273 24723 292 24757
rect 318 24764 324 24833
rect 318 24754 335 24764
rect 303 24732 316 24748
rect 28 24711 64 24719
rect 127 24718 161 24719
rect 127 24711 182 24718
rect 62 24702 64 24711
rect 282 24665 292 24723
rect 303 24714 316 24730
rect 318 24701 324 24754
rect 346 24748 348 24833
rect 400 24825 430 24833
rect 476 24831 480 24899
rect 511 24868 582 24902
rect 544 24861 548 24868
rect 400 24821 434 24825
rect 400 24791 408 24821
rect 420 24791 434 24821
rect 544 24823 548 24831
rect 333 24714 353 24748
rect 428 24744 430 24791
rect 476 24751 480 24819
rect 544 24789 552 24823
rect 578 24789 582 24823
rect 544 24781 548 24789
rect 346 24701 348 24714
rect 367 24710 380 24744
rect 396 24710 408 24744
rect 420 24710 434 24744
rect 544 24741 553 24769
rect 319 24698 335 24700
rect 120 24649 170 24651
rect 76 24643 92 24649
rect 94 24643 110 24649
rect 76 24633 99 24642
rect 60 24623 67 24633
rect 76 24613 77 24633
rect 96 24608 99 24633
rect 109 24613 110 24633
rect 119 24623 126 24633
rect 76 24599 110 24603
rect 170 24599 172 24649
rect 186 24631 190 24665
rect 216 24631 220 24665
rect 182 24593 224 24594
rect 186 24552 220 24586
rect 223 24552 257 24586
rect 160 24545 182 24551
rect 224 24545 246 24551
rect 288 24545 292 24665
rect 296 24663 368 24671
rect 428 24663 430 24710
rect 476 24673 480 24741
rect 485 24697 495 24731
rect 505 24697 519 24731
rect 544 24697 555 24741
rect 485 24673 492 24697
rect 579 24682 582 24772
rect 599 24752 649 24754
rect 610 24744 624 24745
rect 607 24743 624 24744
rect 586 24736 644 24743
rect 607 24735 644 24736
rect 607 24719 610 24735
rect 616 24719 644 24735
rect 607 24718 644 24719
rect 586 24711 644 24718
rect 607 24710 610 24711
rect 649 24702 651 24752
rect 544 24665 548 24673
rect 400 24633 408 24663
rect 420 24633 434 24663
rect 400 24629 434 24633
rect 400 24621 430 24629
rect 428 24605 430 24621
rect 476 24593 480 24661
rect 544 24631 552 24665
rect 578 24631 582 24665
rect 544 24623 548 24631
rect 295 24552 300 24586
rect 324 24552 329 24586
rect 378 24583 450 24591
rect 544 24588 548 24593
rect 544 24584 582 24588
rect 544 24554 552 24584
rect 578 24554 582 24584
rect 544 24551 548 24554
rect 522 24545 548 24551
rect 586 24545 608 24551
rect 182 24529 224 24545
rect 544 24529 586 24545
rect 17 24515 67 24517
rect 119 24515 169 24517
rect 599 24515 649 24517
rect 42 24473 59 24507
rect 67 24465 69 24515
rect 160 24507 246 24515
rect 522 24507 608 24515
rect 76 24473 110 24507
rect 127 24473 144 24507
rect 152 24473 161 24507
rect 162 24505 195 24507
rect 224 24505 244 24507
rect 162 24473 244 24505
rect 524 24505 548 24507
rect 573 24505 582 24507
rect 586 24505 606 24507
rect 160 24465 246 24473
rect 186 24449 220 24451
rect 182 24435 224 24436
rect 160 24429 182 24435
rect 224 24429 246 24435
rect 186 24394 220 24428
rect 223 24394 257 24428
rect 120 24381 170 24383
rect 76 24377 130 24381
rect 110 24372 130 24377
rect 60 24347 67 24357
rect 76 24347 77 24367
rect 96 24338 99 24372
rect 109 24347 110 24367
rect 119 24347 126 24357
rect 76 24331 92 24337
rect 94 24331 110 24337
rect 170 24331 172 24381
rect 186 24315 190 24349
rect 216 24315 220 24349
rect 288 24315 292 24503
rect 476 24435 480 24503
rect 524 24473 606 24505
rect 607 24473 616 24507
rect 522 24465 608 24473
rect 649 24465 651 24515
rect 548 24449 582 24451
rect 522 24430 548 24435
rect 522 24429 582 24430
rect 586 24429 608 24435
rect 295 24394 300 24428
rect 324 24394 329 24428
rect 544 24426 582 24429
rect 378 24389 450 24397
rect 428 24359 430 24375
rect 400 24351 430 24359
rect 476 24357 480 24425
rect 544 24396 552 24426
rect 578 24396 582 24426
rect 544 24387 548 24396
rect 400 24347 434 24351
rect 400 24317 408 24347
rect 420 24317 434 24347
rect 544 24349 548 24357
rect 12 24278 62 24280
rect 28 24269 59 24271
rect 62 24269 64 24278
rect 28 24261 64 24269
rect 127 24269 158 24271
rect 127 24262 182 24269
rect 215 24267 224 24295
rect 127 24261 161 24262
rect 59 24245 64 24261
rect 158 24245 161 24261
rect 28 24237 64 24245
rect 127 24244 161 24245
rect 127 24237 182 24244
rect 62 24228 64 24237
rect 213 24229 224 24267
rect 282 24257 292 24315
rect 296 24309 368 24317
rect 319 24280 335 24282
rect 251 24223 263 24257
rect 273 24223 292 24257
rect 303 24250 316 24266
rect 303 24232 316 24248
rect 120 24175 170 24177
rect 76 24169 92 24175
rect 94 24169 110 24175
rect 76 24159 99 24168
rect 60 24149 67 24159
rect 76 24139 77 24159
rect 96 24134 99 24159
rect 109 24139 110 24159
rect 119 24149 126 24159
rect 76 24125 110 24129
rect 170 24125 172 24175
rect 186 24157 190 24191
rect 216 24157 220 24191
rect 186 24080 220 24114
rect 282 24111 292 24223
rect 318 24226 324 24279
rect 346 24266 348 24279
rect 428 24270 430 24317
rect 443 24307 450 24309
rect 476 24277 480 24345
rect 544 24315 552 24349
rect 578 24315 582 24349
rect 481 24283 517 24311
rect 481 24277 495 24283
rect 333 24232 353 24266
rect 367 24236 380 24270
rect 396 24236 408 24270
rect 420 24236 434 24270
rect 318 24216 335 24226
rect 318 24147 324 24216
rect 346 24147 348 24232
rect 428 24189 430 24236
rect 476 24199 480 24267
rect 485 24249 495 24277
rect 505 24249 519 24283
rect 544 24277 555 24315
rect 544 24249 553 24277
rect 544 24229 548 24249
rect 579 24208 582 24298
rect 599 24278 649 24280
rect 610 24270 624 24271
rect 607 24269 624 24270
rect 586 24262 644 24269
rect 607 24261 644 24262
rect 607 24245 610 24261
rect 616 24245 644 24261
rect 607 24244 644 24245
rect 586 24237 644 24244
rect 607 24236 610 24237
rect 649 24228 651 24278
rect 544 24191 548 24199
rect 400 24159 408 24189
rect 420 24159 434 24189
rect 400 24155 434 24159
rect 400 24147 430 24155
rect 428 24131 430 24147
rect 476 24119 480 24187
rect 544 24157 552 24191
rect 578 24157 582 24191
rect 544 24149 548 24157
rect 544 24119 586 24120
rect 288 24079 292 24111
rect 296 24109 368 24117
rect 378 24109 450 24117
rect 544 24112 548 24119
rect 439 24081 444 24109
rect 120 24065 170 24067
rect 76 24061 130 24065
rect 110 24056 130 24061
rect 60 24031 67 24041
rect 76 24031 77 24051
rect 96 24022 99 24056
rect 109 24031 110 24051
rect 119 24031 126 24041
rect 76 24015 92 24021
rect 94 24015 110 24021
rect 170 24015 172 24065
rect 186 23999 190 24033
rect 216 23999 220 24033
rect 213 23967 224 23999
rect 282 23995 292 24079
rect 296 24073 368 24081
rect 378 24073 450 24081
rect 468 24078 473 24112
rect 428 24043 430 24059
rect 251 23967 292 23995
rect 12 23962 62 23964
rect 28 23953 59 23955
rect 62 23953 64 23962
rect 251 23961 263 23967
rect 28 23945 64 23953
rect 127 23953 158 23955
rect 127 23946 182 23953
rect 127 23945 161 23946
rect 59 23929 64 23945
rect 158 23929 161 23945
rect 253 23933 263 23961
rect 273 23933 292 23967
rect 318 23974 324 24043
rect 318 23964 335 23974
rect 303 23942 316 23958
rect 28 23921 64 23929
rect 127 23928 161 23929
rect 127 23921 182 23928
rect 62 23912 64 23921
rect 282 23875 292 23933
rect 303 23924 316 23940
rect 318 23911 324 23964
rect 346 23958 348 24043
rect 400 24035 430 24043
rect 476 24041 480 24109
rect 511 24078 582 24112
rect 544 24071 548 24078
rect 400 24031 434 24035
rect 400 24001 408 24031
rect 420 24001 434 24031
rect 544 24033 548 24041
rect 333 23924 353 23958
rect 428 23954 430 24001
rect 476 23961 480 24029
rect 544 23999 552 24033
rect 578 23999 582 24033
rect 544 23991 548 23999
rect 346 23911 348 23924
rect 367 23920 380 23954
rect 396 23920 408 23954
rect 420 23920 434 23954
rect 544 23951 553 23979
rect 319 23908 335 23910
rect 120 23859 170 23861
rect 76 23853 92 23859
rect 94 23853 110 23859
rect 76 23843 99 23852
rect 60 23833 67 23843
rect 76 23823 77 23843
rect 96 23818 99 23843
rect 109 23823 110 23843
rect 119 23833 126 23843
rect 76 23809 110 23813
rect 170 23809 172 23859
rect 186 23841 190 23875
rect 216 23841 220 23875
rect 182 23803 224 23804
rect 186 23762 220 23796
rect 223 23762 257 23796
rect 160 23755 182 23761
rect 224 23755 246 23761
rect 288 23755 292 23875
rect 296 23873 368 23881
rect 428 23873 430 23920
rect 476 23883 480 23951
rect 485 23907 495 23941
rect 505 23907 519 23941
rect 544 23907 555 23951
rect 485 23883 492 23907
rect 579 23892 582 23982
rect 599 23962 649 23964
rect 610 23954 624 23955
rect 607 23953 624 23954
rect 586 23946 644 23953
rect 607 23945 644 23946
rect 607 23929 610 23945
rect 616 23929 644 23945
rect 607 23928 644 23929
rect 586 23921 644 23928
rect 607 23920 610 23921
rect 649 23912 651 23962
rect 544 23875 548 23883
rect 400 23843 408 23873
rect 420 23843 434 23873
rect 400 23839 434 23843
rect 400 23831 430 23839
rect 428 23815 430 23831
rect 476 23803 480 23871
rect 544 23841 552 23875
rect 578 23841 582 23875
rect 544 23833 548 23841
rect 295 23762 300 23796
rect 324 23762 329 23796
rect 378 23793 450 23801
rect 544 23798 548 23803
rect 544 23794 582 23798
rect 544 23764 552 23794
rect 578 23764 582 23794
rect 544 23761 548 23764
rect 522 23755 548 23761
rect 586 23755 608 23761
rect 182 23739 224 23755
rect 544 23739 586 23755
rect 17 23725 67 23727
rect 119 23725 169 23727
rect 599 23725 649 23727
rect 42 23683 59 23717
rect 67 23675 69 23725
rect 160 23717 246 23725
rect 522 23717 608 23725
rect 76 23683 110 23717
rect 127 23683 144 23717
rect 152 23683 161 23717
rect 162 23715 195 23717
rect 224 23715 244 23717
rect 162 23683 244 23715
rect 524 23715 548 23717
rect 573 23715 582 23717
rect 586 23715 606 23717
rect 160 23675 246 23683
rect 186 23659 220 23661
rect 182 23645 224 23646
rect 160 23639 182 23645
rect 224 23639 246 23645
rect 186 23604 220 23638
rect 223 23604 257 23638
rect 120 23591 170 23593
rect 76 23587 130 23591
rect 110 23582 130 23587
rect 60 23557 67 23567
rect 76 23557 77 23577
rect 96 23548 99 23582
rect 109 23557 110 23577
rect 119 23557 126 23567
rect 76 23541 92 23547
rect 94 23541 110 23547
rect 170 23541 172 23591
rect 186 23525 190 23559
rect 216 23525 220 23559
rect 288 23525 292 23713
rect 476 23645 480 23713
rect 524 23683 606 23715
rect 607 23683 616 23717
rect 522 23675 608 23683
rect 649 23675 651 23725
rect 548 23659 582 23661
rect 522 23640 548 23645
rect 522 23639 582 23640
rect 586 23639 608 23645
rect 295 23604 300 23638
rect 324 23604 329 23638
rect 544 23636 582 23639
rect 378 23599 450 23607
rect 428 23569 430 23585
rect 400 23561 430 23569
rect 476 23567 480 23635
rect 544 23606 552 23636
rect 578 23606 582 23636
rect 544 23597 548 23606
rect 400 23557 434 23561
rect 400 23527 408 23557
rect 420 23527 434 23557
rect 544 23559 548 23567
rect 12 23488 62 23490
rect 28 23479 59 23481
rect 62 23479 64 23488
rect 28 23471 64 23479
rect 127 23479 158 23481
rect 127 23472 182 23479
rect 215 23477 224 23505
rect 127 23471 161 23472
rect 59 23455 64 23471
rect 158 23455 161 23471
rect 28 23447 64 23455
rect 127 23454 161 23455
rect 127 23447 182 23454
rect 62 23438 64 23447
rect 213 23439 224 23477
rect 282 23467 292 23525
rect 296 23519 368 23527
rect 319 23490 335 23492
rect 251 23433 263 23467
rect 273 23433 292 23467
rect 303 23460 316 23476
rect 303 23442 316 23458
rect 120 23385 170 23387
rect 76 23379 92 23385
rect 94 23379 110 23385
rect 76 23369 99 23378
rect 60 23359 67 23369
rect 76 23349 77 23369
rect 96 23344 99 23369
rect 109 23349 110 23369
rect 119 23359 126 23369
rect 76 23335 110 23339
rect 170 23335 172 23385
rect 186 23367 190 23401
rect 216 23367 220 23401
rect 186 23290 220 23324
rect 282 23321 292 23433
rect 318 23436 324 23489
rect 346 23476 348 23489
rect 428 23480 430 23527
rect 443 23517 450 23519
rect 476 23487 480 23555
rect 544 23525 552 23559
rect 578 23525 582 23559
rect 481 23493 517 23521
rect 481 23487 495 23493
rect 333 23442 353 23476
rect 367 23446 380 23480
rect 396 23446 408 23480
rect 420 23446 434 23480
rect 318 23426 335 23436
rect 318 23357 324 23426
rect 346 23357 348 23442
rect 428 23399 430 23446
rect 476 23409 480 23477
rect 485 23459 495 23487
rect 505 23459 519 23493
rect 544 23487 555 23525
rect 544 23459 553 23487
rect 544 23439 548 23459
rect 579 23418 582 23508
rect 599 23488 649 23490
rect 610 23480 624 23481
rect 607 23479 624 23480
rect 586 23472 644 23479
rect 607 23471 644 23472
rect 607 23455 610 23471
rect 616 23455 644 23471
rect 607 23454 644 23455
rect 586 23447 644 23454
rect 607 23446 610 23447
rect 649 23438 651 23488
rect 544 23401 548 23409
rect 400 23369 408 23399
rect 420 23369 434 23399
rect 400 23365 434 23369
rect 400 23357 430 23365
rect 428 23341 430 23357
rect 476 23329 480 23397
rect 544 23367 552 23401
rect 578 23367 582 23401
rect 544 23359 548 23367
rect 544 23329 586 23330
rect 288 23289 292 23321
rect 296 23319 368 23327
rect 378 23319 450 23327
rect 544 23322 548 23329
rect 439 23291 444 23319
rect 120 23275 170 23277
rect 76 23271 130 23275
rect 110 23266 130 23271
rect 60 23241 67 23251
rect 76 23241 77 23261
rect 96 23232 99 23266
rect 109 23241 110 23261
rect 119 23241 126 23251
rect 76 23225 92 23231
rect 94 23225 110 23231
rect 170 23225 172 23275
rect 186 23209 190 23243
rect 216 23209 220 23243
rect 213 23177 224 23209
rect 282 23205 292 23289
rect 296 23283 368 23291
rect 378 23283 450 23291
rect 468 23288 473 23322
rect 428 23253 430 23269
rect 251 23177 292 23205
rect 12 23172 62 23174
rect 28 23163 59 23165
rect 62 23163 64 23172
rect 251 23171 263 23177
rect 28 23155 64 23163
rect 127 23163 158 23165
rect 127 23156 182 23163
rect 127 23155 161 23156
rect 59 23139 64 23155
rect 158 23139 161 23155
rect 253 23143 263 23171
rect 273 23143 292 23177
rect 318 23184 324 23253
rect 318 23174 335 23184
rect 303 23152 316 23168
rect 28 23131 64 23139
rect 127 23138 161 23139
rect 127 23131 182 23138
rect 62 23122 64 23131
rect 282 23085 292 23143
rect 303 23134 316 23150
rect 318 23121 324 23174
rect 346 23168 348 23253
rect 400 23245 430 23253
rect 476 23251 480 23319
rect 511 23288 582 23322
rect 544 23281 548 23288
rect 400 23241 434 23245
rect 400 23211 408 23241
rect 420 23211 434 23241
rect 544 23243 548 23251
rect 333 23134 353 23168
rect 428 23164 430 23211
rect 476 23171 480 23239
rect 544 23209 552 23243
rect 578 23209 582 23243
rect 544 23201 548 23209
rect 346 23121 348 23134
rect 367 23130 380 23164
rect 396 23130 408 23164
rect 420 23130 434 23164
rect 544 23161 553 23189
rect 319 23118 335 23120
rect 120 23069 170 23071
rect 76 23063 92 23069
rect 94 23063 110 23069
rect 76 23053 99 23062
rect 60 23043 67 23053
rect 76 23033 77 23053
rect 96 23028 99 23053
rect 109 23033 110 23053
rect 119 23043 126 23053
rect 76 23019 110 23023
rect 170 23019 172 23069
rect 186 23051 190 23085
rect 216 23051 220 23085
rect 182 23013 224 23014
rect 186 22972 220 23006
rect 223 22972 257 23006
rect 160 22965 182 22971
rect 224 22965 246 22971
rect 288 22965 292 23085
rect 296 23083 368 23091
rect 428 23083 430 23130
rect 476 23093 480 23161
rect 485 23117 495 23151
rect 505 23117 519 23151
rect 544 23117 555 23161
rect 485 23093 492 23117
rect 579 23102 582 23192
rect 599 23172 649 23174
rect 610 23164 624 23165
rect 607 23163 624 23164
rect 586 23156 644 23163
rect 607 23155 644 23156
rect 607 23139 610 23155
rect 616 23139 644 23155
rect 607 23138 644 23139
rect 586 23131 644 23138
rect 607 23130 610 23131
rect 649 23122 651 23172
rect 544 23085 548 23093
rect 400 23053 408 23083
rect 420 23053 434 23083
rect 400 23049 434 23053
rect 400 23041 430 23049
rect 428 23025 430 23041
rect 476 23013 480 23081
rect 544 23051 552 23085
rect 578 23051 582 23085
rect 544 23043 548 23051
rect 295 22972 300 23006
rect 324 22972 329 23006
rect 378 23003 450 23011
rect 544 23008 548 23013
rect 544 23004 582 23008
rect 544 22974 552 23004
rect 578 22974 582 23004
rect 544 22971 548 22974
rect 522 22965 548 22971
rect 586 22965 608 22971
rect 182 22949 224 22965
rect 544 22949 586 22965
rect 17 22935 67 22937
rect 119 22935 169 22937
rect 599 22935 649 22937
rect 42 22893 59 22927
rect 67 22885 69 22935
rect 160 22927 246 22935
rect 522 22927 608 22935
rect 76 22893 110 22927
rect 127 22893 144 22927
rect 152 22893 161 22927
rect 162 22925 195 22927
rect 224 22925 244 22927
rect 162 22893 244 22925
rect 524 22925 548 22927
rect 573 22925 582 22927
rect 586 22925 606 22927
rect 160 22885 246 22893
rect 186 22869 220 22871
rect 182 22855 224 22856
rect 160 22849 182 22855
rect 224 22849 246 22855
rect 186 22814 220 22848
rect 223 22814 257 22848
rect 120 22801 170 22803
rect 76 22797 130 22801
rect 110 22792 130 22797
rect 60 22767 67 22777
rect 76 22767 77 22787
rect 96 22758 99 22792
rect 109 22767 110 22787
rect 119 22767 126 22777
rect 76 22751 92 22757
rect 94 22751 110 22757
rect 170 22751 172 22801
rect 186 22735 190 22769
rect 216 22735 220 22769
rect 288 22735 292 22923
rect 476 22855 480 22923
rect 524 22893 606 22925
rect 607 22893 616 22927
rect 522 22885 608 22893
rect 649 22885 651 22935
rect 548 22869 582 22871
rect 522 22850 548 22855
rect 522 22849 582 22850
rect 586 22849 608 22855
rect 295 22814 300 22848
rect 324 22814 329 22848
rect 544 22846 582 22849
rect 378 22809 450 22817
rect 428 22779 430 22795
rect 400 22771 430 22779
rect 476 22777 480 22845
rect 544 22816 552 22846
rect 578 22816 582 22846
rect 544 22807 548 22816
rect 400 22767 434 22771
rect 400 22737 408 22767
rect 420 22737 434 22767
rect 544 22769 548 22777
rect 12 22698 62 22700
rect 28 22689 59 22691
rect 62 22689 64 22698
rect 28 22681 64 22689
rect 127 22689 158 22691
rect 127 22682 182 22689
rect 215 22687 224 22715
rect 127 22681 161 22682
rect 59 22665 64 22681
rect 158 22665 161 22681
rect 28 22657 64 22665
rect 127 22664 161 22665
rect 127 22657 182 22664
rect 62 22648 64 22657
rect 213 22649 224 22687
rect 282 22677 292 22735
rect 296 22729 368 22737
rect 319 22700 335 22702
rect 251 22643 263 22677
rect 273 22643 292 22677
rect 303 22670 316 22686
rect 303 22652 316 22668
rect 120 22595 170 22597
rect 76 22589 92 22595
rect 94 22589 110 22595
rect 76 22579 99 22588
rect 60 22569 67 22579
rect 76 22559 77 22579
rect 96 22554 99 22579
rect 109 22559 110 22579
rect 119 22569 126 22579
rect 76 22545 110 22549
rect 170 22545 172 22595
rect 186 22577 190 22611
rect 216 22577 220 22611
rect 186 22500 220 22534
rect 282 22531 292 22643
rect 318 22646 324 22699
rect 346 22686 348 22699
rect 428 22690 430 22737
rect 443 22727 450 22729
rect 476 22697 480 22765
rect 544 22735 552 22769
rect 578 22735 582 22769
rect 481 22703 517 22731
rect 481 22697 495 22703
rect 333 22652 353 22686
rect 367 22656 380 22690
rect 396 22656 408 22690
rect 420 22656 434 22690
rect 318 22636 335 22646
rect 318 22567 324 22636
rect 346 22567 348 22652
rect 428 22609 430 22656
rect 476 22619 480 22687
rect 485 22669 495 22697
rect 505 22669 519 22703
rect 544 22697 555 22735
rect 544 22669 553 22697
rect 544 22649 548 22669
rect 579 22628 582 22718
rect 599 22698 649 22700
rect 610 22690 624 22691
rect 607 22689 624 22690
rect 586 22682 644 22689
rect 607 22681 644 22682
rect 607 22665 610 22681
rect 616 22665 644 22681
rect 607 22664 644 22665
rect 586 22657 644 22664
rect 607 22656 610 22657
rect 649 22648 651 22698
rect 544 22611 548 22619
rect 400 22579 408 22609
rect 420 22579 434 22609
rect 400 22575 434 22579
rect 400 22567 430 22575
rect 428 22551 430 22567
rect 476 22539 480 22607
rect 544 22577 552 22611
rect 578 22577 582 22611
rect 544 22569 548 22577
rect 544 22539 586 22540
rect 288 22499 292 22531
rect 296 22529 368 22537
rect 378 22529 450 22537
rect 544 22532 548 22539
rect 439 22501 444 22529
rect 120 22485 170 22487
rect 76 22481 130 22485
rect 110 22476 130 22481
rect 60 22451 67 22461
rect 76 22451 77 22471
rect 96 22442 99 22476
rect 109 22451 110 22471
rect 119 22451 126 22461
rect 76 22435 92 22441
rect 94 22435 110 22441
rect 170 22435 172 22485
rect 186 22419 190 22453
rect 216 22419 220 22453
rect 213 22387 224 22419
rect 282 22415 292 22499
rect 296 22493 368 22501
rect 378 22493 450 22501
rect 468 22498 473 22532
rect 428 22463 430 22479
rect 251 22387 292 22415
rect 12 22382 62 22384
rect 28 22373 59 22375
rect 62 22373 64 22382
rect 251 22381 263 22387
rect 28 22365 64 22373
rect 127 22373 158 22375
rect 127 22366 182 22373
rect 127 22365 161 22366
rect 59 22349 64 22365
rect 158 22349 161 22365
rect 253 22353 263 22381
rect 273 22353 292 22387
rect 318 22394 324 22463
rect 318 22384 335 22394
rect 303 22362 316 22378
rect 28 22341 64 22349
rect 127 22348 161 22349
rect 127 22341 182 22348
rect 62 22332 64 22341
rect 282 22295 292 22353
rect 303 22344 316 22360
rect 318 22331 324 22384
rect 346 22378 348 22463
rect 400 22455 430 22463
rect 476 22461 480 22529
rect 511 22498 582 22532
rect 544 22491 548 22498
rect 400 22451 434 22455
rect 400 22421 408 22451
rect 420 22421 434 22451
rect 544 22453 548 22461
rect 333 22344 353 22378
rect 428 22374 430 22421
rect 476 22381 480 22449
rect 544 22419 552 22453
rect 578 22419 582 22453
rect 544 22411 548 22419
rect 346 22331 348 22344
rect 367 22340 380 22374
rect 396 22340 408 22374
rect 420 22340 434 22374
rect 544 22371 553 22399
rect 319 22328 335 22330
rect 120 22279 170 22281
rect 76 22273 92 22279
rect 94 22273 110 22279
rect 76 22263 99 22272
rect 60 22253 67 22263
rect 76 22243 77 22263
rect 96 22238 99 22263
rect 109 22243 110 22263
rect 119 22253 126 22263
rect 76 22229 110 22233
rect 170 22229 172 22279
rect 186 22261 190 22295
rect 216 22261 220 22295
rect 182 22223 224 22224
rect 186 22182 220 22216
rect 223 22182 257 22216
rect 160 22175 182 22181
rect 224 22175 246 22181
rect 288 22175 292 22295
rect 296 22293 368 22301
rect 428 22293 430 22340
rect 476 22303 480 22371
rect 485 22327 495 22361
rect 505 22327 519 22361
rect 544 22327 555 22371
rect 485 22303 492 22327
rect 579 22312 582 22402
rect 599 22382 649 22384
rect 610 22374 624 22375
rect 607 22373 624 22374
rect 586 22366 644 22373
rect 607 22365 644 22366
rect 607 22349 610 22365
rect 616 22349 644 22365
rect 607 22348 644 22349
rect 586 22341 644 22348
rect 607 22340 610 22341
rect 649 22332 651 22382
rect 544 22295 548 22303
rect 400 22263 408 22293
rect 420 22263 434 22293
rect 400 22259 434 22263
rect 400 22251 430 22259
rect 428 22235 430 22251
rect 476 22223 480 22291
rect 544 22261 552 22295
rect 578 22261 582 22295
rect 544 22253 548 22261
rect 295 22182 300 22216
rect 324 22182 329 22216
rect 378 22213 450 22221
rect 544 22218 548 22223
rect 544 22214 582 22218
rect 544 22184 552 22214
rect 578 22184 582 22214
rect 544 22181 548 22184
rect 522 22175 548 22181
rect 586 22175 608 22181
rect 182 22159 224 22175
rect 544 22159 586 22175
rect 17 22145 67 22147
rect 119 22145 169 22147
rect 599 22145 649 22147
rect 42 22103 59 22137
rect 67 22095 69 22145
rect 160 22137 246 22145
rect 522 22137 608 22145
rect 76 22103 110 22137
rect 127 22103 144 22137
rect 152 22103 161 22137
rect 162 22135 195 22137
rect 224 22135 244 22137
rect 162 22103 244 22135
rect 524 22135 548 22137
rect 573 22135 582 22137
rect 586 22135 606 22137
rect 160 22095 246 22103
rect 186 22079 220 22081
rect 182 22065 224 22066
rect 160 22059 182 22065
rect 224 22059 246 22065
rect 186 22024 220 22058
rect 223 22024 257 22058
rect 120 22011 170 22013
rect 76 22007 130 22011
rect 110 22002 130 22007
rect 60 21977 67 21987
rect 76 21977 77 21997
rect 96 21968 99 22002
rect 109 21977 110 21997
rect 119 21977 126 21987
rect 76 21961 92 21967
rect 94 21961 110 21967
rect 170 21961 172 22011
rect 186 21945 190 21979
rect 216 21945 220 21979
rect 288 21945 292 22133
rect 476 22065 480 22133
rect 524 22103 606 22135
rect 607 22103 616 22137
rect 522 22095 608 22103
rect 649 22095 651 22145
rect 548 22079 582 22081
rect 522 22060 548 22065
rect 522 22059 582 22060
rect 586 22059 608 22065
rect 295 22024 300 22058
rect 324 22024 329 22058
rect 544 22056 582 22059
rect 378 22019 450 22027
rect 428 21989 430 22005
rect 400 21981 430 21989
rect 476 21987 480 22055
rect 544 22026 552 22056
rect 578 22026 582 22056
rect 544 22017 548 22026
rect 400 21977 434 21981
rect 400 21947 408 21977
rect 420 21947 434 21977
rect 544 21979 548 21987
rect 12 21908 62 21910
rect 28 21899 59 21901
rect 62 21899 64 21908
rect 28 21891 64 21899
rect 127 21899 158 21901
rect 127 21892 182 21899
rect 215 21897 224 21925
rect 127 21891 161 21892
rect 59 21875 64 21891
rect 158 21875 161 21891
rect 28 21867 64 21875
rect 127 21874 161 21875
rect 127 21867 182 21874
rect 62 21858 64 21867
rect 213 21859 224 21897
rect 282 21887 292 21945
rect 296 21939 368 21947
rect 319 21910 335 21912
rect 251 21853 263 21887
rect 273 21853 292 21887
rect 303 21880 316 21896
rect 303 21862 316 21878
rect 120 21805 170 21807
rect 76 21799 92 21805
rect 94 21799 110 21805
rect 76 21789 99 21798
rect 60 21779 67 21789
rect 76 21769 77 21789
rect 96 21764 99 21789
rect 109 21769 110 21789
rect 119 21779 126 21789
rect 76 21755 110 21759
rect 170 21755 172 21805
rect 186 21787 190 21821
rect 216 21787 220 21821
rect 186 21710 220 21744
rect 282 21741 292 21853
rect 318 21856 324 21909
rect 346 21896 348 21909
rect 428 21900 430 21947
rect 443 21937 450 21939
rect 476 21907 480 21975
rect 544 21945 552 21979
rect 578 21945 582 21979
rect 481 21913 517 21941
rect 481 21907 495 21913
rect 333 21862 353 21896
rect 367 21866 380 21900
rect 396 21866 408 21900
rect 420 21866 434 21900
rect 318 21846 335 21856
rect 318 21777 324 21846
rect 346 21777 348 21862
rect 428 21819 430 21866
rect 476 21829 480 21897
rect 485 21879 495 21907
rect 505 21879 519 21913
rect 544 21907 555 21945
rect 544 21879 553 21907
rect 544 21859 548 21879
rect 579 21838 582 21928
rect 599 21908 649 21910
rect 610 21900 624 21901
rect 607 21899 624 21900
rect 586 21892 644 21899
rect 607 21891 644 21892
rect 607 21875 610 21891
rect 616 21875 644 21891
rect 607 21874 644 21875
rect 586 21867 644 21874
rect 607 21866 610 21867
rect 649 21858 651 21908
rect 544 21821 548 21829
rect 400 21789 408 21819
rect 420 21789 434 21819
rect 400 21785 434 21789
rect 400 21777 430 21785
rect 428 21761 430 21777
rect 476 21749 480 21817
rect 544 21787 552 21821
rect 578 21787 582 21821
rect 544 21779 548 21787
rect 544 21749 586 21750
rect 288 21709 292 21741
rect 296 21739 368 21747
rect 378 21739 450 21747
rect 544 21742 548 21749
rect 439 21711 444 21739
rect 120 21695 170 21697
rect 76 21691 130 21695
rect 110 21686 130 21691
rect 60 21661 67 21671
rect 76 21661 77 21681
rect 96 21652 99 21686
rect 109 21661 110 21681
rect 119 21661 126 21671
rect 76 21645 92 21651
rect 94 21645 110 21651
rect 170 21645 172 21695
rect 186 21629 190 21663
rect 216 21629 220 21663
rect 213 21597 224 21629
rect 282 21625 292 21709
rect 296 21703 368 21711
rect 378 21703 450 21711
rect 468 21708 473 21742
rect 428 21673 430 21689
rect 251 21597 292 21625
rect 12 21592 62 21594
rect 28 21583 59 21585
rect 62 21583 64 21592
rect 251 21591 263 21597
rect 28 21575 64 21583
rect 127 21583 158 21585
rect 127 21576 182 21583
rect 127 21575 161 21576
rect 59 21559 64 21575
rect 158 21559 161 21575
rect 253 21563 263 21591
rect 273 21563 292 21597
rect 318 21604 324 21673
rect 318 21594 335 21604
rect 303 21572 316 21588
rect 28 21551 64 21559
rect 127 21558 161 21559
rect 127 21551 182 21558
rect 62 21542 64 21551
rect 282 21505 292 21563
rect 303 21554 316 21570
rect 318 21541 324 21594
rect 346 21588 348 21673
rect 400 21665 430 21673
rect 476 21671 480 21739
rect 511 21708 582 21742
rect 544 21701 548 21708
rect 400 21661 434 21665
rect 400 21631 408 21661
rect 420 21631 434 21661
rect 544 21663 548 21671
rect 333 21554 353 21588
rect 428 21584 430 21631
rect 476 21591 480 21659
rect 544 21629 552 21663
rect 578 21629 582 21663
rect 544 21621 548 21629
rect 346 21541 348 21554
rect 367 21550 380 21584
rect 396 21550 408 21584
rect 420 21550 434 21584
rect 544 21581 553 21609
rect 319 21538 335 21540
rect 120 21489 170 21491
rect 76 21483 92 21489
rect 94 21483 110 21489
rect 76 21473 99 21482
rect 60 21463 67 21473
rect 76 21453 77 21473
rect 96 21448 99 21473
rect 109 21453 110 21473
rect 119 21463 126 21473
rect 76 21439 110 21443
rect 170 21439 172 21489
rect 186 21471 190 21505
rect 216 21471 220 21505
rect 182 21433 224 21434
rect 186 21392 220 21426
rect 223 21392 257 21426
rect 160 21385 182 21391
rect 224 21385 246 21391
rect 288 21385 292 21505
rect 296 21503 368 21511
rect 428 21503 430 21550
rect 476 21513 480 21581
rect 485 21537 495 21571
rect 505 21537 519 21571
rect 544 21537 555 21581
rect 485 21513 492 21537
rect 579 21522 582 21612
rect 599 21592 649 21594
rect 610 21584 624 21585
rect 607 21583 624 21584
rect 586 21576 644 21583
rect 607 21575 644 21576
rect 607 21559 610 21575
rect 616 21559 644 21575
rect 607 21558 644 21559
rect 586 21551 644 21558
rect 607 21550 610 21551
rect 649 21542 651 21592
rect 544 21505 548 21513
rect 400 21473 408 21503
rect 420 21473 434 21503
rect 400 21469 434 21473
rect 400 21461 430 21469
rect 428 21445 430 21461
rect 476 21433 480 21501
rect 544 21471 552 21505
rect 578 21471 582 21505
rect 544 21463 548 21471
rect 295 21392 300 21426
rect 324 21392 329 21426
rect 378 21423 450 21431
rect 544 21428 548 21433
rect 544 21424 582 21428
rect 544 21394 552 21424
rect 578 21394 582 21424
rect 544 21391 548 21394
rect 522 21385 548 21391
rect 586 21385 608 21391
rect 182 21369 224 21385
rect 544 21369 586 21385
rect 17 21355 67 21357
rect 119 21355 169 21357
rect 599 21355 649 21357
rect 42 21313 59 21347
rect 67 21305 69 21355
rect 160 21347 246 21355
rect 522 21347 608 21355
rect 76 21313 110 21347
rect 127 21313 144 21347
rect 152 21313 161 21347
rect 162 21345 195 21347
rect 224 21345 244 21347
rect 162 21313 244 21345
rect 524 21345 548 21347
rect 573 21345 582 21347
rect 586 21345 606 21347
rect 160 21305 246 21313
rect 186 21289 220 21291
rect 182 21275 224 21276
rect 160 21269 182 21275
rect 224 21269 246 21275
rect 186 21234 220 21268
rect 223 21234 257 21268
rect 120 21221 170 21223
rect 76 21217 130 21221
rect 110 21212 130 21217
rect 60 21187 67 21197
rect 76 21187 77 21207
rect 96 21178 99 21212
rect 109 21187 110 21207
rect 119 21187 126 21197
rect 76 21171 92 21177
rect 94 21171 110 21177
rect 170 21171 172 21221
rect 186 21155 190 21189
rect 216 21155 220 21189
rect 288 21155 292 21343
rect 476 21275 480 21343
rect 524 21313 606 21345
rect 607 21313 616 21347
rect 522 21305 608 21313
rect 649 21305 651 21355
rect 548 21289 582 21291
rect 522 21270 548 21275
rect 522 21269 582 21270
rect 586 21269 608 21275
rect 295 21234 300 21268
rect 324 21234 329 21268
rect 544 21266 582 21269
rect 378 21229 450 21237
rect 428 21199 430 21215
rect 400 21191 430 21199
rect 476 21197 480 21265
rect 544 21236 552 21266
rect 578 21236 582 21266
rect 544 21227 548 21236
rect 400 21187 434 21191
rect 400 21157 408 21187
rect 420 21157 434 21187
rect 544 21189 548 21197
rect 12 21118 62 21120
rect 28 21109 59 21111
rect 62 21109 64 21118
rect 28 21101 64 21109
rect 127 21109 158 21111
rect 127 21102 182 21109
rect 215 21107 224 21135
rect 127 21101 161 21102
rect 59 21085 64 21101
rect 158 21085 161 21101
rect 28 21077 64 21085
rect 127 21084 161 21085
rect 127 21077 182 21084
rect 62 21068 64 21077
rect 213 21069 224 21107
rect 282 21097 292 21155
rect 296 21149 368 21157
rect 319 21120 335 21122
rect 251 21063 263 21097
rect 273 21063 292 21097
rect 303 21090 316 21106
rect 303 21072 316 21088
rect 120 21015 170 21017
rect 76 21009 92 21015
rect 94 21009 110 21015
rect 76 20999 99 21008
rect 60 20989 67 20999
rect 76 20979 77 20999
rect 96 20974 99 20999
rect 109 20979 110 20999
rect 119 20989 126 20999
rect 76 20965 110 20969
rect 170 20965 172 21015
rect 186 20997 190 21031
rect 216 20997 220 21031
rect 186 20920 220 20954
rect 282 20951 292 21063
rect 318 21066 324 21119
rect 346 21106 348 21119
rect 428 21110 430 21157
rect 443 21147 450 21149
rect 476 21117 480 21185
rect 544 21155 552 21189
rect 578 21155 582 21189
rect 481 21123 517 21151
rect 481 21117 495 21123
rect 333 21072 353 21106
rect 367 21076 380 21110
rect 396 21076 408 21110
rect 420 21076 434 21110
rect 318 21056 335 21066
rect 318 20987 324 21056
rect 346 20987 348 21072
rect 428 21029 430 21076
rect 476 21039 480 21107
rect 485 21089 495 21117
rect 505 21089 519 21123
rect 544 21117 555 21155
rect 544 21089 553 21117
rect 544 21069 548 21089
rect 579 21048 582 21138
rect 599 21118 649 21120
rect 610 21110 624 21111
rect 607 21109 624 21110
rect 586 21102 644 21109
rect 607 21101 644 21102
rect 607 21085 610 21101
rect 616 21085 644 21101
rect 607 21084 644 21085
rect 586 21077 644 21084
rect 607 21076 610 21077
rect 649 21068 651 21118
rect 544 21031 548 21039
rect 400 20999 408 21029
rect 420 20999 434 21029
rect 400 20995 434 20999
rect 400 20987 430 20995
rect 428 20971 430 20987
rect 476 20959 480 21027
rect 544 20997 552 21031
rect 578 20997 582 21031
rect 544 20989 548 20997
rect 544 20959 586 20960
rect 288 20919 292 20951
rect 296 20949 368 20957
rect 378 20949 450 20957
rect 544 20952 548 20959
rect 439 20921 444 20949
rect 120 20905 170 20907
rect 76 20901 130 20905
rect 110 20896 130 20901
rect 60 20871 67 20881
rect 76 20871 77 20891
rect 96 20862 99 20896
rect 109 20871 110 20891
rect 119 20871 126 20881
rect 76 20855 92 20861
rect 94 20855 110 20861
rect 170 20855 172 20905
rect 186 20839 190 20873
rect 216 20839 220 20873
rect 213 20807 224 20839
rect 282 20835 292 20919
rect 296 20913 368 20921
rect 378 20913 450 20921
rect 468 20918 473 20952
rect 428 20883 430 20899
rect 251 20807 292 20835
rect 12 20802 62 20804
rect 28 20793 59 20795
rect 62 20793 64 20802
rect 251 20801 263 20807
rect 28 20785 64 20793
rect 127 20793 158 20795
rect 127 20786 182 20793
rect 127 20785 161 20786
rect 59 20769 64 20785
rect 158 20769 161 20785
rect 253 20773 263 20801
rect 273 20773 292 20807
rect 318 20814 324 20883
rect 318 20804 335 20814
rect 303 20782 316 20798
rect 28 20761 64 20769
rect 127 20768 161 20769
rect 127 20761 182 20768
rect 62 20752 64 20761
rect 282 20715 292 20773
rect 303 20764 316 20780
rect 318 20751 324 20804
rect 346 20798 348 20883
rect 400 20875 430 20883
rect 476 20881 480 20949
rect 511 20918 582 20952
rect 544 20911 548 20918
rect 400 20871 434 20875
rect 400 20841 408 20871
rect 420 20841 434 20871
rect 544 20873 548 20881
rect 333 20764 353 20798
rect 428 20794 430 20841
rect 476 20801 480 20869
rect 544 20839 552 20873
rect 578 20839 582 20873
rect 544 20831 548 20839
rect 346 20751 348 20764
rect 367 20760 380 20794
rect 396 20760 408 20794
rect 420 20760 434 20794
rect 544 20791 553 20819
rect 319 20748 335 20750
rect 120 20699 170 20701
rect 76 20693 92 20699
rect 94 20693 110 20699
rect 76 20683 99 20692
rect 60 20673 67 20683
rect 76 20663 77 20683
rect 96 20658 99 20683
rect 109 20663 110 20683
rect 119 20673 126 20683
rect 76 20649 110 20653
rect 170 20649 172 20699
rect 186 20681 190 20715
rect 216 20681 220 20715
rect 182 20643 224 20644
rect 186 20602 220 20636
rect 223 20602 257 20636
rect 160 20595 182 20601
rect 224 20595 246 20601
rect 288 20595 292 20715
rect 296 20713 368 20721
rect 428 20713 430 20760
rect 476 20723 480 20791
rect 485 20747 495 20781
rect 505 20747 519 20781
rect 544 20747 555 20791
rect 485 20723 492 20747
rect 579 20732 582 20822
rect 599 20802 649 20804
rect 610 20794 624 20795
rect 607 20793 624 20794
rect 586 20786 644 20793
rect 607 20785 644 20786
rect 607 20769 610 20785
rect 616 20769 644 20785
rect 607 20768 644 20769
rect 586 20761 644 20768
rect 607 20760 610 20761
rect 649 20752 651 20802
rect 544 20715 548 20723
rect 400 20683 408 20713
rect 420 20683 434 20713
rect 400 20679 434 20683
rect 400 20671 430 20679
rect 428 20655 430 20671
rect 476 20643 480 20711
rect 544 20681 552 20715
rect 578 20681 582 20715
rect 544 20673 548 20681
rect 295 20602 300 20636
rect 324 20602 329 20636
rect 378 20633 450 20641
rect 544 20638 548 20643
rect 544 20634 582 20638
rect 544 20604 552 20634
rect 578 20604 582 20634
rect 544 20601 548 20604
rect 522 20595 548 20601
rect 586 20595 608 20601
rect 182 20579 224 20595
rect 544 20579 586 20595
rect 17 20565 67 20567
rect 119 20565 169 20567
rect 599 20565 649 20567
rect 42 20523 59 20557
rect 67 20515 69 20565
rect 160 20557 246 20565
rect 522 20557 608 20565
rect 76 20523 110 20557
rect 127 20523 144 20557
rect 152 20523 161 20557
rect 162 20555 195 20557
rect 224 20555 244 20557
rect 162 20523 244 20555
rect 524 20555 548 20557
rect 573 20555 582 20557
rect 586 20555 606 20557
rect 160 20515 246 20523
rect 186 20499 220 20501
rect 182 20485 224 20486
rect 160 20479 182 20485
rect 224 20479 246 20485
rect 186 20444 220 20478
rect 223 20444 257 20478
rect 120 20431 170 20433
rect 76 20427 130 20431
rect 110 20422 130 20427
rect 60 20397 67 20407
rect 76 20397 77 20417
rect 96 20388 99 20422
rect 109 20397 110 20417
rect 119 20397 126 20407
rect 76 20381 92 20387
rect 94 20381 110 20387
rect 170 20381 172 20431
rect 186 20365 190 20399
rect 216 20365 220 20399
rect 288 20365 292 20553
rect 476 20485 480 20553
rect 524 20523 606 20555
rect 607 20523 616 20557
rect 522 20515 608 20523
rect 649 20515 651 20565
rect 548 20499 582 20501
rect 522 20480 548 20485
rect 522 20479 582 20480
rect 586 20479 608 20485
rect 295 20444 300 20478
rect 324 20444 329 20478
rect 544 20476 582 20479
rect 378 20439 450 20447
rect 428 20409 430 20425
rect 400 20401 430 20409
rect 476 20407 480 20475
rect 544 20446 552 20476
rect 578 20446 582 20476
rect 544 20437 548 20446
rect 400 20397 434 20401
rect 400 20367 408 20397
rect 420 20367 434 20397
rect 544 20399 548 20407
rect 12 20328 62 20330
rect 28 20319 59 20321
rect 62 20319 64 20328
rect 28 20311 64 20319
rect 127 20319 158 20321
rect 127 20312 182 20319
rect 215 20317 224 20345
rect 127 20311 161 20312
rect 59 20295 64 20311
rect 158 20295 161 20311
rect 28 20287 64 20295
rect 127 20294 161 20295
rect 127 20287 182 20294
rect 62 20278 64 20287
rect 213 20279 224 20317
rect 282 20307 292 20365
rect 296 20359 368 20367
rect 319 20330 335 20332
rect 251 20273 263 20307
rect 273 20273 292 20307
rect 303 20300 316 20316
rect 303 20282 316 20298
rect 120 20225 170 20227
rect 76 20219 92 20225
rect 94 20219 110 20225
rect 76 20209 99 20218
rect 60 20199 67 20209
rect 76 20189 77 20209
rect 96 20184 99 20209
rect 109 20189 110 20209
rect 119 20199 126 20209
rect 76 20175 110 20179
rect 170 20175 172 20225
rect 186 20207 190 20241
rect 216 20207 220 20241
rect 186 20130 220 20164
rect 282 20161 292 20273
rect 318 20276 324 20329
rect 346 20316 348 20329
rect 428 20320 430 20367
rect 443 20357 450 20359
rect 476 20327 480 20395
rect 544 20365 552 20399
rect 578 20365 582 20399
rect 481 20333 517 20361
rect 481 20327 495 20333
rect 333 20282 353 20316
rect 367 20286 380 20320
rect 396 20286 408 20320
rect 420 20286 434 20320
rect 318 20266 335 20276
rect 318 20197 324 20266
rect 346 20197 348 20282
rect 428 20239 430 20286
rect 476 20249 480 20317
rect 485 20299 495 20327
rect 505 20299 519 20333
rect 544 20327 555 20365
rect 544 20299 553 20327
rect 544 20279 548 20299
rect 579 20258 582 20348
rect 599 20328 649 20330
rect 610 20320 624 20321
rect 607 20319 624 20320
rect 586 20312 644 20319
rect 607 20311 644 20312
rect 607 20295 610 20311
rect 616 20295 644 20311
rect 607 20294 644 20295
rect 586 20287 644 20294
rect 607 20286 610 20287
rect 649 20278 651 20328
rect 544 20241 548 20249
rect 400 20209 408 20239
rect 420 20209 434 20239
rect 400 20205 434 20209
rect 400 20197 430 20205
rect 428 20181 430 20197
rect 476 20169 480 20237
rect 544 20207 552 20241
rect 578 20207 582 20241
rect 544 20199 548 20207
rect 544 20169 586 20170
rect 288 20129 292 20161
rect 296 20159 368 20167
rect 378 20159 450 20167
rect 544 20162 548 20169
rect 439 20131 444 20159
rect 120 20115 170 20117
rect 76 20111 130 20115
rect 110 20106 130 20111
rect 60 20081 67 20091
rect 76 20081 77 20101
rect 96 20072 99 20106
rect 109 20081 110 20101
rect 119 20081 126 20091
rect 76 20065 92 20071
rect 94 20065 110 20071
rect 170 20065 172 20115
rect 186 20049 190 20083
rect 216 20049 220 20083
rect 213 20017 224 20049
rect 282 20045 292 20129
rect 296 20123 368 20131
rect 378 20123 450 20131
rect 468 20128 473 20162
rect 428 20093 430 20109
rect 251 20017 292 20045
rect 12 20012 62 20014
rect 28 20003 59 20005
rect 62 20003 64 20012
rect 251 20011 263 20017
rect 28 19995 64 20003
rect 127 20003 158 20005
rect 127 19996 182 20003
rect 127 19995 161 19996
rect 59 19979 64 19995
rect 158 19979 161 19995
rect 253 19983 263 20011
rect 273 19983 292 20017
rect 318 20024 324 20093
rect 318 20014 335 20024
rect 303 19992 316 20008
rect 28 19971 64 19979
rect 127 19978 161 19979
rect 127 19971 182 19978
rect 62 19962 64 19971
rect 282 19925 292 19983
rect 303 19974 316 19990
rect 318 19961 324 20014
rect 346 20008 348 20093
rect 400 20085 430 20093
rect 476 20091 480 20159
rect 511 20128 582 20162
rect 544 20121 548 20128
rect 400 20081 434 20085
rect 400 20051 408 20081
rect 420 20051 434 20081
rect 544 20083 548 20091
rect 333 19974 353 20008
rect 428 20004 430 20051
rect 476 20011 480 20079
rect 544 20049 552 20083
rect 578 20049 582 20083
rect 544 20041 548 20049
rect 346 19961 348 19974
rect 367 19970 380 20004
rect 396 19970 408 20004
rect 420 19970 434 20004
rect 544 20001 553 20029
rect 319 19958 335 19960
rect 120 19909 170 19911
rect 76 19903 92 19909
rect 94 19903 110 19909
rect 76 19893 99 19902
rect 60 19883 67 19893
rect 76 19873 77 19893
rect 96 19868 99 19893
rect 109 19873 110 19893
rect 119 19883 126 19893
rect 76 19859 110 19863
rect 170 19859 172 19909
rect 186 19891 190 19925
rect 216 19891 220 19925
rect 182 19853 224 19854
rect 186 19812 220 19846
rect 223 19812 257 19846
rect 160 19805 182 19811
rect 224 19805 246 19811
rect 288 19805 292 19925
rect 296 19923 368 19931
rect 428 19923 430 19970
rect 476 19933 480 20001
rect 485 19957 495 19991
rect 505 19957 519 19991
rect 544 19957 555 20001
rect 485 19933 492 19957
rect 579 19942 582 20032
rect 599 20012 649 20014
rect 610 20004 624 20005
rect 607 20003 624 20004
rect 586 19996 644 20003
rect 607 19995 644 19996
rect 607 19979 610 19995
rect 616 19979 644 19995
rect 607 19978 644 19979
rect 586 19971 644 19978
rect 607 19970 610 19971
rect 649 19962 651 20012
rect 544 19925 548 19933
rect 400 19893 408 19923
rect 420 19893 434 19923
rect 400 19889 434 19893
rect 400 19881 430 19889
rect 428 19865 430 19881
rect 476 19853 480 19921
rect 544 19891 552 19925
rect 578 19891 582 19925
rect 544 19883 548 19891
rect 295 19812 300 19846
rect 324 19812 329 19846
rect 378 19843 450 19851
rect 544 19848 548 19853
rect 544 19844 582 19848
rect 544 19814 552 19844
rect 578 19814 582 19844
rect 544 19811 548 19814
rect 522 19805 548 19811
rect 586 19805 608 19811
rect 182 19789 224 19805
rect 544 19789 586 19805
rect 17 19775 67 19777
rect 119 19775 169 19777
rect 599 19775 649 19777
rect 42 19733 59 19767
rect 67 19725 69 19775
rect 160 19767 246 19775
rect 522 19767 608 19775
rect 76 19733 110 19767
rect 127 19733 144 19767
rect 152 19733 161 19767
rect 162 19765 195 19767
rect 224 19765 244 19767
rect 162 19733 244 19765
rect 524 19765 548 19767
rect 573 19765 582 19767
rect 586 19765 606 19767
rect 160 19725 246 19733
rect 186 19709 220 19711
rect 182 19695 224 19696
rect 160 19689 182 19695
rect 224 19689 246 19695
rect 186 19654 220 19688
rect 223 19654 257 19688
rect 120 19641 170 19643
rect 76 19637 130 19641
rect 110 19632 130 19637
rect 60 19607 67 19617
rect 76 19607 77 19627
rect 96 19598 99 19632
rect 109 19607 110 19627
rect 119 19607 126 19617
rect 76 19591 92 19597
rect 94 19591 110 19597
rect 170 19591 172 19641
rect 186 19575 190 19609
rect 216 19575 220 19609
rect 288 19575 292 19763
rect 476 19695 480 19763
rect 524 19733 606 19765
rect 607 19733 616 19767
rect 522 19725 608 19733
rect 649 19725 651 19775
rect 548 19709 582 19711
rect 522 19690 548 19695
rect 522 19689 582 19690
rect 586 19689 608 19695
rect 295 19654 300 19688
rect 324 19654 329 19688
rect 544 19686 582 19689
rect 378 19649 450 19657
rect 428 19619 430 19635
rect 400 19611 430 19619
rect 476 19617 480 19685
rect 544 19656 552 19686
rect 578 19656 582 19686
rect 544 19647 548 19656
rect 400 19607 434 19611
rect 400 19577 408 19607
rect 420 19577 434 19607
rect 544 19609 548 19617
rect 12 19538 62 19540
rect 28 19529 59 19531
rect 62 19529 64 19538
rect 28 19521 64 19529
rect 127 19529 158 19531
rect 127 19522 182 19529
rect 215 19527 224 19555
rect 127 19521 161 19522
rect 59 19505 64 19521
rect 158 19505 161 19521
rect 28 19497 64 19505
rect 127 19504 161 19505
rect 127 19497 182 19504
rect 62 19488 64 19497
rect 213 19489 224 19527
rect 282 19517 292 19575
rect 296 19569 368 19577
rect 319 19540 335 19542
rect 251 19483 263 19517
rect 273 19483 292 19517
rect 303 19510 316 19526
rect 303 19492 316 19508
rect 120 19435 170 19437
rect 76 19429 92 19435
rect 94 19429 110 19435
rect 76 19419 99 19428
rect 60 19409 67 19419
rect 76 19399 77 19419
rect 96 19394 99 19419
rect 109 19399 110 19419
rect 119 19409 126 19419
rect 76 19385 110 19389
rect 170 19385 172 19435
rect 186 19417 190 19451
rect 216 19417 220 19451
rect 186 19340 220 19374
rect 282 19371 292 19483
rect 318 19486 324 19539
rect 346 19526 348 19539
rect 428 19530 430 19577
rect 443 19567 450 19569
rect 476 19537 480 19605
rect 544 19575 552 19609
rect 578 19575 582 19609
rect 481 19543 517 19571
rect 481 19537 495 19543
rect 333 19492 353 19526
rect 367 19496 380 19530
rect 396 19496 408 19530
rect 420 19496 434 19530
rect 318 19476 335 19486
rect 318 19407 324 19476
rect 346 19407 348 19492
rect 428 19449 430 19496
rect 476 19459 480 19527
rect 485 19509 495 19537
rect 505 19509 519 19543
rect 544 19537 555 19575
rect 544 19509 553 19537
rect 544 19489 548 19509
rect 579 19468 582 19558
rect 599 19538 649 19540
rect 610 19530 624 19531
rect 607 19529 624 19530
rect 586 19522 644 19529
rect 607 19521 644 19522
rect 607 19505 610 19521
rect 616 19505 644 19521
rect 607 19504 644 19505
rect 586 19497 644 19504
rect 607 19496 610 19497
rect 649 19488 651 19538
rect 544 19451 548 19459
rect 400 19419 408 19449
rect 420 19419 434 19449
rect 400 19415 434 19419
rect 400 19407 430 19415
rect 428 19391 430 19407
rect 476 19379 480 19447
rect 544 19417 552 19451
rect 578 19417 582 19451
rect 544 19409 548 19417
rect 544 19379 586 19380
rect 288 19339 292 19371
rect 296 19369 368 19377
rect 378 19369 450 19377
rect 544 19372 548 19379
rect 439 19341 444 19369
rect 120 19325 170 19327
rect 76 19321 130 19325
rect 110 19316 130 19321
rect 60 19291 67 19301
rect 76 19291 77 19311
rect 96 19282 99 19316
rect 109 19291 110 19311
rect 119 19291 126 19301
rect 76 19275 92 19281
rect 94 19275 110 19281
rect 170 19275 172 19325
rect 186 19259 190 19293
rect 216 19259 220 19293
rect 213 19227 224 19259
rect 282 19255 292 19339
rect 296 19333 368 19341
rect 378 19333 450 19341
rect 468 19338 473 19372
rect 428 19303 430 19319
rect 251 19227 292 19255
rect 12 19222 62 19224
rect 28 19213 59 19215
rect 62 19213 64 19222
rect 251 19221 263 19227
rect 28 19205 64 19213
rect 127 19213 158 19215
rect 127 19206 182 19213
rect 127 19205 161 19206
rect 59 19189 64 19205
rect 158 19189 161 19205
rect 253 19193 263 19221
rect 273 19193 292 19227
rect 318 19234 324 19303
rect 318 19224 335 19234
rect 303 19202 316 19218
rect 28 19181 64 19189
rect 127 19188 161 19189
rect 127 19181 182 19188
rect 62 19172 64 19181
rect 282 19135 292 19193
rect 303 19184 316 19200
rect 318 19171 324 19224
rect 346 19218 348 19303
rect 400 19295 430 19303
rect 476 19301 480 19369
rect 511 19338 582 19372
rect 544 19331 548 19338
rect 400 19291 434 19295
rect 400 19261 408 19291
rect 420 19261 434 19291
rect 544 19293 548 19301
rect 333 19184 353 19218
rect 428 19214 430 19261
rect 476 19221 480 19289
rect 544 19259 552 19293
rect 578 19259 582 19293
rect 544 19251 548 19259
rect 346 19171 348 19184
rect 367 19180 380 19214
rect 396 19180 408 19214
rect 420 19180 434 19214
rect 544 19211 553 19239
rect 319 19168 335 19170
rect 120 19119 170 19121
rect 76 19113 92 19119
rect 94 19113 110 19119
rect 76 19103 99 19112
rect 60 19093 67 19103
rect 76 19083 77 19103
rect 96 19078 99 19103
rect 109 19083 110 19103
rect 119 19093 126 19103
rect 76 19069 110 19073
rect 170 19069 172 19119
rect 186 19101 190 19135
rect 216 19101 220 19135
rect 182 19063 224 19064
rect 186 19022 220 19056
rect 223 19022 257 19056
rect 160 19015 182 19021
rect 224 19015 246 19021
rect 288 19015 292 19135
rect 296 19133 368 19141
rect 428 19133 430 19180
rect 476 19143 480 19211
rect 485 19167 495 19201
rect 505 19167 519 19201
rect 544 19167 555 19211
rect 485 19143 492 19167
rect 579 19152 582 19242
rect 599 19222 649 19224
rect 610 19214 624 19215
rect 607 19213 624 19214
rect 586 19206 644 19213
rect 607 19205 644 19206
rect 607 19189 610 19205
rect 616 19189 644 19205
rect 607 19188 644 19189
rect 586 19181 644 19188
rect 607 19180 610 19181
rect 649 19172 651 19222
rect 544 19135 548 19143
rect 400 19103 408 19133
rect 420 19103 434 19133
rect 400 19099 434 19103
rect 400 19091 430 19099
rect 428 19075 430 19091
rect 476 19063 480 19131
rect 544 19101 552 19135
rect 578 19101 582 19135
rect 544 19093 548 19101
rect 295 19022 300 19056
rect 324 19022 329 19056
rect 378 19053 450 19061
rect 544 19058 548 19063
rect 544 19054 582 19058
rect 544 19024 552 19054
rect 578 19024 582 19054
rect 544 19021 548 19024
rect 522 19015 548 19021
rect 586 19015 608 19021
rect 182 18999 224 19015
rect 544 18999 586 19015
rect 17 18985 67 18987
rect 119 18985 169 18987
rect 599 18985 649 18987
rect 42 18943 59 18977
rect 67 18935 69 18985
rect 160 18977 246 18985
rect 522 18977 608 18985
rect 76 18943 110 18977
rect 127 18943 144 18977
rect 152 18943 161 18977
rect 162 18975 195 18977
rect 224 18975 244 18977
rect 162 18943 244 18975
rect 524 18975 548 18977
rect 573 18975 582 18977
rect 586 18975 606 18977
rect 160 18935 246 18943
rect 186 18919 220 18921
rect 182 18905 224 18906
rect 160 18899 182 18905
rect 224 18899 246 18905
rect 186 18864 220 18898
rect 223 18864 257 18898
rect 120 18851 170 18853
rect 76 18847 130 18851
rect 110 18842 130 18847
rect 60 18817 67 18827
rect 76 18817 77 18837
rect 96 18808 99 18842
rect 109 18817 110 18837
rect 119 18817 126 18827
rect 76 18801 92 18807
rect 94 18801 110 18807
rect 170 18801 172 18851
rect 186 18785 190 18819
rect 216 18785 220 18819
rect 288 18785 292 18973
rect 476 18905 480 18973
rect 524 18943 606 18975
rect 607 18943 616 18977
rect 522 18935 608 18943
rect 649 18935 651 18985
rect 548 18919 582 18921
rect 522 18900 548 18905
rect 522 18899 582 18900
rect 586 18899 608 18905
rect 295 18864 300 18898
rect 324 18864 329 18898
rect 544 18896 582 18899
rect 378 18859 450 18867
rect 428 18829 430 18845
rect 400 18821 430 18829
rect 476 18827 480 18895
rect 544 18866 552 18896
rect 578 18866 582 18896
rect 544 18857 548 18866
rect 400 18817 434 18821
rect 400 18787 408 18817
rect 420 18787 434 18817
rect 544 18819 548 18827
rect 12 18748 62 18750
rect 28 18739 59 18741
rect 62 18739 64 18748
rect 28 18731 64 18739
rect 127 18739 158 18741
rect 127 18732 182 18739
rect 215 18737 224 18765
rect 127 18731 161 18732
rect 59 18715 64 18731
rect 158 18715 161 18731
rect 28 18707 64 18715
rect 127 18714 161 18715
rect 127 18707 182 18714
rect 62 18698 64 18707
rect 213 18699 224 18737
rect 282 18727 292 18785
rect 296 18779 368 18787
rect 319 18750 335 18752
rect 251 18693 263 18727
rect 273 18693 292 18727
rect 303 18720 316 18736
rect 303 18702 316 18718
rect 120 18645 170 18647
rect 76 18639 92 18645
rect 94 18639 110 18645
rect 76 18629 99 18638
rect 60 18619 67 18629
rect 76 18609 77 18629
rect 96 18604 99 18629
rect 109 18609 110 18629
rect 119 18619 126 18629
rect 76 18595 110 18599
rect 170 18595 172 18645
rect 186 18627 190 18661
rect 216 18627 220 18661
rect 186 18550 220 18584
rect 282 18581 292 18693
rect 318 18696 324 18749
rect 346 18736 348 18749
rect 428 18740 430 18787
rect 443 18777 450 18779
rect 476 18747 480 18815
rect 544 18785 552 18819
rect 578 18785 582 18819
rect 481 18753 517 18781
rect 481 18747 495 18753
rect 333 18702 353 18736
rect 367 18706 380 18740
rect 396 18706 408 18740
rect 420 18706 434 18740
rect 318 18686 335 18696
rect 318 18617 324 18686
rect 346 18617 348 18702
rect 428 18659 430 18706
rect 476 18669 480 18737
rect 485 18719 495 18747
rect 505 18719 519 18753
rect 544 18747 555 18785
rect 544 18719 553 18747
rect 544 18699 548 18719
rect 579 18678 582 18768
rect 599 18748 649 18750
rect 610 18740 624 18741
rect 607 18739 624 18740
rect 586 18732 644 18739
rect 607 18731 644 18732
rect 607 18715 610 18731
rect 616 18715 644 18731
rect 607 18714 644 18715
rect 586 18707 644 18714
rect 607 18706 610 18707
rect 649 18698 651 18748
rect 544 18661 548 18669
rect 400 18629 408 18659
rect 420 18629 434 18659
rect 400 18625 434 18629
rect 400 18617 430 18625
rect 428 18601 430 18617
rect 476 18589 480 18657
rect 544 18627 552 18661
rect 578 18627 582 18661
rect 544 18619 548 18627
rect 544 18589 586 18590
rect 288 18549 292 18581
rect 296 18579 368 18587
rect 378 18579 450 18587
rect 544 18582 548 18589
rect 439 18551 444 18579
rect 120 18535 170 18537
rect 76 18531 130 18535
rect 110 18526 130 18531
rect 60 18501 67 18511
rect 76 18501 77 18521
rect 96 18492 99 18526
rect 109 18501 110 18521
rect 119 18501 126 18511
rect 76 18485 92 18491
rect 94 18485 110 18491
rect 170 18485 172 18535
rect 186 18469 190 18503
rect 216 18469 220 18503
rect 213 18437 224 18469
rect 282 18465 292 18549
rect 296 18543 368 18551
rect 378 18543 450 18551
rect 468 18548 473 18582
rect 428 18513 430 18529
rect 251 18437 292 18465
rect 12 18432 62 18434
rect 28 18423 59 18425
rect 62 18423 64 18432
rect 251 18431 263 18437
rect 28 18415 64 18423
rect 127 18423 158 18425
rect 127 18416 182 18423
rect 127 18415 161 18416
rect 59 18399 64 18415
rect 158 18399 161 18415
rect 253 18403 263 18431
rect 273 18403 292 18437
rect 318 18444 324 18513
rect 318 18434 335 18444
rect 303 18412 316 18428
rect 28 18391 64 18399
rect 127 18398 161 18399
rect 127 18391 182 18398
rect 62 18382 64 18391
rect 282 18345 292 18403
rect 303 18394 316 18410
rect 318 18381 324 18434
rect 346 18428 348 18513
rect 400 18505 430 18513
rect 476 18511 480 18579
rect 511 18548 582 18582
rect 544 18541 548 18548
rect 400 18501 434 18505
rect 400 18471 408 18501
rect 420 18471 434 18501
rect 544 18503 548 18511
rect 333 18394 353 18428
rect 428 18424 430 18471
rect 476 18431 480 18499
rect 544 18469 552 18503
rect 578 18469 582 18503
rect 544 18461 548 18469
rect 346 18381 348 18394
rect 367 18390 380 18424
rect 396 18390 408 18424
rect 420 18390 434 18424
rect 544 18421 553 18449
rect 319 18378 335 18380
rect 120 18329 170 18331
rect 76 18323 92 18329
rect 94 18323 110 18329
rect 76 18313 99 18322
rect 60 18303 67 18313
rect 76 18293 77 18313
rect 96 18288 99 18313
rect 109 18293 110 18313
rect 119 18303 126 18313
rect 76 18279 110 18283
rect 170 18279 172 18329
rect 186 18311 190 18345
rect 216 18311 220 18345
rect 182 18273 224 18274
rect 186 18232 220 18266
rect 223 18232 257 18266
rect 160 18225 182 18231
rect 224 18225 246 18231
rect 288 18225 292 18345
rect 296 18343 368 18351
rect 428 18343 430 18390
rect 476 18353 480 18421
rect 485 18377 495 18411
rect 505 18377 519 18411
rect 544 18377 555 18421
rect 485 18353 492 18377
rect 579 18362 582 18452
rect 599 18432 649 18434
rect 610 18424 624 18425
rect 607 18423 624 18424
rect 586 18416 644 18423
rect 607 18415 644 18416
rect 607 18399 610 18415
rect 616 18399 644 18415
rect 607 18398 644 18399
rect 586 18391 644 18398
rect 607 18390 610 18391
rect 649 18382 651 18432
rect 544 18345 548 18353
rect 400 18313 408 18343
rect 420 18313 434 18343
rect 400 18309 434 18313
rect 400 18301 430 18309
rect 428 18285 430 18301
rect 476 18273 480 18341
rect 544 18311 552 18345
rect 578 18311 582 18345
rect 544 18303 548 18311
rect 295 18232 300 18266
rect 324 18232 329 18266
rect 378 18263 450 18271
rect 544 18268 548 18273
rect 544 18264 582 18268
rect 544 18234 552 18264
rect 578 18234 582 18264
rect 544 18231 548 18234
rect 522 18225 548 18231
rect 586 18225 608 18231
rect 182 18209 224 18225
rect 544 18209 586 18225
rect 17 18195 67 18197
rect 119 18195 169 18197
rect 599 18195 649 18197
rect 42 18153 59 18187
rect 67 18145 69 18195
rect 160 18187 246 18195
rect 522 18187 608 18195
rect 76 18153 110 18187
rect 127 18153 144 18187
rect 152 18153 161 18187
rect 162 18185 195 18187
rect 224 18185 244 18187
rect 162 18153 244 18185
rect 524 18185 548 18187
rect 573 18185 582 18187
rect 586 18185 606 18187
rect 160 18145 246 18153
rect 186 18129 220 18131
rect 182 18115 224 18116
rect 160 18109 182 18115
rect 224 18109 246 18115
rect 186 18074 220 18108
rect 223 18074 257 18108
rect 120 18061 170 18063
rect 76 18057 130 18061
rect 110 18052 130 18057
rect 60 18027 67 18037
rect 76 18027 77 18047
rect 96 18018 99 18052
rect 109 18027 110 18047
rect 119 18027 126 18037
rect 76 18011 92 18017
rect 94 18011 110 18017
rect 170 18011 172 18061
rect 186 17995 190 18029
rect 216 17995 220 18029
rect 288 17995 292 18183
rect 476 18115 480 18183
rect 524 18153 606 18185
rect 607 18153 616 18187
rect 522 18145 608 18153
rect 649 18145 651 18195
rect 548 18129 582 18131
rect 522 18110 548 18115
rect 522 18109 582 18110
rect 586 18109 608 18115
rect 295 18074 300 18108
rect 324 18074 329 18108
rect 544 18106 582 18109
rect 378 18069 450 18077
rect 428 18039 430 18055
rect 400 18031 430 18039
rect 476 18037 480 18105
rect 544 18076 552 18106
rect 578 18076 582 18106
rect 544 18067 548 18076
rect 400 18027 434 18031
rect 400 17997 408 18027
rect 420 17997 434 18027
rect 544 18029 548 18037
rect 12 17958 62 17960
rect 28 17949 59 17951
rect 62 17949 64 17958
rect 28 17941 64 17949
rect 127 17949 158 17951
rect 127 17942 182 17949
rect 215 17947 224 17975
rect 127 17941 161 17942
rect 59 17925 64 17941
rect 158 17925 161 17941
rect 28 17917 64 17925
rect 127 17924 161 17925
rect 127 17917 182 17924
rect 62 17908 64 17917
rect 213 17909 224 17947
rect 282 17937 292 17995
rect 296 17989 368 17997
rect 319 17960 335 17962
rect 251 17903 263 17937
rect 273 17903 292 17937
rect 303 17930 316 17946
rect 303 17912 316 17928
rect 120 17855 170 17857
rect 76 17849 92 17855
rect 94 17849 110 17855
rect 76 17839 99 17848
rect 60 17829 67 17839
rect 76 17819 77 17839
rect 96 17814 99 17839
rect 109 17819 110 17839
rect 119 17829 126 17839
rect 76 17805 110 17809
rect 170 17805 172 17855
rect 186 17837 190 17871
rect 216 17837 220 17871
rect 186 17760 220 17794
rect 282 17791 292 17903
rect 318 17906 324 17959
rect 346 17946 348 17959
rect 428 17950 430 17997
rect 443 17987 450 17989
rect 476 17957 480 18025
rect 544 17995 552 18029
rect 578 17995 582 18029
rect 481 17963 517 17991
rect 481 17957 495 17963
rect 333 17912 353 17946
rect 367 17916 380 17950
rect 396 17916 408 17950
rect 420 17916 434 17950
rect 318 17896 335 17906
rect 318 17827 324 17896
rect 346 17827 348 17912
rect 428 17869 430 17916
rect 476 17879 480 17947
rect 485 17929 495 17957
rect 505 17929 519 17963
rect 544 17957 555 17995
rect 544 17929 553 17957
rect 544 17909 548 17929
rect 579 17888 582 17978
rect 599 17958 649 17960
rect 610 17950 624 17951
rect 607 17949 624 17950
rect 586 17942 644 17949
rect 607 17941 644 17942
rect 607 17925 610 17941
rect 616 17925 644 17941
rect 607 17924 644 17925
rect 586 17917 644 17924
rect 607 17916 610 17917
rect 649 17908 651 17958
rect 544 17871 548 17879
rect 400 17839 408 17869
rect 420 17839 434 17869
rect 400 17835 434 17839
rect 400 17827 430 17835
rect 428 17811 430 17827
rect 476 17799 480 17867
rect 544 17837 552 17871
rect 578 17837 582 17871
rect 544 17829 548 17837
rect 544 17799 586 17800
rect 288 17759 292 17791
rect 296 17789 368 17797
rect 378 17789 450 17797
rect 544 17792 548 17799
rect 439 17761 444 17789
rect 120 17745 170 17747
rect 76 17741 130 17745
rect 110 17736 130 17741
rect 60 17711 67 17721
rect 76 17711 77 17731
rect 96 17702 99 17736
rect 109 17711 110 17731
rect 119 17711 126 17721
rect 76 17695 92 17701
rect 94 17695 110 17701
rect 170 17695 172 17745
rect 186 17679 190 17713
rect 216 17679 220 17713
rect 213 17647 224 17679
rect 282 17675 292 17759
rect 296 17753 368 17761
rect 378 17753 450 17761
rect 468 17758 473 17792
rect 428 17723 430 17739
rect 251 17647 292 17675
rect 12 17642 62 17644
rect 28 17633 59 17635
rect 62 17633 64 17642
rect 251 17641 263 17647
rect 28 17625 64 17633
rect 127 17633 158 17635
rect 127 17626 182 17633
rect 127 17625 161 17626
rect 59 17609 64 17625
rect 158 17609 161 17625
rect 253 17613 263 17641
rect 273 17613 292 17647
rect 318 17654 324 17723
rect 318 17644 335 17654
rect 303 17622 316 17638
rect 28 17601 64 17609
rect 127 17608 161 17609
rect 127 17601 182 17608
rect 62 17592 64 17601
rect 282 17555 292 17613
rect 303 17604 316 17620
rect 318 17591 324 17644
rect 346 17638 348 17723
rect 400 17715 430 17723
rect 476 17721 480 17789
rect 511 17758 582 17792
rect 544 17751 548 17758
rect 400 17711 434 17715
rect 400 17681 408 17711
rect 420 17681 434 17711
rect 544 17713 548 17721
rect 333 17604 353 17638
rect 428 17634 430 17681
rect 476 17641 480 17709
rect 544 17679 552 17713
rect 578 17679 582 17713
rect 544 17671 548 17679
rect 346 17591 348 17604
rect 367 17600 380 17634
rect 396 17600 408 17634
rect 420 17600 434 17634
rect 544 17631 553 17659
rect 319 17588 335 17590
rect 120 17539 170 17541
rect 76 17533 92 17539
rect 94 17533 110 17539
rect 76 17523 99 17532
rect 60 17513 67 17523
rect 76 17503 77 17523
rect 96 17498 99 17523
rect 109 17503 110 17523
rect 119 17513 126 17523
rect 76 17489 110 17493
rect 170 17489 172 17539
rect 186 17521 190 17555
rect 216 17521 220 17555
rect 182 17483 224 17484
rect 186 17442 220 17476
rect 223 17442 257 17476
rect 160 17435 182 17441
rect 224 17435 246 17441
rect 288 17435 292 17555
rect 296 17553 368 17561
rect 428 17553 430 17600
rect 476 17563 480 17631
rect 485 17587 495 17621
rect 505 17587 519 17621
rect 544 17587 555 17631
rect 485 17563 492 17587
rect 579 17572 582 17662
rect 599 17642 649 17644
rect 610 17634 624 17635
rect 607 17633 624 17634
rect 586 17626 644 17633
rect 607 17625 644 17626
rect 607 17609 610 17625
rect 616 17609 644 17625
rect 607 17608 644 17609
rect 586 17601 644 17608
rect 607 17600 610 17601
rect 649 17592 651 17642
rect 544 17555 548 17563
rect 400 17523 408 17553
rect 420 17523 434 17553
rect 400 17519 434 17523
rect 400 17511 430 17519
rect 428 17495 430 17511
rect 476 17483 480 17551
rect 544 17521 552 17555
rect 578 17521 582 17555
rect 544 17513 548 17521
rect 295 17442 300 17476
rect 324 17442 329 17476
rect 378 17473 450 17481
rect 544 17478 548 17483
rect 544 17474 582 17478
rect 544 17444 552 17474
rect 578 17444 582 17474
rect 544 17441 548 17444
rect 522 17435 548 17441
rect 586 17435 608 17441
rect 182 17419 224 17435
rect 544 17419 586 17435
rect 17 17405 67 17407
rect 119 17405 169 17407
rect 599 17405 649 17407
rect 42 17363 59 17397
rect 67 17355 69 17405
rect 160 17397 246 17405
rect 522 17397 608 17405
rect 76 17363 110 17397
rect 127 17363 144 17397
rect 152 17363 161 17397
rect 162 17395 195 17397
rect 224 17395 244 17397
rect 162 17363 244 17395
rect 524 17395 548 17397
rect 573 17395 582 17397
rect 586 17395 606 17397
rect 160 17355 246 17363
rect 186 17339 220 17341
rect 182 17325 224 17326
rect 160 17319 182 17325
rect 224 17319 246 17325
rect 186 17284 220 17318
rect 223 17284 257 17318
rect 120 17271 170 17273
rect 76 17267 130 17271
rect 110 17262 130 17267
rect 60 17237 67 17247
rect 76 17237 77 17257
rect 96 17228 99 17262
rect 109 17237 110 17257
rect 119 17237 126 17247
rect 76 17221 92 17227
rect 94 17221 110 17227
rect 170 17221 172 17271
rect 186 17205 190 17239
rect 216 17205 220 17239
rect 288 17205 292 17393
rect 476 17325 480 17393
rect 524 17363 606 17395
rect 607 17363 616 17397
rect 522 17355 608 17363
rect 649 17355 651 17405
rect 548 17339 582 17341
rect 522 17320 548 17325
rect 522 17319 582 17320
rect 586 17319 608 17325
rect 295 17284 300 17318
rect 324 17284 329 17318
rect 544 17316 582 17319
rect 378 17279 450 17287
rect 428 17249 430 17265
rect 400 17241 430 17249
rect 476 17247 480 17315
rect 544 17286 552 17316
rect 578 17286 582 17316
rect 544 17277 548 17286
rect 400 17237 434 17241
rect 400 17207 408 17237
rect 420 17207 434 17237
rect 544 17239 548 17247
rect 12 17168 62 17170
rect 28 17159 59 17161
rect 62 17159 64 17168
rect 28 17151 64 17159
rect 127 17159 158 17161
rect 127 17152 182 17159
rect 215 17157 224 17185
rect 127 17151 161 17152
rect 59 17135 64 17151
rect 158 17135 161 17151
rect 28 17127 64 17135
rect 127 17134 161 17135
rect 127 17127 182 17134
rect 62 17118 64 17127
rect 213 17119 224 17157
rect 282 17147 292 17205
rect 296 17199 368 17207
rect 319 17170 335 17172
rect 251 17113 263 17147
rect 273 17113 292 17147
rect 303 17140 316 17156
rect 303 17122 316 17138
rect 120 17065 170 17067
rect 76 17059 92 17065
rect 94 17059 110 17065
rect 76 17049 99 17058
rect 60 17039 67 17049
rect 76 17029 77 17049
rect 96 17024 99 17049
rect 109 17029 110 17049
rect 119 17039 126 17049
rect 76 17015 110 17019
rect 170 17015 172 17065
rect 186 17047 190 17081
rect 216 17047 220 17081
rect 186 16970 220 17004
rect 282 17001 292 17113
rect 318 17116 324 17169
rect 346 17156 348 17169
rect 428 17160 430 17207
rect 443 17197 450 17199
rect 476 17167 480 17235
rect 544 17205 552 17239
rect 578 17205 582 17239
rect 481 17173 517 17201
rect 481 17167 495 17173
rect 333 17122 353 17156
rect 367 17126 380 17160
rect 396 17126 408 17160
rect 420 17126 434 17160
rect 318 17106 335 17116
rect 318 17037 324 17106
rect 346 17037 348 17122
rect 428 17079 430 17126
rect 476 17089 480 17157
rect 485 17139 495 17167
rect 505 17139 519 17173
rect 544 17167 555 17205
rect 544 17139 553 17167
rect 544 17119 548 17139
rect 579 17098 582 17188
rect 599 17168 649 17170
rect 610 17160 624 17161
rect 607 17159 624 17160
rect 586 17152 644 17159
rect 607 17151 644 17152
rect 607 17135 610 17151
rect 616 17135 644 17151
rect 607 17134 644 17135
rect 586 17127 644 17134
rect 607 17126 610 17127
rect 649 17118 651 17168
rect 544 17081 548 17089
rect 400 17049 408 17079
rect 420 17049 434 17079
rect 400 17045 434 17049
rect 400 17037 430 17045
rect 428 17021 430 17037
rect 476 17009 480 17077
rect 544 17047 552 17081
rect 578 17047 582 17081
rect 544 17039 548 17047
rect 544 17009 586 17010
rect 288 16969 292 17001
rect 296 16999 368 17007
rect 378 16999 450 17007
rect 544 17002 548 17009
rect 439 16971 444 16999
rect 120 16955 170 16957
rect 76 16951 130 16955
rect 110 16946 130 16951
rect 60 16921 67 16931
rect 76 16921 77 16941
rect 96 16912 99 16946
rect 109 16921 110 16941
rect 119 16921 126 16931
rect 76 16905 92 16911
rect 94 16905 110 16911
rect 170 16905 172 16955
rect 186 16889 190 16923
rect 216 16889 220 16923
rect 213 16857 224 16889
rect 282 16885 292 16969
rect 296 16963 368 16971
rect 378 16963 450 16971
rect 468 16968 473 17002
rect 428 16933 430 16949
rect 251 16857 292 16885
rect 12 16852 62 16854
rect 28 16843 59 16845
rect 62 16843 64 16852
rect 251 16851 263 16857
rect 28 16835 64 16843
rect 127 16843 158 16845
rect 127 16836 182 16843
rect 127 16835 161 16836
rect 59 16819 64 16835
rect 158 16819 161 16835
rect 253 16823 263 16851
rect 273 16823 292 16857
rect 318 16864 324 16933
rect 318 16854 335 16864
rect 303 16832 316 16848
rect 28 16811 64 16819
rect 127 16818 161 16819
rect 127 16811 182 16818
rect 62 16802 64 16811
rect 282 16765 292 16823
rect 303 16814 316 16830
rect 318 16801 324 16854
rect 346 16848 348 16933
rect 400 16925 430 16933
rect 476 16931 480 16999
rect 511 16968 582 17002
rect 544 16961 548 16968
rect 400 16921 434 16925
rect 400 16891 408 16921
rect 420 16891 434 16921
rect 544 16923 548 16931
rect 333 16814 353 16848
rect 428 16844 430 16891
rect 476 16851 480 16919
rect 544 16889 552 16923
rect 578 16889 582 16923
rect 544 16881 548 16889
rect 346 16801 348 16814
rect 367 16810 380 16844
rect 396 16810 408 16844
rect 420 16810 434 16844
rect 544 16841 553 16869
rect 319 16798 335 16800
rect 120 16749 170 16751
rect 76 16743 92 16749
rect 94 16743 110 16749
rect 76 16733 99 16742
rect 60 16723 67 16733
rect 76 16713 77 16733
rect 96 16708 99 16733
rect 109 16713 110 16733
rect 119 16723 126 16733
rect 76 16699 110 16703
rect 170 16699 172 16749
rect 186 16731 190 16765
rect 216 16731 220 16765
rect 182 16693 224 16694
rect 186 16652 220 16686
rect 223 16652 257 16686
rect 160 16645 182 16651
rect 224 16645 246 16651
rect 288 16645 292 16765
rect 296 16763 368 16771
rect 428 16763 430 16810
rect 476 16773 480 16841
rect 485 16797 495 16831
rect 505 16797 519 16831
rect 544 16797 555 16841
rect 485 16773 492 16797
rect 579 16782 582 16872
rect 599 16852 649 16854
rect 610 16844 624 16845
rect 607 16843 624 16844
rect 586 16836 644 16843
rect 607 16835 644 16836
rect 607 16819 610 16835
rect 616 16819 644 16835
rect 607 16818 644 16819
rect 586 16811 644 16818
rect 607 16810 610 16811
rect 649 16802 651 16852
rect 544 16765 548 16773
rect 400 16733 408 16763
rect 420 16733 434 16763
rect 400 16729 434 16733
rect 400 16721 430 16729
rect 428 16705 430 16721
rect 476 16693 480 16761
rect 544 16731 552 16765
rect 578 16731 582 16765
rect 544 16723 548 16731
rect 295 16652 300 16686
rect 324 16652 329 16686
rect 378 16683 450 16691
rect 544 16688 548 16693
rect 544 16684 582 16688
rect 544 16654 552 16684
rect 578 16654 582 16684
rect 544 16651 548 16654
rect 522 16645 548 16651
rect 586 16645 608 16651
rect 182 16629 224 16645
rect 544 16629 586 16645
rect 17 16615 67 16617
rect 119 16615 169 16617
rect 599 16615 649 16617
rect 42 16573 59 16607
rect 67 16565 69 16615
rect 160 16607 246 16615
rect 522 16607 608 16615
rect 76 16573 110 16607
rect 127 16573 144 16607
rect 152 16573 161 16607
rect 162 16605 195 16607
rect 224 16605 244 16607
rect 162 16573 244 16605
rect 524 16605 548 16607
rect 573 16605 582 16607
rect 586 16605 606 16607
rect 160 16565 246 16573
rect 186 16549 220 16551
rect 182 16535 224 16536
rect 160 16529 182 16535
rect 224 16529 246 16535
rect 186 16494 220 16528
rect 223 16494 257 16528
rect 120 16481 170 16483
rect 76 16477 130 16481
rect 110 16472 130 16477
rect 60 16447 67 16457
rect 76 16447 77 16467
rect 96 16438 99 16472
rect 109 16447 110 16467
rect 119 16447 126 16457
rect 76 16431 92 16437
rect 94 16431 110 16437
rect 170 16431 172 16481
rect 186 16415 190 16449
rect 216 16415 220 16449
rect 288 16415 292 16603
rect 476 16535 480 16603
rect 524 16573 606 16605
rect 607 16573 616 16607
rect 522 16565 608 16573
rect 649 16565 651 16615
rect 548 16549 582 16551
rect 522 16530 548 16535
rect 522 16529 582 16530
rect 586 16529 608 16535
rect 295 16494 300 16528
rect 324 16494 329 16528
rect 544 16526 582 16529
rect 378 16489 450 16497
rect 428 16459 430 16475
rect 400 16451 430 16459
rect 476 16457 480 16525
rect 544 16496 552 16526
rect 578 16496 582 16526
rect 544 16487 548 16496
rect 400 16447 434 16451
rect 400 16417 408 16447
rect 420 16417 434 16447
rect 544 16449 548 16457
rect 12 16378 62 16380
rect 28 16369 59 16371
rect 62 16369 64 16378
rect 28 16361 64 16369
rect 127 16369 158 16371
rect 127 16362 182 16369
rect 215 16367 224 16395
rect 127 16361 161 16362
rect 59 16345 64 16361
rect 158 16345 161 16361
rect 28 16337 64 16345
rect 127 16344 161 16345
rect 127 16337 182 16344
rect 62 16328 64 16337
rect 213 16329 224 16367
rect 282 16357 292 16415
rect 296 16409 368 16417
rect 319 16380 335 16382
rect 251 16323 263 16357
rect 273 16323 292 16357
rect 303 16350 316 16366
rect 303 16332 316 16348
rect 120 16275 170 16277
rect 76 16269 92 16275
rect 94 16269 110 16275
rect 76 16259 99 16268
rect 60 16249 67 16259
rect 76 16239 77 16259
rect 96 16234 99 16259
rect 109 16239 110 16259
rect 119 16249 126 16259
rect 76 16225 110 16229
rect 170 16225 172 16275
rect 186 16257 190 16291
rect 216 16257 220 16291
rect 186 16180 220 16214
rect 282 16211 292 16323
rect 318 16326 324 16379
rect 346 16366 348 16379
rect 428 16370 430 16417
rect 443 16407 450 16409
rect 476 16377 480 16445
rect 544 16415 552 16449
rect 578 16415 582 16449
rect 481 16383 517 16411
rect 481 16377 495 16383
rect 333 16332 353 16366
rect 367 16336 380 16370
rect 396 16336 408 16370
rect 420 16336 434 16370
rect 318 16316 335 16326
rect 318 16247 324 16316
rect 346 16247 348 16332
rect 428 16289 430 16336
rect 476 16299 480 16367
rect 485 16349 495 16377
rect 505 16349 519 16383
rect 544 16377 555 16415
rect 544 16349 553 16377
rect 544 16329 548 16349
rect 579 16308 582 16398
rect 599 16378 649 16380
rect 610 16370 624 16371
rect 607 16369 624 16370
rect 586 16362 644 16369
rect 607 16361 644 16362
rect 607 16345 610 16361
rect 616 16345 644 16361
rect 607 16344 644 16345
rect 586 16337 644 16344
rect 607 16336 610 16337
rect 649 16328 651 16378
rect 544 16291 548 16299
rect 400 16259 408 16289
rect 420 16259 434 16289
rect 400 16255 434 16259
rect 400 16247 430 16255
rect 428 16231 430 16247
rect 476 16219 480 16287
rect 544 16257 552 16291
rect 578 16257 582 16291
rect 544 16249 548 16257
rect 544 16219 586 16220
rect 288 16179 292 16211
rect 296 16209 368 16217
rect 378 16209 450 16217
rect 544 16212 548 16219
rect 439 16181 444 16209
rect 120 16165 170 16167
rect 76 16161 130 16165
rect 110 16156 130 16161
rect 60 16131 67 16141
rect 76 16131 77 16151
rect 96 16122 99 16156
rect 109 16131 110 16151
rect 119 16131 126 16141
rect 76 16115 92 16121
rect 94 16115 110 16121
rect 170 16115 172 16165
rect 186 16099 190 16133
rect 216 16099 220 16133
rect 213 16067 224 16099
rect 282 16095 292 16179
rect 296 16173 368 16181
rect 378 16173 450 16181
rect 468 16178 473 16212
rect 428 16143 430 16159
rect 251 16067 292 16095
rect 12 16062 62 16064
rect 28 16053 59 16055
rect 62 16053 64 16062
rect 251 16061 263 16067
rect 28 16045 64 16053
rect 127 16053 158 16055
rect 127 16046 182 16053
rect 127 16045 161 16046
rect 59 16029 64 16045
rect 158 16029 161 16045
rect 253 16033 263 16061
rect 273 16033 292 16067
rect 318 16074 324 16143
rect 318 16064 335 16074
rect 303 16042 316 16058
rect 28 16021 64 16029
rect 127 16028 161 16029
rect 127 16021 182 16028
rect 62 16012 64 16021
rect 282 15975 292 16033
rect 303 16024 316 16040
rect 318 16011 324 16064
rect 346 16058 348 16143
rect 400 16135 430 16143
rect 476 16141 480 16209
rect 511 16178 582 16212
rect 544 16171 548 16178
rect 400 16131 434 16135
rect 400 16101 408 16131
rect 420 16101 434 16131
rect 544 16133 548 16141
rect 333 16024 353 16058
rect 428 16054 430 16101
rect 476 16061 480 16129
rect 544 16099 552 16133
rect 578 16099 582 16133
rect 544 16091 548 16099
rect 346 16011 348 16024
rect 367 16020 380 16054
rect 396 16020 408 16054
rect 420 16020 434 16054
rect 544 16051 553 16079
rect 319 16008 335 16010
rect 120 15959 170 15961
rect 76 15953 92 15959
rect 94 15953 110 15959
rect 76 15943 99 15952
rect 60 15933 67 15943
rect 76 15923 77 15943
rect 96 15918 99 15943
rect 109 15923 110 15943
rect 119 15933 126 15943
rect 76 15909 110 15913
rect 170 15909 172 15959
rect 186 15941 190 15975
rect 216 15941 220 15975
rect 182 15903 224 15904
rect 186 15862 220 15896
rect 223 15862 257 15896
rect 160 15855 182 15861
rect 224 15855 246 15861
rect 288 15855 292 15975
rect 296 15973 368 15981
rect 428 15973 430 16020
rect 476 15983 480 16051
rect 485 16007 495 16041
rect 505 16007 519 16041
rect 544 16007 555 16051
rect 485 15983 492 16007
rect 579 15992 582 16082
rect 599 16062 649 16064
rect 610 16054 624 16055
rect 607 16053 624 16054
rect 586 16046 644 16053
rect 607 16045 644 16046
rect 607 16029 610 16045
rect 616 16029 644 16045
rect 607 16028 644 16029
rect 586 16021 644 16028
rect 607 16020 610 16021
rect 649 16012 651 16062
rect 544 15975 548 15983
rect 400 15943 408 15973
rect 420 15943 434 15973
rect 400 15939 434 15943
rect 400 15931 430 15939
rect 428 15915 430 15931
rect 476 15903 480 15971
rect 544 15941 552 15975
rect 578 15941 582 15975
rect 544 15933 548 15941
rect 295 15862 300 15896
rect 324 15862 329 15896
rect 378 15893 450 15901
rect 544 15898 548 15903
rect 544 15894 582 15898
rect 544 15864 552 15894
rect 578 15864 582 15894
rect 544 15861 548 15864
rect 522 15855 548 15861
rect 586 15855 608 15861
rect 182 15839 224 15855
rect 544 15839 586 15855
rect 17 15825 67 15827
rect 119 15825 169 15827
rect 599 15825 649 15827
rect 42 15783 59 15817
rect 67 15775 69 15825
rect 160 15817 246 15825
rect 522 15817 608 15825
rect 76 15783 110 15817
rect 127 15783 144 15817
rect 152 15783 161 15817
rect 162 15815 195 15817
rect 224 15815 244 15817
rect 162 15783 244 15815
rect 524 15815 548 15817
rect 573 15815 582 15817
rect 586 15815 606 15817
rect 160 15775 246 15783
rect 186 15759 220 15761
rect 182 15745 224 15746
rect 160 15739 182 15745
rect 224 15739 246 15745
rect 186 15704 220 15738
rect 223 15704 257 15738
rect 120 15691 170 15693
rect 76 15687 130 15691
rect 110 15682 130 15687
rect 60 15657 67 15667
rect 76 15657 77 15677
rect 96 15648 99 15682
rect 109 15657 110 15677
rect 119 15657 126 15667
rect 76 15641 92 15647
rect 94 15641 110 15647
rect 170 15641 172 15691
rect 186 15625 190 15659
rect 216 15625 220 15659
rect 288 15625 292 15813
rect 476 15745 480 15813
rect 524 15783 606 15815
rect 607 15783 616 15817
rect 522 15775 608 15783
rect 649 15775 651 15825
rect 548 15759 582 15761
rect 522 15740 548 15745
rect 522 15739 582 15740
rect 586 15739 608 15745
rect 295 15704 300 15738
rect 324 15704 329 15738
rect 544 15736 582 15739
rect 378 15699 450 15707
rect 428 15669 430 15685
rect 400 15661 430 15669
rect 476 15667 480 15735
rect 544 15706 552 15736
rect 578 15706 582 15736
rect 544 15697 548 15706
rect 400 15657 434 15661
rect 400 15627 408 15657
rect 420 15627 434 15657
rect 544 15659 548 15667
rect 12 15588 62 15590
rect 28 15579 59 15581
rect 62 15579 64 15588
rect 28 15571 64 15579
rect 127 15579 158 15581
rect 127 15572 182 15579
rect 215 15577 224 15605
rect 127 15571 161 15572
rect 59 15555 64 15571
rect 158 15555 161 15571
rect 28 15547 64 15555
rect 127 15554 161 15555
rect 127 15547 182 15554
rect 62 15538 64 15547
rect 213 15539 224 15577
rect 282 15567 292 15625
rect 296 15619 368 15627
rect 319 15590 335 15592
rect 251 15533 263 15567
rect 273 15533 292 15567
rect 303 15560 316 15576
rect 303 15542 316 15558
rect 120 15485 170 15487
rect 76 15479 92 15485
rect 94 15479 110 15485
rect 76 15469 99 15478
rect 60 15459 67 15469
rect 76 15449 77 15469
rect 96 15444 99 15469
rect 109 15449 110 15469
rect 119 15459 126 15469
rect 76 15435 110 15439
rect 170 15435 172 15485
rect 186 15467 190 15501
rect 216 15467 220 15501
rect 186 15390 220 15424
rect 282 15421 292 15533
rect 318 15536 324 15589
rect 346 15576 348 15589
rect 428 15580 430 15627
rect 443 15617 450 15619
rect 476 15587 480 15655
rect 544 15625 552 15659
rect 578 15625 582 15659
rect 481 15593 517 15621
rect 481 15587 495 15593
rect 333 15542 353 15576
rect 367 15546 380 15580
rect 396 15546 408 15580
rect 420 15546 434 15580
rect 318 15526 335 15536
rect 318 15457 324 15526
rect 346 15457 348 15542
rect 428 15499 430 15546
rect 476 15509 480 15577
rect 485 15559 495 15587
rect 505 15559 519 15593
rect 544 15587 555 15625
rect 544 15559 553 15587
rect 544 15539 548 15559
rect 579 15518 582 15608
rect 599 15588 649 15590
rect 610 15580 624 15581
rect 607 15579 624 15580
rect 586 15572 644 15579
rect 607 15571 644 15572
rect 607 15555 610 15571
rect 616 15555 644 15571
rect 607 15554 644 15555
rect 586 15547 644 15554
rect 607 15546 610 15547
rect 649 15538 651 15588
rect 544 15501 548 15509
rect 400 15469 408 15499
rect 420 15469 434 15499
rect 400 15465 434 15469
rect 400 15457 430 15465
rect 428 15441 430 15457
rect 476 15429 480 15497
rect 544 15467 552 15501
rect 578 15467 582 15501
rect 544 15459 548 15467
rect 544 15429 586 15430
rect 288 15389 292 15421
rect 296 15419 368 15427
rect 378 15419 450 15427
rect 544 15422 548 15429
rect 439 15391 444 15419
rect 120 15375 170 15377
rect 76 15371 130 15375
rect 110 15366 130 15371
rect 60 15341 67 15351
rect 76 15341 77 15361
rect 96 15332 99 15366
rect 109 15341 110 15361
rect 119 15341 126 15351
rect 76 15325 92 15331
rect 94 15325 110 15331
rect 170 15325 172 15375
rect 186 15309 190 15343
rect 216 15309 220 15343
rect 213 15277 224 15309
rect 282 15305 292 15389
rect 296 15383 368 15391
rect 378 15383 450 15391
rect 468 15388 473 15422
rect 428 15353 430 15369
rect 251 15277 292 15305
rect 12 15272 62 15274
rect 28 15263 59 15265
rect 62 15263 64 15272
rect 251 15271 263 15277
rect 28 15255 64 15263
rect 127 15263 158 15265
rect 127 15256 182 15263
rect 127 15255 161 15256
rect 59 15239 64 15255
rect 158 15239 161 15255
rect 253 15243 263 15271
rect 273 15243 292 15277
rect 318 15284 324 15353
rect 318 15274 335 15284
rect 303 15252 316 15268
rect 28 15231 64 15239
rect 127 15238 161 15239
rect 127 15231 182 15238
rect 62 15222 64 15231
rect 282 15185 292 15243
rect 303 15234 316 15250
rect 318 15221 324 15274
rect 346 15268 348 15353
rect 400 15345 430 15353
rect 476 15351 480 15419
rect 511 15388 582 15422
rect 544 15381 548 15388
rect 400 15341 434 15345
rect 400 15311 408 15341
rect 420 15311 434 15341
rect 544 15343 548 15351
rect 333 15234 353 15268
rect 428 15264 430 15311
rect 476 15271 480 15339
rect 544 15309 552 15343
rect 578 15309 582 15343
rect 544 15301 548 15309
rect 346 15221 348 15234
rect 367 15230 380 15264
rect 396 15230 408 15264
rect 420 15230 434 15264
rect 544 15261 553 15289
rect 319 15218 335 15220
rect 120 15169 170 15171
rect 76 15163 92 15169
rect 94 15163 110 15169
rect 76 15153 99 15162
rect 60 15143 67 15153
rect 76 15133 77 15153
rect 96 15128 99 15153
rect 109 15133 110 15153
rect 119 15143 126 15153
rect 76 15119 110 15123
rect 170 15119 172 15169
rect 186 15151 190 15185
rect 216 15151 220 15185
rect 182 15113 224 15114
rect 186 15072 220 15106
rect 223 15072 257 15106
rect 160 15065 182 15071
rect 224 15065 246 15071
rect 288 15065 292 15185
rect 296 15183 368 15191
rect 428 15183 430 15230
rect 476 15193 480 15261
rect 485 15217 495 15251
rect 505 15217 519 15251
rect 544 15217 555 15261
rect 485 15193 492 15217
rect 579 15202 582 15292
rect 599 15272 649 15274
rect 610 15264 624 15265
rect 607 15263 624 15264
rect 586 15256 644 15263
rect 607 15255 644 15256
rect 607 15239 610 15255
rect 616 15239 644 15255
rect 607 15238 644 15239
rect 586 15231 644 15238
rect 607 15230 610 15231
rect 649 15222 651 15272
rect 544 15185 548 15193
rect 400 15153 408 15183
rect 420 15153 434 15183
rect 400 15149 434 15153
rect 400 15141 430 15149
rect 428 15125 430 15141
rect 476 15113 480 15181
rect 544 15151 552 15185
rect 578 15151 582 15185
rect 544 15143 548 15151
rect 295 15072 300 15106
rect 324 15072 329 15106
rect 378 15103 450 15111
rect 544 15108 548 15113
rect 544 15104 582 15108
rect 544 15074 552 15104
rect 578 15074 582 15104
rect 544 15071 548 15074
rect 522 15065 548 15071
rect 586 15065 608 15071
rect 182 15049 224 15065
rect 544 15049 586 15065
rect 17 15035 67 15037
rect 119 15035 169 15037
rect 599 15035 649 15037
rect 42 14993 59 15027
rect 67 14985 69 15035
rect 160 15027 246 15035
rect 522 15027 608 15035
rect 76 14993 110 15027
rect 127 14993 144 15027
rect 152 14993 161 15027
rect 162 15025 195 15027
rect 224 15025 244 15027
rect 162 14993 244 15025
rect 524 15025 548 15027
rect 573 15025 582 15027
rect 586 15025 606 15027
rect 160 14985 246 14993
rect 186 14969 220 14971
rect 182 14955 224 14956
rect 160 14949 182 14955
rect 224 14949 246 14955
rect 186 14914 220 14948
rect 223 14914 257 14948
rect 120 14901 170 14903
rect 76 14897 130 14901
rect 110 14892 130 14897
rect 60 14867 67 14877
rect 76 14867 77 14887
rect 96 14858 99 14892
rect 109 14867 110 14887
rect 119 14867 126 14877
rect 76 14851 92 14857
rect 94 14851 110 14857
rect 170 14851 172 14901
rect 186 14835 190 14869
rect 216 14835 220 14869
rect 288 14835 292 15023
rect 476 14955 480 15023
rect 524 14993 606 15025
rect 607 14993 616 15027
rect 522 14985 608 14993
rect 649 14985 651 15035
rect 548 14969 582 14971
rect 522 14950 548 14955
rect 522 14949 582 14950
rect 586 14949 608 14955
rect 295 14914 300 14948
rect 324 14914 329 14948
rect 544 14946 582 14949
rect 378 14909 450 14917
rect 428 14879 430 14895
rect 400 14871 430 14879
rect 476 14877 480 14945
rect 544 14916 552 14946
rect 578 14916 582 14946
rect 544 14907 548 14916
rect 400 14867 434 14871
rect 400 14837 408 14867
rect 420 14837 434 14867
rect 544 14869 548 14877
rect 12 14798 62 14800
rect 28 14789 59 14791
rect 62 14789 64 14798
rect 28 14781 64 14789
rect 127 14789 158 14791
rect 127 14782 182 14789
rect 215 14787 224 14815
rect 127 14781 161 14782
rect 59 14765 64 14781
rect 158 14765 161 14781
rect 28 14757 64 14765
rect 127 14764 161 14765
rect 127 14757 182 14764
rect 62 14748 64 14757
rect 213 14749 224 14787
rect 282 14777 292 14835
rect 296 14829 368 14837
rect 319 14800 335 14802
rect 251 14743 263 14777
rect 273 14743 292 14777
rect 303 14770 316 14786
rect 303 14752 316 14768
rect 120 14695 170 14697
rect 76 14689 92 14695
rect 94 14689 110 14695
rect 76 14679 99 14688
rect 60 14669 67 14679
rect 76 14659 77 14679
rect 96 14654 99 14679
rect 109 14659 110 14679
rect 119 14669 126 14679
rect 76 14645 110 14649
rect 170 14645 172 14695
rect 186 14677 190 14711
rect 216 14677 220 14711
rect 186 14600 220 14634
rect 282 14631 292 14743
rect 318 14746 324 14799
rect 346 14786 348 14799
rect 428 14790 430 14837
rect 443 14827 450 14829
rect 476 14797 480 14865
rect 544 14835 552 14869
rect 578 14835 582 14869
rect 481 14803 517 14831
rect 481 14797 495 14803
rect 333 14752 353 14786
rect 367 14756 380 14790
rect 396 14756 408 14790
rect 420 14756 434 14790
rect 318 14736 335 14746
rect 318 14667 324 14736
rect 346 14667 348 14752
rect 428 14709 430 14756
rect 476 14719 480 14787
rect 485 14769 495 14797
rect 505 14769 519 14803
rect 544 14797 555 14835
rect 544 14769 553 14797
rect 544 14749 548 14769
rect 579 14728 582 14818
rect 599 14798 649 14800
rect 610 14790 624 14791
rect 607 14789 624 14790
rect 586 14782 644 14789
rect 607 14781 644 14782
rect 607 14765 610 14781
rect 616 14765 644 14781
rect 607 14764 644 14765
rect 586 14757 644 14764
rect 607 14756 610 14757
rect 649 14748 651 14798
rect 544 14711 548 14719
rect 400 14679 408 14709
rect 420 14679 434 14709
rect 400 14675 434 14679
rect 400 14667 430 14675
rect 428 14651 430 14667
rect 476 14639 480 14707
rect 544 14677 552 14711
rect 578 14677 582 14711
rect 544 14669 548 14677
rect 544 14639 586 14640
rect 288 14599 292 14631
rect 296 14629 368 14637
rect 378 14629 450 14637
rect 544 14632 548 14639
rect 439 14601 444 14629
rect 120 14585 170 14587
rect 76 14581 130 14585
rect 110 14576 130 14581
rect 60 14551 67 14561
rect 76 14551 77 14571
rect 96 14542 99 14576
rect 109 14551 110 14571
rect 119 14551 126 14561
rect 76 14535 92 14541
rect 94 14535 110 14541
rect 170 14535 172 14585
rect 186 14519 190 14553
rect 216 14519 220 14553
rect 213 14487 224 14519
rect 282 14515 292 14599
rect 296 14593 368 14601
rect 378 14593 450 14601
rect 468 14598 473 14632
rect 428 14563 430 14579
rect 251 14487 292 14515
rect 12 14482 62 14484
rect 28 14473 59 14475
rect 62 14473 64 14482
rect 251 14481 263 14487
rect 28 14465 64 14473
rect 127 14473 158 14475
rect 127 14466 182 14473
rect 127 14465 161 14466
rect 59 14449 64 14465
rect 158 14449 161 14465
rect 253 14453 263 14481
rect 273 14453 292 14487
rect 318 14494 324 14563
rect 318 14484 335 14494
rect 303 14462 316 14478
rect 28 14441 64 14449
rect 127 14448 161 14449
rect 127 14441 182 14448
rect 62 14432 64 14441
rect 282 14395 292 14453
rect 303 14444 316 14460
rect 318 14431 324 14484
rect 346 14478 348 14563
rect 400 14555 430 14563
rect 476 14561 480 14629
rect 511 14598 582 14632
rect 544 14591 548 14598
rect 400 14551 434 14555
rect 400 14521 408 14551
rect 420 14521 434 14551
rect 544 14553 548 14561
rect 333 14444 353 14478
rect 428 14474 430 14521
rect 476 14481 480 14549
rect 544 14519 552 14553
rect 578 14519 582 14553
rect 544 14511 548 14519
rect 346 14431 348 14444
rect 367 14440 380 14474
rect 396 14440 408 14474
rect 420 14440 434 14474
rect 544 14471 553 14499
rect 319 14428 335 14430
rect 120 14379 170 14381
rect 76 14373 92 14379
rect 94 14373 110 14379
rect 76 14363 99 14372
rect 60 14353 67 14363
rect 76 14343 77 14363
rect 96 14338 99 14363
rect 109 14343 110 14363
rect 119 14353 126 14363
rect 76 14329 110 14333
rect 170 14329 172 14379
rect 186 14361 190 14395
rect 216 14361 220 14395
rect 182 14323 224 14324
rect 186 14282 220 14316
rect 223 14282 257 14316
rect 160 14275 182 14281
rect 224 14275 246 14281
rect 288 14275 292 14395
rect 296 14393 368 14401
rect 428 14393 430 14440
rect 476 14403 480 14471
rect 485 14427 495 14461
rect 505 14427 519 14461
rect 544 14427 555 14471
rect 485 14403 492 14427
rect 579 14412 582 14502
rect 599 14482 649 14484
rect 610 14474 624 14475
rect 607 14473 624 14474
rect 586 14466 644 14473
rect 607 14465 644 14466
rect 607 14449 610 14465
rect 616 14449 644 14465
rect 607 14448 644 14449
rect 586 14441 644 14448
rect 607 14440 610 14441
rect 649 14432 651 14482
rect 544 14395 548 14403
rect 400 14363 408 14393
rect 420 14363 434 14393
rect 400 14359 434 14363
rect 400 14351 430 14359
rect 428 14335 430 14351
rect 476 14323 480 14391
rect 544 14361 552 14395
rect 578 14361 582 14395
rect 544 14353 548 14361
rect 295 14282 300 14316
rect 324 14282 329 14316
rect 378 14313 450 14321
rect 544 14318 548 14323
rect 544 14314 582 14318
rect 544 14284 552 14314
rect 578 14284 582 14314
rect 544 14281 548 14284
rect 522 14275 548 14281
rect 586 14275 608 14281
rect 182 14259 224 14275
rect 544 14259 586 14275
rect 17 14245 67 14247
rect 119 14245 169 14247
rect 599 14245 649 14247
rect 42 14203 59 14237
rect 67 14195 69 14245
rect 160 14237 246 14245
rect 522 14237 608 14245
rect 76 14203 110 14237
rect 127 14203 144 14237
rect 152 14203 161 14237
rect 162 14235 195 14237
rect 224 14235 244 14237
rect 162 14203 244 14235
rect 524 14235 548 14237
rect 573 14235 582 14237
rect 586 14235 606 14237
rect 160 14195 246 14203
rect 186 14179 220 14181
rect 182 14165 224 14166
rect 160 14159 182 14165
rect 224 14159 246 14165
rect 186 14124 220 14158
rect 223 14124 257 14158
rect 120 14111 170 14113
rect 76 14107 130 14111
rect 110 14102 130 14107
rect 60 14077 67 14087
rect 76 14077 77 14097
rect 96 14068 99 14102
rect 109 14077 110 14097
rect 119 14077 126 14087
rect 76 14061 92 14067
rect 94 14061 110 14067
rect 170 14061 172 14111
rect 186 14045 190 14079
rect 216 14045 220 14079
rect 288 14045 292 14233
rect 476 14165 480 14233
rect 524 14203 606 14235
rect 607 14203 616 14237
rect 522 14195 608 14203
rect 649 14195 651 14245
rect 548 14179 582 14181
rect 522 14160 548 14165
rect 522 14159 582 14160
rect 586 14159 608 14165
rect 295 14124 300 14158
rect 324 14124 329 14158
rect 544 14156 582 14159
rect 378 14119 450 14127
rect 428 14089 430 14105
rect 400 14081 430 14089
rect 476 14087 480 14155
rect 544 14126 552 14156
rect 578 14126 582 14156
rect 544 14117 548 14126
rect 400 14077 434 14081
rect 400 14047 408 14077
rect 420 14047 434 14077
rect 544 14079 548 14087
rect 12 14008 62 14010
rect 28 13999 59 14001
rect 62 13999 64 14008
rect 28 13991 64 13999
rect 127 13999 158 14001
rect 127 13992 182 13999
rect 215 13997 224 14025
rect 127 13991 161 13992
rect 59 13975 64 13991
rect 158 13975 161 13991
rect 28 13967 64 13975
rect 127 13974 161 13975
rect 127 13967 182 13974
rect 62 13958 64 13967
rect 213 13959 224 13997
rect 282 13987 292 14045
rect 296 14039 368 14047
rect 319 14010 335 14012
rect 251 13953 263 13987
rect 273 13953 292 13987
rect 303 13980 316 13996
rect 303 13962 316 13978
rect 120 13905 170 13907
rect 76 13899 92 13905
rect 94 13899 110 13905
rect 76 13889 99 13898
rect 60 13879 67 13889
rect 76 13869 77 13889
rect 96 13864 99 13889
rect 109 13869 110 13889
rect 119 13879 126 13889
rect 76 13855 110 13859
rect 170 13855 172 13905
rect 186 13887 190 13921
rect 216 13887 220 13921
rect 186 13810 220 13844
rect 282 13841 292 13953
rect 318 13956 324 14009
rect 346 13996 348 14009
rect 428 14000 430 14047
rect 443 14037 450 14039
rect 476 14007 480 14075
rect 544 14045 552 14079
rect 578 14045 582 14079
rect 481 14013 517 14041
rect 481 14007 495 14013
rect 333 13962 353 13996
rect 367 13966 380 14000
rect 396 13966 408 14000
rect 420 13966 434 14000
rect 318 13946 335 13956
rect 318 13877 324 13946
rect 346 13877 348 13962
rect 428 13919 430 13966
rect 476 13929 480 13997
rect 485 13979 495 14007
rect 505 13979 519 14013
rect 544 14007 555 14045
rect 544 13979 553 14007
rect 544 13959 548 13979
rect 579 13938 582 14028
rect 599 14008 649 14010
rect 610 14000 624 14001
rect 607 13999 624 14000
rect 586 13992 644 13999
rect 607 13991 644 13992
rect 607 13975 610 13991
rect 616 13975 644 13991
rect 607 13974 644 13975
rect 586 13967 644 13974
rect 607 13966 610 13967
rect 649 13958 651 14008
rect 544 13921 548 13929
rect 400 13889 408 13919
rect 420 13889 434 13919
rect 400 13885 434 13889
rect 400 13877 430 13885
rect 428 13861 430 13877
rect 476 13849 480 13917
rect 544 13887 552 13921
rect 578 13887 582 13921
rect 544 13879 548 13887
rect 544 13849 586 13850
rect 288 13809 292 13841
rect 296 13839 368 13847
rect 378 13839 450 13847
rect 544 13842 548 13849
rect 439 13811 444 13839
rect 120 13795 170 13797
rect 76 13791 130 13795
rect 110 13786 130 13791
rect 60 13761 67 13771
rect 76 13761 77 13781
rect 96 13752 99 13786
rect 109 13761 110 13781
rect 119 13761 126 13771
rect 76 13745 92 13751
rect 94 13745 110 13751
rect 170 13745 172 13795
rect 186 13729 190 13763
rect 216 13729 220 13763
rect 213 13697 224 13729
rect 282 13725 292 13809
rect 296 13803 368 13811
rect 378 13803 450 13811
rect 468 13808 473 13842
rect 428 13773 430 13789
rect 251 13697 292 13725
rect 12 13692 62 13694
rect 28 13683 59 13685
rect 62 13683 64 13692
rect 251 13691 263 13697
rect 28 13675 64 13683
rect 127 13683 158 13685
rect 127 13676 182 13683
rect 127 13675 161 13676
rect 59 13659 64 13675
rect 158 13659 161 13675
rect 253 13663 263 13691
rect 273 13663 292 13697
rect 318 13704 324 13773
rect 318 13694 335 13704
rect 303 13672 316 13688
rect 28 13651 64 13659
rect 127 13658 161 13659
rect 127 13651 182 13658
rect 62 13642 64 13651
rect 282 13605 292 13663
rect 303 13654 316 13670
rect 318 13641 324 13694
rect 346 13688 348 13773
rect 400 13765 430 13773
rect 476 13771 480 13839
rect 511 13808 582 13842
rect 544 13801 548 13808
rect 400 13761 434 13765
rect 400 13731 408 13761
rect 420 13731 434 13761
rect 544 13763 548 13771
rect 333 13654 353 13688
rect 428 13684 430 13731
rect 476 13691 480 13759
rect 544 13729 552 13763
rect 578 13729 582 13763
rect 544 13721 548 13729
rect 346 13641 348 13654
rect 367 13650 380 13684
rect 396 13650 408 13684
rect 420 13650 434 13684
rect 544 13681 553 13709
rect 319 13638 335 13640
rect 120 13589 170 13591
rect 76 13583 92 13589
rect 94 13583 110 13589
rect 76 13573 99 13582
rect 60 13563 67 13573
rect 76 13553 77 13573
rect 96 13548 99 13573
rect 109 13553 110 13573
rect 119 13563 126 13573
rect 76 13539 110 13543
rect 170 13539 172 13589
rect 186 13571 190 13605
rect 216 13571 220 13605
rect 182 13533 224 13534
rect 186 13492 220 13526
rect 223 13492 257 13526
rect 160 13485 182 13491
rect 224 13485 246 13491
rect 288 13485 292 13605
rect 296 13603 368 13611
rect 428 13603 430 13650
rect 476 13613 480 13681
rect 485 13637 495 13671
rect 505 13637 519 13671
rect 544 13637 555 13681
rect 485 13613 492 13637
rect 579 13622 582 13712
rect 599 13692 649 13694
rect 610 13684 624 13685
rect 607 13683 624 13684
rect 586 13676 644 13683
rect 607 13675 644 13676
rect 607 13659 610 13675
rect 616 13659 644 13675
rect 607 13658 644 13659
rect 586 13651 644 13658
rect 607 13650 610 13651
rect 649 13642 651 13692
rect 544 13605 548 13613
rect 400 13573 408 13603
rect 420 13573 434 13603
rect 400 13569 434 13573
rect 400 13561 430 13569
rect 428 13545 430 13561
rect 476 13533 480 13601
rect 544 13571 552 13605
rect 578 13571 582 13605
rect 544 13563 548 13571
rect 295 13492 300 13526
rect 324 13492 329 13526
rect 378 13523 450 13531
rect 544 13528 548 13533
rect 544 13524 582 13528
rect 544 13494 552 13524
rect 578 13494 582 13524
rect 544 13491 548 13494
rect 522 13485 548 13491
rect 586 13485 608 13491
rect 182 13469 224 13485
rect 544 13469 586 13485
rect 17 13455 67 13457
rect 119 13455 169 13457
rect 599 13455 649 13457
rect 42 13413 59 13447
rect 67 13405 69 13455
rect 160 13447 246 13455
rect 522 13447 608 13455
rect 76 13413 110 13447
rect 127 13413 144 13447
rect 152 13413 161 13447
rect 162 13445 195 13447
rect 224 13445 244 13447
rect 162 13413 244 13445
rect 524 13445 548 13447
rect 573 13445 582 13447
rect 586 13445 606 13447
rect 160 13405 246 13413
rect 186 13389 220 13391
rect 182 13375 224 13376
rect 160 13369 182 13375
rect 224 13369 246 13375
rect 186 13334 220 13368
rect 223 13334 257 13368
rect 120 13321 170 13323
rect 76 13317 130 13321
rect 110 13312 130 13317
rect 60 13287 67 13297
rect 76 13287 77 13307
rect 96 13278 99 13312
rect 109 13287 110 13307
rect 119 13287 126 13297
rect 76 13271 92 13277
rect 94 13271 110 13277
rect 170 13271 172 13321
rect 186 13255 190 13289
rect 216 13255 220 13289
rect 288 13255 292 13443
rect 476 13375 480 13443
rect 524 13413 606 13445
rect 607 13413 616 13447
rect 522 13405 608 13413
rect 649 13405 651 13455
rect 548 13389 582 13391
rect 522 13370 548 13375
rect 522 13369 582 13370
rect 586 13369 608 13375
rect 295 13334 300 13368
rect 324 13334 329 13368
rect 544 13366 582 13369
rect 378 13329 450 13337
rect 428 13299 430 13315
rect 400 13291 430 13299
rect 476 13297 480 13365
rect 544 13336 552 13366
rect 578 13336 582 13366
rect 544 13327 548 13336
rect 400 13287 434 13291
rect 400 13257 408 13287
rect 420 13257 434 13287
rect 544 13289 548 13297
rect 12 13218 62 13220
rect 28 13209 59 13211
rect 62 13209 64 13218
rect 28 13201 64 13209
rect 127 13209 158 13211
rect 127 13202 182 13209
rect 215 13207 224 13235
rect 127 13201 161 13202
rect 59 13185 64 13201
rect 158 13185 161 13201
rect 28 13177 64 13185
rect 127 13184 161 13185
rect 127 13177 182 13184
rect 62 13168 64 13177
rect 213 13169 224 13207
rect 282 13197 292 13255
rect 296 13249 368 13257
rect 319 13220 335 13222
rect 251 13163 263 13197
rect 273 13163 292 13197
rect 303 13190 316 13206
rect 303 13172 316 13188
rect 120 13115 170 13117
rect 76 13109 92 13115
rect 94 13109 110 13115
rect 76 13099 99 13108
rect 60 13089 67 13099
rect 76 13079 77 13099
rect 96 13074 99 13099
rect 109 13079 110 13099
rect 119 13089 126 13099
rect 76 13065 110 13069
rect 170 13065 172 13115
rect 186 13097 190 13131
rect 216 13097 220 13131
rect 186 13020 220 13054
rect 282 13051 292 13163
rect 318 13166 324 13219
rect 346 13206 348 13219
rect 428 13210 430 13257
rect 443 13247 450 13249
rect 476 13217 480 13285
rect 544 13255 552 13289
rect 578 13255 582 13289
rect 481 13223 517 13251
rect 481 13217 495 13223
rect 333 13172 353 13206
rect 367 13176 380 13210
rect 396 13176 408 13210
rect 420 13176 434 13210
rect 318 13156 335 13166
rect 318 13087 324 13156
rect 346 13087 348 13172
rect 428 13129 430 13176
rect 476 13139 480 13207
rect 485 13189 495 13217
rect 505 13189 519 13223
rect 544 13217 555 13255
rect 544 13189 553 13217
rect 544 13169 548 13189
rect 579 13148 582 13238
rect 599 13218 649 13220
rect 610 13210 624 13211
rect 607 13209 624 13210
rect 586 13202 644 13209
rect 607 13201 644 13202
rect 607 13185 610 13201
rect 616 13185 644 13201
rect 607 13184 644 13185
rect 586 13177 644 13184
rect 607 13176 610 13177
rect 649 13168 651 13218
rect 544 13131 548 13139
rect 400 13099 408 13129
rect 420 13099 434 13129
rect 400 13095 434 13099
rect 400 13087 430 13095
rect 428 13071 430 13087
rect 476 13059 480 13127
rect 544 13097 552 13131
rect 578 13097 582 13131
rect 544 13089 548 13097
rect 544 13059 586 13060
rect 288 13019 292 13051
rect 296 13049 368 13057
rect 378 13049 450 13057
rect 544 13052 548 13059
rect 439 13021 444 13049
rect 120 13005 170 13007
rect 76 13001 130 13005
rect 110 12996 130 13001
rect 60 12971 67 12981
rect 76 12971 77 12991
rect 96 12962 99 12996
rect 109 12971 110 12991
rect 119 12971 126 12981
rect 76 12955 92 12961
rect 94 12955 110 12961
rect 170 12955 172 13005
rect 186 12939 190 12973
rect 216 12939 220 12973
rect 213 12907 224 12939
rect 282 12935 292 13019
rect 296 13013 368 13021
rect 378 13013 450 13021
rect 468 13018 473 13052
rect 428 12983 430 12999
rect 251 12907 292 12935
rect 12 12902 62 12904
rect 28 12893 59 12895
rect 62 12893 64 12902
rect 251 12901 263 12907
rect 28 12885 64 12893
rect 127 12893 158 12895
rect 127 12886 182 12893
rect 127 12885 161 12886
rect 59 12869 64 12885
rect 158 12869 161 12885
rect 253 12873 263 12901
rect 273 12873 292 12907
rect 318 12914 324 12983
rect 318 12904 335 12914
rect 303 12882 316 12898
rect 28 12861 64 12869
rect 127 12868 161 12869
rect 127 12861 182 12868
rect 62 12852 64 12861
rect 282 12815 292 12873
rect 303 12864 316 12880
rect 318 12851 324 12904
rect 346 12898 348 12983
rect 400 12975 430 12983
rect 476 12981 480 13049
rect 511 13018 582 13052
rect 544 13011 548 13018
rect 400 12971 434 12975
rect 400 12941 408 12971
rect 420 12941 434 12971
rect 544 12973 548 12981
rect 333 12864 353 12898
rect 428 12894 430 12941
rect 476 12901 480 12969
rect 544 12939 552 12973
rect 578 12939 582 12973
rect 544 12931 548 12939
rect 346 12851 348 12864
rect 367 12860 380 12894
rect 396 12860 408 12894
rect 420 12860 434 12894
rect 544 12891 553 12919
rect 319 12848 335 12850
rect 120 12799 170 12801
rect 76 12793 92 12799
rect 94 12793 110 12799
rect 76 12783 99 12792
rect 60 12773 67 12783
rect 76 12763 77 12783
rect 96 12758 99 12783
rect 109 12763 110 12783
rect 119 12773 126 12783
rect 76 12749 110 12753
rect 170 12749 172 12799
rect 186 12781 190 12815
rect 216 12781 220 12815
rect 182 12743 224 12744
rect 186 12702 220 12736
rect 223 12702 257 12736
rect 160 12695 182 12701
rect 224 12695 246 12701
rect 288 12695 292 12815
rect 296 12813 368 12821
rect 428 12813 430 12860
rect 476 12823 480 12891
rect 485 12847 495 12881
rect 505 12847 519 12881
rect 544 12847 555 12891
rect 485 12823 492 12847
rect 579 12832 582 12922
rect 599 12902 649 12904
rect 610 12894 624 12895
rect 607 12893 624 12894
rect 586 12886 644 12893
rect 607 12885 644 12886
rect 607 12869 610 12885
rect 616 12869 644 12885
rect 607 12868 644 12869
rect 586 12861 644 12868
rect 607 12860 610 12861
rect 649 12852 651 12902
rect 544 12815 548 12823
rect 400 12783 408 12813
rect 420 12783 434 12813
rect 400 12779 434 12783
rect 400 12771 430 12779
rect 428 12755 430 12771
rect 476 12743 480 12811
rect 544 12781 552 12815
rect 578 12781 582 12815
rect 544 12773 548 12781
rect 295 12702 300 12736
rect 324 12702 329 12736
rect 378 12733 450 12741
rect 544 12738 548 12743
rect 544 12734 582 12738
rect 544 12704 552 12734
rect 578 12704 582 12734
rect 544 12701 548 12704
rect 522 12695 548 12701
rect 586 12695 608 12701
rect 182 12679 224 12695
rect 544 12679 586 12695
rect 17 12665 67 12667
rect 119 12665 169 12667
rect 599 12665 649 12667
rect 42 12623 59 12657
rect 67 12615 69 12665
rect 160 12657 246 12665
rect 522 12657 608 12665
rect 76 12623 110 12657
rect 127 12623 144 12657
rect 152 12623 161 12657
rect 162 12655 195 12657
rect 224 12655 244 12657
rect 162 12623 244 12655
rect 524 12655 548 12657
rect 573 12655 582 12657
rect 586 12655 606 12657
rect 160 12615 246 12623
rect 186 12599 220 12601
rect 182 12585 224 12586
rect 160 12579 182 12585
rect 224 12579 246 12585
rect 186 12544 220 12578
rect 223 12544 257 12578
rect 120 12531 170 12533
rect 76 12527 130 12531
rect 110 12522 130 12527
rect 60 12497 67 12507
rect 76 12497 77 12517
rect 96 12488 99 12522
rect 109 12497 110 12517
rect 119 12497 126 12507
rect 76 12481 92 12487
rect 94 12481 110 12487
rect 170 12481 172 12531
rect 186 12465 190 12499
rect 216 12465 220 12499
rect 288 12465 292 12653
rect 476 12585 480 12653
rect 524 12623 606 12655
rect 607 12623 616 12657
rect 522 12615 608 12623
rect 649 12615 651 12665
rect 548 12599 582 12601
rect 522 12580 548 12585
rect 522 12579 582 12580
rect 586 12579 608 12585
rect 295 12544 300 12578
rect 324 12544 329 12578
rect 544 12576 582 12579
rect 378 12539 450 12547
rect 428 12509 430 12525
rect 400 12501 430 12509
rect 476 12507 480 12575
rect 544 12546 552 12576
rect 578 12546 582 12576
rect 544 12537 548 12546
rect 400 12497 434 12501
rect 400 12467 408 12497
rect 420 12467 434 12497
rect 544 12499 548 12507
rect 12 12428 62 12430
rect 28 12419 59 12421
rect 62 12419 64 12428
rect 28 12411 64 12419
rect 127 12419 158 12421
rect 127 12412 182 12419
rect 215 12417 224 12445
rect 127 12411 161 12412
rect 59 12395 64 12411
rect 158 12395 161 12411
rect 28 12387 64 12395
rect 127 12394 161 12395
rect 127 12387 182 12394
rect 62 12378 64 12387
rect 213 12379 224 12417
rect 282 12407 292 12465
rect 296 12459 368 12467
rect 319 12430 335 12432
rect 251 12373 263 12407
rect 273 12373 292 12407
rect 303 12400 316 12416
rect 303 12382 316 12398
rect 120 12325 170 12327
rect 76 12319 92 12325
rect 94 12319 110 12325
rect 76 12309 99 12318
rect 60 12299 67 12309
rect 76 12289 77 12309
rect 96 12284 99 12309
rect 109 12289 110 12309
rect 119 12299 126 12309
rect 76 12275 110 12279
rect 170 12275 172 12325
rect 186 12307 190 12341
rect 216 12307 220 12341
rect 186 12230 220 12264
rect 282 12261 292 12373
rect 318 12376 324 12429
rect 346 12416 348 12429
rect 428 12420 430 12467
rect 443 12457 450 12459
rect 476 12427 480 12495
rect 544 12465 552 12499
rect 578 12465 582 12499
rect 481 12433 517 12461
rect 481 12427 495 12433
rect 333 12382 353 12416
rect 367 12386 380 12420
rect 396 12386 408 12420
rect 420 12386 434 12420
rect 318 12366 335 12376
rect 318 12297 324 12366
rect 346 12297 348 12382
rect 428 12339 430 12386
rect 476 12349 480 12417
rect 485 12399 495 12427
rect 505 12399 519 12433
rect 544 12427 555 12465
rect 544 12399 553 12427
rect 544 12379 548 12399
rect 579 12358 582 12448
rect 599 12428 649 12430
rect 610 12420 624 12421
rect 607 12419 624 12420
rect 586 12412 644 12419
rect 607 12411 644 12412
rect 607 12395 610 12411
rect 616 12395 644 12411
rect 607 12394 644 12395
rect 586 12387 644 12394
rect 607 12386 610 12387
rect 649 12378 651 12428
rect 544 12341 548 12349
rect 400 12309 408 12339
rect 420 12309 434 12339
rect 400 12305 434 12309
rect 400 12297 430 12305
rect 428 12281 430 12297
rect 476 12269 480 12337
rect 544 12307 552 12341
rect 578 12307 582 12341
rect 544 12299 548 12307
rect 544 12269 586 12270
rect 288 12229 292 12261
rect 296 12259 368 12267
rect 378 12259 450 12267
rect 544 12262 548 12269
rect 439 12231 444 12259
rect 120 12215 170 12217
rect 76 12211 130 12215
rect 110 12206 130 12211
rect 60 12181 67 12191
rect 76 12181 77 12201
rect 96 12172 99 12206
rect 109 12181 110 12201
rect 119 12181 126 12191
rect 76 12165 92 12171
rect 94 12165 110 12171
rect 170 12165 172 12215
rect 186 12149 190 12183
rect 216 12149 220 12183
rect 213 12117 224 12149
rect 282 12145 292 12229
rect 296 12223 368 12231
rect 378 12223 450 12231
rect 468 12228 473 12262
rect 428 12193 430 12209
rect 251 12117 292 12145
rect 12 12112 62 12114
rect 28 12103 59 12105
rect 62 12103 64 12112
rect 251 12111 263 12117
rect 28 12095 64 12103
rect 127 12103 158 12105
rect 127 12096 182 12103
rect 127 12095 161 12096
rect 59 12079 64 12095
rect 158 12079 161 12095
rect 253 12083 263 12111
rect 273 12083 292 12117
rect 318 12124 324 12193
rect 318 12114 335 12124
rect 303 12092 316 12108
rect 28 12071 64 12079
rect 127 12078 161 12079
rect 127 12071 182 12078
rect 62 12062 64 12071
rect 282 12025 292 12083
rect 303 12074 316 12090
rect 318 12061 324 12114
rect 346 12108 348 12193
rect 400 12185 430 12193
rect 476 12191 480 12259
rect 511 12228 582 12262
rect 544 12221 548 12228
rect 400 12181 434 12185
rect 400 12151 408 12181
rect 420 12151 434 12181
rect 544 12183 548 12191
rect 333 12074 353 12108
rect 428 12104 430 12151
rect 476 12111 480 12179
rect 544 12149 552 12183
rect 578 12149 582 12183
rect 544 12141 548 12149
rect 346 12061 348 12074
rect 367 12070 380 12104
rect 396 12070 408 12104
rect 420 12070 434 12104
rect 544 12101 553 12129
rect 319 12058 335 12060
rect 120 12009 170 12011
rect 76 12003 92 12009
rect 94 12003 110 12009
rect 76 11993 99 12002
rect 60 11983 67 11993
rect 76 11973 77 11993
rect 96 11968 99 11993
rect 109 11973 110 11993
rect 119 11983 126 11993
rect 76 11959 110 11963
rect 170 11959 172 12009
rect 186 11991 190 12025
rect 216 11991 220 12025
rect 182 11953 224 11954
rect 186 11912 220 11946
rect 223 11912 257 11946
rect 160 11905 182 11911
rect 224 11905 246 11911
rect 288 11905 292 12025
rect 296 12023 368 12031
rect 428 12023 430 12070
rect 476 12033 480 12101
rect 485 12057 495 12091
rect 505 12057 519 12091
rect 544 12057 555 12101
rect 485 12033 492 12057
rect 579 12042 582 12132
rect 599 12112 649 12114
rect 610 12104 624 12105
rect 607 12103 624 12104
rect 586 12096 644 12103
rect 607 12095 644 12096
rect 607 12079 610 12095
rect 616 12079 644 12095
rect 607 12078 644 12079
rect 586 12071 644 12078
rect 607 12070 610 12071
rect 649 12062 651 12112
rect 544 12025 548 12033
rect 400 11993 408 12023
rect 420 11993 434 12023
rect 400 11989 434 11993
rect 400 11981 430 11989
rect 428 11965 430 11981
rect 476 11953 480 12021
rect 544 11991 552 12025
rect 578 11991 582 12025
rect 544 11983 548 11991
rect 295 11912 300 11946
rect 324 11912 329 11946
rect 378 11943 450 11951
rect 544 11948 548 11953
rect 544 11944 582 11948
rect 544 11914 552 11944
rect 578 11914 582 11944
rect 544 11911 548 11914
rect 522 11905 548 11911
rect 586 11905 608 11911
rect 182 11889 224 11905
rect 544 11889 586 11905
rect 17 11875 67 11877
rect 119 11875 169 11877
rect 599 11875 649 11877
rect 42 11833 59 11867
rect 67 11825 69 11875
rect 160 11867 246 11875
rect 522 11867 608 11875
rect 76 11833 110 11867
rect 127 11833 144 11867
rect 152 11833 161 11867
rect 162 11865 195 11867
rect 224 11865 244 11867
rect 162 11833 244 11865
rect 524 11865 548 11867
rect 573 11865 582 11867
rect 586 11865 606 11867
rect 160 11825 246 11833
rect 186 11809 220 11811
rect 182 11795 224 11796
rect 160 11789 182 11795
rect 224 11789 246 11795
rect 186 11754 220 11788
rect 223 11754 257 11788
rect 120 11741 170 11743
rect 76 11737 130 11741
rect 110 11732 130 11737
rect 60 11707 67 11717
rect 76 11707 77 11727
rect 96 11698 99 11732
rect 109 11707 110 11727
rect 119 11707 126 11717
rect 76 11691 92 11697
rect 94 11691 110 11697
rect 170 11691 172 11741
rect 186 11675 190 11709
rect 216 11675 220 11709
rect 288 11675 292 11863
rect 476 11795 480 11863
rect 524 11833 606 11865
rect 607 11833 616 11867
rect 522 11825 608 11833
rect 649 11825 651 11875
rect 548 11809 582 11811
rect 522 11790 548 11795
rect 522 11789 582 11790
rect 586 11789 608 11795
rect 295 11754 300 11788
rect 324 11754 329 11788
rect 544 11786 582 11789
rect 378 11749 450 11757
rect 428 11719 430 11735
rect 400 11711 430 11719
rect 476 11717 480 11785
rect 544 11756 552 11786
rect 578 11756 582 11786
rect 544 11747 548 11756
rect 400 11707 434 11711
rect 400 11677 408 11707
rect 420 11677 434 11707
rect 544 11709 548 11717
rect 12 11638 62 11640
rect 28 11629 59 11631
rect 62 11629 64 11638
rect 28 11621 64 11629
rect 127 11629 158 11631
rect 127 11622 182 11629
rect 215 11627 224 11655
rect 127 11621 161 11622
rect 59 11605 64 11621
rect 158 11605 161 11621
rect 28 11597 64 11605
rect 127 11604 161 11605
rect 127 11597 182 11604
rect 62 11588 64 11597
rect 213 11589 224 11627
rect 282 11617 292 11675
rect 296 11669 368 11677
rect 319 11640 335 11642
rect 251 11583 263 11617
rect 273 11583 292 11617
rect 303 11610 316 11626
rect 303 11592 316 11608
rect 120 11535 170 11537
rect 76 11529 92 11535
rect 94 11529 110 11535
rect 76 11519 99 11528
rect 60 11509 67 11519
rect 76 11499 77 11519
rect 96 11494 99 11519
rect 109 11499 110 11519
rect 119 11509 126 11519
rect 76 11485 110 11489
rect 170 11485 172 11535
rect 186 11517 190 11551
rect 216 11517 220 11551
rect 186 11440 220 11474
rect 282 11471 292 11583
rect 318 11586 324 11639
rect 346 11626 348 11639
rect 428 11630 430 11677
rect 443 11667 450 11669
rect 476 11637 480 11705
rect 544 11675 552 11709
rect 578 11675 582 11709
rect 481 11643 517 11671
rect 481 11637 495 11643
rect 333 11592 353 11626
rect 367 11596 380 11630
rect 396 11596 408 11630
rect 420 11596 434 11630
rect 318 11576 335 11586
rect 318 11507 324 11576
rect 346 11507 348 11592
rect 428 11549 430 11596
rect 476 11559 480 11627
rect 485 11609 495 11637
rect 505 11609 519 11643
rect 544 11637 555 11675
rect 544 11609 553 11637
rect 544 11589 548 11609
rect 579 11568 582 11658
rect 599 11638 649 11640
rect 610 11630 624 11631
rect 607 11629 624 11630
rect 586 11622 644 11629
rect 607 11621 644 11622
rect 607 11605 610 11621
rect 616 11605 644 11621
rect 607 11604 644 11605
rect 586 11597 644 11604
rect 607 11596 610 11597
rect 649 11588 651 11638
rect 544 11551 548 11559
rect 400 11519 408 11549
rect 420 11519 434 11549
rect 400 11515 434 11519
rect 400 11507 430 11515
rect 428 11491 430 11507
rect 476 11479 480 11547
rect 544 11517 552 11551
rect 578 11517 582 11551
rect 544 11509 548 11517
rect 544 11479 586 11480
rect 288 11439 292 11471
rect 296 11469 368 11477
rect 378 11469 450 11477
rect 544 11472 548 11479
rect 439 11441 444 11469
rect 120 11425 170 11427
rect 76 11421 130 11425
rect 110 11416 130 11421
rect 60 11391 67 11401
rect 76 11391 77 11411
rect 96 11382 99 11416
rect 109 11391 110 11411
rect 119 11391 126 11401
rect 76 11375 92 11381
rect 94 11375 110 11381
rect 170 11375 172 11425
rect 186 11359 190 11393
rect 216 11359 220 11393
rect 213 11327 224 11359
rect 282 11355 292 11439
rect 296 11433 368 11441
rect 378 11433 450 11441
rect 468 11438 473 11472
rect 428 11403 430 11419
rect 251 11327 292 11355
rect 12 11322 62 11324
rect 28 11313 59 11315
rect 62 11313 64 11322
rect 251 11321 263 11327
rect 28 11305 64 11313
rect 127 11313 158 11315
rect 127 11306 182 11313
rect 127 11305 161 11306
rect 59 11289 64 11305
rect 158 11289 161 11305
rect 253 11293 263 11321
rect 273 11293 292 11327
rect 318 11334 324 11403
rect 318 11324 335 11334
rect 303 11302 316 11318
rect 28 11281 64 11289
rect 127 11288 161 11289
rect 127 11281 182 11288
rect 62 11272 64 11281
rect 282 11235 292 11293
rect 303 11284 316 11300
rect 318 11271 324 11324
rect 346 11318 348 11403
rect 400 11395 430 11403
rect 476 11401 480 11469
rect 511 11438 582 11472
rect 544 11431 548 11438
rect 400 11391 434 11395
rect 400 11361 408 11391
rect 420 11361 434 11391
rect 544 11393 548 11401
rect 333 11284 353 11318
rect 428 11314 430 11361
rect 476 11321 480 11389
rect 544 11359 552 11393
rect 578 11359 582 11393
rect 544 11351 548 11359
rect 346 11271 348 11284
rect 367 11280 380 11314
rect 396 11280 408 11314
rect 420 11280 434 11314
rect 544 11311 553 11339
rect 319 11268 335 11270
rect 120 11219 170 11221
rect 76 11213 92 11219
rect 94 11213 110 11219
rect 76 11203 99 11212
rect 60 11193 67 11203
rect 76 11183 77 11203
rect 96 11178 99 11203
rect 109 11183 110 11203
rect 119 11193 126 11203
rect 76 11169 110 11173
rect 170 11169 172 11219
rect 186 11201 190 11235
rect 216 11201 220 11235
rect 182 11163 224 11164
rect 186 11122 220 11156
rect 223 11122 257 11156
rect 160 11115 182 11121
rect 224 11115 246 11121
rect 288 11115 292 11235
rect 296 11233 368 11241
rect 428 11233 430 11280
rect 476 11243 480 11311
rect 485 11267 495 11301
rect 505 11267 519 11301
rect 544 11267 555 11311
rect 485 11243 492 11267
rect 579 11252 582 11342
rect 599 11322 649 11324
rect 610 11314 624 11315
rect 607 11313 624 11314
rect 586 11306 644 11313
rect 607 11305 644 11306
rect 607 11289 610 11305
rect 616 11289 644 11305
rect 607 11288 644 11289
rect 586 11281 644 11288
rect 607 11280 610 11281
rect 649 11272 651 11322
rect 544 11235 548 11243
rect 400 11203 408 11233
rect 420 11203 434 11233
rect 400 11199 434 11203
rect 400 11191 430 11199
rect 428 11175 430 11191
rect 476 11163 480 11231
rect 544 11201 552 11235
rect 578 11201 582 11235
rect 544 11193 548 11201
rect 295 11122 300 11156
rect 324 11122 329 11156
rect 378 11153 450 11161
rect 544 11158 548 11163
rect 544 11154 582 11158
rect 544 11124 552 11154
rect 578 11124 582 11154
rect 544 11121 548 11124
rect 522 11115 548 11121
rect 586 11115 608 11121
rect 182 11099 224 11115
rect 544 11099 586 11115
rect 17 11085 67 11087
rect 119 11085 169 11087
rect 599 11085 649 11087
rect 42 11043 59 11077
rect 67 11035 69 11085
rect 160 11077 246 11085
rect 522 11077 608 11085
rect 76 11043 110 11077
rect 127 11043 144 11077
rect 152 11043 161 11077
rect 162 11075 195 11077
rect 224 11075 244 11077
rect 162 11043 244 11075
rect 524 11075 548 11077
rect 573 11075 582 11077
rect 586 11075 606 11077
rect 160 11035 246 11043
rect 186 11019 220 11021
rect 182 11005 224 11006
rect 160 10999 182 11005
rect 224 10999 246 11005
rect 186 10964 220 10998
rect 223 10964 257 10998
rect 120 10951 170 10953
rect 76 10947 130 10951
rect 110 10942 130 10947
rect 60 10917 67 10927
rect 76 10917 77 10937
rect 96 10908 99 10942
rect 109 10917 110 10937
rect 119 10917 126 10927
rect 76 10901 92 10907
rect 94 10901 110 10907
rect 170 10901 172 10951
rect 186 10885 190 10919
rect 216 10885 220 10919
rect 288 10885 292 11073
rect 476 11005 480 11073
rect 524 11043 606 11075
rect 607 11043 616 11077
rect 522 11035 608 11043
rect 649 11035 651 11085
rect 548 11019 582 11021
rect 522 11000 548 11005
rect 522 10999 582 11000
rect 586 10999 608 11005
rect 295 10964 300 10998
rect 324 10964 329 10998
rect 544 10996 582 10999
rect 378 10959 450 10967
rect 428 10929 430 10945
rect 400 10921 430 10929
rect 476 10927 480 10995
rect 544 10966 552 10996
rect 578 10966 582 10996
rect 544 10957 548 10966
rect 400 10917 434 10921
rect 400 10887 408 10917
rect 420 10887 434 10917
rect 544 10919 548 10927
rect 12 10848 62 10850
rect 28 10839 59 10841
rect 62 10839 64 10848
rect 28 10831 64 10839
rect 127 10839 158 10841
rect 127 10832 182 10839
rect 215 10837 224 10865
rect 127 10831 161 10832
rect 59 10815 64 10831
rect 158 10815 161 10831
rect 28 10807 64 10815
rect 127 10814 161 10815
rect 127 10807 182 10814
rect 62 10798 64 10807
rect 213 10799 224 10837
rect 282 10827 292 10885
rect 296 10879 368 10887
rect 319 10850 335 10852
rect 251 10793 263 10827
rect 273 10793 292 10827
rect 303 10820 316 10836
rect 303 10802 316 10818
rect 120 10745 170 10747
rect 76 10739 92 10745
rect 94 10739 110 10745
rect 76 10729 99 10738
rect 60 10719 67 10729
rect 76 10709 77 10729
rect 96 10704 99 10729
rect 109 10709 110 10729
rect 119 10719 126 10729
rect 76 10695 110 10699
rect 170 10695 172 10745
rect 186 10727 190 10761
rect 216 10727 220 10761
rect 186 10650 220 10684
rect 282 10681 292 10793
rect 318 10796 324 10849
rect 346 10836 348 10849
rect 428 10840 430 10887
rect 443 10877 450 10879
rect 476 10847 480 10915
rect 544 10885 552 10919
rect 578 10885 582 10919
rect 481 10853 517 10881
rect 481 10847 495 10853
rect 333 10802 353 10836
rect 367 10806 380 10840
rect 396 10806 408 10840
rect 420 10806 434 10840
rect 318 10786 335 10796
rect 318 10717 324 10786
rect 346 10717 348 10802
rect 428 10759 430 10806
rect 476 10769 480 10837
rect 485 10819 495 10847
rect 505 10819 519 10853
rect 544 10847 555 10885
rect 544 10819 553 10847
rect 544 10799 548 10819
rect 579 10778 582 10868
rect 599 10848 649 10850
rect 610 10840 624 10841
rect 607 10839 624 10840
rect 586 10832 644 10839
rect 607 10831 644 10832
rect 607 10815 610 10831
rect 616 10815 644 10831
rect 607 10814 644 10815
rect 586 10807 644 10814
rect 607 10806 610 10807
rect 649 10798 651 10848
rect 544 10761 548 10769
rect 400 10729 408 10759
rect 420 10729 434 10759
rect 400 10725 434 10729
rect 400 10717 430 10725
rect 428 10701 430 10717
rect 476 10689 480 10757
rect 544 10727 552 10761
rect 578 10727 582 10761
rect 544 10719 548 10727
rect 544 10689 586 10690
rect 288 10649 292 10681
rect 296 10679 368 10687
rect 378 10679 450 10687
rect 544 10682 548 10689
rect 439 10651 444 10679
rect 120 10635 170 10637
rect 76 10631 130 10635
rect 110 10626 130 10631
rect 60 10601 67 10611
rect 76 10601 77 10621
rect 96 10592 99 10626
rect 109 10601 110 10621
rect 119 10601 126 10611
rect 76 10585 92 10591
rect 94 10585 110 10591
rect 170 10585 172 10635
rect 186 10569 190 10603
rect 216 10569 220 10603
rect 213 10537 224 10569
rect 282 10565 292 10649
rect 296 10643 368 10651
rect 378 10643 450 10651
rect 468 10648 473 10682
rect 428 10613 430 10629
rect 251 10537 292 10565
rect 12 10532 62 10534
rect 28 10523 59 10525
rect 62 10523 64 10532
rect 251 10531 263 10537
rect 28 10515 64 10523
rect 127 10523 158 10525
rect 127 10516 182 10523
rect 127 10515 161 10516
rect 59 10499 64 10515
rect 158 10499 161 10515
rect 253 10503 263 10531
rect 273 10503 292 10537
rect 318 10544 324 10613
rect 318 10534 335 10544
rect 303 10512 316 10528
rect 28 10491 64 10499
rect 127 10498 161 10499
rect 127 10491 182 10498
rect 62 10482 64 10491
rect 282 10445 292 10503
rect 303 10494 316 10510
rect 318 10481 324 10534
rect 346 10528 348 10613
rect 400 10605 430 10613
rect 476 10611 480 10679
rect 511 10648 582 10682
rect 544 10641 548 10648
rect 400 10601 434 10605
rect 400 10571 408 10601
rect 420 10571 434 10601
rect 544 10603 548 10611
rect 333 10494 353 10528
rect 428 10524 430 10571
rect 476 10531 480 10599
rect 544 10569 552 10603
rect 578 10569 582 10603
rect 544 10561 548 10569
rect 346 10481 348 10494
rect 367 10490 380 10524
rect 396 10490 408 10524
rect 420 10490 434 10524
rect 544 10521 553 10549
rect 319 10478 335 10480
rect 120 10429 170 10431
rect 76 10423 92 10429
rect 94 10423 110 10429
rect 76 10413 99 10422
rect 60 10403 67 10413
rect 76 10393 77 10413
rect 96 10388 99 10413
rect 109 10393 110 10413
rect 119 10403 126 10413
rect 76 10379 110 10383
rect 170 10379 172 10429
rect 186 10411 190 10445
rect 216 10411 220 10445
rect 182 10373 224 10374
rect 186 10332 220 10366
rect 223 10332 257 10366
rect 160 10325 182 10331
rect 224 10325 246 10331
rect 288 10325 292 10445
rect 296 10443 368 10451
rect 428 10443 430 10490
rect 476 10453 480 10521
rect 485 10477 495 10511
rect 505 10477 519 10511
rect 544 10477 555 10521
rect 485 10453 492 10477
rect 579 10462 582 10552
rect 599 10532 649 10534
rect 610 10524 624 10525
rect 607 10523 624 10524
rect 586 10516 644 10523
rect 607 10515 644 10516
rect 607 10499 610 10515
rect 616 10499 644 10515
rect 607 10498 644 10499
rect 586 10491 644 10498
rect 607 10490 610 10491
rect 649 10482 651 10532
rect 544 10445 548 10453
rect 400 10413 408 10443
rect 420 10413 434 10443
rect 400 10409 434 10413
rect 400 10401 430 10409
rect 428 10385 430 10401
rect 476 10373 480 10441
rect 544 10411 552 10445
rect 578 10411 582 10445
rect 544 10403 548 10411
rect 295 10332 300 10366
rect 324 10332 329 10366
rect 378 10363 450 10371
rect 544 10368 548 10373
rect 544 10364 582 10368
rect 544 10334 552 10364
rect 578 10334 582 10364
rect 544 10331 548 10334
rect 522 10325 548 10331
rect 586 10325 608 10331
rect 182 10309 224 10325
rect 544 10309 586 10325
rect 17 10295 67 10297
rect 119 10295 169 10297
rect 599 10295 649 10297
rect 42 10253 59 10287
rect 67 10245 69 10295
rect 160 10287 246 10295
rect 522 10287 608 10295
rect 76 10253 110 10287
rect 127 10253 144 10287
rect 152 10253 161 10287
rect 162 10285 195 10287
rect 224 10285 244 10287
rect 162 10253 244 10285
rect 524 10285 548 10287
rect 573 10285 582 10287
rect 586 10285 606 10287
rect 160 10245 246 10253
rect 186 10229 220 10231
rect 182 10215 224 10216
rect 160 10209 182 10215
rect 224 10209 246 10215
rect 186 10174 220 10208
rect 223 10174 257 10208
rect 120 10161 170 10163
rect 76 10157 130 10161
rect 110 10152 130 10157
rect 60 10127 67 10137
rect 76 10127 77 10147
rect 96 10118 99 10152
rect 109 10127 110 10147
rect 119 10127 126 10137
rect 76 10111 92 10117
rect 94 10111 110 10117
rect 170 10111 172 10161
rect 186 10095 190 10129
rect 216 10095 220 10129
rect 288 10095 292 10283
rect 476 10215 480 10283
rect 524 10253 606 10285
rect 607 10253 616 10287
rect 522 10245 608 10253
rect 649 10245 651 10295
rect 548 10229 582 10231
rect 522 10210 548 10215
rect 522 10209 582 10210
rect 586 10209 608 10215
rect 295 10174 300 10208
rect 324 10174 329 10208
rect 544 10206 582 10209
rect 378 10169 450 10177
rect 428 10139 430 10155
rect 400 10131 430 10139
rect 476 10137 480 10205
rect 544 10176 552 10206
rect 578 10176 582 10206
rect 544 10167 548 10176
rect 400 10127 434 10131
rect 400 10097 408 10127
rect 420 10097 434 10127
rect 544 10129 548 10137
rect 12 10058 62 10060
rect 28 10049 59 10051
rect 62 10049 64 10058
rect 28 10041 64 10049
rect 127 10049 158 10051
rect 127 10042 182 10049
rect 215 10047 224 10075
rect 127 10041 161 10042
rect 59 10025 64 10041
rect 158 10025 161 10041
rect 28 10017 64 10025
rect 127 10024 161 10025
rect 127 10017 182 10024
rect 62 10008 64 10017
rect 213 10009 224 10047
rect 282 10037 292 10095
rect 296 10089 368 10097
rect 319 10060 335 10062
rect 251 10003 263 10037
rect 273 10003 292 10037
rect 303 10030 316 10046
rect 303 10012 316 10028
rect 120 9955 170 9957
rect 76 9949 92 9955
rect 94 9949 110 9955
rect 76 9939 99 9948
rect 60 9929 67 9939
rect 76 9919 77 9939
rect 96 9914 99 9939
rect 109 9919 110 9939
rect 119 9929 126 9939
rect 76 9905 110 9909
rect 170 9905 172 9955
rect 186 9937 190 9971
rect 216 9937 220 9971
rect 186 9860 220 9894
rect 282 9891 292 10003
rect 318 10006 324 10059
rect 346 10046 348 10059
rect 428 10050 430 10097
rect 443 10087 450 10089
rect 476 10057 480 10125
rect 544 10095 552 10129
rect 578 10095 582 10129
rect 481 10063 517 10091
rect 481 10057 495 10063
rect 333 10012 353 10046
rect 367 10016 380 10050
rect 396 10016 408 10050
rect 420 10016 434 10050
rect 318 9996 335 10006
rect 318 9927 324 9996
rect 346 9927 348 10012
rect 428 9969 430 10016
rect 476 9979 480 10047
rect 485 10029 495 10057
rect 505 10029 519 10063
rect 544 10057 555 10095
rect 544 10029 553 10057
rect 544 10009 548 10029
rect 579 9988 582 10078
rect 599 10058 649 10060
rect 610 10050 624 10051
rect 607 10049 624 10050
rect 586 10042 644 10049
rect 607 10041 644 10042
rect 607 10025 610 10041
rect 616 10025 644 10041
rect 607 10024 644 10025
rect 586 10017 644 10024
rect 607 10016 610 10017
rect 649 10008 651 10058
rect 544 9971 548 9979
rect 400 9939 408 9969
rect 420 9939 434 9969
rect 400 9935 434 9939
rect 400 9927 430 9935
rect 428 9911 430 9927
rect 476 9899 480 9967
rect 544 9937 552 9971
rect 578 9937 582 9971
rect 544 9929 548 9937
rect 544 9899 586 9900
rect 288 9859 292 9891
rect 296 9889 368 9897
rect 378 9889 450 9897
rect 544 9892 548 9899
rect 439 9861 444 9889
rect 120 9845 170 9847
rect 76 9841 130 9845
rect 110 9836 130 9841
rect 60 9811 67 9821
rect 76 9811 77 9831
rect 96 9802 99 9836
rect 109 9811 110 9831
rect 119 9811 126 9821
rect 76 9795 92 9801
rect 94 9795 110 9801
rect 170 9795 172 9845
rect 186 9779 190 9813
rect 216 9779 220 9813
rect 213 9747 224 9779
rect 282 9775 292 9859
rect 296 9853 368 9861
rect 378 9853 450 9861
rect 468 9858 473 9892
rect 428 9823 430 9839
rect 251 9747 292 9775
rect 12 9742 62 9744
rect 28 9733 59 9735
rect 62 9733 64 9742
rect 251 9741 263 9747
rect 28 9725 64 9733
rect 127 9733 158 9735
rect 127 9726 182 9733
rect 127 9725 161 9726
rect 59 9709 64 9725
rect 158 9709 161 9725
rect 253 9713 263 9741
rect 273 9713 292 9747
rect 318 9754 324 9823
rect 318 9744 335 9754
rect 303 9722 316 9738
rect 28 9701 64 9709
rect 127 9708 161 9709
rect 127 9701 182 9708
rect 62 9692 64 9701
rect 282 9655 292 9713
rect 303 9704 316 9720
rect 318 9691 324 9744
rect 346 9738 348 9823
rect 400 9815 430 9823
rect 476 9821 480 9889
rect 511 9858 582 9892
rect 544 9851 548 9858
rect 400 9811 434 9815
rect 400 9781 408 9811
rect 420 9781 434 9811
rect 544 9813 548 9821
rect 333 9704 353 9738
rect 428 9734 430 9781
rect 476 9741 480 9809
rect 544 9779 552 9813
rect 578 9779 582 9813
rect 544 9771 548 9779
rect 346 9691 348 9704
rect 367 9700 380 9734
rect 396 9700 408 9734
rect 420 9700 434 9734
rect 544 9731 553 9759
rect 319 9688 335 9690
rect 120 9639 170 9641
rect 76 9633 92 9639
rect 94 9633 110 9639
rect 76 9623 99 9632
rect 60 9613 67 9623
rect 76 9603 77 9623
rect 96 9598 99 9623
rect 109 9603 110 9623
rect 119 9613 126 9623
rect 76 9589 110 9593
rect 170 9589 172 9639
rect 186 9621 190 9655
rect 216 9621 220 9655
rect 182 9583 224 9584
rect 186 9542 220 9576
rect 223 9542 257 9576
rect 160 9535 182 9541
rect 224 9535 246 9541
rect 288 9535 292 9655
rect 296 9653 368 9661
rect 428 9653 430 9700
rect 476 9663 480 9731
rect 485 9687 495 9721
rect 505 9687 519 9721
rect 544 9687 555 9731
rect 485 9663 492 9687
rect 579 9672 582 9762
rect 599 9742 649 9744
rect 610 9734 624 9735
rect 607 9733 624 9734
rect 586 9726 644 9733
rect 607 9725 644 9726
rect 607 9709 610 9725
rect 616 9709 644 9725
rect 607 9708 644 9709
rect 586 9701 644 9708
rect 607 9700 610 9701
rect 649 9692 651 9742
rect 544 9655 548 9663
rect 400 9623 408 9653
rect 420 9623 434 9653
rect 400 9619 434 9623
rect 400 9611 430 9619
rect 428 9595 430 9611
rect 476 9583 480 9651
rect 544 9621 552 9655
rect 578 9621 582 9655
rect 544 9613 548 9621
rect 295 9542 300 9576
rect 324 9542 329 9576
rect 378 9573 450 9581
rect 544 9578 548 9583
rect 544 9574 582 9578
rect 544 9544 552 9574
rect 578 9544 582 9574
rect 544 9541 548 9544
rect 522 9535 548 9541
rect 586 9535 608 9541
rect 182 9519 224 9535
rect 544 9519 586 9535
rect 17 9505 67 9507
rect 119 9505 169 9507
rect 599 9505 649 9507
rect 42 9463 59 9497
rect 67 9455 69 9505
rect 160 9497 246 9505
rect 522 9497 608 9505
rect 76 9463 110 9497
rect 127 9463 144 9497
rect 152 9463 161 9497
rect 162 9495 195 9497
rect 224 9495 244 9497
rect 162 9463 244 9495
rect 524 9495 548 9497
rect 573 9495 582 9497
rect 586 9495 606 9497
rect 160 9455 246 9463
rect 186 9439 220 9441
rect 182 9425 224 9426
rect 160 9419 182 9425
rect 224 9419 246 9425
rect 186 9384 220 9418
rect 223 9384 257 9418
rect 120 9371 170 9373
rect 76 9367 130 9371
rect 110 9362 130 9367
rect 60 9337 67 9347
rect 76 9337 77 9357
rect 96 9328 99 9362
rect 109 9337 110 9357
rect 119 9337 126 9347
rect 76 9321 92 9327
rect 94 9321 110 9327
rect 170 9321 172 9371
rect 186 9305 190 9339
rect 216 9305 220 9339
rect 288 9305 292 9493
rect 476 9425 480 9493
rect 524 9463 606 9495
rect 607 9463 616 9497
rect 522 9455 608 9463
rect 649 9455 651 9505
rect 548 9439 582 9441
rect 522 9420 548 9425
rect 522 9419 582 9420
rect 586 9419 608 9425
rect 295 9384 300 9418
rect 324 9384 329 9418
rect 544 9416 582 9419
rect 378 9379 450 9387
rect 428 9349 430 9365
rect 400 9341 430 9349
rect 476 9347 480 9415
rect 544 9386 552 9416
rect 578 9386 582 9416
rect 544 9377 548 9386
rect 400 9337 434 9341
rect 400 9307 408 9337
rect 420 9307 434 9337
rect 544 9339 548 9347
rect 12 9268 62 9270
rect 28 9259 59 9261
rect 62 9259 64 9268
rect 28 9251 64 9259
rect 127 9259 158 9261
rect 127 9252 182 9259
rect 215 9257 224 9285
rect 127 9251 161 9252
rect 59 9235 64 9251
rect 158 9235 161 9251
rect 28 9227 64 9235
rect 127 9234 161 9235
rect 127 9227 182 9234
rect 62 9218 64 9227
rect 213 9219 224 9257
rect 282 9247 292 9305
rect 296 9299 368 9307
rect 319 9270 335 9272
rect 251 9213 263 9247
rect 273 9213 292 9247
rect 303 9240 316 9256
rect 303 9222 316 9238
rect 120 9165 170 9167
rect 76 9159 92 9165
rect 94 9159 110 9165
rect 76 9149 99 9158
rect 60 9139 67 9149
rect 76 9129 77 9149
rect 96 9124 99 9149
rect 109 9129 110 9149
rect 119 9139 126 9149
rect 76 9115 110 9119
rect 170 9115 172 9165
rect 186 9147 190 9181
rect 216 9147 220 9181
rect 186 9070 220 9104
rect 282 9101 292 9213
rect 318 9216 324 9269
rect 346 9256 348 9269
rect 428 9260 430 9307
rect 443 9297 450 9299
rect 476 9267 480 9335
rect 544 9305 552 9339
rect 578 9305 582 9339
rect 481 9273 517 9301
rect 481 9267 495 9273
rect 333 9222 353 9256
rect 367 9226 380 9260
rect 396 9226 408 9260
rect 420 9226 434 9260
rect 318 9206 335 9216
rect 318 9137 324 9206
rect 346 9137 348 9222
rect 428 9179 430 9226
rect 476 9189 480 9257
rect 485 9239 495 9267
rect 505 9239 519 9273
rect 544 9267 555 9305
rect 544 9239 553 9267
rect 544 9219 548 9239
rect 579 9198 582 9288
rect 599 9268 649 9270
rect 610 9260 624 9261
rect 607 9259 624 9260
rect 586 9252 644 9259
rect 607 9251 644 9252
rect 607 9235 610 9251
rect 616 9235 644 9251
rect 607 9234 644 9235
rect 586 9227 644 9234
rect 607 9226 610 9227
rect 649 9218 651 9268
rect 544 9181 548 9189
rect 400 9149 408 9179
rect 420 9149 434 9179
rect 400 9145 434 9149
rect 400 9137 430 9145
rect 428 9121 430 9137
rect 476 9109 480 9177
rect 544 9147 552 9181
rect 578 9147 582 9181
rect 544 9139 548 9147
rect 544 9109 586 9110
rect 288 9069 292 9101
rect 296 9099 368 9107
rect 378 9099 450 9107
rect 544 9102 548 9109
rect 439 9071 444 9099
rect 120 9055 170 9057
rect 76 9051 130 9055
rect 110 9046 130 9051
rect 60 9021 67 9031
rect 76 9021 77 9041
rect 96 9012 99 9046
rect 109 9021 110 9041
rect 119 9021 126 9031
rect 76 9005 92 9011
rect 94 9005 110 9011
rect 170 9005 172 9055
rect 186 8989 190 9023
rect 216 8989 220 9023
rect 213 8957 224 8989
rect 282 8985 292 9069
rect 296 9063 368 9071
rect 378 9063 450 9071
rect 468 9068 473 9102
rect 428 9033 430 9049
rect 251 8957 292 8985
rect 12 8952 62 8954
rect 28 8943 59 8945
rect 62 8943 64 8952
rect 251 8951 263 8957
rect 28 8935 64 8943
rect 127 8943 158 8945
rect 127 8936 182 8943
rect 127 8935 161 8936
rect 59 8919 64 8935
rect 158 8919 161 8935
rect 253 8923 263 8951
rect 273 8923 292 8957
rect 318 8964 324 9033
rect 318 8954 335 8964
rect 303 8932 316 8948
rect 28 8911 64 8919
rect 127 8918 161 8919
rect 127 8911 182 8918
rect 62 8902 64 8911
rect 282 8865 292 8923
rect 303 8914 316 8930
rect 318 8901 324 8954
rect 346 8948 348 9033
rect 400 9025 430 9033
rect 476 9031 480 9099
rect 511 9068 582 9102
rect 544 9061 548 9068
rect 400 9021 434 9025
rect 400 8991 408 9021
rect 420 8991 434 9021
rect 544 9023 548 9031
rect 333 8914 353 8948
rect 428 8944 430 8991
rect 476 8951 480 9019
rect 544 8989 552 9023
rect 578 8989 582 9023
rect 544 8981 548 8989
rect 346 8901 348 8914
rect 367 8910 380 8944
rect 396 8910 408 8944
rect 420 8910 434 8944
rect 544 8941 553 8969
rect 319 8898 335 8900
rect 120 8849 170 8851
rect 76 8843 92 8849
rect 94 8843 110 8849
rect 76 8833 99 8842
rect 60 8823 67 8833
rect 76 8813 77 8833
rect 96 8808 99 8833
rect 109 8813 110 8833
rect 119 8823 126 8833
rect 76 8799 110 8803
rect 170 8799 172 8849
rect 186 8831 190 8865
rect 216 8831 220 8865
rect 182 8793 224 8794
rect 186 8752 220 8786
rect 223 8752 257 8786
rect 160 8745 182 8751
rect 224 8745 246 8751
rect 288 8745 292 8865
rect 296 8863 368 8871
rect 428 8863 430 8910
rect 476 8873 480 8941
rect 485 8897 495 8931
rect 505 8897 519 8931
rect 544 8897 555 8941
rect 485 8873 492 8897
rect 579 8882 582 8972
rect 599 8952 649 8954
rect 610 8944 624 8945
rect 607 8943 624 8944
rect 586 8936 644 8943
rect 607 8935 644 8936
rect 607 8919 610 8935
rect 616 8919 644 8935
rect 607 8918 644 8919
rect 586 8911 644 8918
rect 607 8910 610 8911
rect 649 8902 651 8952
rect 544 8865 548 8873
rect 400 8833 408 8863
rect 420 8833 434 8863
rect 400 8829 434 8833
rect 400 8821 430 8829
rect 428 8805 430 8821
rect 476 8793 480 8861
rect 544 8831 552 8865
rect 578 8831 582 8865
rect 544 8823 548 8831
rect 295 8752 300 8786
rect 324 8752 329 8786
rect 378 8783 450 8791
rect 544 8788 548 8793
rect 544 8784 582 8788
rect 544 8754 552 8784
rect 578 8754 582 8784
rect 544 8751 548 8754
rect 522 8745 548 8751
rect 586 8745 608 8751
rect 182 8729 224 8745
rect 544 8729 586 8745
rect 17 8715 67 8717
rect 119 8715 169 8717
rect 599 8715 649 8717
rect 42 8673 59 8707
rect 67 8665 69 8715
rect 160 8707 246 8715
rect 522 8707 608 8715
rect 76 8673 110 8707
rect 127 8673 144 8707
rect 152 8673 161 8707
rect 162 8705 195 8707
rect 224 8705 244 8707
rect 162 8673 244 8705
rect 524 8705 548 8707
rect 573 8705 582 8707
rect 586 8705 606 8707
rect 160 8665 246 8673
rect 186 8649 220 8651
rect 182 8635 224 8636
rect 160 8629 182 8635
rect 224 8629 246 8635
rect 186 8594 220 8628
rect 223 8594 257 8628
rect 120 8581 170 8583
rect 76 8577 130 8581
rect 110 8572 130 8577
rect 60 8547 67 8557
rect 76 8547 77 8567
rect 96 8538 99 8572
rect 109 8547 110 8567
rect 119 8547 126 8557
rect 76 8531 92 8537
rect 94 8531 110 8537
rect 170 8531 172 8581
rect 186 8515 190 8549
rect 216 8515 220 8549
rect 288 8515 292 8703
rect 476 8635 480 8703
rect 524 8673 606 8705
rect 607 8673 616 8707
rect 522 8665 608 8673
rect 649 8665 651 8715
rect 548 8649 582 8651
rect 522 8630 548 8635
rect 522 8629 582 8630
rect 586 8629 608 8635
rect 295 8594 300 8628
rect 324 8594 329 8628
rect 544 8626 582 8629
rect 378 8589 450 8597
rect 428 8559 430 8575
rect 400 8551 430 8559
rect 476 8557 480 8625
rect 544 8596 552 8626
rect 578 8596 582 8626
rect 544 8587 548 8596
rect 400 8547 434 8551
rect 400 8517 408 8547
rect 420 8517 434 8547
rect 544 8549 548 8557
rect 12 8478 62 8480
rect 28 8469 59 8471
rect 62 8469 64 8478
rect 28 8461 64 8469
rect 127 8469 158 8471
rect 127 8462 182 8469
rect 215 8467 224 8495
rect 127 8461 161 8462
rect 59 8445 64 8461
rect 158 8445 161 8461
rect 28 8437 64 8445
rect 127 8444 161 8445
rect 127 8437 182 8444
rect 62 8428 64 8437
rect 213 8429 224 8467
rect 282 8457 292 8515
rect 296 8509 368 8517
rect 319 8480 335 8482
rect 251 8423 263 8457
rect 273 8423 292 8457
rect 303 8450 316 8466
rect 303 8432 316 8448
rect 120 8375 170 8377
rect 76 8369 92 8375
rect 94 8369 110 8375
rect 76 8359 99 8368
rect 60 8349 67 8359
rect 76 8339 77 8359
rect 96 8334 99 8359
rect 109 8339 110 8359
rect 119 8349 126 8359
rect 76 8325 110 8329
rect 170 8325 172 8375
rect 186 8357 190 8391
rect 216 8357 220 8391
rect 186 8280 220 8314
rect 282 8311 292 8423
rect 318 8426 324 8479
rect 346 8466 348 8479
rect 428 8470 430 8517
rect 443 8507 450 8509
rect 476 8477 480 8545
rect 544 8515 552 8549
rect 578 8515 582 8549
rect 481 8483 517 8511
rect 481 8477 495 8483
rect 333 8432 353 8466
rect 367 8436 380 8470
rect 396 8436 408 8470
rect 420 8436 434 8470
rect 318 8416 335 8426
rect 318 8347 324 8416
rect 346 8347 348 8432
rect 428 8389 430 8436
rect 476 8399 480 8467
rect 485 8449 495 8477
rect 505 8449 519 8483
rect 544 8477 555 8515
rect 544 8449 553 8477
rect 544 8429 548 8449
rect 579 8408 582 8498
rect 599 8478 649 8480
rect 610 8470 624 8471
rect 607 8469 624 8470
rect 586 8462 644 8469
rect 607 8461 644 8462
rect 607 8445 610 8461
rect 616 8445 644 8461
rect 607 8444 644 8445
rect 586 8437 644 8444
rect 607 8436 610 8437
rect 649 8428 651 8478
rect 544 8391 548 8399
rect 400 8359 408 8389
rect 420 8359 434 8389
rect 400 8355 434 8359
rect 400 8347 430 8355
rect 428 8331 430 8347
rect 476 8319 480 8387
rect 544 8357 552 8391
rect 578 8357 582 8391
rect 544 8349 548 8357
rect 544 8319 586 8320
rect 288 8279 292 8311
rect 296 8309 368 8317
rect 378 8309 450 8317
rect 544 8312 548 8319
rect 439 8281 444 8309
rect 120 8265 170 8267
rect 76 8261 130 8265
rect 110 8256 130 8261
rect 60 8231 67 8241
rect 76 8231 77 8251
rect 96 8222 99 8256
rect 109 8231 110 8251
rect 119 8231 126 8241
rect 76 8215 92 8221
rect 94 8215 110 8221
rect 170 8215 172 8265
rect 186 8199 190 8233
rect 216 8199 220 8233
rect 213 8167 224 8199
rect 282 8195 292 8279
rect 296 8273 368 8281
rect 378 8273 450 8281
rect 468 8278 473 8312
rect 428 8243 430 8259
rect 251 8167 292 8195
rect 12 8162 62 8164
rect 28 8153 59 8155
rect 62 8153 64 8162
rect 251 8161 263 8167
rect 28 8145 64 8153
rect 127 8153 158 8155
rect 127 8146 182 8153
rect 127 8145 161 8146
rect 59 8129 64 8145
rect 158 8129 161 8145
rect 253 8133 263 8161
rect 273 8133 292 8167
rect 318 8174 324 8243
rect 318 8164 335 8174
rect 303 8142 316 8158
rect 28 8121 64 8129
rect 127 8128 161 8129
rect 127 8121 182 8128
rect 62 8112 64 8121
rect 282 8075 292 8133
rect 303 8124 316 8140
rect 318 8111 324 8164
rect 346 8158 348 8243
rect 400 8235 430 8243
rect 476 8241 480 8309
rect 511 8278 582 8312
rect 544 8271 548 8278
rect 400 8231 434 8235
rect 400 8201 408 8231
rect 420 8201 434 8231
rect 544 8233 548 8241
rect 333 8124 353 8158
rect 428 8154 430 8201
rect 476 8161 480 8229
rect 544 8199 552 8233
rect 578 8199 582 8233
rect 544 8191 548 8199
rect 346 8111 348 8124
rect 367 8120 380 8154
rect 396 8120 408 8154
rect 420 8120 434 8154
rect 544 8151 553 8179
rect 319 8108 335 8110
rect 120 8059 170 8061
rect 76 8053 92 8059
rect 94 8053 110 8059
rect 76 8043 99 8052
rect 60 8033 67 8043
rect 76 8023 77 8043
rect 96 8018 99 8043
rect 109 8023 110 8043
rect 119 8033 126 8043
rect 76 8009 110 8013
rect 170 8009 172 8059
rect 186 8041 190 8075
rect 216 8041 220 8075
rect 182 8003 224 8004
rect 186 7962 220 7996
rect 223 7962 257 7996
rect 160 7955 182 7961
rect 224 7955 246 7961
rect 288 7955 292 8075
rect 296 8073 368 8081
rect 428 8073 430 8120
rect 476 8083 480 8151
rect 485 8107 495 8141
rect 505 8107 519 8141
rect 544 8107 555 8151
rect 485 8083 492 8107
rect 579 8092 582 8182
rect 599 8162 649 8164
rect 610 8154 624 8155
rect 607 8153 624 8154
rect 586 8146 644 8153
rect 607 8145 644 8146
rect 607 8129 610 8145
rect 616 8129 644 8145
rect 607 8128 644 8129
rect 586 8121 644 8128
rect 607 8120 610 8121
rect 649 8112 651 8162
rect 544 8075 548 8083
rect 400 8043 408 8073
rect 420 8043 434 8073
rect 400 8039 434 8043
rect 400 8031 430 8039
rect 428 8015 430 8031
rect 476 8003 480 8071
rect 544 8041 552 8075
rect 578 8041 582 8075
rect 544 8033 548 8041
rect 295 7962 300 7996
rect 324 7962 329 7996
rect 378 7993 450 8001
rect 544 7998 548 8003
rect 544 7994 582 7998
rect 544 7964 552 7994
rect 578 7964 582 7994
rect 544 7961 548 7964
rect 522 7955 548 7961
rect 586 7955 608 7961
rect 182 7939 224 7955
rect 544 7939 586 7955
rect 17 7925 67 7927
rect 119 7925 169 7927
rect 599 7925 649 7927
rect 42 7883 59 7917
rect 67 7875 69 7925
rect 160 7917 246 7925
rect 522 7917 608 7925
rect 76 7883 110 7917
rect 127 7883 144 7917
rect 152 7883 161 7917
rect 162 7915 195 7917
rect 224 7915 244 7917
rect 162 7883 244 7915
rect 524 7915 548 7917
rect 573 7915 582 7917
rect 586 7915 606 7917
rect 160 7875 246 7883
rect 186 7859 220 7861
rect 182 7845 224 7846
rect 160 7839 182 7845
rect 224 7839 246 7845
rect 186 7804 220 7838
rect 223 7804 257 7838
rect 120 7791 170 7793
rect 76 7787 130 7791
rect 110 7782 130 7787
rect 60 7757 67 7767
rect 76 7757 77 7777
rect 96 7748 99 7782
rect 109 7757 110 7777
rect 119 7757 126 7767
rect 76 7741 92 7747
rect 94 7741 110 7747
rect 170 7741 172 7791
rect 186 7725 190 7759
rect 216 7725 220 7759
rect 288 7725 292 7913
rect 476 7845 480 7913
rect 524 7883 606 7915
rect 607 7883 616 7917
rect 522 7875 608 7883
rect 649 7875 651 7925
rect 548 7859 582 7861
rect 522 7840 548 7845
rect 522 7839 582 7840
rect 586 7839 608 7845
rect 295 7804 300 7838
rect 324 7804 329 7838
rect 544 7836 582 7839
rect 378 7799 450 7807
rect 428 7769 430 7785
rect 400 7761 430 7769
rect 476 7767 480 7835
rect 544 7806 552 7836
rect 578 7806 582 7836
rect 544 7797 548 7806
rect 400 7757 434 7761
rect 400 7727 408 7757
rect 420 7727 434 7757
rect 544 7759 548 7767
rect 12 7688 62 7690
rect 28 7679 59 7681
rect 62 7679 64 7688
rect 28 7671 64 7679
rect 127 7679 158 7681
rect 127 7672 182 7679
rect 215 7677 224 7705
rect 127 7671 161 7672
rect 59 7655 64 7671
rect 158 7655 161 7671
rect 28 7647 64 7655
rect 127 7654 161 7655
rect 127 7647 182 7654
rect 62 7638 64 7647
rect 213 7639 224 7677
rect 282 7667 292 7725
rect 296 7719 368 7727
rect 319 7690 335 7692
rect 251 7633 263 7667
rect 273 7633 292 7667
rect 303 7660 316 7676
rect 303 7642 316 7658
rect 120 7585 170 7587
rect 76 7579 92 7585
rect 94 7579 110 7585
rect 76 7569 99 7578
rect 60 7559 67 7569
rect 76 7549 77 7569
rect 96 7544 99 7569
rect 109 7549 110 7569
rect 119 7559 126 7569
rect 76 7535 110 7539
rect 170 7535 172 7585
rect 186 7567 190 7601
rect 216 7567 220 7601
rect 186 7490 220 7524
rect 282 7521 292 7633
rect 318 7636 324 7689
rect 346 7676 348 7689
rect 428 7680 430 7727
rect 443 7717 450 7719
rect 476 7687 480 7755
rect 544 7725 552 7759
rect 578 7725 582 7759
rect 481 7693 517 7721
rect 481 7687 495 7693
rect 333 7642 353 7676
rect 367 7646 380 7680
rect 396 7646 408 7680
rect 420 7646 434 7680
rect 318 7626 335 7636
rect 318 7557 324 7626
rect 346 7557 348 7642
rect 428 7599 430 7646
rect 476 7609 480 7677
rect 485 7659 495 7687
rect 505 7659 519 7693
rect 544 7687 555 7725
rect 544 7659 553 7687
rect 544 7639 548 7659
rect 579 7618 582 7708
rect 599 7688 649 7690
rect 610 7680 624 7681
rect 607 7679 624 7680
rect 586 7672 644 7679
rect 607 7671 644 7672
rect 607 7655 610 7671
rect 616 7655 644 7671
rect 607 7654 644 7655
rect 586 7647 644 7654
rect 607 7646 610 7647
rect 649 7638 651 7688
rect 544 7601 548 7609
rect 400 7569 408 7599
rect 420 7569 434 7599
rect 400 7565 434 7569
rect 400 7557 430 7565
rect 428 7541 430 7557
rect 476 7529 480 7597
rect 544 7567 552 7601
rect 578 7567 582 7601
rect 544 7559 548 7567
rect 544 7529 586 7530
rect 288 7489 292 7521
rect 296 7519 368 7527
rect 378 7519 450 7527
rect 544 7522 548 7529
rect 439 7491 444 7519
rect 120 7475 170 7477
rect 76 7471 130 7475
rect 110 7466 130 7471
rect 60 7441 67 7451
rect 76 7441 77 7461
rect 96 7432 99 7466
rect 109 7441 110 7461
rect 119 7441 126 7451
rect 76 7425 92 7431
rect 94 7425 110 7431
rect 170 7425 172 7475
rect 186 7409 190 7443
rect 216 7409 220 7443
rect 213 7377 224 7409
rect 282 7405 292 7489
rect 296 7483 368 7491
rect 378 7483 450 7491
rect 468 7488 473 7522
rect 428 7453 430 7469
rect 251 7377 292 7405
rect 12 7372 62 7374
rect 28 7363 59 7365
rect 62 7363 64 7372
rect 251 7371 263 7377
rect 28 7355 64 7363
rect 127 7363 158 7365
rect 127 7356 182 7363
rect 127 7355 161 7356
rect 59 7339 64 7355
rect 158 7339 161 7355
rect 253 7343 263 7371
rect 273 7343 292 7377
rect 318 7384 324 7453
rect 318 7374 335 7384
rect 303 7352 316 7368
rect 28 7331 64 7339
rect 127 7338 161 7339
rect 127 7331 182 7338
rect 62 7322 64 7331
rect 282 7285 292 7343
rect 303 7334 316 7350
rect 318 7321 324 7374
rect 346 7368 348 7453
rect 400 7445 430 7453
rect 476 7451 480 7519
rect 511 7488 582 7522
rect 544 7481 548 7488
rect 400 7441 434 7445
rect 400 7411 408 7441
rect 420 7411 434 7441
rect 544 7443 548 7451
rect 333 7334 353 7368
rect 428 7364 430 7411
rect 476 7371 480 7439
rect 544 7409 552 7443
rect 578 7409 582 7443
rect 544 7401 548 7409
rect 346 7321 348 7334
rect 367 7330 380 7364
rect 396 7330 408 7364
rect 420 7330 434 7364
rect 544 7361 553 7389
rect 319 7318 335 7320
rect 120 7269 170 7271
rect 76 7263 92 7269
rect 94 7263 110 7269
rect 76 7253 99 7262
rect 60 7243 67 7253
rect 76 7233 77 7253
rect 96 7228 99 7253
rect 109 7233 110 7253
rect 119 7243 126 7253
rect 76 7219 110 7223
rect 170 7219 172 7269
rect 186 7251 190 7285
rect 216 7251 220 7285
rect 182 7213 224 7214
rect 186 7172 220 7206
rect 223 7172 257 7206
rect 160 7165 182 7171
rect 224 7165 246 7171
rect 288 7165 292 7285
rect 296 7283 368 7291
rect 428 7283 430 7330
rect 476 7293 480 7361
rect 485 7317 495 7351
rect 505 7317 519 7351
rect 544 7317 555 7361
rect 485 7293 492 7317
rect 579 7302 582 7392
rect 599 7372 649 7374
rect 610 7364 624 7365
rect 607 7363 624 7364
rect 586 7356 644 7363
rect 607 7355 644 7356
rect 607 7339 610 7355
rect 616 7339 644 7355
rect 607 7338 644 7339
rect 586 7331 644 7338
rect 607 7330 610 7331
rect 649 7322 651 7372
rect 544 7285 548 7293
rect 400 7253 408 7283
rect 420 7253 434 7283
rect 400 7249 434 7253
rect 400 7241 430 7249
rect 428 7225 430 7241
rect 476 7213 480 7281
rect 544 7251 552 7285
rect 578 7251 582 7285
rect 544 7243 548 7251
rect 295 7172 300 7206
rect 324 7172 329 7206
rect 378 7203 450 7211
rect 544 7208 548 7213
rect 544 7204 582 7208
rect 544 7174 552 7204
rect 578 7174 582 7204
rect 544 7171 548 7174
rect 522 7165 548 7171
rect 586 7165 608 7171
rect 182 7149 224 7165
rect 544 7149 586 7165
rect 17 7135 67 7137
rect 119 7135 169 7137
rect 599 7135 649 7137
rect 42 7093 59 7127
rect 67 7085 69 7135
rect 160 7127 246 7135
rect 522 7127 608 7135
rect 76 7093 110 7127
rect 127 7093 144 7127
rect 152 7093 161 7127
rect 162 7125 195 7127
rect 224 7125 244 7127
rect 162 7093 244 7125
rect 524 7125 548 7127
rect 573 7125 582 7127
rect 586 7125 606 7127
rect 160 7085 246 7093
rect 186 7069 220 7071
rect 182 7055 224 7056
rect 160 7049 182 7055
rect 224 7049 246 7055
rect 186 7014 220 7048
rect 223 7014 257 7048
rect 120 7001 170 7003
rect 76 6997 130 7001
rect 110 6992 130 6997
rect 60 6967 67 6977
rect 76 6967 77 6987
rect 96 6958 99 6992
rect 109 6967 110 6987
rect 119 6967 126 6977
rect 76 6951 92 6957
rect 94 6951 110 6957
rect 170 6951 172 7001
rect 186 6935 190 6969
rect 216 6935 220 6969
rect 288 6935 292 7123
rect 476 7055 480 7123
rect 524 7093 606 7125
rect 607 7093 616 7127
rect 522 7085 608 7093
rect 649 7085 651 7135
rect 548 7069 582 7071
rect 522 7050 548 7055
rect 522 7049 582 7050
rect 586 7049 608 7055
rect 295 7014 300 7048
rect 324 7014 329 7048
rect 544 7046 582 7049
rect 378 7009 450 7017
rect 428 6979 430 6995
rect 400 6971 430 6979
rect 476 6977 480 7045
rect 544 7016 552 7046
rect 578 7016 582 7046
rect 544 7007 548 7016
rect 400 6967 434 6971
rect 400 6937 408 6967
rect 420 6937 434 6967
rect 544 6969 548 6977
rect 12 6898 62 6900
rect 28 6889 59 6891
rect 62 6889 64 6898
rect 28 6881 64 6889
rect 127 6889 158 6891
rect 127 6882 182 6889
rect 215 6887 224 6915
rect 127 6881 161 6882
rect 59 6865 64 6881
rect 158 6865 161 6881
rect 28 6857 64 6865
rect 127 6864 161 6865
rect 127 6857 182 6864
rect 62 6848 64 6857
rect 213 6849 224 6887
rect 282 6877 292 6935
rect 296 6929 368 6937
rect 319 6900 335 6902
rect 251 6843 263 6877
rect 273 6843 292 6877
rect 303 6870 316 6886
rect 303 6852 316 6868
rect 120 6795 170 6797
rect 76 6789 92 6795
rect 94 6789 110 6795
rect 76 6779 99 6788
rect 60 6769 67 6779
rect 76 6759 77 6779
rect 96 6754 99 6779
rect 109 6759 110 6779
rect 119 6769 126 6779
rect 76 6745 110 6749
rect 170 6745 172 6795
rect 186 6777 190 6811
rect 216 6777 220 6811
rect 186 6700 220 6734
rect 282 6731 292 6843
rect 318 6846 324 6899
rect 346 6886 348 6899
rect 428 6890 430 6937
rect 443 6927 450 6929
rect 476 6897 480 6965
rect 544 6935 552 6969
rect 578 6935 582 6969
rect 481 6903 517 6931
rect 481 6897 495 6903
rect 333 6852 353 6886
rect 367 6856 380 6890
rect 396 6856 408 6890
rect 420 6856 434 6890
rect 318 6836 335 6846
rect 318 6767 324 6836
rect 346 6767 348 6852
rect 428 6809 430 6856
rect 476 6819 480 6887
rect 485 6869 495 6897
rect 505 6869 519 6903
rect 544 6897 555 6935
rect 544 6869 553 6897
rect 544 6849 548 6869
rect 579 6828 582 6918
rect 599 6898 649 6900
rect 610 6890 624 6891
rect 607 6889 624 6890
rect 586 6882 644 6889
rect 607 6881 644 6882
rect 607 6865 610 6881
rect 616 6865 644 6881
rect 607 6864 644 6865
rect 586 6857 644 6864
rect 607 6856 610 6857
rect 649 6848 651 6898
rect 544 6811 548 6819
rect 400 6779 408 6809
rect 420 6779 434 6809
rect 400 6775 434 6779
rect 400 6767 430 6775
rect 428 6751 430 6767
rect 476 6739 480 6807
rect 544 6777 552 6811
rect 578 6777 582 6811
rect 544 6769 548 6777
rect 544 6739 586 6740
rect 288 6699 292 6731
rect 296 6729 368 6737
rect 378 6729 450 6737
rect 544 6732 548 6739
rect 439 6701 444 6729
rect 120 6685 170 6687
rect 76 6681 130 6685
rect 110 6676 130 6681
rect 60 6651 67 6661
rect 76 6651 77 6671
rect 96 6642 99 6676
rect 109 6651 110 6671
rect 119 6651 126 6661
rect 76 6635 92 6641
rect 94 6635 110 6641
rect 170 6635 172 6685
rect 186 6619 190 6653
rect 216 6619 220 6653
rect 213 6587 224 6619
rect 282 6615 292 6699
rect 296 6693 368 6701
rect 378 6693 450 6701
rect 468 6698 473 6732
rect 428 6663 430 6679
rect 251 6587 292 6615
rect 12 6582 62 6584
rect 28 6573 59 6575
rect 62 6573 64 6582
rect 251 6581 263 6587
rect 28 6565 64 6573
rect 127 6573 158 6575
rect 127 6566 182 6573
rect 127 6565 161 6566
rect 59 6549 64 6565
rect 158 6549 161 6565
rect 253 6553 263 6581
rect 273 6553 292 6587
rect 318 6594 324 6663
rect 318 6584 335 6594
rect 303 6562 316 6578
rect 28 6541 64 6549
rect 127 6548 161 6549
rect 127 6541 182 6548
rect 62 6532 64 6541
rect 282 6495 292 6553
rect 303 6544 316 6560
rect 318 6531 324 6584
rect 346 6578 348 6663
rect 400 6655 430 6663
rect 476 6661 480 6729
rect 511 6698 582 6732
rect 544 6691 548 6698
rect 400 6651 434 6655
rect 400 6621 408 6651
rect 420 6621 434 6651
rect 544 6653 548 6661
rect 333 6544 353 6578
rect 428 6574 430 6621
rect 476 6581 480 6649
rect 544 6619 552 6653
rect 578 6619 582 6653
rect 544 6611 548 6619
rect 346 6531 348 6544
rect 367 6540 380 6574
rect 396 6540 408 6574
rect 420 6540 434 6574
rect 544 6571 553 6599
rect 319 6528 335 6530
rect 120 6479 170 6481
rect 76 6473 92 6479
rect 94 6473 110 6479
rect 76 6463 99 6472
rect 60 6453 67 6463
rect 76 6443 77 6463
rect 96 6438 99 6463
rect 109 6443 110 6463
rect 119 6453 126 6463
rect 76 6429 110 6433
rect 170 6429 172 6479
rect 186 6461 190 6495
rect 216 6461 220 6495
rect 182 6423 224 6424
rect 186 6382 220 6416
rect 223 6382 257 6416
rect 160 6375 182 6381
rect 224 6375 246 6381
rect 288 6375 292 6495
rect 296 6493 368 6501
rect 428 6493 430 6540
rect 476 6503 480 6571
rect 485 6527 495 6561
rect 505 6527 519 6561
rect 544 6527 555 6571
rect 485 6503 492 6527
rect 579 6512 582 6602
rect 599 6582 649 6584
rect 610 6574 624 6575
rect 607 6573 624 6574
rect 586 6566 644 6573
rect 607 6565 644 6566
rect 607 6549 610 6565
rect 616 6549 644 6565
rect 607 6548 644 6549
rect 586 6541 644 6548
rect 607 6540 610 6541
rect 649 6532 651 6582
rect 544 6495 548 6503
rect 400 6463 408 6493
rect 420 6463 434 6493
rect 400 6459 434 6463
rect 400 6451 430 6459
rect 428 6435 430 6451
rect 476 6423 480 6491
rect 544 6461 552 6495
rect 578 6461 582 6495
rect 544 6453 548 6461
rect 295 6382 300 6416
rect 324 6382 329 6416
rect 378 6413 450 6421
rect 544 6418 548 6423
rect 544 6414 582 6418
rect 544 6384 552 6414
rect 578 6384 582 6414
rect 544 6381 548 6384
rect 522 6375 548 6381
rect 586 6375 608 6381
rect 182 6359 224 6375
rect 544 6359 586 6375
rect 17 6345 67 6347
rect 119 6345 169 6347
rect 599 6345 649 6347
rect 42 6303 59 6337
rect 67 6295 69 6345
rect 160 6337 246 6345
rect 522 6337 608 6345
rect 76 6303 110 6337
rect 127 6303 144 6337
rect 152 6303 161 6337
rect 162 6335 195 6337
rect 224 6335 244 6337
rect 162 6303 244 6335
rect 524 6335 548 6337
rect 573 6335 582 6337
rect 586 6335 606 6337
rect 160 6295 246 6303
rect 186 6279 220 6281
rect 182 6265 224 6266
rect 160 6259 182 6265
rect 224 6259 246 6265
rect 186 6224 220 6258
rect 223 6224 257 6258
rect 120 6211 170 6213
rect 76 6207 130 6211
rect 110 6202 130 6207
rect 60 6177 67 6187
rect 76 6177 77 6197
rect 96 6168 99 6202
rect 109 6177 110 6197
rect 119 6177 126 6187
rect 76 6161 92 6167
rect 94 6161 110 6167
rect 170 6161 172 6211
rect 186 6145 190 6179
rect 216 6145 220 6179
rect 288 6145 292 6333
rect 476 6265 480 6333
rect 524 6303 606 6335
rect 607 6303 616 6337
rect 522 6295 608 6303
rect 649 6295 651 6345
rect 548 6279 582 6281
rect 522 6260 548 6265
rect 522 6259 582 6260
rect 586 6259 608 6265
rect 295 6224 300 6258
rect 324 6224 329 6258
rect 544 6256 582 6259
rect 378 6219 450 6227
rect 428 6189 430 6205
rect 400 6181 430 6189
rect 476 6187 480 6255
rect 544 6226 552 6256
rect 578 6226 582 6256
rect 544 6217 548 6226
rect 400 6177 434 6181
rect 400 6147 408 6177
rect 420 6147 434 6177
rect 544 6179 548 6187
rect 12 6108 62 6110
rect 28 6099 59 6101
rect 62 6099 64 6108
rect 28 6091 64 6099
rect 127 6099 158 6101
rect 127 6092 182 6099
rect 215 6097 224 6125
rect 127 6091 161 6092
rect 59 6075 64 6091
rect 158 6075 161 6091
rect 28 6067 64 6075
rect 127 6074 161 6075
rect 127 6067 182 6074
rect 62 6058 64 6067
rect 213 6059 224 6097
rect 282 6087 292 6145
rect 296 6139 368 6147
rect 319 6110 335 6112
rect 251 6053 263 6087
rect 273 6053 292 6087
rect 303 6080 316 6096
rect 303 6062 316 6078
rect 120 6005 170 6007
rect 76 5999 92 6005
rect 94 5999 110 6005
rect 76 5989 99 5998
rect 60 5979 67 5989
rect 76 5969 77 5989
rect 96 5964 99 5989
rect 109 5969 110 5989
rect 119 5979 126 5989
rect 76 5955 110 5959
rect 170 5955 172 6005
rect 186 5987 190 6021
rect 216 5987 220 6021
rect 186 5910 220 5944
rect 282 5941 292 6053
rect 318 6056 324 6109
rect 346 6096 348 6109
rect 428 6100 430 6147
rect 443 6137 450 6139
rect 476 6107 480 6175
rect 544 6145 552 6179
rect 578 6145 582 6179
rect 481 6113 517 6141
rect 481 6107 495 6113
rect 333 6062 353 6096
rect 367 6066 380 6100
rect 396 6066 408 6100
rect 420 6066 434 6100
rect 318 6046 335 6056
rect 318 5977 324 6046
rect 346 5977 348 6062
rect 428 6019 430 6066
rect 476 6029 480 6097
rect 485 6079 495 6107
rect 505 6079 519 6113
rect 544 6107 555 6145
rect 544 6079 553 6107
rect 544 6059 548 6079
rect 579 6038 582 6128
rect 599 6108 649 6110
rect 610 6100 624 6101
rect 607 6099 624 6100
rect 586 6092 644 6099
rect 607 6091 644 6092
rect 607 6075 610 6091
rect 616 6075 644 6091
rect 607 6074 644 6075
rect 586 6067 644 6074
rect 607 6066 610 6067
rect 649 6058 651 6108
rect 544 6021 548 6029
rect 400 5989 408 6019
rect 420 5989 434 6019
rect 400 5985 434 5989
rect 400 5977 430 5985
rect 428 5961 430 5977
rect 476 5949 480 6017
rect 544 5987 552 6021
rect 578 5987 582 6021
rect 544 5979 548 5987
rect 544 5949 586 5950
rect 288 5909 292 5941
rect 296 5939 368 5947
rect 378 5939 450 5947
rect 544 5942 548 5949
rect 439 5911 444 5939
rect 120 5895 170 5897
rect 76 5891 130 5895
rect 110 5886 130 5891
rect 60 5861 67 5871
rect 76 5861 77 5881
rect 96 5852 99 5886
rect 109 5861 110 5881
rect 119 5861 126 5871
rect 76 5845 92 5851
rect 94 5845 110 5851
rect 170 5845 172 5895
rect 186 5829 190 5863
rect 216 5829 220 5863
rect 213 5797 224 5829
rect 282 5825 292 5909
rect 296 5903 368 5911
rect 378 5903 450 5911
rect 468 5908 473 5942
rect 428 5873 430 5889
rect 251 5797 292 5825
rect 12 5792 62 5794
rect 28 5783 59 5785
rect 62 5783 64 5792
rect 251 5791 263 5797
rect 28 5775 64 5783
rect 127 5783 158 5785
rect 127 5776 182 5783
rect 127 5775 161 5776
rect 59 5759 64 5775
rect 158 5759 161 5775
rect 253 5763 263 5791
rect 273 5763 292 5797
rect 318 5804 324 5873
rect 318 5794 335 5804
rect 303 5772 316 5788
rect 28 5751 64 5759
rect 127 5758 161 5759
rect 127 5751 182 5758
rect 62 5742 64 5751
rect 282 5705 292 5763
rect 303 5754 316 5770
rect 318 5741 324 5794
rect 346 5788 348 5873
rect 400 5865 430 5873
rect 476 5871 480 5939
rect 511 5908 582 5942
rect 544 5901 548 5908
rect 400 5861 434 5865
rect 400 5831 408 5861
rect 420 5831 434 5861
rect 544 5863 548 5871
rect 333 5754 353 5788
rect 428 5784 430 5831
rect 476 5791 480 5859
rect 544 5829 552 5863
rect 578 5829 582 5863
rect 544 5821 548 5829
rect 346 5741 348 5754
rect 367 5750 380 5784
rect 396 5750 408 5784
rect 420 5750 434 5784
rect 544 5781 553 5809
rect 319 5738 335 5740
rect 120 5689 170 5691
rect 76 5683 92 5689
rect 94 5683 110 5689
rect 76 5673 99 5682
rect 60 5663 67 5673
rect 76 5653 77 5673
rect 96 5648 99 5673
rect 109 5653 110 5673
rect 119 5663 126 5673
rect 76 5639 110 5643
rect 170 5639 172 5689
rect 186 5671 190 5705
rect 216 5671 220 5705
rect 182 5633 224 5634
rect 186 5592 220 5626
rect 223 5592 257 5626
rect 160 5585 182 5591
rect 224 5585 246 5591
rect 288 5585 292 5705
rect 296 5703 368 5711
rect 428 5703 430 5750
rect 476 5713 480 5781
rect 485 5737 495 5771
rect 505 5737 519 5771
rect 544 5737 555 5781
rect 485 5713 492 5737
rect 579 5722 582 5812
rect 599 5792 649 5794
rect 610 5784 624 5785
rect 607 5783 624 5784
rect 586 5776 644 5783
rect 607 5775 644 5776
rect 607 5759 610 5775
rect 616 5759 644 5775
rect 607 5758 644 5759
rect 586 5751 644 5758
rect 607 5750 610 5751
rect 649 5742 651 5792
rect 544 5705 548 5713
rect 400 5673 408 5703
rect 420 5673 434 5703
rect 400 5669 434 5673
rect 400 5661 430 5669
rect 428 5645 430 5661
rect 476 5633 480 5701
rect 544 5671 552 5705
rect 578 5671 582 5705
rect 544 5663 548 5671
rect 295 5592 300 5626
rect 324 5592 329 5626
rect 378 5623 450 5631
rect 544 5628 548 5633
rect 544 5624 582 5628
rect 544 5594 552 5624
rect 578 5594 582 5624
rect 544 5591 548 5594
rect 522 5585 548 5591
rect 586 5585 608 5591
rect 182 5569 224 5585
rect 544 5569 586 5585
rect 17 5555 67 5557
rect 119 5555 169 5557
rect 599 5555 649 5557
rect 42 5513 59 5547
rect 67 5505 69 5555
rect 160 5547 246 5555
rect 522 5547 608 5555
rect 76 5513 110 5547
rect 127 5513 144 5547
rect 152 5513 161 5547
rect 162 5545 195 5547
rect 224 5545 244 5547
rect 162 5513 244 5545
rect 524 5545 548 5547
rect 573 5545 582 5547
rect 586 5545 606 5547
rect 160 5505 246 5513
rect 186 5489 220 5491
rect 182 5475 224 5476
rect 160 5469 182 5475
rect 224 5469 246 5475
rect 186 5434 220 5468
rect 223 5434 257 5468
rect 120 5421 170 5423
rect 76 5417 130 5421
rect 110 5412 130 5417
rect 60 5387 67 5397
rect 76 5387 77 5407
rect 96 5378 99 5412
rect 109 5387 110 5407
rect 119 5387 126 5397
rect 76 5371 92 5377
rect 94 5371 110 5377
rect 170 5371 172 5421
rect 186 5355 190 5389
rect 216 5355 220 5389
rect 288 5355 292 5543
rect 476 5475 480 5543
rect 524 5513 606 5545
rect 607 5513 616 5547
rect 522 5505 608 5513
rect 649 5505 651 5555
rect 548 5489 582 5491
rect 522 5470 548 5475
rect 522 5469 582 5470
rect 586 5469 608 5475
rect 295 5434 300 5468
rect 324 5434 329 5468
rect 544 5466 582 5469
rect 378 5429 450 5437
rect 428 5399 430 5415
rect 400 5391 430 5399
rect 476 5397 480 5465
rect 544 5436 552 5466
rect 578 5436 582 5466
rect 544 5427 548 5436
rect 400 5387 434 5391
rect 400 5357 408 5387
rect 420 5357 434 5387
rect 544 5389 548 5397
rect 12 5318 62 5320
rect 28 5309 59 5311
rect 62 5309 64 5318
rect 28 5301 64 5309
rect 127 5309 158 5311
rect 127 5302 182 5309
rect 215 5307 224 5335
rect 127 5301 161 5302
rect 59 5285 64 5301
rect 158 5285 161 5301
rect 28 5277 64 5285
rect 127 5284 161 5285
rect 127 5277 182 5284
rect 62 5268 64 5277
rect 213 5269 224 5307
rect 282 5297 292 5355
rect 296 5349 368 5357
rect 319 5320 335 5322
rect 251 5263 263 5297
rect 273 5263 292 5297
rect 303 5290 316 5306
rect 303 5272 316 5288
rect 120 5215 170 5217
rect 76 5209 92 5215
rect 94 5209 110 5215
rect 76 5199 99 5208
rect 60 5189 67 5199
rect 76 5179 77 5199
rect 96 5174 99 5199
rect 109 5179 110 5199
rect 119 5189 126 5199
rect 76 5165 110 5169
rect 170 5165 172 5215
rect 186 5197 190 5231
rect 216 5197 220 5231
rect 186 5120 220 5154
rect 282 5151 292 5263
rect 318 5266 324 5319
rect 346 5306 348 5319
rect 428 5310 430 5357
rect 443 5347 450 5349
rect 476 5317 480 5385
rect 544 5355 552 5389
rect 578 5355 582 5389
rect 481 5323 517 5351
rect 481 5317 495 5323
rect 333 5272 353 5306
rect 367 5276 380 5310
rect 396 5276 408 5310
rect 420 5276 434 5310
rect 318 5256 335 5266
rect 318 5187 324 5256
rect 346 5187 348 5272
rect 428 5229 430 5276
rect 476 5239 480 5307
rect 485 5289 495 5317
rect 505 5289 519 5323
rect 544 5317 555 5355
rect 544 5289 553 5317
rect 544 5269 548 5289
rect 579 5248 582 5338
rect 599 5318 649 5320
rect 610 5310 624 5311
rect 607 5309 624 5310
rect 586 5302 644 5309
rect 607 5301 644 5302
rect 607 5285 610 5301
rect 616 5285 644 5301
rect 607 5284 644 5285
rect 586 5277 644 5284
rect 607 5276 610 5277
rect 649 5268 651 5318
rect 544 5231 548 5239
rect 400 5199 408 5229
rect 420 5199 434 5229
rect 400 5195 434 5199
rect 400 5187 430 5195
rect 428 5171 430 5187
rect 476 5159 480 5227
rect 544 5197 552 5231
rect 578 5197 582 5231
rect 544 5189 548 5197
rect 544 5159 586 5160
rect 288 5119 292 5151
rect 296 5149 368 5157
rect 378 5149 450 5157
rect 544 5152 548 5159
rect 439 5121 444 5149
rect 120 5105 170 5107
rect 76 5101 130 5105
rect 110 5096 130 5101
rect 60 5071 67 5081
rect 76 5071 77 5091
rect 96 5062 99 5096
rect 109 5071 110 5091
rect 119 5071 126 5081
rect 76 5055 92 5061
rect 94 5055 110 5061
rect 170 5055 172 5105
rect 186 5039 190 5073
rect 216 5039 220 5073
rect 213 5007 224 5039
rect 282 5035 292 5119
rect 296 5113 368 5121
rect 378 5113 450 5121
rect 468 5118 473 5152
rect 428 5083 430 5099
rect 251 5007 292 5035
rect 12 5002 62 5004
rect 28 4993 59 4995
rect 62 4993 64 5002
rect 251 5001 263 5007
rect 28 4985 64 4993
rect 127 4993 158 4995
rect 127 4986 182 4993
rect 127 4985 161 4986
rect 59 4969 64 4985
rect 158 4969 161 4985
rect 253 4973 263 5001
rect 273 4973 292 5007
rect 318 5014 324 5083
rect 318 5004 335 5014
rect 303 4982 316 4998
rect 28 4961 64 4969
rect 127 4968 161 4969
rect 127 4961 182 4968
rect 62 4952 64 4961
rect 282 4915 292 4973
rect 303 4964 316 4980
rect 318 4951 324 5004
rect 346 4998 348 5083
rect 400 5075 430 5083
rect 476 5081 480 5149
rect 511 5118 582 5152
rect 544 5111 548 5118
rect 400 5071 434 5075
rect 400 5041 408 5071
rect 420 5041 434 5071
rect 544 5073 548 5081
rect 333 4964 353 4998
rect 428 4994 430 5041
rect 476 5001 480 5069
rect 544 5039 552 5073
rect 578 5039 582 5073
rect 544 5031 548 5039
rect 346 4951 348 4964
rect 367 4960 380 4994
rect 396 4960 408 4994
rect 420 4960 434 4994
rect 544 4991 553 5019
rect 319 4948 335 4950
rect 120 4899 170 4901
rect 76 4893 92 4899
rect 94 4893 110 4899
rect 76 4883 99 4892
rect 60 4873 67 4883
rect 76 4863 77 4883
rect 96 4858 99 4883
rect 109 4863 110 4883
rect 119 4873 126 4883
rect 76 4849 110 4853
rect 170 4849 172 4899
rect 186 4881 190 4915
rect 216 4881 220 4915
rect 182 4843 224 4844
rect 186 4802 220 4836
rect 223 4802 257 4836
rect 160 4795 182 4801
rect 224 4795 246 4801
rect 288 4795 292 4915
rect 296 4913 368 4921
rect 428 4913 430 4960
rect 476 4923 480 4991
rect 485 4947 495 4981
rect 505 4947 519 4981
rect 544 4947 555 4991
rect 485 4923 492 4947
rect 579 4932 582 5022
rect 599 5002 649 5004
rect 610 4994 624 4995
rect 607 4993 624 4994
rect 586 4986 644 4993
rect 607 4985 644 4986
rect 607 4969 610 4985
rect 616 4969 644 4985
rect 607 4968 644 4969
rect 586 4961 644 4968
rect 607 4960 610 4961
rect 649 4952 651 5002
rect 544 4915 548 4923
rect 400 4883 408 4913
rect 420 4883 434 4913
rect 400 4879 434 4883
rect 400 4871 430 4879
rect 428 4855 430 4871
rect 476 4843 480 4911
rect 544 4881 552 4915
rect 578 4881 582 4915
rect 544 4873 548 4881
rect 295 4802 300 4836
rect 324 4802 329 4836
rect 378 4833 450 4841
rect 544 4838 548 4843
rect 544 4834 582 4838
rect 544 4804 552 4834
rect 578 4804 582 4834
rect 544 4801 548 4804
rect 522 4795 548 4801
rect 586 4795 608 4801
rect 182 4779 224 4795
rect 544 4779 586 4795
rect 17 4765 67 4767
rect 119 4765 169 4767
rect 599 4765 649 4767
rect 42 4723 59 4757
rect 67 4715 69 4765
rect 160 4757 246 4765
rect 522 4757 608 4765
rect 76 4723 110 4757
rect 127 4723 144 4757
rect 152 4723 161 4757
rect 162 4755 195 4757
rect 224 4755 244 4757
rect 162 4723 244 4755
rect 524 4755 548 4757
rect 573 4755 582 4757
rect 586 4755 606 4757
rect 160 4715 246 4723
rect 186 4699 220 4701
rect 182 4685 224 4686
rect 160 4679 182 4685
rect 224 4679 246 4685
rect 186 4644 220 4678
rect 223 4644 257 4678
rect 120 4631 170 4633
rect 76 4627 130 4631
rect 110 4622 130 4627
rect 60 4597 67 4607
rect 76 4597 77 4617
rect 96 4588 99 4622
rect 109 4597 110 4617
rect 119 4597 126 4607
rect 76 4581 92 4587
rect 94 4581 110 4587
rect 170 4581 172 4631
rect 186 4565 190 4599
rect 216 4565 220 4599
rect 288 4565 292 4753
rect 476 4685 480 4753
rect 524 4723 606 4755
rect 607 4723 616 4757
rect 522 4715 608 4723
rect 649 4715 651 4765
rect 548 4699 582 4701
rect 522 4680 548 4685
rect 522 4679 582 4680
rect 586 4679 608 4685
rect 295 4644 300 4678
rect 324 4644 329 4678
rect 544 4676 582 4679
rect 378 4639 450 4647
rect 428 4609 430 4625
rect 400 4601 430 4609
rect 476 4607 480 4675
rect 544 4646 552 4676
rect 578 4646 582 4676
rect 544 4637 548 4646
rect 400 4597 434 4601
rect 400 4567 408 4597
rect 420 4567 434 4597
rect 544 4599 548 4607
rect 12 4528 62 4530
rect 28 4519 59 4521
rect 62 4519 64 4528
rect 28 4511 64 4519
rect 127 4519 158 4521
rect 127 4512 182 4519
rect 215 4517 224 4545
rect 127 4511 161 4512
rect 59 4495 64 4511
rect 158 4495 161 4511
rect 28 4487 64 4495
rect 127 4494 161 4495
rect 127 4487 182 4494
rect 62 4478 64 4487
rect 213 4479 224 4517
rect 282 4507 292 4565
rect 296 4559 368 4567
rect 319 4530 335 4532
rect 251 4473 263 4507
rect 273 4473 292 4507
rect 303 4500 316 4516
rect 303 4482 316 4498
rect 120 4425 170 4427
rect 76 4419 92 4425
rect 94 4419 110 4425
rect 76 4409 99 4418
rect 60 4399 67 4409
rect 76 4389 77 4409
rect 96 4384 99 4409
rect 109 4389 110 4409
rect 119 4399 126 4409
rect 76 4375 110 4379
rect 170 4375 172 4425
rect 186 4407 190 4441
rect 216 4407 220 4441
rect 186 4330 220 4364
rect 282 4361 292 4473
rect 318 4476 324 4529
rect 346 4516 348 4529
rect 428 4520 430 4567
rect 443 4557 450 4559
rect 476 4527 480 4595
rect 544 4565 552 4599
rect 578 4565 582 4599
rect 481 4533 517 4561
rect 481 4527 495 4533
rect 333 4482 353 4516
rect 367 4486 380 4520
rect 396 4486 408 4520
rect 420 4486 434 4520
rect 318 4466 335 4476
rect 318 4397 324 4466
rect 346 4397 348 4482
rect 428 4439 430 4486
rect 476 4449 480 4517
rect 485 4499 495 4527
rect 505 4499 519 4533
rect 544 4527 555 4565
rect 544 4499 553 4527
rect 544 4479 548 4499
rect 579 4458 582 4548
rect 599 4528 649 4530
rect 610 4520 624 4521
rect 607 4519 624 4520
rect 586 4512 644 4519
rect 607 4511 644 4512
rect 607 4495 610 4511
rect 616 4495 644 4511
rect 607 4494 644 4495
rect 586 4487 644 4494
rect 607 4486 610 4487
rect 649 4478 651 4528
rect 544 4441 548 4449
rect 400 4409 408 4439
rect 420 4409 434 4439
rect 400 4405 434 4409
rect 400 4397 430 4405
rect 428 4381 430 4397
rect 476 4369 480 4437
rect 544 4407 552 4441
rect 578 4407 582 4441
rect 544 4399 548 4407
rect 544 4369 586 4370
rect 288 4329 292 4361
rect 296 4359 368 4367
rect 378 4359 450 4367
rect 544 4362 548 4369
rect 439 4331 444 4359
rect 120 4315 170 4317
rect 76 4311 130 4315
rect 110 4306 130 4311
rect 60 4281 67 4291
rect 76 4281 77 4301
rect 96 4272 99 4306
rect 109 4281 110 4301
rect 119 4281 126 4291
rect 76 4265 92 4271
rect 94 4265 110 4271
rect 170 4265 172 4315
rect 186 4249 190 4283
rect 216 4249 220 4283
rect 213 4217 224 4249
rect 282 4245 292 4329
rect 296 4323 368 4331
rect 378 4323 450 4331
rect 468 4328 473 4362
rect 428 4293 430 4309
rect 251 4217 292 4245
rect 12 4212 62 4214
rect 28 4203 59 4205
rect 62 4203 64 4212
rect 251 4211 263 4217
rect 28 4195 64 4203
rect 127 4203 158 4205
rect 127 4196 182 4203
rect 127 4195 161 4196
rect 59 4179 64 4195
rect 158 4179 161 4195
rect 253 4183 263 4211
rect 273 4183 292 4217
rect 318 4224 324 4293
rect 318 4214 335 4224
rect 303 4192 316 4208
rect 28 4171 64 4179
rect 127 4178 161 4179
rect 127 4171 182 4178
rect 62 4162 64 4171
rect 282 4125 292 4183
rect 303 4174 316 4190
rect 318 4161 324 4214
rect 346 4208 348 4293
rect 400 4285 430 4293
rect 476 4291 480 4359
rect 511 4328 582 4362
rect 544 4321 548 4328
rect 400 4281 434 4285
rect 400 4251 408 4281
rect 420 4251 434 4281
rect 544 4283 548 4291
rect 333 4174 353 4208
rect 428 4204 430 4251
rect 476 4211 480 4279
rect 544 4249 552 4283
rect 578 4249 582 4283
rect 544 4241 548 4249
rect 346 4161 348 4174
rect 367 4170 380 4204
rect 396 4170 408 4204
rect 420 4170 434 4204
rect 544 4201 553 4229
rect 319 4158 335 4160
rect 120 4109 170 4111
rect 76 4103 92 4109
rect 94 4103 110 4109
rect 76 4093 99 4102
rect 60 4083 67 4093
rect 76 4073 77 4093
rect 96 4068 99 4093
rect 109 4073 110 4093
rect 119 4083 126 4093
rect 76 4059 110 4063
rect 170 4059 172 4109
rect 186 4091 190 4125
rect 216 4091 220 4125
rect 182 4053 224 4054
rect 186 4012 220 4046
rect 223 4012 257 4046
rect 160 4005 182 4011
rect 224 4005 246 4011
rect 288 4005 292 4125
rect 296 4123 368 4131
rect 428 4123 430 4170
rect 476 4133 480 4201
rect 485 4157 495 4191
rect 505 4157 519 4191
rect 544 4157 555 4201
rect 485 4133 492 4157
rect 579 4142 582 4232
rect 599 4212 649 4214
rect 610 4204 624 4205
rect 607 4203 624 4204
rect 586 4196 644 4203
rect 607 4195 644 4196
rect 607 4179 610 4195
rect 616 4179 644 4195
rect 607 4178 644 4179
rect 586 4171 644 4178
rect 607 4170 610 4171
rect 649 4162 651 4212
rect 544 4125 548 4133
rect 400 4093 408 4123
rect 420 4093 434 4123
rect 400 4089 434 4093
rect 400 4081 430 4089
rect 428 4065 430 4081
rect 476 4053 480 4121
rect 544 4091 552 4125
rect 578 4091 582 4125
rect 544 4083 548 4091
rect 295 4012 300 4046
rect 324 4012 329 4046
rect 378 4043 450 4051
rect 544 4048 548 4053
rect 544 4044 582 4048
rect 544 4014 552 4044
rect 578 4014 582 4044
rect 544 4011 548 4014
rect 522 4005 548 4011
rect 586 4005 608 4011
rect 182 3989 224 4005
rect 544 3989 586 4005
rect 17 3975 67 3977
rect 119 3975 169 3977
rect 599 3975 649 3977
rect 42 3933 59 3967
rect 67 3925 69 3975
rect 160 3967 246 3975
rect 522 3967 608 3975
rect 76 3933 110 3967
rect 127 3933 144 3967
rect 152 3933 161 3967
rect 162 3965 195 3967
rect 224 3965 244 3967
rect 162 3933 244 3965
rect 524 3965 548 3967
rect 573 3965 582 3967
rect 586 3965 606 3967
rect 160 3925 246 3933
rect 186 3909 220 3911
rect 182 3895 224 3896
rect 160 3889 182 3895
rect 224 3889 246 3895
rect 186 3854 220 3888
rect 223 3854 257 3888
rect 120 3841 170 3843
rect 76 3837 130 3841
rect 110 3832 130 3837
rect 60 3807 67 3817
rect 76 3807 77 3827
rect 96 3798 99 3832
rect 109 3807 110 3827
rect 119 3807 126 3817
rect 76 3791 92 3797
rect 94 3791 110 3797
rect 170 3791 172 3841
rect 186 3775 190 3809
rect 216 3775 220 3809
rect 288 3775 292 3963
rect 476 3895 480 3963
rect 524 3933 606 3965
rect 607 3933 616 3967
rect 522 3925 608 3933
rect 649 3925 651 3975
rect 548 3909 582 3911
rect 522 3890 548 3895
rect 522 3889 582 3890
rect 586 3889 608 3895
rect 295 3854 300 3888
rect 324 3854 329 3888
rect 544 3886 582 3889
rect 378 3849 450 3857
rect 428 3819 430 3835
rect 400 3811 430 3819
rect 476 3817 480 3885
rect 544 3856 552 3886
rect 578 3856 582 3886
rect 544 3847 548 3856
rect 400 3807 434 3811
rect 400 3777 408 3807
rect 420 3777 434 3807
rect 544 3809 548 3817
rect 12 3738 62 3740
rect 28 3729 59 3731
rect 62 3729 64 3738
rect 28 3721 64 3729
rect 127 3729 158 3731
rect 127 3722 182 3729
rect 215 3727 224 3755
rect 127 3721 161 3722
rect 59 3705 64 3721
rect 158 3705 161 3721
rect 28 3697 64 3705
rect 127 3704 161 3705
rect 127 3697 182 3704
rect 62 3688 64 3697
rect 213 3689 224 3727
rect 282 3717 292 3775
rect 296 3769 368 3777
rect 319 3740 335 3742
rect 251 3683 263 3717
rect 273 3683 292 3717
rect 303 3710 316 3726
rect 303 3692 316 3708
rect 120 3635 170 3637
rect 76 3629 92 3635
rect 94 3629 110 3635
rect 76 3619 99 3628
rect 60 3609 67 3619
rect 76 3599 77 3619
rect 96 3594 99 3619
rect 109 3599 110 3619
rect 119 3609 126 3619
rect 76 3585 110 3589
rect 170 3585 172 3635
rect 186 3617 190 3651
rect 216 3617 220 3651
rect 186 3540 220 3574
rect 282 3571 292 3683
rect 318 3686 324 3739
rect 346 3726 348 3739
rect 428 3730 430 3777
rect 443 3767 450 3769
rect 476 3737 480 3805
rect 544 3775 552 3809
rect 578 3775 582 3809
rect 481 3743 517 3771
rect 481 3737 495 3743
rect 333 3692 353 3726
rect 367 3696 380 3730
rect 396 3696 408 3730
rect 420 3696 434 3730
rect 318 3676 335 3686
rect 318 3607 324 3676
rect 346 3607 348 3692
rect 428 3649 430 3696
rect 476 3659 480 3727
rect 485 3709 495 3737
rect 505 3709 519 3743
rect 544 3737 555 3775
rect 544 3709 553 3737
rect 544 3689 548 3709
rect 579 3668 582 3758
rect 599 3738 649 3740
rect 610 3730 624 3731
rect 607 3729 624 3730
rect 586 3722 644 3729
rect 607 3721 644 3722
rect 607 3705 610 3721
rect 616 3705 644 3721
rect 607 3704 644 3705
rect 586 3697 644 3704
rect 607 3696 610 3697
rect 649 3688 651 3738
rect 544 3651 548 3659
rect 400 3619 408 3649
rect 420 3619 434 3649
rect 400 3615 434 3619
rect 400 3607 430 3615
rect 428 3591 430 3607
rect 476 3579 480 3647
rect 544 3617 552 3651
rect 578 3617 582 3651
rect 544 3609 548 3617
rect 544 3579 586 3580
rect 288 3539 292 3571
rect 296 3569 368 3577
rect 378 3569 450 3577
rect 544 3572 548 3579
rect 439 3541 444 3569
rect 120 3525 170 3527
rect 76 3521 130 3525
rect 110 3516 130 3521
rect 60 3491 67 3501
rect 76 3491 77 3511
rect 96 3482 99 3516
rect 109 3491 110 3511
rect 119 3491 126 3501
rect 76 3475 92 3481
rect 94 3475 110 3481
rect 170 3475 172 3525
rect 186 3459 190 3493
rect 216 3459 220 3493
rect 213 3427 224 3459
rect 282 3455 292 3539
rect 296 3533 368 3541
rect 378 3533 450 3541
rect 468 3538 473 3572
rect 428 3503 430 3519
rect 251 3427 292 3455
rect 12 3422 62 3424
rect 28 3413 59 3415
rect 62 3413 64 3422
rect 251 3421 263 3427
rect 28 3405 64 3413
rect 127 3413 158 3415
rect 127 3406 182 3413
rect 127 3405 161 3406
rect 59 3389 64 3405
rect 158 3389 161 3405
rect 253 3393 263 3421
rect 273 3393 292 3427
rect 318 3434 324 3503
rect 318 3424 335 3434
rect 303 3402 316 3418
rect 28 3381 64 3389
rect 127 3388 161 3389
rect 127 3381 182 3388
rect 62 3372 64 3381
rect 282 3335 292 3393
rect 303 3384 316 3400
rect 318 3371 324 3424
rect 346 3418 348 3503
rect 400 3495 430 3503
rect 476 3501 480 3569
rect 511 3538 582 3572
rect 544 3531 548 3538
rect 400 3491 434 3495
rect 400 3461 408 3491
rect 420 3461 434 3491
rect 544 3493 548 3501
rect 333 3384 353 3418
rect 428 3414 430 3461
rect 476 3421 480 3489
rect 544 3459 552 3493
rect 578 3459 582 3493
rect 544 3451 548 3459
rect 346 3371 348 3384
rect 367 3380 380 3414
rect 396 3380 408 3414
rect 420 3380 434 3414
rect 544 3411 553 3439
rect 319 3368 335 3370
rect 120 3319 170 3321
rect 76 3313 92 3319
rect 94 3313 110 3319
rect 76 3303 99 3312
rect 60 3293 67 3303
rect 76 3283 77 3303
rect 96 3278 99 3303
rect 109 3283 110 3303
rect 119 3293 126 3303
rect 76 3269 110 3273
rect 170 3269 172 3319
rect 186 3301 190 3335
rect 216 3301 220 3335
rect 182 3263 224 3264
rect 186 3222 220 3256
rect 223 3222 257 3256
rect 160 3215 182 3221
rect 224 3215 246 3221
rect 288 3215 292 3335
rect 296 3333 368 3341
rect 428 3333 430 3380
rect 476 3343 480 3411
rect 485 3367 495 3401
rect 505 3367 519 3401
rect 544 3367 555 3411
rect 485 3343 492 3367
rect 579 3352 582 3442
rect 599 3422 649 3424
rect 610 3414 624 3415
rect 607 3413 624 3414
rect 586 3406 644 3413
rect 607 3405 644 3406
rect 607 3389 610 3405
rect 616 3389 644 3405
rect 607 3388 644 3389
rect 586 3381 644 3388
rect 607 3380 610 3381
rect 649 3372 651 3422
rect 544 3335 548 3343
rect 400 3303 408 3333
rect 420 3303 434 3333
rect 400 3299 434 3303
rect 400 3291 430 3299
rect 428 3275 430 3291
rect 476 3263 480 3331
rect 544 3301 552 3335
rect 578 3301 582 3335
rect 544 3293 548 3301
rect 295 3222 300 3256
rect 324 3222 329 3256
rect 378 3253 450 3261
rect 544 3258 548 3263
rect 544 3254 582 3258
rect 544 3224 552 3254
rect 578 3224 582 3254
rect 544 3221 548 3224
rect 522 3215 548 3221
rect 586 3215 608 3221
rect 182 3199 224 3215
rect 544 3199 586 3215
rect 17 3185 67 3187
rect 119 3185 169 3187
rect 599 3185 649 3187
rect 42 3143 59 3177
rect 67 3135 69 3185
rect 160 3177 246 3185
rect 522 3177 608 3185
rect 76 3143 110 3177
rect 127 3143 144 3177
rect 152 3143 161 3177
rect 162 3175 195 3177
rect 224 3175 244 3177
rect 162 3143 244 3175
rect 524 3175 548 3177
rect 573 3175 582 3177
rect 586 3175 606 3177
rect 160 3135 246 3143
rect 186 3119 220 3121
rect 182 3105 224 3106
rect 160 3099 182 3105
rect 224 3099 246 3105
rect 186 3064 220 3098
rect 223 3064 257 3098
rect 120 3051 170 3053
rect 76 3047 130 3051
rect 110 3042 130 3047
rect 60 3017 67 3027
rect 76 3017 77 3037
rect 96 3008 99 3042
rect 109 3017 110 3037
rect 119 3017 126 3027
rect 76 3001 92 3007
rect 94 3001 110 3007
rect 170 3001 172 3051
rect 186 2985 190 3019
rect 216 2985 220 3019
rect 288 2985 292 3173
rect 476 3105 480 3173
rect 524 3143 606 3175
rect 607 3143 616 3177
rect 522 3135 608 3143
rect 649 3135 651 3185
rect 548 3119 582 3121
rect 522 3100 548 3105
rect 522 3099 582 3100
rect 586 3099 608 3105
rect 295 3064 300 3098
rect 324 3064 329 3098
rect 544 3096 582 3099
rect 378 3059 450 3067
rect 428 3029 430 3045
rect 400 3021 430 3029
rect 476 3027 480 3095
rect 544 3066 552 3096
rect 578 3066 582 3096
rect 544 3057 548 3066
rect 400 3017 434 3021
rect 400 2987 408 3017
rect 420 2987 434 3017
rect 544 3019 548 3027
rect 12 2948 62 2950
rect 28 2939 59 2941
rect 62 2939 64 2948
rect 28 2931 64 2939
rect 127 2939 158 2941
rect 127 2932 182 2939
rect 215 2937 224 2965
rect 127 2931 161 2932
rect 59 2915 64 2931
rect 158 2915 161 2931
rect 28 2907 64 2915
rect 127 2914 161 2915
rect 127 2907 182 2914
rect 62 2898 64 2907
rect 213 2899 224 2937
rect 282 2927 292 2985
rect 296 2979 368 2987
rect 319 2950 335 2952
rect 251 2893 263 2927
rect 273 2893 292 2927
rect 303 2920 316 2936
rect 303 2902 316 2918
rect 120 2845 170 2847
rect 76 2839 92 2845
rect 94 2839 110 2845
rect 76 2829 99 2838
rect 60 2819 67 2829
rect 76 2809 77 2829
rect 96 2804 99 2829
rect 109 2809 110 2829
rect 119 2819 126 2829
rect 76 2795 110 2799
rect 170 2795 172 2845
rect 186 2827 190 2861
rect 216 2827 220 2861
rect 186 2750 220 2784
rect 282 2781 292 2893
rect 318 2896 324 2949
rect 346 2936 348 2949
rect 428 2940 430 2987
rect 443 2977 450 2979
rect 476 2947 480 3015
rect 544 2985 552 3019
rect 578 2985 582 3019
rect 481 2953 517 2981
rect 481 2947 495 2953
rect 333 2902 353 2936
rect 367 2906 380 2940
rect 396 2906 408 2940
rect 420 2906 434 2940
rect 318 2886 335 2896
rect 318 2817 324 2886
rect 346 2817 348 2902
rect 428 2859 430 2906
rect 476 2869 480 2937
rect 485 2919 495 2947
rect 505 2919 519 2953
rect 544 2947 555 2985
rect 544 2919 553 2947
rect 544 2899 548 2919
rect 579 2878 582 2968
rect 599 2948 649 2950
rect 610 2940 624 2941
rect 607 2939 624 2940
rect 586 2932 644 2939
rect 607 2931 644 2932
rect 607 2915 610 2931
rect 616 2915 644 2931
rect 607 2914 644 2915
rect 586 2907 644 2914
rect 607 2906 610 2907
rect 649 2898 651 2948
rect 544 2861 548 2869
rect 400 2829 408 2859
rect 420 2829 434 2859
rect 400 2825 434 2829
rect 400 2817 430 2825
rect 428 2801 430 2817
rect 476 2789 480 2857
rect 544 2827 552 2861
rect 578 2827 582 2861
rect 544 2819 548 2827
rect 544 2789 586 2790
rect 288 2749 292 2781
rect 296 2779 368 2787
rect 378 2779 450 2787
rect 544 2782 548 2789
rect 439 2751 444 2779
rect 120 2735 170 2737
rect 76 2731 130 2735
rect 110 2726 130 2731
rect 60 2701 67 2711
rect 76 2701 77 2721
rect 96 2692 99 2726
rect 109 2701 110 2721
rect 119 2701 126 2711
rect 76 2685 92 2691
rect 94 2685 110 2691
rect 170 2685 172 2735
rect 186 2669 190 2703
rect 216 2669 220 2703
rect 213 2637 224 2669
rect 282 2665 292 2749
rect 296 2743 368 2751
rect 378 2743 450 2751
rect 468 2748 473 2782
rect 428 2713 430 2729
rect 251 2637 292 2665
rect 12 2632 62 2634
rect 28 2623 59 2625
rect 62 2623 64 2632
rect 251 2631 263 2637
rect 28 2615 64 2623
rect 127 2623 158 2625
rect 127 2616 182 2623
rect 127 2615 161 2616
rect 59 2599 64 2615
rect 158 2599 161 2615
rect 253 2603 263 2631
rect 273 2603 292 2637
rect 318 2644 324 2713
rect 318 2634 335 2644
rect 303 2612 316 2628
rect 28 2591 64 2599
rect 127 2598 161 2599
rect 127 2591 182 2598
rect 62 2582 64 2591
rect 282 2545 292 2603
rect 303 2594 316 2610
rect 318 2581 324 2634
rect 346 2628 348 2713
rect 400 2705 430 2713
rect 476 2711 480 2779
rect 511 2748 582 2782
rect 544 2741 548 2748
rect 400 2701 434 2705
rect 400 2671 408 2701
rect 420 2671 434 2701
rect 544 2703 548 2711
rect 333 2594 353 2628
rect 428 2624 430 2671
rect 476 2631 480 2699
rect 544 2669 552 2703
rect 578 2669 582 2703
rect 544 2661 548 2669
rect 346 2581 348 2594
rect 367 2590 380 2624
rect 396 2590 408 2624
rect 420 2590 434 2624
rect 544 2621 553 2649
rect 319 2578 335 2580
rect 120 2529 170 2531
rect 76 2523 92 2529
rect 94 2523 110 2529
rect 76 2513 99 2522
rect 60 2503 67 2513
rect 76 2493 77 2513
rect 96 2488 99 2513
rect 109 2493 110 2513
rect 119 2503 126 2513
rect 76 2479 110 2483
rect 170 2479 172 2529
rect 186 2511 190 2545
rect 216 2511 220 2545
rect 182 2473 224 2474
rect 186 2432 220 2466
rect 223 2432 257 2466
rect 160 2425 182 2431
rect 224 2425 246 2431
rect 288 2425 292 2545
rect 296 2543 368 2551
rect 428 2543 430 2590
rect 476 2553 480 2621
rect 485 2577 495 2611
rect 505 2577 519 2611
rect 544 2577 555 2621
rect 485 2553 492 2577
rect 579 2562 582 2652
rect 599 2632 649 2634
rect 610 2624 624 2625
rect 607 2623 624 2624
rect 586 2616 644 2623
rect 607 2615 644 2616
rect 607 2599 610 2615
rect 616 2599 644 2615
rect 607 2598 644 2599
rect 586 2591 644 2598
rect 607 2590 610 2591
rect 649 2582 651 2632
rect 544 2545 548 2553
rect 400 2513 408 2543
rect 420 2513 434 2543
rect 400 2509 434 2513
rect 400 2501 430 2509
rect 428 2485 430 2501
rect 476 2473 480 2541
rect 544 2511 552 2545
rect 578 2511 582 2545
rect 544 2503 548 2511
rect 295 2432 300 2466
rect 324 2432 329 2466
rect 378 2463 450 2471
rect 544 2468 548 2473
rect 544 2464 582 2468
rect 544 2434 552 2464
rect 578 2434 582 2464
rect 544 2431 548 2434
rect 522 2425 548 2431
rect 586 2425 608 2431
rect 182 2409 224 2425
rect 544 2409 586 2425
rect 17 2395 67 2397
rect 119 2395 169 2397
rect 599 2395 649 2397
rect 42 2353 59 2387
rect 67 2345 69 2395
rect 160 2387 246 2395
rect 522 2387 608 2395
rect 76 2353 110 2387
rect 127 2353 144 2387
rect 152 2353 161 2387
rect 162 2385 195 2387
rect 224 2385 244 2387
rect 162 2353 244 2385
rect 524 2385 548 2387
rect 573 2385 582 2387
rect 586 2385 606 2387
rect 160 2345 246 2353
rect 186 2329 220 2331
rect 182 2315 224 2316
rect 160 2309 182 2315
rect 224 2309 246 2315
rect 186 2274 220 2308
rect 223 2274 257 2308
rect 120 2261 170 2263
rect 76 2257 130 2261
rect 110 2252 130 2257
rect 60 2227 67 2237
rect 76 2227 77 2247
rect 96 2218 99 2252
rect 109 2227 110 2247
rect 119 2227 126 2237
rect 76 2211 92 2217
rect 94 2211 110 2217
rect 170 2211 172 2261
rect 186 2195 190 2229
rect 216 2195 220 2229
rect 288 2195 292 2383
rect 476 2315 480 2383
rect 524 2353 606 2385
rect 607 2353 616 2387
rect 522 2345 608 2353
rect 649 2345 651 2395
rect 548 2329 582 2331
rect 522 2310 548 2315
rect 522 2309 582 2310
rect 586 2309 608 2315
rect 295 2274 300 2308
rect 324 2274 329 2308
rect 544 2306 582 2309
rect 378 2269 450 2277
rect 428 2239 430 2255
rect 400 2231 430 2239
rect 476 2237 480 2305
rect 544 2276 552 2306
rect 578 2276 582 2306
rect 544 2267 548 2276
rect 400 2227 434 2231
rect 400 2197 408 2227
rect 420 2197 434 2227
rect 544 2229 548 2237
rect 12 2158 62 2160
rect 28 2149 59 2151
rect 62 2149 64 2158
rect 28 2141 64 2149
rect 127 2149 158 2151
rect 127 2142 182 2149
rect 215 2147 224 2175
rect 127 2141 161 2142
rect 59 2125 64 2141
rect 158 2125 161 2141
rect 28 2117 64 2125
rect 127 2124 161 2125
rect 127 2117 182 2124
rect 62 2108 64 2117
rect 213 2109 224 2147
rect 282 2137 292 2195
rect 296 2189 368 2197
rect 319 2160 335 2162
rect 251 2103 263 2137
rect 273 2103 292 2137
rect 303 2130 316 2146
rect 303 2112 316 2128
rect 120 2055 170 2057
rect 76 2049 92 2055
rect 94 2049 110 2055
rect 76 2039 99 2048
rect 60 2029 67 2039
rect 76 2019 77 2039
rect 96 2014 99 2039
rect 109 2019 110 2039
rect 119 2029 126 2039
rect 76 2005 110 2009
rect 170 2005 172 2055
rect 186 2037 190 2071
rect 216 2037 220 2071
rect 186 1960 220 1994
rect 282 1991 292 2103
rect 318 2106 324 2159
rect 346 2146 348 2159
rect 428 2150 430 2197
rect 443 2187 450 2189
rect 476 2157 480 2225
rect 544 2195 552 2229
rect 578 2195 582 2229
rect 481 2163 517 2191
rect 481 2157 495 2163
rect 333 2112 353 2146
rect 367 2116 380 2150
rect 396 2116 408 2150
rect 420 2116 434 2150
rect 318 2096 335 2106
rect 318 2027 324 2096
rect 346 2027 348 2112
rect 428 2069 430 2116
rect 476 2079 480 2147
rect 485 2129 495 2157
rect 505 2129 519 2163
rect 544 2157 555 2195
rect 544 2129 553 2157
rect 544 2109 548 2129
rect 579 2088 582 2178
rect 599 2158 649 2160
rect 610 2150 624 2151
rect 607 2149 624 2150
rect 586 2142 644 2149
rect 607 2141 644 2142
rect 607 2125 610 2141
rect 616 2125 644 2141
rect 607 2124 644 2125
rect 586 2117 644 2124
rect 607 2116 610 2117
rect 649 2108 651 2158
rect 544 2071 548 2079
rect 400 2039 408 2069
rect 420 2039 434 2069
rect 400 2035 434 2039
rect 400 2027 430 2035
rect 428 2011 430 2027
rect 476 1999 480 2067
rect 544 2037 552 2071
rect 578 2037 582 2071
rect 544 2029 548 2037
rect 544 1999 586 2000
rect 288 1959 292 1991
rect 296 1989 368 1997
rect 378 1989 450 1997
rect 544 1992 548 1999
rect 439 1961 444 1989
rect 120 1945 170 1947
rect 76 1941 130 1945
rect 110 1936 130 1941
rect 60 1911 67 1921
rect 76 1911 77 1931
rect 96 1902 99 1936
rect 109 1911 110 1931
rect 119 1911 126 1921
rect 76 1895 92 1901
rect 94 1895 110 1901
rect 170 1895 172 1945
rect 186 1879 190 1913
rect 216 1879 220 1913
rect 213 1847 224 1879
rect 282 1875 292 1959
rect 296 1953 368 1961
rect 378 1953 450 1961
rect 468 1958 473 1992
rect 428 1923 430 1939
rect 251 1847 292 1875
rect 12 1842 62 1844
rect 28 1833 59 1835
rect 62 1833 64 1842
rect 251 1841 263 1847
rect 28 1825 64 1833
rect 127 1833 158 1835
rect 127 1826 182 1833
rect 127 1825 161 1826
rect 59 1809 64 1825
rect 158 1809 161 1825
rect 253 1813 263 1841
rect 273 1813 292 1847
rect 318 1854 324 1923
rect 318 1844 335 1854
rect 303 1822 316 1838
rect 28 1801 64 1809
rect 127 1808 161 1809
rect 127 1801 182 1808
rect 62 1792 64 1801
rect 282 1755 292 1813
rect 303 1804 316 1820
rect 318 1791 324 1844
rect 346 1838 348 1923
rect 400 1915 430 1923
rect 476 1921 480 1989
rect 511 1958 582 1992
rect 544 1951 548 1958
rect 400 1911 434 1915
rect 400 1881 408 1911
rect 420 1881 434 1911
rect 544 1913 548 1921
rect 333 1804 353 1838
rect 428 1834 430 1881
rect 476 1841 480 1909
rect 544 1879 552 1913
rect 578 1879 582 1913
rect 544 1871 548 1879
rect 346 1791 348 1804
rect 367 1800 380 1834
rect 396 1800 408 1834
rect 420 1800 434 1834
rect 544 1831 553 1859
rect 319 1788 335 1790
rect 120 1739 170 1741
rect 76 1733 92 1739
rect 94 1733 110 1739
rect 76 1723 99 1732
rect 60 1713 67 1723
rect 76 1703 77 1723
rect 96 1698 99 1723
rect 109 1703 110 1723
rect 119 1713 126 1723
rect 76 1689 110 1693
rect 170 1689 172 1739
rect 186 1721 190 1755
rect 216 1721 220 1755
rect 182 1683 224 1684
rect 186 1642 220 1676
rect 223 1642 257 1676
rect 160 1635 182 1641
rect 224 1635 246 1641
rect 288 1635 292 1755
rect 296 1753 368 1761
rect 428 1753 430 1800
rect 476 1763 480 1831
rect 485 1787 495 1821
rect 505 1787 519 1821
rect 544 1787 555 1831
rect 485 1763 492 1787
rect 579 1772 582 1862
rect 599 1842 649 1844
rect 610 1834 624 1835
rect 607 1833 624 1834
rect 586 1826 644 1833
rect 607 1825 644 1826
rect 607 1809 610 1825
rect 616 1809 644 1825
rect 607 1808 644 1809
rect 586 1801 644 1808
rect 607 1800 610 1801
rect 649 1792 651 1842
rect 544 1755 548 1763
rect 400 1723 408 1753
rect 420 1723 434 1753
rect 400 1719 434 1723
rect 400 1711 430 1719
rect 428 1695 430 1711
rect 476 1683 480 1751
rect 544 1721 552 1755
rect 578 1721 582 1755
rect 544 1713 548 1721
rect 295 1642 300 1676
rect 324 1642 329 1676
rect 378 1673 450 1681
rect 544 1678 548 1683
rect 544 1674 582 1678
rect 544 1644 552 1674
rect 578 1644 582 1674
rect 544 1641 548 1644
rect 522 1635 548 1641
rect 586 1635 608 1641
rect 182 1619 224 1635
rect 544 1619 586 1635
rect 17 1605 67 1607
rect 119 1605 169 1607
rect 599 1605 649 1607
rect 42 1563 59 1597
rect 67 1555 69 1605
rect 160 1597 246 1605
rect 522 1597 608 1605
rect 76 1563 110 1597
rect 127 1563 144 1597
rect 152 1563 161 1597
rect 162 1595 195 1597
rect 224 1595 244 1597
rect 162 1563 244 1595
rect 524 1595 548 1597
rect 573 1595 582 1597
rect 586 1595 606 1597
rect 160 1555 246 1563
rect 186 1539 220 1541
rect 182 1525 224 1526
rect 160 1519 182 1525
rect 224 1519 246 1525
rect 186 1484 220 1518
rect 223 1484 257 1518
rect 120 1471 170 1473
rect 76 1467 130 1471
rect 110 1462 130 1467
rect 60 1437 67 1447
rect 76 1437 77 1457
rect 96 1428 99 1462
rect 109 1437 110 1457
rect 119 1437 126 1447
rect 76 1421 92 1427
rect 94 1421 110 1427
rect 170 1421 172 1471
rect 186 1405 190 1439
rect 216 1405 220 1439
rect 288 1405 292 1593
rect 476 1525 480 1593
rect 524 1563 606 1595
rect 607 1563 616 1597
rect 522 1555 608 1563
rect 649 1555 651 1605
rect 548 1539 582 1541
rect 522 1520 548 1525
rect 522 1519 582 1520
rect 586 1519 608 1525
rect 295 1484 300 1518
rect 324 1484 329 1518
rect 544 1516 582 1519
rect 378 1479 450 1487
rect 428 1449 430 1465
rect 400 1441 430 1449
rect 476 1447 480 1515
rect 544 1486 552 1516
rect 578 1486 582 1516
rect 544 1477 548 1486
rect 400 1437 434 1441
rect 400 1407 408 1437
rect 420 1407 434 1437
rect 544 1439 548 1447
rect 12 1368 62 1370
rect 28 1359 59 1361
rect 62 1359 64 1368
rect 28 1351 64 1359
rect 127 1359 158 1361
rect 127 1352 182 1359
rect 215 1357 224 1385
rect 127 1351 161 1352
rect 59 1335 64 1351
rect 158 1335 161 1351
rect 28 1327 64 1335
rect 127 1334 161 1335
rect 127 1327 182 1334
rect 62 1318 64 1327
rect 213 1319 224 1357
rect 282 1347 292 1405
rect 296 1399 368 1407
rect 319 1370 335 1372
rect 251 1313 263 1347
rect 273 1313 292 1347
rect 303 1340 316 1356
rect 303 1322 316 1338
rect 120 1265 170 1267
rect 76 1259 92 1265
rect 94 1259 110 1265
rect 76 1249 99 1258
rect 60 1239 67 1249
rect 76 1229 77 1249
rect 96 1224 99 1249
rect 109 1229 110 1249
rect 119 1239 126 1249
rect 76 1215 110 1219
rect 170 1215 172 1265
rect 186 1247 190 1281
rect 216 1247 220 1281
rect 186 1170 220 1204
rect 282 1201 292 1313
rect 318 1316 324 1369
rect 346 1356 348 1369
rect 428 1360 430 1407
rect 443 1397 450 1399
rect 476 1367 480 1435
rect 544 1405 552 1439
rect 578 1405 582 1439
rect 481 1373 517 1401
rect 481 1367 495 1373
rect 333 1322 353 1356
rect 367 1326 380 1360
rect 396 1326 408 1360
rect 420 1326 434 1360
rect 318 1306 335 1316
rect 318 1237 324 1306
rect 346 1237 348 1322
rect 428 1279 430 1326
rect 476 1289 480 1357
rect 485 1339 495 1367
rect 505 1339 519 1373
rect 544 1367 555 1405
rect 544 1339 553 1367
rect 544 1319 548 1339
rect 579 1298 582 1388
rect 599 1368 649 1370
rect 610 1360 624 1361
rect 607 1359 624 1360
rect 586 1352 644 1359
rect 607 1351 644 1352
rect 607 1335 610 1351
rect 616 1335 644 1351
rect 607 1334 644 1335
rect 586 1327 644 1334
rect 607 1326 610 1327
rect 649 1318 651 1368
rect 544 1281 548 1289
rect 400 1249 408 1279
rect 420 1249 434 1279
rect 400 1245 434 1249
rect 400 1237 430 1245
rect 428 1221 430 1237
rect 476 1209 480 1277
rect 544 1247 552 1281
rect 578 1247 582 1281
rect 544 1239 548 1247
rect 544 1209 586 1210
rect 288 1169 292 1201
rect 296 1199 368 1207
rect 378 1199 450 1207
rect 544 1202 548 1209
rect 439 1171 444 1199
rect 120 1155 170 1157
rect 76 1151 130 1155
rect 110 1146 130 1151
rect 60 1121 67 1131
rect 76 1121 77 1141
rect 96 1112 99 1146
rect 109 1121 110 1141
rect 119 1121 126 1131
rect 76 1105 92 1111
rect 94 1105 110 1111
rect 170 1105 172 1155
rect 186 1089 190 1123
rect 216 1089 220 1123
rect 213 1057 224 1089
rect 282 1085 292 1169
rect 296 1163 368 1171
rect 378 1163 450 1171
rect 468 1168 473 1202
rect 428 1133 430 1149
rect 251 1057 292 1085
rect 12 1052 62 1054
rect 28 1043 59 1045
rect 62 1043 64 1052
rect 251 1051 263 1057
rect 28 1035 64 1043
rect 127 1043 158 1045
rect 127 1036 182 1043
rect 127 1035 161 1036
rect 59 1019 64 1035
rect 158 1019 161 1035
rect 253 1023 263 1051
rect 273 1023 292 1057
rect 318 1064 324 1133
rect 318 1054 335 1064
rect 303 1032 316 1048
rect 28 1011 64 1019
rect 127 1018 161 1019
rect 127 1011 182 1018
rect 62 1002 64 1011
rect 282 965 292 1023
rect 303 1014 316 1030
rect 318 1001 324 1054
rect 346 1048 348 1133
rect 400 1125 430 1133
rect 476 1131 480 1199
rect 511 1168 582 1202
rect 544 1161 548 1168
rect 400 1121 434 1125
rect 400 1091 408 1121
rect 420 1091 434 1121
rect 544 1123 548 1131
rect 333 1014 353 1048
rect 428 1044 430 1091
rect 476 1051 480 1119
rect 544 1089 552 1123
rect 578 1089 582 1123
rect 544 1081 548 1089
rect 346 1001 348 1014
rect 367 1010 380 1044
rect 396 1010 408 1044
rect 420 1010 434 1044
rect 544 1041 553 1069
rect 319 998 335 1000
rect 120 949 170 951
rect 76 943 92 949
rect 94 943 110 949
rect 76 933 99 942
rect 60 923 67 933
rect 76 913 77 933
rect 96 908 99 933
rect 109 913 110 933
rect 119 923 126 933
rect 76 899 110 903
rect 170 899 172 949
rect 186 931 190 965
rect 216 931 220 965
rect 182 893 224 894
rect 186 852 220 886
rect 223 852 257 886
rect 160 845 182 851
rect 224 845 246 851
rect 288 845 292 965
rect 296 963 368 971
rect 428 963 430 1010
rect 476 973 480 1041
rect 485 997 495 1031
rect 505 997 519 1031
rect 544 997 555 1041
rect 485 973 492 997
rect 579 982 582 1072
rect 599 1052 649 1054
rect 610 1044 624 1045
rect 607 1043 624 1044
rect 586 1036 644 1043
rect 607 1035 644 1036
rect 607 1019 610 1035
rect 616 1019 644 1035
rect 607 1018 644 1019
rect 586 1011 644 1018
rect 607 1010 610 1011
rect 649 1002 651 1052
rect 544 965 548 973
rect 400 933 408 963
rect 420 933 434 963
rect 400 929 434 933
rect 400 921 430 929
rect 428 905 430 921
rect 476 893 480 961
rect 544 931 552 965
rect 578 931 582 965
rect 544 923 548 931
rect 295 852 300 886
rect 324 852 329 886
rect 378 883 450 891
rect 544 888 548 893
rect 544 884 582 888
rect 544 854 552 884
rect 578 854 582 884
rect 544 851 548 854
rect 522 845 548 851
rect 586 845 608 851
rect 182 829 224 845
rect 544 829 586 845
rect 17 815 67 817
rect 119 815 169 817
rect 599 815 649 817
rect 42 773 59 807
rect 67 765 69 815
rect 160 807 246 815
rect 522 807 608 815
rect 76 773 110 807
rect 127 773 144 807
rect 152 773 161 807
rect 162 805 195 807
rect 224 805 244 807
rect 162 773 244 805
rect 524 805 548 807
rect 573 805 582 807
rect 586 805 606 807
rect 160 765 246 773
rect 186 749 220 751
rect 182 735 224 736
rect 160 729 182 735
rect 224 729 246 735
rect 186 694 220 728
rect 223 694 257 728
rect 120 681 170 683
rect 76 677 130 681
rect 110 672 130 677
rect 60 647 67 657
rect 76 647 77 667
rect 96 638 99 672
rect 109 647 110 667
rect 119 647 126 657
rect 76 631 92 637
rect 94 631 110 637
rect 170 631 172 681
rect 186 615 190 649
rect 216 615 220 649
rect 288 615 292 803
rect 476 735 480 803
rect 524 773 606 805
rect 607 773 616 807
rect 522 765 608 773
rect 649 765 651 815
rect 548 749 582 751
rect 522 730 548 735
rect 522 729 582 730
rect 586 729 608 735
rect 295 694 300 728
rect 324 694 329 728
rect 544 726 582 729
rect 378 689 450 697
rect 428 659 430 675
rect 400 651 430 659
rect 476 657 480 725
rect 544 696 552 726
rect 578 696 582 726
rect 544 687 548 696
rect 400 647 434 651
rect 400 617 408 647
rect 420 617 434 647
rect 544 649 548 657
rect 12 578 62 580
rect 28 569 59 571
rect 62 569 64 578
rect 28 561 64 569
rect 127 569 158 571
rect 127 562 182 569
rect 215 567 224 595
rect 127 561 161 562
rect 59 545 64 561
rect 158 545 161 561
rect 28 537 64 545
rect 127 544 161 545
rect 127 537 182 544
rect 62 528 64 537
rect 213 529 224 567
rect 282 557 292 615
rect 296 609 368 617
rect 319 580 335 582
rect 251 523 263 557
rect 273 523 292 557
rect 303 550 316 566
rect 303 532 316 548
rect 120 475 170 477
rect 76 469 92 475
rect 94 469 110 475
rect 76 459 99 468
rect 60 449 67 459
rect 76 439 77 459
rect 96 434 99 459
rect 109 439 110 459
rect 119 449 126 459
rect 76 425 110 429
rect 170 425 172 475
rect 186 457 190 491
rect 216 457 220 491
rect 186 411 220 429
rect 282 411 292 523
rect 318 526 324 579
rect 346 566 348 579
rect 428 570 430 617
rect 443 607 450 609
rect 476 577 480 645
rect 544 615 552 649
rect 578 615 582 649
rect 481 583 517 611
rect 481 577 495 583
rect 333 532 353 566
rect 367 536 380 570
rect 396 536 408 570
rect 420 536 434 570
rect 318 516 335 526
rect 318 447 324 516
rect 346 447 348 532
rect 428 489 430 536
rect 476 499 480 567
rect 485 549 495 577
rect 505 549 519 583
rect 544 577 555 615
rect 544 549 553 577
rect 544 529 548 549
rect 579 508 582 598
rect 599 578 649 580
rect 610 570 624 571
rect 607 569 624 570
rect 586 562 644 569
rect 607 561 644 562
rect 607 545 610 561
rect 616 545 644 561
rect 607 544 644 545
rect 586 537 644 544
rect 607 536 610 537
rect 649 528 651 578
rect 544 491 548 499
rect 400 459 408 489
rect 420 459 434 489
rect 400 455 434 459
rect 400 447 430 455
rect 428 431 430 447
rect 476 419 480 487
rect 544 457 552 491
rect 578 457 582 491
rect 544 449 548 457
rect 548 420 582 429
rect 544 419 586 420
rect 170 410 236 411
rect 186 403 190 410
rect 216 403 220 410
rect 186 395 220 403
rect 288 395 292 411
rect 296 409 368 417
rect 378 409 450 417
rect 544 412 582 419
rect 182 369 224 395
rect 439 378 444 409
rect 468 378 473 412
rect 511 395 582 412
rect 511 378 586 395
rect 544 369 586 378
<< metal1 >>
rect 222 0 258 26860
rect 294 0 330 26860
rect 366 26149 402 26490
rect 366 25359 402 25991
rect 366 24569 402 25201
rect 366 23779 402 24411
rect 366 22989 402 23621
rect 366 22199 402 22831
rect 366 21409 402 22041
rect 366 20619 402 21251
rect 366 19829 402 20461
rect 366 19039 402 19671
rect 366 18249 402 18881
rect 366 17459 402 18091
rect 366 16669 402 17301
rect 366 15879 402 16511
rect 366 15089 402 15721
rect 366 14299 402 14931
rect 366 13509 402 14141
rect 366 12719 402 13351
rect 366 11929 402 12561
rect 366 11139 402 11771
rect 366 10349 402 10981
rect 366 9559 402 10191
rect 366 8769 402 9401
rect 366 7979 402 8611
rect 366 7189 402 7821
rect 366 6399 402 7031
rect 366 5609 402 6241
rect 366 4819 402 5451
rect 366 4029 402 4661
rect 366 3239 402 3871
rect 366 2449 402 3081
rect 366 1659 402 2291
rect 366 869 402 1501
rect 366 370 402 711
rect 438 0 474 26860
rect 510 0 546 26860
<< metal2 >>
rect 0 26576 624 26686
rect 0 26393 624 26441
rect 330 26269 438 26345
rect 0 26173 624 26221
rect 330 26015 438 26125
rect 0 25919 624 25967
rect 330 25795 438 25871
rect 0 25699 624 25747
rect 0 25603 624 25651
rect 330 25479 438 25555
rect 0 25383 624 25431
rect 330 25225 438 25335
rect 0 25129 624 25177
rect 330 25005 438 25081
rect 0 24909 624 24957
rect 0 24813 624 24861
rect 330 24689 438 24765
rect 0 24593 624 24641
rect 330 24435 438 24545
rect 0 24339 624 24387
rect 330 24215 438 24291
rect 0 24119 624 24167
rect 0 24023 624 24071
rect 330 23899 438 23975
rect 0 23803 624 23851
rect 330 23645 438 23755
rect 0 23549 624 23597
rect 330 23425 438 23501
rect 0 23329 624 23377
rect 0 23233 624 23281
rect 330 23109 438 23185
rect 0 23013 624 23061
rect 330 22855 438 22965
rect 0 22759 624 22807
rect 330 22635 438 22711
rect 0 22539 624 22587
rect 0 22443 624 22491
rect 330 22319 438 22395
rect 0 22223 624 22271
rect 330 22065 438 22175
rect 0 21969 624 22017
rect 330 21845 438 21921
rect 0 21749 624 21797
rect 0 21653 624 21701
rect 330 21529 438 21605
rect 0 21433 624 21481
rect 330 21275 438 21385
rect 0 21179 624 21227
rect 330 21055 438 21131
rect 0 20959 624 21007
rect 0 20863 624 20911
rect 330 20739 438 20815
rect 0 20643 624 20691
rect 330 20485 438 20595
rect 0 20389 624 20437
rect 330 20265 438 20341
rect 0 20169 624 20217
rect 0 20073 624 20121
rect 330 19949 438 20025
rect 0 19853 624 19901
rect 330 19695 438 19805
rect 0 19599 624 19647
rect 330 19475 438 19551
rect 0 19379 624 19427
rect 0 19283 624 19331
rect 330 19159 438 19235
rect 0 19063 624 19111
rect 330 18905 438 19015
rect 0 18809 624 18857
rect 330 18685 438 18761
rect 0 18589 624 18637
rect 0 18493 624 18541
rect 330 18369 438 18445
rect 0 18273 624 18321
rect 330 18115 438 18225
rect 0 18019 624 18067
rect 330 17895 438 17971
rect 0 17799 624 17847
rect 0 17703 624 17751
rect 330 17579 438 17655
rect 0 17483 624 17531
rect 330 17325 438 17435
rect 0 17229 624 17277
rect 330 17105 438 17181
rect 0 17009 624 17057
rect 0 16913 624 16961
rect 330 16789 438 16865
rect 0 16693 624 16741
rect 330 16535 438 16645
rect 0 16439 624 16487
rect 330 16315 438 16391
rect 0 16219 624 16267
rect 0 16123 624 16171
rect 330 15999 438 16075
rect 0 15903 624 15951
rect 330 15745 438 15855
rect 0 15649 624 15697
rect 330 15525 438 15601
rect 0 15429 624 15477
rect 0 15333 624 15381
rect 330 15209 438 15285
rect 0 15113 624 15161
rect 330 14955 438 15065
rect 0 14859 624 14907
rect 330 14735 438 14811
rect 0 14639 624 14687
rect 0 14543 624 14591
rect 330 14419 438 14495
rect 0 14323 624 14371
rect 330 14165 438 14275
rect 0 14069 624 14117
rect 330 13945 438 14021
rect 0 13849 624 13897
rect 0 13753 624 13801
rect 330 13629 438 13705
rect 0 13533 624 13581
rect 330 13375 438 13485
rect 0 13279 624 13327
rect 330 13155 438 13231
rect 0 13059 624 13107
rect 0 12963 624 13011
rect 330 12839 438 12915
rect 0 12743 624 12791
rect 330 12585 438 12695
rect 0 12489 624 12537
rect 330 12365 438 12441
rect 0 12269 624 12317
rect 0 12173 624 12221
rect 330 12049 438 12125
rect 0 11953 624 12001
rect 330 11795 438 11905
rect 0 11699 624 11747
rect 330 11575 438 11651
rect 0 11479 624 11527
rect 0 11383 624 11431
rect 330 11259 438 11335
rect 0 11163 624 11211
rect 330 11005 438 11115
rect 0 10909 624 10957
rect 330 10785 438 10861
rect 0 10689 624 10737
rect 0 10593 624 10641
rect 330 10469 438 10545
rect 0 10373 624 10421
rect 330 10215 438 10325
rect 0 10119 624 10167
rect 330 9995 438 10071
rect 0 9899 624 9947
rect 0 9803 624 9851
rect 330 9679 438 9755
rect 0 9583 624 9631
rect 330 9425 438 9535
rect 0 9329 624 9377
rect 330 9205 438 9281
rect 0 9109 624 9157
rect 0 9013 624 9061
rect 330 8889 438 8965
rect 0 8793 624 8841
rect 330 8635 438 8745
rect 0 8539 624 8587
rect 330 8415 438 8491
rect 0 8319 624 8367
rect 0 8223 624 8271
rect 330 8099 438 8175
rect 0 8003 624 8051
rect 330 7845 438 7955
rect 0 7749 624 7797
rect 330 7625 438 7701
rect 0 7529 624 7577
rect 0 7433 624 7481
rect 330 7309 438 7385
rect 0 7213 624 7261
rect 330 7055 438 7165
rect 0 6959 624 7007
rect 330 6835 438 6911
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 330 6519 438 6595
rect 0 6423 624 6471
rect 330 6265 438 6375
rect 0 6169 624 6217
rect 330 6045 438 6121
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 330 5729 438 5805
rect 0 5633 624 5681
rect 330 5475 438 5585
rect 0 5379 624 5427
rect 330 5255 438 5331
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 330 4939 438 5015
rect 0 4843 624 4891
rect 330 4685 438 4795
rect 0 4589 624 4637
rect 330 4465 438 4541
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 330 4149 438 4225
rect 0 4053 624 4101
rect 330 3895 438 4005
rect 0 3799 624 3847
rect 330 3675 438 3751
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 330 3359 438 3435
rect 0 3263 624 3311
rect 330 3105 438 3215
rect 0 3009 624 3057
rect 330 2885 438 2961
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 330 2569 438 2645
rect 0 2473 624 2521
rect 330 2315 438 2425
rect 0 2219 624 2267
rect 330 2095 438 2171
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 330 1779 438 1855
rect 0 1683 624 1731
rect 330 1525 438 1635
rect 0 1429 624 1477
rect 330 1305 438 1381
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 330 989 438 1065
rect 0 893 624 941
rect 330 735 438 845
rect 0 639 624 687
rect 330 515 438 591
rect 0 419 624 467
rect 0 174 624 284
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_0
timestamp 1661296025
transform -1 0 624 0 -1 26860
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_cap_col  sky130_fd_bd_sram__openram_dp_cell_cap_col_1
timestamp 1661296025
transform -1 0 624 0 1 0
box 0 0 624 474
use sky130_fd_bd_sram__openram_dp_cell_dummy  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1661296025
transform -1 0 624 0 1 26070
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_0
timestamp 1661296025
transform -1 0 624 0 -1 26070
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_1
timestamp 1661296025
transform -1 0 624 0 1 25280
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_2
timestamp 1661296025
transform -1 0 624 0 -1 25280
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_3
timestamp 1661296025
transform -1 0 624 0 1 24490
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_4
timestamp 1661296025
transform -1 0 624 0 -1 24490
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_5
timestamp 1661296025
transform -1 0 624 0 1 23700
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_6
timestamp 1661296025
transform -1 0 624 0 -1 23700
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_7
timestamp 1661296025
transform -1 0 624 0 1 22910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_8
timestamp 1661296025
transform -1 0 624 0 -1 22910
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_9
timestamp 1661296025
transform -1 0 624 0 1 22120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_10
timestamp 1661296025
transform -1 0 624 0 -1 22120
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_11
timestamp 1661296025
transform -1 0 624 0 1 21330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_12
timestamp 1661296025
transform -1 0 624 0 -1 21330
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_13
timestamp 1661296025
transform -1 0 624 0 1 20540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_14
timestamp 1661296025
transform -1 0 624 0 -1 20540
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_15
timestamp 1661296025
transform -1 0 624 0 1 19750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_16
timestamp 1661296025
transform -1 0 624 0 -1 19750
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_17
timestamp 1661296025
transform -1 0 624 0 1 18960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_18
timestamp 1661296025
transform -1 0 624 0 -1 18960
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_19
timestamp 1661296025
transform -1 0 624 0 1 18170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_20
timestamp 1661296025
transform -1 0 624 0 -1 18170
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_21
timestamp 1661296025
transform -1 0 624 0 1 17380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_22
timestamp 1661296025
transform -1 0 624 0 -1 17380
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_23
timestamp 1661296025
transform -1 0 624 0 1 16590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_24
timestamp 1661296025
transform -1 0 624 0 -1 16590
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_25
timestamp 1661296025
transform -1 0 624 0 1 15800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_26
timestamp 1661296025
transform -1 0 624 0 -1 15800
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_27
timestamp 1661296025
transform -1 0 624 0 1 15010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_28
timestamp 1661296025
transform -1 0 624 0 -1 15010
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_29
timestamp 1661296025
transform -1 0 624 0 1 14220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_30
timestamp 1661296025
transform -1 0 624 0 -1 14220
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_31
timestamp 1661296025
transform -1 0 624 0 1 13430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_32
timestamp 1661296025
transform -1 0 624 0 -1 13430
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_33
timestamp 1661296025
transform -1 0 624 0 1 12640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_34
timestamp 1661296025
transform -1 0 624 0 -1 12640
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_35
timestamp 1661296025
transform -1 0 624 0 1 11850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_36
timestamp 1661296025
transform -1 0 624 0 -1 11850
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_37
timestamp 1661296025
transform -1 0 624 0 1 11060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_38
timestamp 1661296025
transform -1 0 624 0 -1 11060
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_39
timestamp 1661296025
transform -1 0 624 0 1 10270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_40
timestamp 1661296025
transform -1 0 624 0 -1 10270
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_41
timestamp 1661296025
transform -1 0 624 0 1 9480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_42
timestamp 1661296025
transform -1 0 624 0 -1 9480
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_43
timestamp 1661296025
transform -1 0 624 0 1 8690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_44
timestamp 1661296025
transform -1 0 624 0 -1 8690
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_45
timestamp 1661296025
transform -1 0 624 0 1 7900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_46
timestamp 1661296025
transform -1 0 624 0 -1 7900
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_47
timestamp 1661296025
transform -1 0 624 0 1 7110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_48
timestamp 1661296025
transform -1 0 624 0 -1 7110
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_49
timestamp 1661296025
transform -1 0 624 0 1 6320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_50
timestamp 1661296025
transform -1 0 624 0 -1 6320
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_51
timestamp 1661296025
transform -1 0 624 0 1 5530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_52
timestamp 1661296025
transform -1 0 624 0 -1 5530
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_53
timestamp 1661296025
transform -1 0 624 0 1 4740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_54
timestamp 1661296025
transform -1 0 624 0 -1 4740
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_55
timestamp 1661296025
transform -1 0 624 0 1 3950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_56
timestamp 1661296025
transform -1 0 624 0 -1 3950
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_57
timestamp 1661296025
transform -1 0 624 0 1 3160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_58
timestamp 1661296025
transform -1 0 624 0 -1 3160
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_59
timestamp 1661296025
transform -1 0 624 0 1 2370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_60
timestamp 1661296025
transform -1 0 624 0 -1 2370
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_61
timestamp 1661296025
transform -1 0 624 0 1 1580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_62
timestamp 1661296025
transform -1 0 624 0 -1 1580
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_63
timestamp 1661296025
transform -1 0 624 0 1 790
box -42 -105 650 424
use sky130_fd_bd_sram__openram_dp_cell_replica  sky130_fd_bd_sram__openram_dp_cell_replica_64
timestamp 1661296025
transform -1 0 624 0 -1 790
box -42 -105 650 424
<< labels >>
rlabel metal1 s 510 0 546 26860 4 bl_0_0
port 1 nsew
rlabel metal1 s 438 0 474 26860 4 br_0_0
port 2 nsew
rlabel metal1 s 294 0 330 26860 4 bl_1_0
port 3 nsew
rlabel metal1 s 222 0 258 26860 4 br_1_0
port 4 nsew
rlabel metal2 s 0 419 624 467 4 wl_0_0
port 5 nsew
rlabel metal2 s 0 1113 624 1161 4 wl_0_1
port 6 nsew
rlabel metal2 s 0 1209 624 1257 4 wl_0_2
port 7 nsew
rlabel metal2 s 0 1903 624 1951 4 wl_0_3
port 8 nsew
rlabel metal2 s 0 1999 624 2047 4 wl_0_4
port 9 nsew
rlabel metal2 s 0 2693 624 2741 4 wl_0_5
port 10 nsew
rlabel metal2 s 0 2789 624 2837 4 wl_0_6
port 11 nsew
rlabel metal2 s 0 3483 624 3531 4 wl_0_7
port 12 nsew
rlabel metal2 s 0 3579 624 3627 4 wl_0_8
port 13 nsew
rlabel metal2 s 0 4273 624 4321 4 wl_0_9
port 14 nsew
rlabel metal2 s 0 4369 624 4417 4 wl_0_10
port 15 nsew
rlabel metal2 s 0 5063 624 5111 4 wl_0_11
port 16 nsew
rlabel metal2 s 0 5159 624 5207 4 wl_0_12
port 17 nsew
rlabel metal2 s 0 5853 624 5901 4 wl_0_13
port 18 nsew
rlabel metal2 s 0 5949 624 5997 4 wl_0_14
port 19 nsew
rlabel metal2 s 0 6643 624 6691 4 wl_0_15
port 20 nsew
rlabel metal2 s 0 6739 624 6787 4 wl_0_16
port 21 nsew
rlabel metal2 s 0 7433 624 7481 4 wl_0_17
port 22 nsew
rlabel metal2 s 0 7529 624 7577 4 wl_0_18
port 23 nsew
rlabel metal2 s 0 8223 624 8271 4 wl_0_19
port 24 nsew
rlabel metal2 s 0 8319 624 8367 4 wl_0_20
port 25 nsew
rlabel metal2 s 0 9013 624 9061 4 wl_0_21
port 26 nsew
rlabel metal2 s 0 9109 624 9157 4 wl_0_22
port 27 nsew
rlabel metal2 s 0 9803 624 9851 4 wl_0_23
port 28 nsew
rlabel metal2 s 0 9899 624 9947 4 wl_0_24
port 29 nsew
rlabel metal2 s 0 10593 624 10641 4 wl_0_25
port 30 nsew
rlabel metal2 s 0 10689 624 10737 4 wl_0_26
port 31 nsew
rlabel metal2 s 0 11383 624 11431 4 wl_0_27
port 32 nsew
rlabel metal2 s 0 11479 624 11527 4 wl_0_28
port 33 nsew
rlabel metal2 s 0 12173 624 12221 4 wl_0_29
port 34 nsew
rlabel metal2 s 0 12269 624 12317 4 wl_0_30
port 35 nsew
rlabel metal2 s 0 12963 624 13011 4 wl_0_31
port 36 nsew
rlabel metal2 s 0 13059 624 13107 4 wl_0_32
port 37 nsew
rlabel metal2 s 0 13753 624 13801 4 wl_0_33
port 38 nsew
rlabel metal2 s 0 13849 624 13897 4 wl_0_34
port 39 nsew
rlabel metal2 s 0 14543 624 14591 4 wl_0_35
port 40 nsew
rlabel metal2 s 0 14639 624 14687 4 wl_0_36
port 41 nsew
rlabel metal2 s 0 15333 624 15381 4 wl_0_37
port 42 nsew
rlabel metal2 s 0 15429 624 15477 4 wl_0_38
port 43 nsew
rlabel metal2 s 0 16123 624 16171 4 wl_0_39
port 44 nsew
rlabel metal2 s 0 16219 624 16267 4 wl_0_40
port 45 nsew
rlabel metal2 s 0 16913 624 16961 4 wl_0_41
port 46 nsew
rlabel metal2 s 0 17009 624 17057 4 wl_0_42
port 47 nsew
rlabel metal2 s 0 17703 624 17751 4 wl_0_43
port 48 nsew
rlabel metal2 s 0 17799 624 17847 4 wl_0_44
port 49 nsew
rlabel metal2 s 0 18493 624 18541 4 wl_0_45
port 50 nsew
rlabel metal2 s 0 18589 624 18637 4 wl_0_46
port 51 nsew
rlabel metal2 s 0 19283 624 19331 4 wl_0_47
port 52 nsew
rlabel metal2 s 0 19379 624 19427 4 wl_0_48
port 53 nsew
rlabel metal2 s 0 20073 624 20121 4 wl_0_49
port 54 nsew
rlabel metal2 s 0 20169 624 20217 4 wl_0_50
port 55 nsew
rlabel metal2 s 0 20863 624 20911 4 wl_0_51
port 56 nsew
rlabel metal2 s 0 20959 624 21007 4 wl_0_52
port 57 nsew
rlabel metal2 s 0 21653 624 21701 4 wl_0_53
port 58 nsew
rlabel metal2 s 0 21749 624 21797 4 wl_0_54
port 59 nsew
rlabel metal2 s 0 22443 624 22491 4 wl_0_55
port 60 nsew
rlabel metal2 s 0 22539 624 22587 4 wl_0_56
port 61 nsew
rlabel metal2 s 0 23233 624 23281 4 wl_0_57
port 62 nsew
rlabel metal2 s 0 23329 624 23377 4 wl_0_58
port 63 nsew
rlabel metal2 s 0 24023 624 24071 4 wl_0_59
port 64 nsew
rlabel metal2 s 0 24119 624 24167 4 wl_0_60
port 65 nsew
rlabel metal2 s 0 24813 624 24861 4 wl_0_61
port 66 nsew
rlabel metal2 s 0 24909 624 24957 4 wl_0_62
port 67 nsew
rlabel metal2 s 0 25603 624 25651 4 wl_0_63
port 68 nsew
rlabel metal2 s 0 25699 624 25747 4 wl_0_64
port 69 nsew
rlabel metal2 s 0 26393 624 26441 4 wl_0_65
port 70 nsew
rlabel metal2 s 0 639 624 687 4 wl_1_0
port 71 nsew
rlabel metal2 s 0 893 624 941 4 wl_1_1
port 72 nsew
rlabel metal2 s 0 1429 624 1477 4 wl_1_2
port 73 nsew
rlabel metal2 s 0 1683 624 1731 4 wl_1_3
port 74 nsew
rlabel metal2 s 0 2219 624 2267 4 wl_1_4
port 75 nsew
rlabel metal2 s 0 2473 624 2521 4 wl_1_5
port 76 nsew
rlabel metal2 s 0 3009 624 3057 4 wl_1_6
port 77 nsew
rlabel metal2 s 0 3263 624 3311 4 wl_1_7
port 78 nsew
rlabel metal2 s 0 3799 624 3847 4 wl_1_8
port 79 nsew
rlabel metal2 s 0 4053 624 4101 4 wl_1_9
port 80 nsew
rlabel metal2 s 0 4589 624 4637 4 wl_1_10
port 81 nsew
rlabel metal2 s 0 4843 624 4891 4 wl_1_11
port 82 nsew
rlabel metal2 s 0 5379 624 5427 4 wl_1_12
port 83 nsew
rlabel metal2 s 0 5633 624 5681 4 wl_1_13
port 84 nsew
rlabel metal2 s 0 6169 624 6217 4 wl_1_14
port 85 nsew
rlabel metal2 s 0 6423 624 6471 4 wl_1_15
port 86 nsew
rlabel metal2 s 0 6959 624 7007 4 wl_1_16
port 87 nsew
rlabel metal2 s 0 7213 624 7261 4 wl_1_17
port 88 nsew
rlabel metal2 s 0 7749 624 7797 4 wl_1_18
port 89 nsew
rlabel metal2 s 0 8003 624 8051 4 wl_1_19
port 90 nsew
rlabel metal2 s 0 8539 624 8587 4 wl_1_20
port 91 nsew
rlabel metal2 s 0 8793 624 8841 4 wl_1_21
port 92 nsew
rlabel metal2 s 0 9329 624 9377 4 wl_1_22
port 93 nsew
rlabel metal2 s 0 9583 624 9631 4 wl_1_23
port 94 nsew
rlabel metal2 s 0 10119 624 10167 4 wl_1_24
port 95 nsew
rlabel metal2 s 0 10373 624 10421 4 wl_1_25
port 96 nsew
rlabel metal2 s 0 10909 624 10957 4 wl_1_26
port 97 nsew
rlabel metal2 s 0 11163 624 11211 4 wl_1_27
port 98 nsew
rlabel metal2 s 0 11699 624 11747 4 wl_1_28
port 99 nsew
rlabel metal2 s 0 11953 624 12001 4 wl_1_29
port 100 nsew
rlabel metal2 s 0 12489 624 12537 4 wl_1_30
port 101 nsew
rlabel metal2 s 0 12743 624 12791 4 wl_1_31
port 102 nsew
rlabel metal2 s 0 13279 624 13327 4 wl_1_32
port 103 nsew
rlabel metal2 s 0 13533 624 13581 4 wl_1_33
port 104 nsew
rlabel metal2 s 0 14069 624 14117 4 wl_1_34
port 105 nsew
rlabel metal2 s 0 14323 624 14371 4 wl_1_35
port 106 nsew
rlabel metal2 s 0 14859 624 14907 4 wl_1_36
port 107 nsew
rlabel metal2 s 0 15113 624 15161 4 wl_1_37
port 108 nsew
rlabel metal2 s 0 15649 624 15697 4 wl_1_38
port 109 nsew
rlabel metal2 s 0 15903 624 15951 4 wl_1_39
port 110 nsew
rlabel metal2 s 0 16439 624 16487 4 wl_1_40
port 111 nsew
rlabel metal2 s 0 16693 624 16741 4 wl_1_41
port 112 nsew
rlabel metal2 s 0 17229 624 17277 4 wl_1_42
port 113 nsew
rlabel metal2 s 0 17483 624 17531 4 wl_1_43
port 114 nsew
rlabel metal2 s 0 18019 624 18067 4 wl_1_44
port 115 nsew
rlabel metal2 s 0 18273 624 18321 4 wl_1_45
port 116 nsew
rlabel metal2 s 0 18809 624 18857 4 wl_1_46
port 117 nsew
rlabel metal2 s 0 19063 624 19111 4 wl_1_47
port 118 nsew
rlabel metal2 s 0 19599 624 19647 4 wl_1_48
port 119 nsew
rlabel metal2 s 0 19853 624 19901 4 wl_1_49
port 120 nsew
rlabel metal2 s 0 20389 624 20437 4 wl_1_50
port 121 nsew
rlabel metal2 s 0 20643 624 20691 4 wl_1_51
port 122 nsew
rlabel metal2 s 0 21179 624 21227 4 wl_1_52
port 123 nsew
rlabel metal2 s 0 21433 624 21481 4 wl_1_53
port 124 nsew
rlabel metal2 s 0 21969 624 22017 4 wl_1_54
port 125 nsew
rlabel metal2 s 0 22223 624 22271 4 wl_1_55
port 126 nsew
rlabel metal2 s 0 22759 624 22807 4 wl_1_56
port 127 nsew
rlabel metal2 s 0 23013 624 23061 4 wl_1_57
port 128 nsew
rlabel metal2 s 0 23549 624 23597 4 wl_1_58
port 129 nsew
rlabel metal2 s 0 23803 624 23851 4 wl_1_59
port 130 nsew
rlabel metal2 s 0 24339 624 24387 4 wl_1_60
port 131 nsew
rlabel metal2 s 0 24593 624 24641 4 wl_1_61
port 132 nsew
rlabel metal2 s 0 25129 624 25177 4 wl_1_62
port 133 nsew
rlabel metal2 s 0 25383 624 25431 4 wl_1_63
port 134 nsew
rlabel metal2 s 0 25919 624 25967 4 wl_1_64
port 135 nsew
rlabel metal2 s 0 26173 624 26221 4 wl_1_65
port 136 nsew
rlabel metal1 s 366 16960 402 17301 4 vdd
port 137 nsew
rlabel metal1 s 366 9060 402 9401 4 vdd
port 137 nsew
rlabel metal1 s 366 21409 402 21750 4 vdd
port 137 nsew
rlabel metal1 s 366 26149 402 26490 4 vdd
port 137 nsew
rlabel metal1 s 366 1950 402 2291 4 vdd
port 137 nsew
rlabel metal1 s 366 10349 402 10690 4 vdd
port 137 nsew
rlabel metal1 s 366 23779 402 24120 4 vdd
port 137 nsew
rlabel metal1 s 366 12719 402 13060 4 vdd
port 137 nsew
rlabel metal1 s 366 5609 402 5950 4 vdd
port 137 nsew
rlabel metal1 s 366 6399 402 6740 4 vdd
port 137 nsew
rlabel metal1 s 366 9559 402 9900 4 vdd
port 137 nsew
rlabel metal1 s 366 869 402 1210 4 vdd
port 137 nsew
rlabel metal2 s 0 174 624 284 4 vdd
port 137 nsew
rlabel metal1 s 366 3530 402 3871 4 vdd
port 137 nsew
rlabel metal1 s 366 14590 402 14931 4 vdd
port 137 nsew
rlabel metal1 s 366 11929 402 12270 4 vdd
port 137 nsew
rlabel metal1 s 366 17459 402 17800 4 vdd
port 137 nsew
rlabel metal1 s 366 11139 402 11480 4 vdd
port 137 nsew
rlabel metal1 s 366 1659 402 2000 4 vdd
port 137 nsew
rlabel metal1 s 366 18249 402 18590 4 vdd
port 137 nsew
rlabel metal1 s 366 4320 402 4661 4 vdd
port 137 nsew
rlabel metal1 s 366 18540 402 18881 4 vdd
port 137 nsew
rlabel metal1 s 366 24569 402 24910 4 vdd
port 137 nsew
rlabel metal1 s 366 16669 402 17010 4 vdd
port 137 nsew
rlabel metal1 s 366 25359 402 25700 4 vdd
port 137 nsew
rlabel metal1 s 366 5110 402 5451 4 vdd
port 137 nsew
rlabel metal1 s 366 2740 402 3081 4 vdd
port 137 nsew
rlabel metal1 s 366 20120 402 20461 4 vdd
port 137 nsew
rlabel metal1 s 366 10640 402 10981 4 vdd
port 137 nsew
rlabel metal1 s 366 13010 402 13351 4 vdd
port 137 nsew
rlabel metal1 s 366 19330 402 19671 4 vdd
port 137 nsew
rlabel metal1 s 366 20619 402 20960 4 vdd
port 137 nsew
rlabel metal1 s 366 11430 402 11771 4 vdd
port 137 nsew
rlabel metal1 s 366 7189 402 7530 4 vdd
port 137 nsew
rlabel metal1 s 366 15879 402 16220 4 vdd
port 137 nsew
rlabel metal1 s 366 25650 402 25991 4 vdd
port 137 nsew
rlabel metal1 s 366 4029 402 4370 4 vdd
port 137 nsew
rlabel metal1 s 366 9850 402 10191 4 vdd
port 137 nsew
rlabel metal1 s 366 4819 402 5160 4 vdd
port 137 nsew
rlabel metal1 s 366 21700 402 22041 4 vdd
port 137 nsew
rlabel metal1 s 366 17750 402 18091 4 vdd
port 137 nsew
rlabel metal1 s 366 7480 402 7821 4 vdd
port 137 nsew
rlabel metal1 s 366 15380 402 15721 4 vdd
port 137 nsew
rlabel metal1 s 366 2449 402 2790 4 vdd
port 137 nsew
rlabel metal1 s 366 8270 402 8611 4 vdd
port 137 nsew
rlabel metal1 s 366 14299 402 14640 4 vdd
port 137 nsew
rlabel metal1 s 366 23280 402 23621 4 vdd
port 137 nsew
rlabel metal1 s 366 15089 402 15430 4 vdd
port 137 nsew
rlabel metal1 s 366 20910 402 21251 4 vdd
port 137 nsew
rlabel metal2 s 0 26576 624 26686 4 vdd
port 137 nsew
rlabel metal1 s 366 22989 402 23330 4 vdd
port 137 nsew
rlabel metal1 s 366 12220 402 12561 4 vdd
port 137 nsew
rlabel metal1 s 366 370 402 711 4 vdd
port 137 nsew
rlabel metal1 s 366 16170 402 16511 4 vdd
port 137 nsew
rlabel metal1 s 366 19829 402 20170 4 vdd
port 137 nsew
rlabel metal1 s 366 22490 402 22831 4 vdd
port 137 nsew
rlabel metal1 s 366 5900 402 6241 4 vdd
port 137 nsew
rlabel metal1 s 366 8769 402 9110 4 vdd
port 137 nsew
rlabel metal1 s 366 13800 402 14141 4 vdd
port 137 nsew
rlabel metal1 s 366 13509 402 13850 4 vdd
port 137 nsew
rlabel metal1 s 366 3239 402 3580 4 vdd
port 137 nsew
rlabel metal1 s 366 19039 402 19380 4 vdd
port 137 nsew
rlabel metal1 s 366 22199 402 22540 4 vdd
port 137 nsew
rlabel metal1 s 366 24070 402 24411 4 vdd
port 137 nsew
rlabel metal1 s 366 7979 402 8320 4 vdd
port 137 nsew
rlabel metal1 s 366 1160 402 1501 4 vdd
port 137 nsew
rlabel metal1 s 366 6690 402 7031 4 vdd
port 137 nsew
rlabel metal1 s 366 24860 402 25201 4 vdd
port 137 nsew
rlabel metal2 s 330 26015 438 26125 4 gnd
port 138 nsew
rlabel metal2 s 330 989 438 1065 4 gnd
port 138 nsew
rlabel metal2 s 330 17325 438 17435 4 gnd
port 138 nsew
rlabel metal2 s 330 18115 438 18225 4 gnd
port 138 nsew
rlabel metal2 s 330 21529 438 21605 4 gnd
port 138 nsew
rlabel metal2 s 330 4939 438 5015 4 gnd
port 138 nsew
rlabel metal2 s 330 11575 438 11651 4 gnd
port 138 nsew
rlabel metal2 s 330 19695 438 19805 4 gnd
port 138 nsew
rlabel metal2 s 330 22635 438 22711 4 gnd
port 138 nsew
rlabel metal2 s 330 8099 438 8175 4 gnd
port 138 nsew
rlabel metal2 s 330 14165 438 14275 4 gnd
port 138 nsew
rlabel metal2 s 330 21845 438 21921 4 gnd
port 138 nsew
rlabel metal2 s 330 2885 438 2961 4 gnd
port 138 nsew
rlabel metal2 s 330 18685 438 18761 4 gnd
port 138 nsew
rlabel metal2 s 330 4149 438 4225 4 gnd
port 138 nsew
rlabel metal2 s 330 13155 438 13231 4 gnd
port 138 nsew
rlabel metal2 s 330 16315 438 16391 4 gnd
port 138 nsew
rlabel metal2 s 330 23109 438 23185 4 gnd
port 138 nsew
rlabel metal2 s 330 6835 438 6911 4 gnd
port 138 nsew
rlabel metal2 s 330 23645 438 23755 4 gnd
port 138 nsew
rlabel metal2 s 330 14419 438 14495 4 gnd
port 138 nsew
rlabel metal2 s 330 15525 438 15601 4 gnd
port 138 nsew
rlabel metal2 s 330 17105 438 17181 4 gnd
port 138 nsew
rlabel metal2 s 330 5255 438 5331 4 gnd
port 138 nsew
rlabel metal2 s 330 5475 438 5585 4 gnd
port 138 nsew
rlabel metal2 s 330 19475 438 19551 4 gnd
port 138 nsew
rlabel metal2 s 330 11259 438 11335 4 gnd
port 138 nsew
rlabel metal2 s 330 515 438 591 4 gnd
port 138 nsew
rlabel metal2 s 330 25005 438 25081 4 gnd
port 138 nsew
rlabel metal2 s 330 11795 438 11905 4 gnd
port 138 nsew
rlabel metal2 s 330 24435 438 24545 4 gnd
port 138 nsew
rlabel metal2 s 330 15745 438 15855 4 gnd
port 138 nsew
rlabel metal2 s 330 1305 438 1381 4 gnd
port 138 nsew
rlabel metal2 s 330 12049 438 12125 4 gnd
port 138 nsew
rlabel metal2 s 330 10785 438 10861 4 gnd
port 138 nsew
rlabel metal2 s 330 12585 438 12695 4 gnd
port 138 nsew
rlabel metal2 s 330 7845 438 7955 4 gnd
port 138 nsew
rlabel metal2 s 330 13629 438 13705 4 gnd
port 138 nsew
rlabel metal2 s 330 3895 438 4005 4 gnd
port 138 nsew
rlabel metal2 s 330 9205 438 9281 4 gnd
port 138 nsew
rlabel metal2 s 330 9425 438 9535 4 gnd
port 138 nsew
rlabel metal2 s 330 20485 438 20595 4 gnd
port 138 nsew
rlabel metal2 s 330 19949 438 20025 4 gnd
port 138 nsew
rlabel metal2 s 330 13375 438 13485 4 gnd
port 138 nsew
rlabel metal2 s 330 3105 438 3215 4 gnd
port 138 nsew
rlabel metal2 s 330 14735 438 14811 4 gnd
port 138 nsew
rlabel metal2 s 330 2095 438 2171 4 gnd
port 138 nsew
rlabel metal2 s 330 8415 438 8491 4 gnd
port 138 nsew
rlabel metal2 s 330 25479 438 25555 4 gnd
port 138 nsew
rlabel metal2 s 330 6045 438 6121 4 gnd
port 138 nsew
rlabel metal2 s 330 16789 438 16865 4 gnd
port 138 nsew
rlabel metal2 s 330 25225 438 25335 4 gnd
port 138 nsew
rlabel metal2 s 330 3359 438 3435 4 gnd
port 138 nsew
rlabel metal2 s 330 15999 438 16075 4 gnd
port 138 nsew
rlabel metal2 s 330 4685 438 4795 4 gnd
port 138 nsew
rlabel metal2 s 330 4465 438 4541 4 gnd
port 138 nsew
rlabel metal2 s 330 11005 438 11115 4 gnd
port 138 nsew
rlabel metal2 s 330 20739 438 20815 4 gnd
port 138 nsew
rlabel metal2 s 330 1779 438 1855 4 gnd
port 138 nsew
rlabel metal2 s 330 12365 438 12441 4 gnd
port 138 nsew
rlabel metal2 s 330 13945 438 14021 4 gnd
port 138 nsew
rlabel metal2 s 330 7055 438 7165 4 gnd
port 138 nsew
rlabel metal2 s 330 18369 438 18445 4 gnd
port 138 nsew
rlabel metal2 s 330 22065 438 22175 4 gnd
port 138 nsew
rlabel metal2 s 330 14955 438 15065 4 gnd
port 138 nsew
rlabel metal2 s 330 17895 438 17971 4 gnd
port 138 nsew
rlabel metal2 s 330 9679 438 9755 4 gnd
port 138 nsew
rlabel metal2 s 330 10215 438 10325 4 gnd
port 138 nsew
rlabel metal2 s 330 23425 438 23501 4 gnd
port 138 nsew
rlabel metal2 s 330 17579 438 17655 4 gnd
port 138 nsew
rlabel metal2 s 330 21275 438 21385 4 gnd
port 138 nsew
rlabel metal2 s 330 21055 438 21131 4 gnd
port 138 nsew
rlabel metal2 s 330 10469 438 10545 4 gnd
port 138 nsew
rlabel metal2 s 330 20265 438 20341 4 gnd
port 138 nsew
rlabel metal2 s 330 16535 438 16645 4 gnd
port 138 nsew
rlabel metal2 s 330 2569 438 2645 4 gnd
port 138 nsew
rlabel metal2 s 330 26269 438 26345 4 gnd
port 138 nsew
rlabel metal2 s 330 24689 438 24765 4 gnd
port 138 nsew
rlabel metal2 s 330 24215 438 24291 4 gnd
port 138 nsew
rlabel metal2 s 330 7309 438 7385 4 gnd
port 138 nsew
rlabel metal2 s 330 3675 438 3751 4 gnd
port 138 nsew
rlabel metal2 s 330 12839 438 12915 4 gnd
port 138 nsew
rlabel metal2 s 330 6265 438 6375 4 gnd
port 138 nsew
rlabel metal2 s 330 19159 438 19235 4 gnd
port 138 nsew
rlabel metal2 s 330 8889 438 8965 4 gnd
port 138 nsew
rlabel metal2 s 330 2315 438 2425 4 gnd
port 138 nsew
rlabel metal2 s 330 25795 438 25871 4 gnd
port 138 nsew
rlabel metal2 s 330 1525 438 1635 4 gnd
port 138 nsew
rlabel metal2 s 330 735 438 845 4 gnd
port 138 nsew
rlabel metal2 s 330 22855 438 22965 4 gnd
port 138 nsew
rlabel metal2 s 330 5729 438 5805 4 gnd
port 138 nsew
rlabel metal2 s 330 15209 438 15285 4 gnd
port 138 nsew
rlabel metal2 s 330 8635 438 8745 4 gnd
port 138 nsew
rlabel metal2 s 330 23899 438 23975 4 gnd
port 138 nsew
rlabel metal2 s 330 6519 438 6595 4 gnd
port 138 nsew
rlabel metal2 s 330 7625 438 7701 4 gnd
port 138 nsew
rlabel metal2 s 330 9995 438 10071 4 gnd
port 138 nsew
rlabel metal2 s 330 18905 438 19015 4 gnd
port 138 nsew
rlabel metal2 s 330 22319 438 22395 4 gnd
port 138 nsew
<< properties >>
string FIXED_BBOX 0 0 624 26860
<< end >>
