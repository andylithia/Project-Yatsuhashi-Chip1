* NGSPICE file created from captune_flat.ext - technology: sky130B

.subckt captune_flat
X0 BOT_C1 G1 BOT SUB sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=5.656e+12p ps=4.264e+07u w=5.05e+06u l=150000u
X1 BOT G4 BOT_C4 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.828e+12p ps=2.132e+07u w=5.05e+06u l=150000u
X2 BOT G1 BOT_C1 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 TOP BOT_C4 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=4e+06u
X4 BOT_C2 G2 BOT SUB sky130_fd_pr__nfet_01v8 ad=2.828e+12p pd=2.132e+07u as=0p ps=0u w=5.05e+06u l=150000u
X5 TOP BOT_C8 sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=8e+06u
X6 BOT G8 BOT_C8 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.828e+12p ps=2.132e+07u w=5.05e+06u l=150000u
X7 TOP BOT_C2 sky130_fd_pr__cap_mim_m3_1 l=4e+06u w=2.5e+06u
X8 TOP BOT_C1 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2.5e+06u
X9 BOT_C8 G8 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X10 BOT G2 BOT_C2 SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X11 BOT_C4 G4 BOT SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
C0 BOT BOT_C4 3.59fF
C1 TOP BOT_C4 2.51fF
C2 BOT_C2 BOT 3.54fF
C3 BOT_C2 TOP 1.67fF
C4 BOT BOT_C1 3.56fF
C5 BOT BOT_C8 4.38fF
C6 TOP BOT_C1 1.07fF
C7 BOT_C8 TOP 4.54fF
C8 TOP SUB 2.43fF
C9 BOT_C4 SUB 3.66fF
C10 BOT_C8 SUB 3.70fF
C11 BOT_C1 SUB 3.00fF
C12 BOT_C2 SUB 3.19fF
.ends

