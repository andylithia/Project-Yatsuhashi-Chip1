magic
tech sky130B
timestamp 1662579390
<< nwell >>
rect -569 -718 569 718
<< pwell >>
rect -638 718 638 787
rect -638 -718 -569 718
rect 569 -718 638 718
rect -638 -787 638 -718
<< psubdiff >>
rect -620 752 -572 769
rect 572 752 620 769
rect -620 721 -603 752
rect 603 721 620 752
rect -620 -752 -603 -721
rect 603 -752 620 -721
rect -620 -769 -572 -752
rect 572 -769 620 -752
<< nsubdiff >>
rect -551 683 -503 700
rect 503 683 551 700
rect -551 652 -534 683
rect 534 652 551 683
rect -551 415 -534 446
rect 534 415 551 446
rect -551 398 -503 415
rect 503 398 551 415
rect -551 317 -503 334
rect 503 317 551 334
rect -551 286 -534 317
rect 534 286 551 317
rect -551 49 -534 80
rect 534 49 551 80
rect -551 32 -503 49
rect 503 32 551 49
rect -551 -49 -503 -32
rect 503 -49 551 -32
rect -551 -80 -534 -49
rect 534 -80 551 -49
rect -551 -317 -534 -286
rect 534 -317 551 -286
rect -551 -334 -503 -317
rect 503 -334 551 -317
rect -551 -415 -503 -398
rect 503 -415 551 -398
rect -551 -446 -534 -415
rect 534 -446 551 -415
rect -551 -683 -534 -652
rect 534 -683 551 -652
rect -551 -700 -503 -683
rect 503 -700 551 -683
<< psubdiffcont >>
rect -572 752 572 769
rect -620 -721 -603 721
rect 603 -721 620 721
rect -572 -769 572 -752
<< nsubdiffcont >>
rect -503 683 503 700
rect -551 446 -534 652
rect 534 446 551 652
rect -503 398 503 415
rect -503 317 503 334
rect -551 80 -534 286
rect 534 80 551 286
rect -503 32 503 49
rect -503 -49 503 -32
rect -551 -286 -534 -80
rect 534 -286 551 -80
rect -503 -334 503 -317
rect -503 -415 503 -398
rect -551 -652 -534 -446
rect 534 -652 551 -446
rect -503 -700 503 -683
<< pdiode >>
rect -500 643 500 649
rect -500 455 -494 643
rect 494 455 500 643
rect -500 449 500 455
rect -500 277 500 283
rect -500 89 -494 277
rect 494 89 500 277
rect -500 83 500 89
rect -500 -89 500 -83
rect -500 -277 -494 -89
rect 494 -277 500 -89
rect -500 -283 500 -277
rect -500 -455 500 -449
rect -500 -643 -494 -455
rect 494 -643 500 -455
rect -500 -649 500 -643
<< pdiodec >>
rect -494 455 494 643
rect -494 89 494 277
rect -494 -277 494 -89
rect -494 -643 494 -455
<< locali >>
rect -620 752 -572 769
rect 572 752 620 769
rect -620 721 -603 752
rect 603 721 620 752
rect -551 683 -503 700
rect 503 683 551 700
rect -551 652 -534 683
rect 534 652 551 683
rect -502 455 -494 643
rect 494 455 502 643
rect -551 415 -534 446
rect 534 415 551 446
rect -551 398 -503 415
rect 503 398 551 415
rect -551 317 -503 334
rect 503 317 551 334
rect -551 286 -534 317
rect 534 286 551 317
rect -502 89 -494 277
rect 494 89 502 277
rect -551 49 -534 80
rect 534 49 551 80
rect -551 32 -503 49
rect 503 32 551 49
rect -551 -49 -503 -32
rect 503 -49 551 -32
rect -551 -80 -534 -49
rect 534 -80 551 -49
rect -502 -277 -494 -89
rect 494 -277 502 -89
rect -551 -317 -534 -286
rect 534 -317 551 -286
rect -551 -334 -503 -317
rect 503 -334 551 -317
rect -551 -415 -503 -398
rect 503 -415 551 -398
rect -551 -446 -534 -415
rect 534 -446 551 -415
rect -502 -643 -494 -455
rect 494 -643 502 -455
rect -551 -683 -534 -652
rect 534 -683 551 -652
rect -551 -700 -503 -683
rect 503 -700 551 -683
rect -620 -752 -603 -721
rect 603 -752 620 -721
rect -620 -769 -572 -752
rect 572 -769 620 -752
<< viali >>
rect -494 455 494 643
rect -494 89 494 277
rect -494 -277 494 -89
rect -494 -643 494 -455
<< metal1 >>
rect -500 643 500 646
rect -500 455 -494 643
rect 494 455 500 643
rect -500 452 500 455
rect -500 277 500 280
rect -500 89 -494 277
rect 494 89 500 277
rect -500 86 500 89
rect -500 -89 500 -86
rect -500 -277 -494 -89
rect 494 -277 500 -89
rect -500 -280 500 -277
rect -500 -455 500 -452
rect -500 -643 -494 -455
rect 494 -643 500 -455
rect -500 -646 500 -643
<< properties >>
string FIXED_BBOX -542 406 542 691
string gencell sky130_fd_pr__diode_pd2nw_05v5
string library sky130
string parameters w 10 l 2 area 20.0 peri 24.0 nx 1 ny 4 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
