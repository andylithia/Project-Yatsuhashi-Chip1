magic
tech sky130B
magscale 1 2
timestamp 1659629293
<< locali >>
rect -20 -2 1780 20
rect -20 -48 -8 -2
rect 1768 -48 1780 -2
rect -20 -50 1780 -48
<< viali >>
rect -8 -48 1768 -2
<< metal1 >>
rect 268 1055 342 1064
rect 268 1040 277 1055
rect 220 999 277 1040
rect 333 1040 342 1055
rect 463 1055 531 1061
rect 463 1040 469 1055
rect 333 999 469 1040
rect 525 1040 531 1055
rect 655 1055 723 1061
rect 655 1040 661 1055
rect 525 999 661 1040
rect 717 1040 723 1055
rect 847 1055 915 1061
rect 847 1040 853 1055
rect 717 999 853 1040
rect 909 1040 915 1055
rect 1039 1055 1107 1061
rect 1039 1040 1045 1055
rect 909 999 1045 1040
rect 1101 1040 1107 1055
rect 1231 1055 1299 1061
rect 1231 1040 1237 1055
rect 1101 999 1237 1040
rect 1293 1040 1299 1055
rect 1423 1055 1491 1061
rect 1423 1040 1429 1055
rect 1293 999 1429 1040
rect 1485 1040 1491 1055
rect 1615 1055 1683 1061
rect 1615 1040 1621 1055
rect 1485 999 1621 1040
rect 1677 999 1683 1055
rect 220 990 1640 999
rect 82 951 146 957
rect 82 163 88 951
rect 140 163 146 951
rect 82 157 146 163
rect 178 951 242 957
rect 178 163 184 951
rect 236 163 242 951
rect 178 157 242 163
rect 274 951 338 957
rect 274 163 280 951
rect 332 163 338 951
rect 274 157 338 163
rect 370 951 434 957
rect 370 163 376 951
rect 428 163 434 951
rect 370 157 434 163
rect 466 951 530 957
rect 466 163 472 951
rect 524 163 530 951
rect 466 157 530 163
rect 562 951 626 957
rect 562 163 568 951
rect 620 163 626 951
rect 562 157 626 163
rect 658 951 722 957
rect 658 163 664 951
rect 716 163 722 951
rect 658 157 722 163
rect 754 951 818 957
rect 754 163 760 951
rect 812 163 818 951
rect 754 157 818 163
rect 850 951 914 957
rect 850 163 856 951
rect 908 163 914 951
rect 850 157 914 163
rect 946 951 1010 957
rect 946 163 952 951
rect 1004 163 1010 951
rect 946 157 1010 163
rect 1042 951 1106 957
rect 1042 163 1048 951
rect 1100 163 1106 951
rect 1042 157 1106 163
rect 1138 951 1202 957
rect 1138 163 1144 951
rect 1196 163 1202 951
rect 1138 157 1202 163
rect 1234 951 1298 957
rect 1234 163 1240 951
rect 1292 163 1298 951
rect 1234 157 1298 163
rect 1330 951 1394 957
rect 1330 163 1336 951
rect 1388 163 1394 951
rect 1330 157 1394 163
rect 1426 951 1490 957
rect 1426 163 1432 951
rect 1484 163 1490 951
rect 1426 157 1490 163
rect 1522 951 1586 957
rect 1522 163 1528 951
rect 1580 163 1586 951
rect 1522 157 1586 163
rect 1618 951 1682 957
rect 1618 163 1624 951
rect 1676 163 1682 951
rect 1618 157 1682 163
rect 129 106 1600 120
rect 129 60 180 106
rect 170 50 180 60
rect 236 60 380 106
rect 236 50 245 60
rect 370 50 380 60
rect 436 60 570 106
rect 436 50 445 60
rect 560 50 570 60
rect 626 60 760 106
rect 626 50 635 60
rect 750 50 760 60
rect 816 60 950 106
rect 816 50 825 60
rect 940 50 950 60
rect 1006 60 1140 106
rect 1006 50 1015 60
rect 1130 50 1140 60
rect 1196 60 1330 106
rect 1196 50 1205 60
rect 1320 50 1330 60
rect 1386 60 1530 106
rect 1386 50 1395 60
rect 1520 50 1530 60
rect 1586 60 1600 106
rect 1586 50 1595 60
rect 171 41 245 50
rect 371 41 445 50
rect 561 41 635 50
rect 751 41 825 50
rect 941 41 1015 50
rect 1131 41 1205 50
rect 1321 41 1395 50
rect 1521 41 1595 50
rect -20 -2 1780 10
rect -20 -54 -8 -2
rect 1768 -54 1780 -2
rect -20 -60 1780 -54
<< via1 >>
rect 277 999 333 1055
rect 469 999 525 1055
rect 661 999 717 1055
rect 853 999 909 1055
rect 1045 999 1101 1055
rect 1237 999 1293 1055
rect 1429 999 1485 1055
rect 1621 999 1677 1055
rect 88 163 140 951
rect 184 163 236 951
rect 280 163 332 951
rect 376 163 428 951
rect 472 163 524 951
rect 568 163 620 951
rect 664 163 716 951
rect 760 163 812 951
rect 856 163 908 951
rect 952 163 1004 951
rect 1048 163 1100 951
rect 1144 163 1196 951
rect 1240 163 1292 951
rect 1336 163 1388 951
rect 1432 163 1484 951
rect 1528 163 1580 951
rect 1624 163 1676 951
rect 180 50 236 106
rect 380 50 436 106
rect 570 50 626 106
rect 760 50 816 106
rect 950 50 1006 106
rect 1140 50 1196 106
rect 1330 50 1386 106
rect 1530 50 1586 106
rect -8 -48 1768 -2
rect -8 -54 1768 -48
<< metal2 >>
rect 178 1092 242 1122
rect 370 1092 434 1122
rect 562 1092 626 1122
rect 754 1092 818 1122
rect 946 1092 1010 1122
rect 1138 1092 1202 1122
rect 1330 1092 1394 1122
rect 178 962 240 1092
rect 268 1055 342 1064
rect 268 999 277 1055
rect 333 999 342 1055
rect 268 990 342 999
rect 370 962 432 1092
rect 460 1055 534 1064
rect 460 999 469 1055
rect 525 999 534 1055
rect 460 990 534 999
rect 562 962 624 1092
rect 652 1055 726 1064
rect 652 999 661 1055
rect 717 999 726 1055
rect 652 990 726 999
rect 754 962 816 1092
rect 844 1055 918 1064
rect 844 999 853 1055
rect 909 999 918 1055
rect 844 990 918 999
rect 946 962 1008 1092
rect 1036 1055 1110 1064
rect 1036 999 1045 1055
rect 1101 999 1110 1055
rect 1036 990 1110 999
rect 1138 962 1200 1092
rect 1228 1055 1302 1064
rect 1228 999 1237 1055
rect 1293 999 1302 1055
rect 1228 990 1302 999
rect 1330 962 1392 1092
rect 1420 1055 1494 1064
rect 1420 999 1429 1055
rect 1485 999 1494 1055
rect 1420 990 1494 999
rect 1612 1055 1686 1064
rect 1612 999 1621 1055
rect 1677 999 1686 1055
rect 1612 990 1686 999
rect 82 951 146 957
rect 82 163 88 951
rect 140 163 146 951
rect 82 160 146 163
rect 178 951 242 962
rect 178 163 184 951
rect 236 163 242 951
rect 82 10 140 160
rect 178 157 242 163
rect 274 951 338 957
rect 274 163 280 951
rect 332 163 338 951
rect 171 106 245 115
rect 171 50 180 106
rect 236 50 245 106
rect 171 41 245 50
rect 274 10 338 163
rect 370 951 434 962
rect 370 163 376 951
rect 428 163 434 951
rect 370 157 434 163
rect 466 951 530 957
rect 466 163 472 951
rect 524 163 530 951
rect 466 150 530 163
rect 562 951 626 962
rect 562 163 568 951
rect 620 163 626 951
rect 562 157 626 163
rect 658 951 722 957
rect 658 163 664 951
rect 716 163 722 951
rect 658 150 722 163
rect 754 951 818 962
rect 754 163 760 951
rect 812 163 818 951
rect 754 157 818 163
rect 850 951 914 957
rect 850 163 856 951
rect 908 163 914 951
rect 850 150 914 163
rect 946 951 1010 962
rect 946 163 952 951
rect 1004 163 1010 951
rect 946 157 1010 163
rect 1042 951 1106 957
rect 1042 163 1048 951
rect 1100 163 1106 951
rect 1042 150 1106 163
rect 1138 951 1202 962
rect 1138 163 1144 951
rect 1196 163 1202 951
rect 1138 157 1202 163
rect 1234 951 1298 957
rect 1234 163 1240 951
rect 1292 163 1298 951
rect 1234 150 1298 163
rect 1330 951 1394 962
rect 1330 163 1336 951
rect 1388 163 1394 951
rect 1330 157 1394 163
rect 1426 951 1490 957
rect 1426 163 1432 951
rect 1484 163 1490 951
rect 371 106 445 115
rect 371 50 380 106
rect 436 50 445 106
rect 371 41 445 50
rect 473 10 530 150
rect 561 106 635 115
rect 561 50 570 106
rect 626 50 635 106
rect 561 41 635 50
rect 670 10 722 150
rect 751 106 825 115
rect 751 50 760 106
rect 816 50 825 106
rect 751 41 825 50
rect 860 10 910 150
rect 941 106 1015 115
rect 941 50 950 106
rect 1006 50 1015 106
rect 941 41 1015 50
rect 1050 10 1100 150
rect 1131 106 1205 115
rect 1131 50 1140 106
rect 1196 50 1205 106
rect 1131 41 1205 50
rect 1234 10 1290 150
rect 1321 106 1395 115
rect 1321 50 1330 106
rect 1386 50 1395 106
rect 1321 41 1395 50
rect 1426 10 1490 163
rect 1522 951 1586 957
rect 1522 163 1528 951
rect 1580 163 1586 951
rect 1522 157 1586 163
rect 1618 951 1682 957
rect 1618 163 1624 951
rect 1676 163 1682 951
rect 1618 150 1682 163
rect 1521 106 1595 115
rect 1521 50 1530 106
rect 1586 50 1595 106
rect 1521 41 1595 50
rect 1630 10 1682 150
rect -20 -2 1780 10
rect -20 -54 -8 -2
rect 1768 -54 1780 -2
rect -20 -60 1780 -54
<< via2 >>
rect 277 999 333 1055
rect 469 999 525 1055
rect 661 999 717 1055
rect 853 999 909 1055
rect 1045 999 1101 1055
rect 1237 999 1293 1055
rect 1429 999 1485 1055
rect 1621 999 1677 1055
rect 180 50 236 106
rect 380 50 436 106
rect 570 50 626 106
rect 760 50 816 106
rect 950 50 1006 106
rect 1140 50 1196 106
rect 1330 50 1386 106
rect 1530 50 1586 106
<< metal3 >>
rect 268 1055 1686 1064
rect 268 999 277 1055
rect 333 999 469 1055
rect 525 999 661 1055
rect 717 999 853 1055
rect 909 999 1045 1055
rect 1101 999 1237 1055
rect 1293 999 1429 1055
rect 1485 999 1621 1055
rect 1677 999 1686 1055
rect 268 990 1686 999
rect 170 106 1600 120
rect 170 50 180 106
rect 236 50 380 106
rect 436 50 570 106
rect 626 50 760 106
rect 816 50 950 106
rect 1006 50 1140 106
rect 1196 50 1330 106
rect 1386 50 1530 106
rect 1586 50 1600 106
rect 170 40 1600 50
use sky130_fd_pr__nfet_01v8_7RL2PV  sky130_fd_pr__nfet_01v8_7RL2PV_0
timestamp 1659585137
transform 1 0 882 0 1 557
box -935 -610 935 610
<< end >>
