magic
tech sky130A
magscale 1 2
timestamp 1664325575
<< error_s >>
rect 5100 5789 5191 5800
rect 3020 800 3145 820
rect 3215 800 3461 820
rect 3531 800 3777 820
rect 3847 800 4093 820
rect 4163 800 4409 820
rect 4479 800 4725 820
rect 4795 800 5041 820
rect 15620 800 15657 820
rect 15903 800 15973 820
rect 16219 800 16289 820
rect 16535 800 16606 820
rect 16851 800 16921 820
rect 17167 800 17237 820
rect 17483 800 17553 820
rect 1560 720 1565 740
rect 1635 720 1881 740
rect 1951 720 2197 740
rect 2267 720 2513 740
rect 2583 720 2829 740
rect 2899 720 3145 740
rect 3215 720 3461 740
rect 3531 720 3777 740
rect 3847 720 4093 740
rect 4163 720 4409 740
rect 4479 720 4725 740
rect 4795 720 5041 740
rect 11419 720 11657 740
rect 11727 720 11973 740
rect 12043 720 12289 740
rect 12359 720 12605 740
rect 12675 720 12680 740
rect 14160 720 14165 740
rect 14235 720 14481 740
rect 14551 720 14797 740
rect 14867 720 15113 740
rect 15183 720 15429 740
rect 15499 720 15580 740
rect 24019 720 24257 740
rect 24327 720 24573 740
rect 24643 720 24889 740
rect 24959 720 25205 740
rect 25275 720 25280 740
rect 1560 340 3100 360
rect 5000 340 6380 360
rect 7860 340 12680 360
rect 14160 340 15700 360
rect 17600 340 18980 360
rect 20460 340 25280 360
rect 1500 280 3100 300
rect 5000 280 6440 300
rect 7800 280 12740 300
rect 14100 280 15700 300
rect 17600 280 19040 300
rect 20400 280 25340 300
rect 7780 -750 8023 -731
rect 8093 -750 8339 -731
rect 8409 -750 8655 -731
rect 8725 -750 8971 -731
rect 9041 -750 9280 -731
rect 20380 -750 20623 -731
rect 20693 -750 20939 -731
rect 21009 -750 21255 -731
rect 21325 -750 21571 -731
rect 21641 -750 21880 -731
rect 1663 -751 1853 -750
rect 1979 -751 2169 -750
rect 2295 -751 2485 -750
rect 2611 -751 2801 -750
rect 2927 -751 3117 -750
rect 5139 -751 5329 -750
rect 5455 -751 5645 -750
rect 5771 -751 5961 -750
rect 6087 -751 6277 -750
rect 7780 -751 9417 -750
rect 9543 -751 9733 -750
rect 9859 -751 10049 -750
rect 10175 -751 10365 -750
rect 10491 -751 10681 -750
rect 10807 -751 10997 -750
rect 11123 -751 11313 -750
rect 11439 -751 11629 -750
rect 11755 -751 11945 -750
rect 12071 -751 12261 -750
rect 12387 -751 12577 -750
rect 14263 -751 14453 -750
rect 14579 -751 14769 -750
rect 14895 -751 15085 -750
rect 15211 -751 15401 -750
rect 15527 -751 15717 -750
rect 17739 -751 17929 -750
rect 18055 -751 18245 -750
rect 18371 -751 18561 -750
rect 18687 -751 18877 -750
rect 20380 -751 22017 -750
rect 22143 -751 22333 -750
rect 22459 -751 22649 -750
rect 22775 -751 22965 -750
rect 23091 -751 23281 -750
rect 23407 -751 23597 -750
rect 23723 -751 23913 -750
rect 24039 -751 24229 -750
rect 24355 -751 24545 -750
rect 24671 -751 24861 -750
rect 24987 -751 25177 -750
rect 1500 -800 3117 -751
rect 5000 -800 6440 -751
rect 7780 -800 12740 -751
rect 14100 -800 15717 -751
rect 17600 -800 19040 -751
rect 20380 -800 25340 -751
rect 1723 -811 1793 -810
rect 2039 -811 2109 -810
rect 2355 -811 2425 -810
rect 2671 -811 2741 -810
rect 2987 -811 3057 -810
rect 3100 -811 3117 -800
rect 5199 -811 5269 -810
rect 5515 -811 5585 -810
rect 5831 -811 5901 -810
rect 6147 -811 6217 -810
rect 8023 -811 8093 -810
rect 8339 -811 8409 -810
rect 8655 -811 8725 -810
rect 8971 -811 9041 -810
rect 9287 -811 9357 -810
rect 9603 -811 9673 -810
rect 9919 -811 9989 -810
rect 10235 -811 10305 -810
rect 10551 -811 10621 -810
rect 10867 -811 10937 -810
rect 11183 -811 11253 -810
rect 11499 -811 11569 -810
rect 11815 -811 11885 -810
rect 12131 -811 12201 -810
rect 12447 -811 12517 -810
rect 14323 -811 14393 -810
rect 14639 -811 14709 -810
rect 14955 -811 15025 -810
rect 15271 -811 15341 -810
rect 15587 -811 15657 -810
rect 15700 -811 15717 -800
rect 17799 -811 17869 -810
rect 18115 -811 18185 -810
rect 18431 -811 18501 -810
rect 18747 -811 18817 -810
rect 20623 -811 20693 -810
rect 20939 -811 21009 -810
rect 21255 -811 21325 -810
rect 21571 -811 21641 -810
rect 21887 -811 21957 -810
rect 22203 -811 22273 -810
rect 22519 -811 22589 -810
rect 22835 -811 22905 -810
rect 23151 -811 23221 -810
rect 23467 -811 23537 -810
rect 23783 -811 23853 -810
rect 24099 -811 24169 -810
rect 24415 -811 24485 -810
rect 24731 -811 24801 -810
rect 25047 -811 25117 -810
rect 1560 -860 3100 -811
rect 5000 -860 6380 -811
rect 7860 -860 12680 -811
rect 14160 -860 15700 -811
rect 17600 -860 18980 -811
rect 20460 -860 25280 -811
rect 3145 -1291 3215 -1280
rect 5041 -1291 5080 -1280
rect 15745 -1291 15815 -1280
rect 17641 -1291 17680 -1280
rect 1635 -6280 1881 -6260
rect 1951 -6280 2197 -6260
rect 2267 -6280 2513 -6260
rect 2583 -6280 2829 -6260
rect 2899 -6280 3145 -6260
rect 3215 -6280 3461 -6260
rect 3531 -6280 3777 -6260
rect 3847 -6280 4093 -6260
rect 4163 -6280 4409 -6260
rect 4479 -6280 4725 -6260
rect 4795 -6280 5041 -6260
rect 5111 -6280 5357 -6260
rect 5427 -6280 5673 -6260
rect 5743 -6280 5989 -6260
rect 6059 -6280 6305 -6260
rect 6375 -6280 6380 -6260
rect 7935 -6280 8181 -6260
rect 8251 -6280 8497 -6260
rect 8567 -6280 8813 -6260
rect 8883 -6280 9129 -6260
rect 9199 -6280 9445 -6260
rect 9515 -6280 9761 -6260
rect 9831 -6280 10077 -6260
rect 10147 -6280 10393 -6260
rect 10463 -6280 10709 -6260
rect 10779 -6280 11025 -6260
rect 11095 -6280 11341 -6260
rect 11411 -6280 11657 -6260
rect 11727 -6280 11973 -6260
rect 12043 -6280 12289 -6260
rect 12359 -6280 12605 -6260
rect 12675 -6280 12680 -6260
rect 17719 -6280 17957 -6260
rect 18027 -6280 18273 -6260
rect 18343 -6280 18589 -6260
rect 18659 -6280 18905 -6260
rect 18975 -6280 18980 -6260
rect 20460 -6280 20465 -6260
rect 20535 -6280 20781 -6260
rect 20851 -6280 21097 -6260
rect 21167 -6280 21413 -6260
rect 21483 -6280 21729 -6260
rect 21799 -6280 22045 -6260
rect 22115 -6280 22361 -6260
rect 22431 -6280 22677 -6260
rect 22747 -6280 22993 -6260
rect 23063 -6280 23309 -6260
rect 23379 -6280 23625 -6260
rect 23695 -6280 23941 -6260
rect 24011 -6280 24257 -6260
rect 24327 -6280 24573 -6260
rect 24643 -6280 24889 -6260
rect 24959 -6280 25205 -6260
rect 25275 -6280 25280 -6260
<< metal2 >>
rect 6500 6100 7800 6500
rect 12800 6200 14100 6600
rect 19100 6100 20400 6500
rect 6500 5500 7800 5900
rect 12800 5600 14100 6000
rect 19100 5500 20400 5900
rect 6500 4900 7800 5300
rect 12800 5000 14100 5400
rect 19100 4900 20400 5300
rect 6500 4300 7800 4700
rect 12800 4400 14100 4800
rect 19100 4300 20400 4700
rect 6500 3700 7800 4100
rect 12800 3800 14100 4200
rect 19100 3700 20400 4100
rect 6500 3100 7800 3500
rect 12800 3200 14100 3600
rect 19100 3100 20400 3500
rect 6500 2500 7800 2900
rect 12800 2600 14100 3000
rect 19100 2500 20400 2900
rect 6500 1900 7800 2300
rect 12800 2000 14100 2400
rect 19100 1900 20400 2300
rect 6500 1300 7800 1700
rect 12800 1400 14100 1800
rect 19100 1300 20400 1700
rect 6500 700 7800 1100
rect 12800 800 14100 1200
rect 19100 700 20400 1100
rect 6500 100 7800 500
rect 12800 200 14100 600
rect 6900 -500 7400 100
rect 13200 -500 13700 200
rect 19100 100 20400 500
rect 19500 -500 20000 100
rect 6500 -900 7800 -500
rect 12800 -900 14100 -500
rect 19100 -900 20400 -500
rect 6500 -1500 7800 -1100
rect 12800 -1500 14100 -1100
rect 19100 -1500 20400 -1100
rect 6500 -2100 7800 -1700
rect 12800 -2100 14100 -1700
rect 19100 -2100 20400 -1700
rect 6500 -2700 7800 -2300
rect 12800 -2700 14100 -2300
rect 19100 -2700 20400 -2300
rect 6500 -3300 7800 -2900
rect 12800 -3300 14100 -2900
rect 19100 -3300 20400 -2900
rect 6500 -3900 7800 -3500
rect 12800 -3900 14100 -3500
rect 19100 -3900 20400 -3500
rect 6500 -4500 7800 -4100
rect 12800 -4500 14100 -4100
rect 19100 -4500 20400 -4100
rect 6500 -5100 7800 -4700
rect 12800 -5100 14100 -4700
rect 19100 -5100 20400 -4700
rect 6500 -5700 7800 -5300
rect 12800 -5700 14100 -5300
rect 19100 -5700 20400 -5300
rect 6500 -6300 7800 -5900
rect 12800 -6300 14100 -5900
rect 19100 -6300 20400 -5900
rect 6500 -6900 7800 -6500
rect 12800 -6900 14100 -6500
rect 19100 -6900 20400 -6500
<< metal3 >>
rect 1400 5700 5100 5800
rect 1400 3900 1500 5700
rect 2800 3900 5100 5700
rect 1400 3800 5100 3900
rect 7700 5700 9200 5800
rect 7700 3900 7800 5700
rect 9000 3900 9200 5700
rect 7700 3800 9200 3900
rect 14000 5700 15500 5800
rect 14000 3900 14100 5700
rect 15400 3900 15500 5700
rect 14000 3800 15500 3900
rect 20300 5700 21800 5800
rect 20300 3900 20400 5700
rect 21600 3900 21800 5700
rect 20300 3800 21800 3900
rect 1400 2700 5100 2800
rect 1400 900 1500 2700
rect 2800 900 5100 2700
rect 1400 800 5100 900
rect 11500 2700 13000 2800
rect 11500 900 11600 2700
rect 12900 900 13000 2700
rect 11500 800 13000 900
rect 14000 2700 15500 2800
rect 14000 900 14100 2700
rect 15400 900 15500 2700
rect 14000 800 15500 900
rect 24100 2700 25600 2800
rect 24100 900 24200 2700
rect 25500 900 25600 2700
rect 24100 800 25600 900
rect 3100 400 5000 500
rect 3100 300 3300 400
rect 1400 100 3300 300
rect 4800 300 5000 400
rect 15700 400 17600 500
rect 15700 300 15900 400
rect 4800 180 7400 300
rect 4800 100 7020 180
rect 1400 20 7020 100
rect 7380 20 7400 180
rect 1400 0 7400 20
rect 7600 180 13700 300
rect 7600 20 13320 180
rect 13680 20 13700 180
rect 7600 0 13700 20
rect 13900 100 15900 300
rect 17400 300 17600 400
rect 17400 180 20000 300
rect 17400 100 19620 180
rect 13900 20 19620 100
rect 19980 20 20000 180
rect 13900 0 20000 20
rect 20200 0 25400 300
rect 7600 -200 7900 0
rect 9400 -100 12000 0
rect 13900 -100 14100 0
rect 20200 -100 20500 0
rect 22000 -100 24600 0
rect 6500 -400 7900 -200
rect 12800 -300 14100 -100
rect 19100 -300 20500 -100
rect 3100 -500 5000 -400
rect 6500 -500 6800 -400
rect 9400 -500 12000 -400
rect 12800 -500 13100 -300
rect 15700 -500 17600 -400
rect 19100 -500 19400 -300
rect 22000 -500 24600 -400
rect 1400 -800 3300 -500
rect 4800 -800 6800 -500
rect 7000 -520 13100 -500
rect 7000 -680 7020 -520
rect 7380 -680 13100 -520
rect 7000 -800 13100 -680
rect 13300 -520 15900 -500
rect 13300 -680 13320 -520
rect 13680 -680 15900 -520
rect 13300 -800 15900 -680
rect 17400 -800 19400 -500
rect 19600 -520 25400 -500
rect 19600 -680 19620 -520
rect 19980 -680 25400 -520
rect 19600 -800 25400 -680
rect 3100 -900 5000 -800
rect 15700 -900 17600 -800
rect 3300 -1300 4800 -1200
rect 3300 -3100 3400 -1300
rect 4700 -3100 4800 -1300
rect 3300 -3200 4800 -3100
rect 7700 -1300 9200 -1200
rect 7700 -3100 7800 -1300
rect 9100 -3100 9200 -1300
rect 7700 -3200 9200 -3100
rect 15900 -1300 17400 -1200
rect 15900 -3100 16000 -1300
rect 17300 -3100 17400 -1300
rect 15900 -3200 17400 -3100
rect 20300 -1300 21800 -1200
rect 20300 -3100 20400 -1300
rect 21700 -3100 21800 -1300
rect 20300 -3200 21800 -3100
rect 1600 -4300 6700 -4200
rect 1600 -6100 5300 -4300
rect 6600 -6100 6700 -4300
rect 1600 -6200 6700 -6100
rect 7900 -4300 12800 -4200
rect 7900 -6100 9700 -4300
rect 11000 -6100 12800 -4300
rect 7900 -6200 12800 -6100
rect 17800 -4300 19300 -4200
rect 17800 -6100 17900 -4300
rect 19200 -6100 19300 -4300
rect 17800 -6200 19300 -6100
rect 20300 -4300 25600 -4200
rect 20300 -6100 22300 -4300
rect 23600 -6100 25600 -4300
rect 20300 -6200 25600 -6100
<< via3 >>
rect 1500 3900 2800 5700
rect 7800 3900 9000 5700
rect 14100 3900 15400 5700
rect 20400 3900 21600 5700
rect 1500 900 2800 2700
rect 11600 900 12900 2700
rect 14100 900 15400 2700
rect 24200 900 25500 2700
rect 3300 100 4800 400
rect 7020 20 7380 180
rect 13320 20 13680 180
rect 15900 100 17400 400
rect 19620 20 19980 180
rect 3300 -800 4800 -500
rect 7020 -680 7380 -520
rect 13320 -680 13680 -520
rect 15900 -800 17400 -500
rect 19620 -680 19980 -520
rect 3400 -3100 4700 -1300
rect 7800 -3100 9100 -1300
rect 16000 -3100 17300 -1300
rect 20400 -3100 21700 -1300
rect 5300 -6100 6600 -4300
rect 9700 -6100 11000 -4300
rect 17900 -6100 19200 -4300
rect 22300 -6100 23600 -4300
<< metal4 >>
rect 5200 11100 6700 11200
rect 5200 9500 5300 11100
rect 6600 9500 6700 11100
rect 1400 8000 2900 8200
rect 1400 6600 1600 8000
rect 2800 6600 2900 8000
rect 1400 5700 2900 6600
rect 1400 3900 1500 5700
rect 2800 3900 2900 5700
rect 1400 3800 2900 3900
rect 1400 2700 2900 2800
rect 1400 900 1500 2700
rect 2800 900 2900 2700
rect 1400 -9900 2900 900
rect 3200 400 4900 500
rect 3200 100 3300 400
rect 4800 100 4900 400
rect 3200 0 4900 100
rect 3200 -500 4900 -400
rect 3200 -800 3300 -500
rect 4800 -800 4900 -500
rect 3200 -900 4900 -800
rect 3300 -1300 4800 -1200
rect 3300 -3100 3400 -1300
rect 4700 -3100 4800 -1300
rect 3300 -6900 4800 -3100
rect 5200 -4300 6700 9500
rect 7700 11100 9200 11200
rect 7700 9500 7800 11100
rect 9100 9500 9200 11100
rect 7700 5700 9200 9500
rect 17800 11100 19300 11200
rect 17800 9500 17900 11100
rect 19200 9500 19300 11100
rect 7700 3900 7800 5700
rect 9000 3900 9200 5700
rect 7700 3800 9200 3900
rect 9600 8100 11100 8200
rect 9600 6500 9800 8100
rect 11000 6500 11100 8100
rect 7000 180 7400 200
rect 7000 20 7020 180
rect 7380 20 7400 180
rect 7000 -520 7400 20
rect 7000 -680 7020 -520
rect 7380 -680 7400 -520
rect 7000 -700 7400 -680
rect 5200 -6100 5300 -4300
rect 6600 -6100 6700 -4300
rect 5200 -6200 6700 -6100
rect 7700 -1300 9200 -1200
rect 7700 -3100 7800 -1300
rect 9100 -3100 9200 -1300
rect 3300 -8500 3400 -6900
rect 4700 -8500 4800 -6900
rect 3300 -8600 4800 -8500
rect 1400 -11500 1500 -9900
rect 2800 -11500 2900 -9900
rect 1400 -11600 2900 -11500
rect 7700 -9900 9200 -3100
rect 9600 -4300 11100 6500
rect 14000 8000 15500 8200
rect 14000 6600 14200 8000
rect 15400 6600 15500 8000
rect 14000 5700 15500 6600
rect 14000 3900 14100 5700
rect 15400 3900 15500 5700
rect 14000 3800 15500 3900
rect 9600 -6100 9700 -4300
rect 11000 -6100 11100 -4300
rect 9600 -6200 11100 -6100
rect 11500 2700 13000 2800
rect 11500 900 11600 2700
rect 12900 900 13000 2700
rect 11500 -6900 13000 900
rect 14000 2700 15500 2800
rect 14000 900 14100 2700
rect 15400 900 15500 2700
rect 13300 180 13700 200
rect 13300 20 13320 180
rect 13680 20 13700 180
rect 13300 -520 13700 20
rect 13300 -680 13320 -520
rect 13680 -680 13700 -520
rect 13300 -700 13700 -680
rect 11500 -8500 11600 -6900
rect 12900 -8500 13000 -6900
rect 11500 -8600 13000 -8500
rect 14000 -9900 15500 900
rect 15800 400 17500 500
rect 15800 100 15900 400
rect 17400 100 17500 400
rect 15800 0 17500 100
rect 15800 -500 17500 -400
rect 15800 -800 15900 -500
rect 17400 -800 17500 -500
rect 15800 -900 17500 -800
rect 15900 -1300 17400 -1200
rect 15900 -3100 16000 -1300
rect 17300 -3100 17400 -1300
rect 15900 -6900 17400 -3100
rect 17800 -4300 19300 9500
rect 20300 11100 21800 11200
rect 20300 9500 20400 11100
rect 21700 9500 21800 11100
rect 20300 8200 21800 9500
rect 20300 6600 21900 8200
rect 22200 8100 23700 8200
rect 20300 5700 21800 6600
rect 20300 3900 20400 5700
rect 21600 3900 21800 5700
rect 20300 3800 21800 3900
rect 22200 6500 22400 8100
rect 23600 6500 23700 8100
rect 19600 180 20000 200
rect 19600 20 19620 180
rect 19980 20 20000 180
rect 19600 -520 20000 20
rect 19600 -680 19620 -520
rect 19980 -680 20000 -520
rect 19600 -700 20000 -680
rect 17800 -6100 17900 -4300
rect 19200 -6100 19300 -4300
rect 17800 -6200 19300 -6100
rect 20300 -1300 21800 -1200
rect 20300 -3100 20400 -1300
rect 21700 -3100 21800 -1300
rect 15900 -8500 16000 -6900
rect 17300 -8500 17400 -6900
rect 15900 -8600 17400 -8500
rect 7700 -11500 7800 -9900
rect 9100 -11500 9200 -9900
rect 7700 -11600 9200 -11500
rect 11500 -11500 11600 -9900
rect 12800 -11500 13000 -9900
rect 11500 -11600 13000 -11500
rect 14000 -11500 14100 -9900
rect 15400 -11500 15500 -9900
rect 14000 -11600 15500 -11500
rect 20300 -9900 21800 -3100
rect 22200 -4300 23700 6500
rect 22200 -6100 22300 -4300
rect 23600 -6100 23700 -4300
rect 22200 -6200 23700 -6100
rect 24100 2700 25600 2800
rect 24100 900 24200 2700
rect 25500 900 25600 2700
rect 24100 -6900 25600 900
rect 24100 -8500 24200 -6900
rect 25500 -8500 25600 -6900
rect 24100 -8600 25600 -8500
rect 20300 -11500 20400 -9900
rect 21700 -11500 21800 -9900
rect 20300 -11600 21800 -11500
<< via4 >>
rect 5300 9500 6600 11100
rect 1600 6600 2800 8000
rect 3300 100 4800 400
rect 3300 -800 4800 -500
rect 7800 9500 9100 11100
rect 17900 9500 19200 11100
rect 9800 6500 11000 8100
rect 3400 -8500 4700 -6900
rect 1500 -11500 2800 -9900
rect 14200 6600 15400 8000
rect 11600 -8500 12900 -6900
rect 15900 100 17400 400
rect 15900 -800 17400 -500
rect 20400 9500 21700 11100
rect 22400 6500 23600 8100
rect 16000 -8500 17300 -6900
rect 7800 -11500 9100 -9900
rect 14100 -11500 15400 -9900
rect 24200 -8500 25500 -6900
rect 20400 -11500 21700 -9900
<< metal5 >>
rect 1400 8200 4200 11400
rect 22800 11200 25600 11400
rect 5200 11100 25600 11200
rect 5200 9500 5300 11100
rect 6600 9500 7800 11100
rect 9100 9500 17900 11100
rect 19200 9500 20400 11100
rect 21700 9500 25600 11100
rect 5200 9400 25600 9500
rect 1400 8100 23700 8200
rect 1400 8000 9800 8100
rect 1400 6600 1600 8000
rect 2800 6600 9800 8000
rect 1400 6500 9800 6600
rect 11000 8000 22400 8100
rect 11000 6600 14200 8000
rect 15400 6600 22400 8000
rect 11000 6500 22400 6600
rect 23600 6500 23700 8100
rect 1400 6400 23700 6500
rect 1300 400 25500 500
rect 1300 100 3300 400
rect 4800 100 15900 400
rect 17400 100 25500 400
rect 1300 0 25500 100
rect 1300 -500 25500 -400
rect 1300 -800 3300 -500
rect 4800 -800 15900 -500
rect 17400 -800 25500 -500
rect 1300 -900 25500 -800
rect 3300 -6900 25600 -6800
rect 3300 -8500 3400 -6900
rect 4700 -8500 11600 -6900
rect 12900 -8500 16000 -6900
rect 17300 -8500 24200 -6900
rect 25500 -8500 25600 -6900
rect 3300 -8600 25600 -8500
rect 1400 -9900 21800 -9800
rect 1400 -11500 1500 -9900
rect 2800 -11500 7800 -9900
rect 9100 -11500 14100 -9900
rect 15400 -11500 20400 -9900
rect 21700 -11500 21800 -9900
rect 1400 -11600 21800 -11500
rect 1400 -11800 4200 -11600
rect 22800 -11800 25600 -8600
use ./CLASSE/NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_0 CLASSE
timestamp 1664325575
transform 1 0 1400 0 1 0
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_1
timestamp 1664325575
transform 1 0 7700 0 1 0
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_2
timestamp 1664325575
transform 1 0 14000 0 1 0
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_3
timestamp 1664325575
transform 1 0 20300 0 1 0
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_4
timestamp 1664325575
transform 1 0 20300 0 1 -7000
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_5
timestamp 1664325575
transform 1 0 14000 0 1 -7000
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_6
timestamp 1664325575
transform 1 0 7700 0 1 -7000
box 0 0 5138 6516
use ./CLASSE/NMOS_30_0p5_30_1  NMOS_30_0p5_30_1_7
timestamp 1664325575
transform 1 0 1400 0 1 -7000
box 0 0 5138 6516
<< labels >>
rlabel metal5 1300 0 1400 500 1 GL
rlabel metal5 1300 -900 1400 -400 1 GR
rlabel metal5 1400 -11800 4200 -11600 1 SD2L
rlabel metal5 22800 -11800 25600 -11600 1 SD2R
rlabel metal5 22800 11200 25600 11400 1 SD1R
rlabel metal5 1400 11200 4200 11400 1 SD1L
rlabel metal2 14030 -580 14100 -520 1 SUB
<< end >>
