magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< metal1 >>
rect 2092 5397 2152 5453
rect 3340 5397 3400 5453
rect 4588 5397 4648 5453
rect 5836 5397 5896 5453
rect 7084 5397 7144 5453
rect 8332 5397 8392 5453
rect 9580 5397 9640 5453
rect 10828 5397 10888 5453
rect 12076 5397 12136 5453
rect 13324 5397 13384 5453
rect 14572 5397 14632 5453
rect 15820 5397 15880 5453
rect 17068 5397 17128 5453
rect 18316 5397 18376 5453
rect 19564 5397 19624 5453
rect 20812 5397 20872 5453
rect 22060 5397 22120 5453
rect 23308 5397 23368 5453
rect 24556 5397 24616 5453
rect 25804 5397 25864 5453
rect 27052 5397 27112 5453
rect 28300 5397 28360 5453
rect 29548 5397 29608 5453
rect 30796 5397 30856 5453
rect 0 5335 31073 5363
rect 1996 3380 2024 3446
rect 1949 3352 2024 3380
rect 1949 2946 1977 3352
rect 2198 3300 2226 3446
rect 3244 3380 3272 3446
rect 3197 3352 3272 3380
rect 2198 3272 2441 3300
rect 2413 3070 2441 3272
rect 3197 2946 3225 3352
rect 3446 3300 3474 3446
rect 4492 3380 4520 3446
rect 4445 3352 4520 3380
rect 3446 3272 3689 3300
rect 3661 3070 3689 3272
rect 4445 2946 4473 3352
rect 4694 3300 4722 3446
rect 5740 3380 5768 3446
rect 5693 3352 5768 3380
rect 4694 3272 4937 3300
rect 4909 3070 4937 3272
rect 5693 2946 5721 3352
rect 5942 3300 5970 3446
rect 6988 3380 7016 3446
rect 6941 3352 7016 3380
rect 5942 3272 6185 3300
rect 6157 3070 6185 3272
rect 6941 2946 6969 3352
rect 7190 3300 7218 3446
rect 8236 3380 8264 3446
rect 8189 3352 8264 3380
rect 7190 3272 7433 3300
rect 7405 3070 7433 3272
rect 8189 2946 8217 3352
rect 8438 3300 8466 3446
rect 9484 3380 9512 3446
rect 9437 3352 9512 3380
rect 8438 3272 8681 3300
rect 8653 3070 8681 3272
rect 9437 2946 9465 3352
rect 9686 3300 9714 3446
rect 10732 3380 10760 3446
rect 10685 3352 10760 3380
rect 9686 3272 9929 3300
rect 9901 3070 9929 3272
rect 10685 2946 10713 3352
rect 10934 3300 10962 3446
rect 11980 3380 12008 3446
rect 11933 3352 12008 3380
rect 10934 3272 11177 3300
rect 11149 3070 11177 3272
rect 11933 2946 11961 3352
rect 12182 3300 12210 3446
rect 13228 3380 13256 3446
rect 13181 3352 13256 3380
rect 12182 3272 12425 3300
rect 12397 3070 12425 3272
rect 13181 2946 13209 3352
rect 13430 3300 13458 3446
rect 14476 3380 14504 3446
rect 14429 3352 14504 3380
rect 13430 3272 13673 3300
rect 13645 3070 13673 3272
rect 14429 2946 14457 3352
rect 14678 3300 14706 3446
rect 15724 3380 15752 3446
rect 15677 3352 15752 3380
rect 14678 3272 14921 3300
rect 14893 3070 14921 3272
rect 15677 2946 15705 3352
rect 15926 3300 15954 3446
rect 16972 3380 17000 3446
rect 16925 3352 17000 3380
rect 15926 3272 16169 3300
rect 16141 3070 16169 3272
rect 16925 2946 16953 3352
rect 17174 3300 17202 3446
rect 18220 3380 18248 3446
rect 18173 3352 18248 3380
rect 17174 3272 17417 3300
rect 17389 3070 17417 3272
rect 18173 2946 18201 3352
rect 18422 3300 18450 3446
rect 19468 3380 19496 3446
rect 19421 3352 19496 3380
rect 18422 3272 18665 3300
rect 18637 3070 18665 3272
rect 19421 2946 19449 3352
rect 19670 3300 19698 3446
rect 20716 3380 20744 3446
rect 20669 3352 20744 3380
rect 19670 3272 19913 3300
rect 19885 3070 19913 3272
rect 20669 2946 20697 3352
rect 20918 3300 20946 3446
rect 21964 3380 21992 3446
rect 21917 3352 21992 3380
rect 20918 3272 21161 3300
rect 21133 3070 21161 3272
rect 21917 2946 21945 3352
rect 22166 3300 22194 3446
rect 23212 3380 23240 3446
rect 23165 3352 23240 3380
rect 22166 3272 22409 3300
rect 22381 3070 22409 3272
rect 23165 2946 23193 3352
rect 23414 3300 23442 3446
rect 24460 3380 24488 3446
rect 24413 3352 24488 3380
rect 23414 3272 23657 3300
rect 23629 3070 23657 3272
rect 24413 2946 24441 3352
rect 24662 3300 24690 3446
rect 25708 3380 25736 3446
rect 25661 3352 25736 3380
rect 24662 3272 24905 3300
rect 24877 3070 24905 3272
rect 25661 2946 25689 3352
rect 25910 3300 25938 3446
rect 26956 3380 26984 3446
rect 26909 3352 26984 3380
rect 25910 3272 26153 3300
rect 26125 3070 26153 3272
rect 26909 2946 26937 3352
rect 27158 3300 27186 3446
rect 28204 3380 28232 3446
rect 28157 3352 28232 3380
rect 27158 3272 27401 3300
rect 27373 3070 27401 3272
rect 28157 2946 28185 3352
rect 28406 3300 28434 3446
rect 29452 3380 29480 3446
rect 29405 3352 29480 3380
rect 28406 3272 28649 3300
rect 28621 3070 28649 3272
rect 29405 2946 29433 3352
rect 29654 3300 29682 3446
rect 30700 3380 30728 3446
rect 30653 3352 30728 3380
rect 29654 3272 29897 3300
rect 29869 3070 29897 3272
rect 30653 2946 30681 3352
rect 30902 3300 30930 3446
rect 30902 3272 31145 3300
rect 31117 3070 31145 3272
rect 1949 1192 1977 1258
rect 1935 1164 1977 1192
rect 1311 252 1339 1006
rect 1775 252 1803 1006
rect 1935 252 1963 1164
rect 2413 1112 2441 1258
rect 2399 1084 2441 1112
rect 2545 1112 2573 1258
rect 3009 1192 3037 1258
rect 3197 1192 3225 1258
rect 3009 1164 3051 1192
rect 2545 1084 2587 1112
rect 2399 252 2427 1084
rect 2559 252 2587 1084
rect 3023 252 3051 1164
rect 3183 1164 3225 1192
rect 3183 252 3211 1164
rect 3661 1112 3689 1258
rect 3647 1084 3689 1112
rect 3793 1112 3821 1258
rect 4257 1192 4285 1258
rect 4445 1192 4473 1258
rect 4257 1164 4299 1192
rect 3793 1084 3835 1112
rect 3647 252 3675 1084
rect 3807 252 3835 1084
rect 4271 252 4299 1164
rect 4431 1164 4473 1192
rect 4431 252 4459 1164
rect 4909 1112 4937 1258
rect 4895 1084 4937 1112
rect 5041 1112 5069 1258
rect 5505 1192 5533 1258
rect 5693 1192 5721 1258
rect 5505 1164 5547 1192
rect 5041 1084 5083 1112
rect 4895 252 4923 1084
rect 5055 252 5083 1084
rect 5519 252 5547 1164
rect 5679 1164 5721 1192
rect 5679 252 5707 1164
rect 6157 1112 6185 1258
rect 6143 1084 6185 1112
rect 6289 1112 6317 1258
rect 6753 1192 6781 1258
rect 6941 1192 6969 1258
rect 6753 1164 6795 1192
rect 6289 1084 6331 1112
rect 6143 252 6171 1084
rect 6303 252 6331 1084
rect 6767 252 6795 1164
rect 6927 1164 6969 1192
rect 6927 252 6955 1164
rect 7405 1112 7433 1258
rect 7391 1084 7433 1112
rect 7537 1112 7565 1258
rect 8001 1192 8029 1258
rect 8189 1192 8217 1258
rect 8001 1164 8043 1192
rect 7537 1084 7579 1112
rect 7391 252 7419 1084
rect 7551 252 7579 1084
rect 8015 252 8043 1164
rect 8175 1164 8217 1192
rect 8175 252 8203 1164
rect 8653 1112 8681 1258
rect 8639 1084 8681 1112
rect 8785 1112 8813 1258
rect 9249 1192 9277 1258
rect 9437 1192 9465 1258
rect 9249 1164 9291 1192
rect 8785 1084 8827 1112
rect 8639 252 8667 1084
rect 8799 252 8827 1084
rect 9263 252 9291 1164
rect 9423 1164 9465 1192
rect 9423 252 9451 1164
rect 9901 1112 9929 1258
rect 9887 1084 9929 1112
rect 10033 1112 10061 1258
rect 10497 1192 10525 1258
rect 10685 1192 10713 1258
rect 10497 1164 10539 1192
rect 10033 1084 10075 1112
rect 9887 252 9915 1084
rect 10047 252 10075 1084
rect 10511 252 10539 1164
rect 10671 1164 10713 1192
rect 10671 252 10699 1164
rect 11149 1112 11177 1258
rect 11135 1084 11177 1112
rect 11281 1112 11309 1258
rect 11745 1192 11773 1258
rect 11933 1192 11961 1258
rect 11745 1164 11787 1192
rect 11281 1084 11323 1112
rect 11135 252 11163 1084
rect 11295 252 11323 1084
rect 11759 252 11787 1164
rect 11919 1164 11961 1192
rect 11919 252 11947 1164
rect 12397 1112 12425 1258
rect 12383 1084 12425 1112
rect 12529 1112 12557 1258
rect 12993 1192 13021 1258
rect 13181 1192 13209 1258
rect 12993 1164 13035 1192
rect 12529 1084 12571 1112
rect 12383 252 12411 1084
rect 12543 252 12571 1084
rect 13007 252 13035 1164
rect 13167 1164 13209 1192
rect 13167 252 13195 1164
rect 13645 1112 13673 1258
rect 13631 1084 13673 1112
rect 13777 1112 13805 1258
rect 14241 1192 14269 1258
rect 14429 1192 14457 1258
rect 14241 1164 14283 1192
rect 13777 1084 13819 1112
rect 13631 252 13659 1084
rect 13791 252 13819 1084
rect 14255 252 14283 1164
rect 14415 1164 14457 1192
rect 14415 252 14443 1164
rect 14893 1112 14921 1258
rect 14879 1084 14921 1112
rect 15025 1112 15053 1258
rect 15489 1192 15517 1258
rect 15677 1192 15705 1258
rect 15489 1164 15531 1192
rect 15025 1084 15067 1112
rect 14879 252 14907 1084
rect 15039 252 15067 1084
rect 15503 252 15531 1164
rect 15663 1164 15705 1192
rect 15663 252 15691 1164
rect 16141 1112 16169 1258
rect 16127 1084 16169 1112
rect 16273 1112 16301 1258
rect 16737 1192 16765 1258
rect 16925 1192 16953 1258
rect 16737 1164 16779 1192
rect 16273 1084 16315 1112
rect 16127 252 16155 1084
rect 16287 252 16315 1084
rect 16751 252 16779 1164
rect 16911 1164 16953 1192
rect 16911 252 16939 1164
rect 17389 1112 17417 1258
rect 17375 1084 17417 1112
rect 17521 1112 17549 1258
rect 17985 1192 18013 1258
rect 18173 1192 18201 1258
rect 17985 1164 18027 1192
rect 17521 1084 17563 1112
rect 17375 252 17403 1084
rect 17535 252 17563 1084
rect 17999 252 18027 1164
rect 18159 1164 18201 1192
rect 18159 252 18187 1164
rect 18637 1112 18665 1258
rect 18623 1084 18665 1112
rect 18769 1112 18797 1258
rect 19233 1192 19261 1258
rect 19421 1192 19449 1258
rect 19233 1164 19275 1192
rect 18769 1084 18811 1112
rect 18623 252 18651 1084
rect 18783 252 18811 1084
rect 19247 252 19275 1164
rect 19407 1164 19449 1192
rect 19407 252 19435 1164
rect 19885 1112 19913 1258
rect 19871 1084 19913 1112
rect 20017 1112 20045 1258
rect 20481 1192 20509 1258
rect 20669 1192 20697 1258
rect 20481 1164 20523 1192
rect 20017 1084 20059 1112
rect 19871 252 19899 1084
rect 20031 252 20059 1084
rect 20495 252 20523 1164
rect 20655 1164 20697 1192
rect 20655 252 20683 1164
rect 21133 1112 21161 1258
rect 21119 1084 21161 1112
rect 21265 1112 21293 1258
rect 21729 1192 21757 1258
rect 21917 1192 21945 1258
rect 21729 1164 21771 1192
rect 21265 1084 21307 1112
rect 21119 252 21147 1084
rect 21279 252 21307 1084
rect 21743 252 21771 1164
rect 21903 1164 21945 1192
rect 21903 252 21931 1164
rect 22381 1112 22409 1258
rect 22367 1084 22409 1112
rect 22513 1112 22541 1258
rect 22977 1192 23005 1258
rect 23165 1192 23193 1258
rect 22977 1164 23019 1192
rect 22513 1084 22555 1112
rect 22367 252 22395 1084
rect 22527 252 22555 1084
rect 22991 252 23019 1164
rect 23151 1164 23193 1192
rect 23151 252 23179 1164
rect 23629 1112 23657 1258
rect 23615 1084 23657 1112
rect 23761 1112 23789 1258
rect 24225 1192 24253 1258
rect 24413 1192 24441 1258
rect 24225 1164 24267 1192
rect 23761 1084 23803 1112
rect 23615 252 23643 1084
rect 23775 252 23803 1084
rect 24239 252 24267 1164
rect 24399 1164 24441 1192
rect 24399 252 24427 1164
rect 24877 1112 24905 1258
rect 24863 1084 24905 1112
rect 25009 1112 25037 1258
rect 25473 1192 25501 1258
rect 25661 1192 25689 1258
rect 25473 1164 25515 1192
rect 25009 1084 25051 1112
rect 24863 252 24891 1084
rect 25023 252 25051 1084
rect 25487 252 25515 1164
rect 25647 1164 25689 1192
rect 25647 252 25675 1164
rect 26125 1112 26153 1258
rect 26111 1084 26153 1112
rect 26257 1112 26285 1258
rect 26721 1192 26749 1258
rect 26909 1192 26937 1258
rect 26721 1164 26763 1192
rect 26257 1084 26299 1112
rect 26111 252 26139 1084
rect 26271 252 26299 1084
rect 26735 252 26763 1164
rect 26895 1164 26937 1192
rect 26895 252 26923 1164
rect 27373 1112 27401 1258
rect 27359 1084 27401 1112
rect 27505 1112 27533 1258
rect 27969 1192 27997 1258
rect 28157 1192 28185 1258
rect 27969 1164 28011 1192
rect 27505 1084 27547 1112
rect 27359 252 27387 1084
rect 27519 252 27547 1084
rect 27983 252 28011 1164
rect 28143 1164 28185 1192
rect 28143 252 28171 1164
rect 28621 1112 28649 1258
rect 28607 1084 28649 1112
rect 28753 1112 28781 1258
rect 29217 1192 29245 1258
rect 29405 1192 29433 1258
rect 29217 1164 29259 1192
rect 28753 1084 28795 1112
rect 28607 252 28635 1084
rect 28767 252 28795 1084
rect 29231 252 29259 1164
rect 29391 1164 29433 1192
rect 29391 252 29419 1164
rect 29869 1112 29897 1258
rect 29855 1084 29897 1112
rect 30001 1112 30029 1258
rect 30465 1192 30493 1258
rect 30653 1192 30681 1258
rect 30465 1164 30507 1192
rect 30001 1084 30043 1112
rect 29855 252 29883 1084
rect 30015 252 30043 1084
rect 30479 252 30507 1164
rect 30639 1164 30681 1192
rect 30639 252 30667 1164
rect 31117 1112 31145 1258
rect 31103 1084 31145 1112
rect 31249 1112 31277 1258
rect 31713 1192 31741 1258
rect 31713 1164 31755 1192
rect 31249 1084 31291 1112
rect 31103 252 31131 1084
rect 31263 252 31291 1084
rect 31727 252 31755 1164
<< metal3 >>
rect 33 5107 31106 5173
rect 33 4615 31106 4681
rect 33 4283 31106 4349
rect 33 3846 31106 3912
rect 0 2762 31821 2822
rect 0 2638 31821 2698
rect 33 1878 31244 1944
rect 33 948 31854 1014
rect 33 329 31854 395
use sky130_sram_1r1w_24x128_8_column_mux_array  sky130_sram_1r1w_24x128_8_column_mux_array_0
timestamp 1661296025
transform 1 0 0 0 -1 3194
box 0 87 31821 1936
use sky130_sram_1r1w_24x128_8_precharge_array  sky130_sram_1r1w_24x128_8_precharge_array_0
timestamp 1661296025
transform 1 0 0 0 -1 1006
box 33 -12 31854 754
use sky130_sram_1r1w_24x128_8_write_driver_array  sky130_sram_1r1w_24x128_8_write_driver_array_0
timestamp 1661296025
transform 1 0 0 0 -1 5457
box 0 4 31453 2011
<< labels >>
rlabel metal1 s 2092 5397 2152 5453 4 din_0
port 1 nsew
rlabel metal1 s 3340 5397 3400 5453 4 din_1
port 2 nsew
rlabel metal1 s 4588 5397 4648 5453 4 din_2
port 3 nsew
rlabel metal1 s 5836 5397 5896 5453 4 din_3
port 4 nsew
rlabel metal1 s 7084 5397 7144 5453 4 din_4
port 5 nsew
rlabel metal1 s 8332 5397 8392 5453 4 din_5
port 6 nsew
rlabel metal1 s 9580 5397 9640 5453 4 din_6
port 7 nsew
rlabel metal1 s 10828 5397 10888 5453 4 din_7
port 8 nsew
rlabel metal1 s 12076 5397 12136 5453 4 din_8
port 9 nsew
rlabel metal1 s 13324 5397 13384 5453 4 din_9
port 10 nsew
rlabel metal1 s 14572 5397 14632 5453 4 din_10
port 11 nsew
rlabel metal1 s 15820 5397 15880 5453 4 din_11
port 12 nsew
rlabel metal1 s 17068 5397 17128 5453 4 din_12
port 13 nsew
rlabel metal1 s 18316 5397 18376 5453 4 din_13
port 14 nsew
rlabel metal1 s 19564 5397 19624 5453 4 din_14
port 15 nsew
rlabel metal1 s 20812 5397 20872 5453 4 din_15
port 16 nsew
rlabel metal1 s 22060 5397 22120 5453 4 din_16
port 17 nsew
rlabel metal1 s 23308 5397 23368 5453 4 din_17
port 18 nsew
rlabel metal1 s 24556 5397 24616 5453 4 din_18
port 19 nsew
rlabel metal1 s 25804 5397 25864 5453 4 din_19
port 20 nsew
rlabel metal1 s 27052 5397 27112 5453 4 din_20
port 21 nsew
rlabel metal1 s 28300 5397 28360 5453 4 din_21
port 22 nsew
rlabel metal1 s 29548 5397 29608 5453 4 din_22
port 23 nsew
rlabel metal1 s 30796 5397 30856 5453 4 din_23
port 24 nsew
rlabel metal1 s 1775 252 1803 1006 4 rbl_bl
port 25 nsew
rlabel metal1 s 1311 252 1339 1006 4 rbl_br
port 26 nsew
rlabel metal1 s 1935 252 1963 1006 4 bl_0
port 27 nsew
rlabel metal1 s 2399 252 2427 1006 4 br_0
port 28 nsew
rlabel metal1 s 3023 252 3051 1006 4 bl_1
port 29 nsew
rlabel metal1 s 2559 252 2587 1006 4 br_1
port 30 nsew
rlabel metal1 s 3183 252 3211 1006 4 bl_2
port 31 nsew
rlabel metal1 s 3647 252 3675 1006 4 br_2
port 32 nsew
rlabel metal1 s 4271 252 4299 1006 4 bl_3
port 33 nsew
rlabel metal1 s 3807 252 3835 1006 4 br_3
port 34 nsew
rlabel metal1 s 4431 252 4459 1006 4 bl_4
port 35 nsew
rlabel metal1 s 4895 252 4923 1006 4 br_4
port 36 nsew
rlabel metal1 s 5519 252 5547 1006 4 bl_5
port 37 nsew
rlabel metal1 s 5055 252 5083 1006 4 br_5
port 38 nsew
rlabel metal1 s 5679 252 5707 1006 4 bl_6
port 39 nsew
rlabel metal1 s 6143 252 6171 1006 4 br_6
port 40 nsew
rlabel metal1 s 6767 252 6795 1006 4 bl_7
port 41 nsew
rlabel metal1 s 6303 252 6331 1006 4 br_7
port 42 nsew
rlabel metal1 s 6927 252 6955 1006 4 bl_8
port 43 nsew
rlabel metal1 s 7391 252 7419 1006 4 br_8
port 44 nsew
rlabel metal1 s 8015 252 8043 1006 4 bl_9
port 45 nsew
rlabel metal1 s 7551 252 7579 1006 4 br_9
port 46 nsew
rlabel metal1 s 8175 252 8203 1006 4 bl_10
port 47 nsew
rlabel metal1 s 8639 252 8667 1006 4 br_10
port 48 nsew
rlabel metal1 s 9263 252 9291 1006 4 bl_11
port 49 nsew
rlabel metal1 s 8799 252 8827 1006 4 br_11
port 50 nsew
rlabel metal1 s 9423 252 9451 1006 4 bl_12
port 51 nsew
rlabel metal1 s 9887 252 9915 1006 4 br_12
port 52 nsew
rlabel metal1 s 10511 252 10539 1006 4 bl_13
port 53 nsew
rlabel metal1 s 10047 252 10075 1006 4 br_13
port 54 nsew
rlabel metal1 s 10671 252 10699 1006 4 bl_14
port 55 nsew
rlabel metal1 s 11135 252 11163 1006 4 br_14
port 56 nsew
rlabel metal1 s 11759 252 11787 1006 4 bl_15
port 57 nsew
rlabel metal1 s 11295 252 11323 1006 4 br_15
port 58 nsew
rlabel metal1 s 11919 252 11947 1006 4 bl_16
port 59 nsew
rlabel metal1 s 12383 252 12411 1006 4 br_16
port 60 nsew
rlabel metal1 s 13007 252 13035 1006 4 bl_17
port 61 nsew
rlabel metal1 s 12543 252 12571 1006 4 br_17
port 62 nsew
rlabel metal1 s 13167 252 13195 1006 4 bl_18
port 63 nsew
rlabel metal1 s 13631 252 13659 1006 4 br_18
port 64 nsew
rlabel metal1 s 14255 252 14283 1006 4 bl_19
port 65 nsew
rlabel metal1 s 13791 252 13819 1006 4 br_19
port 66 nsew
rlabel metal1 s 14415 252 14443 1006 4 bl_20
port 67 nsew
rlabel metal1 s 14879 252 14907 1006 4 br_20
port 68 nsew
rlabel metal1 s 15503 252 15531 1006 4 bl_21
port 69 nsew
rlabel metal1 s 15039 252 15067 1006 4 br_21
port 70 nsew
rlabel metal1 s 15663 252 15691 1006 4 bl_22
port 71 nsew
rlabel metal1 s 16127 252 16155 1006 4 br_22
port 72 nsew
rlabel metal1 s 16751 252 16779 1006 4 bl_23
port 73 nsew
rlabel metal1 s 16287 252 16315 1006 4 br_23
port 74 nsew
rlabel metal1 s 16911 252 16939 1006 4 bl_24
port 75 nsew
rlabel metal1 s 17375 252 17403 1006 4 br_24
port 76 nsew
rlabel metal1 s 17999 252 18027 1006 4 bl_25
port 77 nsew
rlabel metal1 s 17535 252 17563 1006 4 br_25
port 78 nsew
rlabel metal1 s 18159 252 18187 1006 4 bl_26
port 79 nsew
rlabel metal1 s 18623 252 18651 1006 4 br_26
port 80 nsew
rlabel metal1 s 19247 252 19275 1006 4 bl_27
port 81 nsew
rlabel metal1 s 18783 252 18811 1006 4 br_27
port 82 nsew
rlabel metal1 s 19407 252 19435 1006 4 bl_28
port 83 nsew
rlabel metal1 s 19871 252 19899 1006 4 br_28
port 84 nsew
rlabel metal1 s 20495 252 20523 1006 4 bl_29
port 85 nsew
rlabel metal1 s 20031 252 20059 1006 4 br_29
port 86 nsew
rlabel metal1 s 20655 252 20683 1006 4 bl_30
port 87 nsew
rlabel metal1 s 21119 252 21147 1006 4 br_30
port 88 nsew
rlabel metal1 s 21743 252 21771 1006 4 bl_31
port 89 nsew
rlabel metal1 s 21279 252 21307 1006 4 br_31
port 90 nsew
rlabel metal1 s 21903 252 21931 1006 4 bl_32
port 91 nsew
rlabel metal1 s 22367 252 22395 1006 4 br_32
port 92 nsew
rlabel metal1 s 22991 252 23019 1006 4 bl_33
port 93 nsew
rlabel metal1 s 22527 252 22555 1006 4 br_33
port 94 nsew
rlabel metal1 s 23151 252 23179 1006 4 bl_34
port 95 nsew
rlabel metal1 s 23615 252 23643 1006 4 br_34
port 96 nsew
rlabel metal1 s 24239 252 24267 1006 4 bl_35
port 97 nsew
rlabel metal1 s 23775 252 23803 1006 4 br_35
port 98 nsew
rlabel metal1 s 24399 252 24427 1006 4 bl_36
port 99 nsew
rlabel metal1 s 24863 252 24891 1006 4 br_36
port 100 nsew
rlabel metal1 s 25487 252 25515 1006 4 bl_37
port 101 nsew
rlabel metal1 s 25023 252 25051 1006 4 br_37
port 102 nsew
rlabel metal1 s 25647 252 25675 1006 4 bl_38
port 103 nsew
rlabel metal1 s 26111 252 26139 1006 4 br_38
port 104 nsew
rlabel metal1 s 26735 252 26763 1006 4 bl_39
port 105 nsew
rlabel metal1 s 26271 252 26299 1006 4 br_39
port 106 nsew
rlabel metal1 s 26895 252 26923 1006 4 bl_40
port 107 nsew
rlabel metal1 s 27359 252 27387 1006 4 br_40
port 108 nsew
rlabel metal1 s 27983 252 28011 1006 4 bl_41
port 109 nsew
rlabel metal1 s 27519 252 27547 1006 4 br_41
port 110 nsew
rlabel metal1 s 28143 252 28171 1006 4 bl_42
port 111 nsew
rlabel metal1 s 28607 252 28635 1006 4 br_42
port 112 nsew
rlabel metal1 s 29231 252 29259 1006 4 bl_43
port 113 nsew
rlabel metal1 s 28767 252 28795 1006 4 br_43
port 114 nsew
rlabel metal1 s 29391 252 29419 1006 4 bl_44
port 115 nsew
rlabel metal1 s 29855 252 29883 1006 4 br_44
port 116 nsew
rlabel metal1 s 30479 252 30507 1006 4 bl_45
port 117 nsew
rlabel metal1 s 30015 252 30043 1006 4 br_45
port 118 nsew
rlabel metal1 s 30639 252 30667 1006 4 bl_46
port 119 nsew
rlabel metal1 s 31103 252 31131 1006 4 br_46
port 120 nsew
rlabel metal1 s 31727 252 31755 1006 4 bl_47
port 121 nsew
rlabel metal1 s 31263 252 31291 1006 4 br_47
port 122 nsew
rlabel metal3 s 33 948 31854 1014 4 p_en_bar
port 123 nsew
rlabel metal3 s 0 2762 31821 2822 4 sel_0
port 124 nsew
rlabel metal3 s 0 2638 31821 2698 4 sel_1
port 125 nsew
rlabel metal1 s 0 5335 31073 5363 4 w_en
port 126 nsew
rlabel metal3 s 33 329 31854 395 4 vdd
port 127 nsew
rlabel metal3 s 33 4283 31106 4349 4 vdd
port 127 nsew
rlabel metal3 s 33 5107 31106 5173 4 vdd
port 127 nsew
rlabel metal3 s 33 4615 31106 4681 4 gnd
port 128 nsew
rlabel metal3 s 33 3846 31106 3912 4 gnd
port 128 nsew
rlabel metal3 s 33 1878 31244 1944 4 gnd
port 128 nsew
<< properties >>
string FIXED_BBOX 0 0 31821 5457
<< end >>
