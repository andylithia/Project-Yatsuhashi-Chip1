magic
tech sky130B
timestamp 1662581134
<< pwell >>
rect 1637 870 2775 1906
<< psubdiff >>
rect 1655 1871 1703 1888
rect 2709 1871 2757 1888
rect 1655 1840 1672 1871
rect 2740 1840 2757 1871
rect 1655 1703 1672 1734
rect 2740 1703 2757 1734
rect 1655 1686 1703 1703
rect 2709 1686 2757 1703
rect 1655 1605 1703 1622
rect 2709 1605 2757 1622
rect 1655 1574 1672 1605
rect 2740 1574 2757 1605
rect 1655 1437 1672 1468
rect 2740 1437 2757 1468
rect 1655 1420 1703 1437
rect 2709 1420 2757 1437
rect 1655 1339 1703 1356
rect 2709 1339 2757 1356
rect 1655 1308 1672 1339
rect 2740 1308 2757 1339
rect 1655 1171 1672 1202
rect 2740 1171 2757 1202
rect 1655 1154 1703 1171
rect 2709 1154 2757 1171
rect 1655 1073 1703 1090
rect 2709 1073 2757 1090
rect 1655 1042 1672 1073
rect 2740 1042 2757 1073
rect 1655 905 1672 936
rect 2740 905 2757 936
rect 1655 888 1703 905
rect 2709 888 2757 905
<< psubdiffcont >>
rect 1703 1871 2709 1888
rect 1655 1734 1672 1840
rect 2740 1734 2757 1840
rect 1703 1686 2709 1703
rect 1703 1605 2709 1622
rect 1655 1468 1672 1574
rect 2740 1468 2757 1574
rect 1703 1420 2709 1437
rect 1703 1339 2709 1356
rect 1655 1202 1672 1308
rect 2740 1202 2757 1308
rect 1703 1154 2709 1171
rect 1703 1073 2709 1090
rect 1655 936 1672 1042
rect 2740 936 2757 1042
rect 1703 888 2709 905
<< ndiode >>
rect 1706 1831 2706 1837
rect 1706 1743 1712 1831
rect 2700 1743 2706 1831
rect 1706 1737 2706 1743
rect 1706 1565 2706 1571
rect 1706 1477 1712 1565
rect 2700 1477 2706 1565
rect 1706 1471 2706 1477
rect 1706 1299 2706 1305
rect 1706 1211 1712 1299
rect 2700 1211 2706 1299
rect 1706 1205 2706 1211
rect 1706 1033 2706 1039
rect 1706 945 1712 1033
rect 2700 945 2706 1033
rect 1706 939 2706 945
<< ndiodec >>
rect 1712 1743 2700 1831
rect 1712 1477 2700 1565
rect 1712 1211 2700 1299
rect 1712 945 2700 1033
<< locali >>
rect -85 1935 -40 1960
rect 1120 1935 1165 1960
rect -85 1915 -60 1935
rect 1140 1915 1165 1935
rect -20 1870 30 1900
rect 1060 1870 1100 1900
rect -20 1710 10 1870
rect 1070 1710 1100 1870
rect -20 1680 30 1710
rect 1060 1680 1100 1710
rect -20 1630 10 1680
rect 1070 1630 1100 1680
rect -20 1600 30 1630
rect 1060 1600 1100 1630
rect -20 1440 10 1600
rect 1070 1440 1100 1600
rect -20 1410 30 1440
rect 1060 1410 1100 1440
rect -20 1360 10 1410
rect 1070 1360 1100 1410
rect -20 1330 30 1360
rect 1060 1330 1100 1360
rect -20 1170 10 1330
rect 1070 1170 1100 1330
rect -20 1140 30 1170
rect 1060 1140 1100 1170
rect -20 1100 10 1140
rect 1070 1100 1100 1140
rect -20 1070 30 1100
rect 1060 1070 1100 1100
rect -20 910 10 1070
rect 1070 910 1100 1070
rect -20 880 30 910
rect 1060 880 1100 910
rect -85 840 -60 860
rect 1645 1870 1685 1900
rect 2715 1870 2765 1900
rect 1645 1840 1675 1870
rect 1645 1734 1655 1840
rect 1672 1734 1675 1840
rect 2735 1840 2765 1870
rect 1704 1743 1712 1831
rect 2700 1743 2708 1831
rect 1645 1710 1675 1734
rect 2735 1734 2740 1840
rect 2757 1734 2765 1840
rect 2735 1710 2765 1734
rect 1645 1680 1685 1710
rect 2715 1680 2765 1710
rect 1645 1630 1675 1680
rect 2735 1630 2765 1680
rect 1645 1600 1685 1630
rect 2715 1600 2765 1630
rect 1645 1574 1675 1600
rect 1645 1468 1655 1574
rect 1672 1468 1675 1574
rect 2735 1574 2765 1600
rect 1704 1477 1712 1565
rect 2700 1477 2708 1565
rect 1645 1440 1675 1468
rect 2735 1468 2740 1574
rect 2757 1468 2765 1574
rect 2735 1440 2765 1468
rect 1645 1410 1685 1440
rect 2715 1410 2765 1440
rect 1645 1360 1675 1410
rect 2735 1360 2765 1410
rect 1645 1330 1685 1360
rect 2715 1330 2765 1360
rect 1645 1308 1675 1330
rect 1645 1202 1655 1308
rect 1672 1202 1675 1308
rect 2735 1308 2765 1330
rect 1704 1211 1712 1299
rect 2700 1211 2708 1299
rect 1645 1171 1675 1202
rect 2735 1202 2740 1308
rect 2757 1202 2765 1308
rect 2735 1171 2765 1202
rect 1645 1170 1703 1171
rect 2709 1170 2765 1171
rect 1645 1140 1685 1170
rect 2715 1140 2765 1170
rect 1645 1100 1675 1140
rect 2735 1100 2765 1140
rect 1645 1070 1685 1100
rect 2715 1070 2765 1100
rect 1645 1042 1675 1070
rect 1645 936 1655 1042
rect 1672 936 1675 1042
rect 2735 1042 2765 1070
rect 1704 945 1712 1033
rect 2700 945 2708 1033
rect 1645 910 1675 936
rect 2735 936 2740 1042
rect 2757 936 2765 1042
rect 2735 910 2765 936
rect 1645 880 1685 910
rect 2715 880 2765 910
rect 1140 840 1165 860
rect -85 815 -40 840
rect 1120 815 1165 840
<< viali >>
rect -40 1935 1120 1960
rect -85 860 -60 1915
rect 30 1870 1060 1900
rect 30 1680 1060 1710
rect 30 1600 1060 1630
rect 30 1410 1060 1440
rect 30 1330 1060 1360
rect 30 1140 1060 1170
rect 30 1070 1060 1100
rect 30 880 1060 910
rect 1140 860 1165 1915
rect 1685 1888 2715 1900
rect 1685 1871 1703 1888
rect 1703 1871 2709 1888
rect 2709 1871 2715 1888
rect 1685 1870 2715 1871
rect 1712 1743 2700 1831
rect 1685 1703 2715 1710
rect 1685 1686 1703 1703
rect 1703 1686 2709 1703
rect 2709 1686 2715 1703
rect 1685 1680 2715 1686
rect 1685 1622 2715 1630
rect 1685 1605 1703 1622
rect 1703 1605 2709 1622
rect 2709 1605 2715 1622
rect 1685 1600 2715 1605
rect 1712 1477 2700 1565
rect 1685 1437 2715 1440
rect 1685 1420 1703 1437
rect 1703 1420 2709 1437
rect 2709 1420 2715 1437
rect 1685 1410 2715 1420
rect 1685 1356 2715 1360
rect 1685 1339 1703 1356
rect 1703 1339 2709 1356
rect 2709 1339 2715 1356
rect 1685 1330 2715 1339
rect 1712 1211 2700 1299
rect 1685 1154 1703 1170
rect 1703 1154 2709 1170
rect 2709 1154 2715 1170
rect 1685 1140 2715 1154
rect 1685 1090 2715 1100
rect 1685 1073 1703 1090
rect 1703 1073 2709 1090
rect 2709 1073 2715 1090
rect 1685 1070 2715 1073
rect 1712 945 2700 1033
rect 1685 905 2715 910
rect 1685 888 1703 905
rect 1703 888 2709 905
rect 2709 888 2715 905
rect 1685 880 2715 888
rect -40 815 1120 840
<< metal1 >>
rect -90 1930 -40 1965
rect 1120 1930 1170 1965
rect -90 1915 -55 1930
rect 1135 1915 1170 1930
rect -20 1860 10 1910
rect 1070 1860 1100 1910
rect 35 1825 1040 1840
rect 35 1755 50 1825
rect 1025 1755 1040 1825
rect 35 1740 1040 1755
rect -20 1670 10 1720
rect 1070 1670 1100 1720
rect -20 1590 10 1640
rect 1070 1590 1100 1640
rect 35 1555 1040 1570
rect 35 1485 50 1555
rect 1025 1485 1040 1555
rect 35 1470 1040 1485
rect -20 1400 10 1450
rect 1070 1400 1100 1450
rect -20 1320 10 1370
rect 1070 1320 1100 1370
rect 35 1285 1040 1300
rect 35 1215 50 1285
rect 1025 1215 1040 1285
rect 35 1200 1040 1215
rect -20 1130 10 1180
rect 1070 1130 1100 1180
rect -20 1060 10 1110
rect 1070 1060 1100 1110
rect 35 1025 1040 1040
rect 35 955 50 1025
rect 1025 955 1040 1025
rect 35 940 1040 955
rect -20 870 10 920
rect 1070 870 1100 920
rect -90 845 -55 860
rect 1645 1860 1675 1910
rect 2735 1860 2765 1910
rect 1705 1831 2710 1840
rect 1705 1743 1712 1831
rect 2700 1743 2710 1831
rect 1705 1740 2710 1743
rect 1645 1670 1675 1720
rect 2735 1670 2765 1720
rect 1645 1590 1675 1640
rect 2735 1590 2765 1640
rect 1705 1565 2710 1570
rect 1705 1477 1712 1565
rect 2700 1477 2710 1565
rect 1705 1470 2710 1477
rect 1645 1400 1675 1450
rect 2735 1400 2765 1450
rect 1645 1320 1675 1370
rect 2735 1320 2765 1370
rect 1706 1300 2706 1302
rect 1705 1299 2710 1300
rect 1705 1211 1712 1299
rect 2700 1211 2710 1299
rect 1705 1200 2710 1211
rect 1645 1130 1675 1180
rect 2735 1130 2765 1180
rect 1645 1060 1675 1110
rect 2735 1060 2765 1110
rect 1705 1033 2710 1040
rect 1705 945 1712 1033
rect 2700 945 2710 1033
rect 1705 940 2710 945
rect 1645 870 1675 920
rect 2735 870 2765 920
rect 1135 845 1170 860
rect -90 810 -40 845
rect 1120 810 1170 845
<< via1 >>
rect -40 1960 1120 1965
rect -40 1935 1120 1960
rect -40 1930 1120 1935
rect -90 860 -85 1915
rect -85 860 -60 1915
rect -60 860 -55 1915
rect 10 1900 1070 1910
rect 10 1870 30 1900
rect 30 1870 1060 1900
rect 1060 1870 1070 1900
rect 10 1860 1070 1870
rect 50 1755 1025 1825
rect 10 1710 1070 1720
rect 10 1680 30 1710
rect 30 1680 1060 1710
rect 1060 1680 1070 1710
rect 10 1670 1070 1680
rect 10 1630 1070 1640
rect 10 1600 30 1630
rect 30 1600 1060 1630
rect 1060 1600 1070 1630
rect 10 1590 1070 1600
rect 50 1485 1025 1555
rect 10 1440 1070 1450
rect 10 1410 30 1440
rect 30 1410 1060 1440
rect 1060 1410 1070 1440
rect 10 1400 1070 1410
rect 10 1360 1070 1370
rect 10 1330 30 1360
rect 30 1330 1060 1360
rect 1060 1330 1070 1360
rect 10 1320 1070 1330
rect 50 1215 1025 1285
rect 10 1170 1070 1180
rect 10 1140 30 1170
rect 30 1140 1060 1170
rect 1060 1140 1070 1170
rect 10 1130 1070 1140
rect 10 1100 1070 1110
rect 10 1070 30 1100
rect 30 1070 1060 1100
rect 1060 1070 1070 1100
rect 10 1060 1070 1070
rect 50 955 1025 1025
rect 10 910 1070 920
rect 10 880 30 910
rect 30 880 1060 910
rect 1060 880 1070 910
rect 10 870 1070 880
rect 1135 860 1140 1915
rect 1140 860 1165 1915
rect 1165 860 1170 1915
rect 1675 1900 2735 1910
rect 1675 1870 1685 1900
rect 1685 1870 2715 1900
rect 2715 1870 2735 1900
rect 1675 1860 2735 1870
rect 1720 1755 2695 1825
rect 1675 1710 2735 1720
rect 1675 1680 1685 1710
rect 1685 1680 2715 1710
rect 2715 1680 2735 1710
rect 1675 1670 2735 1680
rect 1675 1630 2735 1640
rect 1675 1600 1685 1630
rect 1685 1600 2715 1630
rect 2715 1600 2735 1630
rect 1675 1590 2735 1600
rect 1720 1485 2695 1555
rect 1675 1440 2735 1450
rect 1675 1410 1685 1440
rect 1685 1410 2715 1440
rect 2715 1410 2735 1440
rect 1675 1400 2735 1410
rect 1675 1360 2735 1370
rect 1675 1330 1685 1360
rect 1685 1330 2715 1360
rect 2715 1330 2735 1360
rect 1675 1320 2735 1330
rect 1720 1215 2695 1285
rect 1675 1170 2735 1180
rect 1675 1140 1685 1170
rect 1685 1140 2715 1170
rect 2715 1140 2735 1170
rect 1675 1130 2735 1140
rect 1675 1100 2735 1110
rect 1675 1070 1685 1100
rect 1685 1070 2715 1100
rect 2715 1070 2735 1100
rect 1675 1060 2735 1070
rect 1720 955 2695 1025
rect 1675 910 2735 920
rect 1675 880 1685 910
rect 1685 880 2715 910
rect 2715 880 2735 910
rect 1675 870 2735 880
rect -40 840 1120 845
rect -40 815 1120 840
rect -40 810 1120 815
<< metal2 >>
rect -90 1930 -40 1965
rect 1120 1930 1170 1965
rect -90 1915 -55 1930
rect -105 1725 -90 1800
rect 1135 1915 1170 1930
rect -20 1905 10 1910
rect 1070 1905 1100 1910
rect -20 1865 -15 1905
rect 1095 1865 1100 1905
rect -20 1860 10 1865
rect 1070 1860 1100 1865
rect 45 1825 1030 1830
rect 45 1755 50 1825
rect 1025 1755 1030 1825
rect 45 1750 1030 1755
rect -20 1715 10 1720
rect 1070 1715 1100 1720
rect -20 1675 -15 1715
rect 1095 1675 1100 1715
rect -20 1670 10 1675
rect 1070 1670 1100 1675
rect -20 1635 10 1640
rect 1070 1635 1100 1640
rect -20 1595 -15 1635
rect 1095 1595 1100 1635
rect -20 1590 10 1595
rect 1070 1590 1100 1595
rect 45 1555 1030 1560
rect 45 1485 50 1555
rect 1025 1485 1030 1555
rect 45 1480 1030 1485
rect -20 1445 10 1450
rect 1070 1445 1100 1450
rect -20 1405 -15 1445
rect 1095 1405 1100 1445
rect -20 1400 10 1405
rect 1070 1400 1100 1405
rect -20 1365 10 1370
rect 1070 1365 1100 1370
rect -20 1325 -15 1365
rect 1095 1325 1100 1365
rect -20 1320 10 1325
rect 1070 1320 1100 1325
rect 45 1285 1030 1290
rect 45 1215 50 1285
rect 1025 1215 1030 1285
rect 45 1210 1030 1215
rect -20 1175 10 1180
rect 1070 1175 1100 1180
rect -20 1135 -15 1175
rect 1095 1135 1100 1175
rect -20 1130 10 1135
rect 1070 1130 1100 1135
rect -20 1105 10 1110
rect 1070 1105 1100 1110
rect -20 1065 -15 1105
rect 1095 1065 1100 1105
rect -20 1060 10 1065
rect 1070 1060 1100 1065
rect 45 1025 1030 1030
rect 45 955 50 1025
rect 1025 955 1030 1025
rect 45 950 1030 955
rect -20 915 10 920
rect 1070 915 1100 920
rect -20 875 -15 915
rect 1095 875 1100 915
rect -20 870 10 875
rect 1070 870 1100 875
rect -90 845 -55 860
rect 1645 1905 1675 1910
rect 2735 1905 2765 1910
rect 1645 1865 1650 1905
rect 2760 1865 2765 1905
rect 1645 1860 1675 1865
rect 2735 1860 2765 1865
rect 1715 1825 2700 1830
rect 1715 1755 1720 1825
rect 2695 1755 2700 1825
rect 1715 1750 2700 1755
rect 1645 1715 1675 1720
rect 2735 1715 2765 1720
rect 1645 1675 1650 1715
rect 2760 1675 2765 1715
rect 1645 1670 1675 1675
rect 2735 1670 2765 1675
rect 1645 1635 1675 1640
rect 2735 1635 2765 1640
rect 1645 1595 1650 1635
rect 2760 1595 2765 1635
rect 1645 1590 1675 1595
rect 2735 1590 2765 1595
rect 1715 1555 2700 1560
rect 1715 1485 1720 1555
rect 2695 1485 2700 1555
rect 1715 1480 2700 1485
rect 1645 1445 1675 1450
rect 2735 1445 2765 1450
rect 1645 1405 1650 1445
rect 2760 1405 2765 1445
rect 1645 1400 1675 1405
rect 2735 1400 2765 1405
rect 1645 1365 1675 1370
rect 2735 1365 2765 1370
rect 1645 1325 1650 1365
rect 2760 1325 2765 1365
rect 1645 1320 1675 1325
rect 2735 1320 2765 1325
rect 1715 1285 2700 1290
rect 1715 1215 1720 1285
rect 2695 1215 2700 1285
rect 1715 1210 2700 1215
rect 1645 1175 1675 1180
rect 2735 1175 2765 1180
rect 1645 1135 1650 1175
rect 2760 1135 2765 1175
rect 1645 1130 1675 1135
rect 2735 1130 2765 1135
rect 1645 1105 1675 1110
rect 2735 1105 2765 1110
rect 1645 1065 1650 1105
rect 2760 1065 2765 1105
rect 1645 1060 1675 1065
rect 2735 1060 2765 1065
rect 1715 1025 2700 1030
rect 1715 955 1720 1025
rect 2695 955 2700 1025
rect 1715 950 2700 955
rect 1645 915 1675 920
rect 2735 915 2765 920
rect 1645 875 1650 915
rect 2760 875 2765 915
rect 1645 870 1675 875
rect 2735 870 2765 875
rect 1135 845 1170 860
rect -90 810 -40 845
rect 1120 810 1170 845
<< via2 >>
rect -15 1865 10 1905
rect 10 1865 1070 1905
rect 1070 1865 1095 1905
rect 50 1755 1025 1825
rect -15 1675 10 1715
rect 10 1675 1070 1715
rect 1070 1675 1095 1715
rect -15 1595 10 1635
rect 10 1595 1070 1635
rect 1070 1595 1095 1635
rect 50 1485 1025 1555
rect -15 1405 10 1445
rect 10 1405 1070 1445
rect 1070 1405 1095 1445
rect -15 1325 10 1365
rect 10 1325 1070 1365
rect 1070 1325 1095 1365
rect 50 1215 1025 1285
rect -15 1135 10 1175
rect 10 1135 1070 1175
rect 1070 1135 1095 1175
rect -15 1065 10 1105
rect 10 1065 1070 1105
rect 1070 1065 1095 1105
rect 50 955 1025 1025
rect -15 875 10 915
rect 10 875 1070 915
rect 1070 875 1095 915
rect 1650 1865 1675 1905
rect 1675 1865 2735 1905
rect 2735 1865 2760 1905
rect 1720 1755 2695 1825
rect 1650 1675 1675 1715
rect 1675 1675 2735 1715
rect 2735 1675 2760 1715
rect 1650 1595 1675 1635
rect 1675 1595 2735 1635
rect 2735 1595 2760 1635
rect 1720 1485 2695 1555
rect 1650 1405 1675 1445
rect 1675 1405 2735 1445
rect 2735 1405 2760 1445
rect 1650 1325 1675 1365
rect 1675 1325 2735 1365
rect 2735 1325 2760 1365
rect 1720 1215 2695 1285
rect 1650 1135 1675 1175
rect 1675 1135 2735 1175
rect 2735 1135 2760 1175
rect 1650 1065 1675 1105
rect 1675 1065 2735 1105
rect 2735 1065 2760 1105
rect 1720 955 2695 1025
rect 1650 875 1675 915
rect 1675 875 2735 915
rect 2735 875 2760 915
<< metal3 >>
rect -105 1905 1100 1910
rect -105 1865 -15 1905
rect 1095 1865 1100 1905
rect 1645 1905 2790 1910
rect -105 1860 1100 1865
rect -105 1815 10 1860
rect 1300 1830 1500 1900
rect 1645 1865 1650 1905
rect 2760 1865 2790 1905
rect 1645 1860 2790 1865
rect -40 1720 10 1815
rect 45 1825 2700 1830
rect 45 1755 50 1825
rect 1025 1755 1720 1825
rect 2695 1755 2700 1825
rect 45 1750 2700 1755
rect 2735 1815 2790 1860
rect -40 1715 1100 1720
rect -40 1675 -15 1715
rect 1095 1675 1100 1715
rect -40 1635 1100 1675
rect -40 1595 -15 1635
rect 1095 1595 1100 1635
rect -40 1590 1100 1595
rect -40 1450 10 1590
rect 1130 1560 1185 1750
rect 1280 1560 1535 1750
rect 1630 1720 1685 1750
rect 2735 1720 2785 1815
rect 1630 1715 2785 1720
rect 1630 1675 1650 1715
rect 2760 1675 2785 1715
rect 1630 1635 2785 1675
rect 1630 1595 1650 1635
rect 2760 1595 2785 1635
rect 1630 1590 2785 1595
rect 1630 1560 1685 1590
rect 45 1555 2700 1560
rect 45 1485 50 1555
rect 1025 1485 1720 1555
rect 2695 1485 2700 1555
rect 45 1480 2700 1485
rect -40 1445 1100 1450
rect -40 1405 -15 1445
rect 1095 1405 1100 1445
rect -40 1365 1100 1405
rect -40 1325 -15 1365
rect 1095 1325 1100 1365
rect -40 1320 1100 1325
rect -40 1180 10 1320
rect 1130 1290 1185 1480
rect 1280 1290 1535 1480
rect 1630 1450 1685 1480
rect 2735 1450 2785 1590
rect 1630 1445 2785 1450
rect 1630 1405 1650 1445
rect 2760 1405 2785 1445
rect 1630 1365 2785 1405
rect 1630 1325 1650 1365
rect 2760 1325 2785 1365
rect 1630 1320 2785 1325
rect 1630 1290 1685 1320
rect 45 1285 2700 1290
rect 45 1215 50 1285
rect 1025 1215 1720 1285
rect 2695 1215 2700 1285
rect 45 1210 2700 1215
rect -40 1175 1100 1180
rect -40 1135 -15 1175
rect 1095 1135 1100 1175
rect -40 1105 1100 1135
rect -40 1065 -15 1105
rect 1095 1065 1100 1105
rect -40 1060 1100 1065
rect -40 920 10 1060
rect 1130 1030 1185 1210
rect 1280 1030 1535 1210
rect 1630 1180 1685 1210
rect 2735 1180 2785 1320
rect 1630 1175 2785 1180
rect 1630 1135 1650 1175
rect 2760 1135 2785 1175
rect 1630 1105 2785 1135
rect 1630 1065 1650 1105
rect 2760 1065 2785 1105
rect 1630 1060 2785 1065
rect 1630 1030 1685 1060
rect 45 1025 2700 1030
rect 45 955 50 1025
rect 1025 955 1720 1025
rect 2695 955 2700 1025
rect 45 950 2700 955
rect -40 915 1100 920
rect -40 875 -15 915
rect 1095 875 1100 915
rect 1300 900 1500 950
rect 2735 920 2785 1060
rect 1645 915 2785 920
rect -40 870 1100 875
rect 1645 875 1650 915
rect 2760 875 2785 915
rect 1645 870 2785 875
use sky130_fd_pr__diode_pd2nw_05v5_PZH3ZX  sky130_fd_pr__diode_pd2nw_05v5_PZH3ZX_0
timestamp 1662579390
transform 1 0 538 0 1 1387
box -638 -587 638 587
<< labels >>
rlabel metal3 -105 1815 -100 1910 3 VHI
rlabel metal3 1185 1750 1190 1830 7 IO
rlabel metal2 -105 1725 -100 1800 3 VLO
<< end >>
