magic
tech sky130B
magscale 1 2
timestamp 1662263286
<< metal1 >>
rect 1540 9540 2030 9620
rect 1670 9120 1750 9540
rect 1540 9040 2020 9120
rect 1670 8620 1750 9040
rect 1540 8540 2020 8620
rect 1670 8120 1750 8540
rect 1540 8040 2010 8120
rect 1670 7630 1750 8040
rect 0 7580 200 7600
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 10200 7580 10400 7600
rect 10200 7420 10220 7580
rect 10380 7420 10400 7580
rect 10200 7400 10400 7420
rect 0 7100 200 7120
rect 0 6480 200 6500
rect 0 6120 20 6480
rect 180 6120 200 6480
rect 0 6100 200 6120
rect 10200 380 10400 400
rect 10200 220 10220 380
rect 10380 220 10400 380
rect 10200 200 10400 220
<< via1 >>
rect 20 7120 180 7580
rect 10220 7420 10380 7580
rect 20 6120 180 6480
rect 10220 220 10380 380
<< metal2 >>
rect 0 7580 200 7600
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 10200 7580 10400 7600
rect 10200 7420 10220 7580
rect 10380 7420 10400 7580
rect 10200 7400 10400 7420
rect 0 7100 200 7120
rect 0 6480 200 6500
rect 0 6120 20 6480
rect 180 6120 200 6480
rect 0 6100 200 6120
rect 10200 380 10400 400
rect 10200 220 10220 380
rect 10380 220 10400 380
rect 10200 200 10400 220
<< via2 >>
rect 20 7120 180 7580
rect 10220 7420 10380 7580
rect 20 6120 180 6480
rect 10220 220 10380 380
<< metal3 >>
rect -5200 12550 -600 12600
rect -5200 12050 -5150 12550
rect -650 12050 -600 12550
rect -5200 8600 -600 12050
rect 6200 11600 11200 11700
rect -350 11550 2000 11600
rect -350 9950 -300 11550
rect 800 9950 2000 11550
rect -350 9900 2000 9950
rect -9600 8400 -6600 8600
rect -9600 6000 -9400 8400
rect -6800 7200 -6600 8400
rect -5200 8350 -2550 8600
rect -5200 7850 -5150 8350
rect -2650 7850 -2550 8350
rect -5200 7800 -2550 7850
rect -1800 8150 -600 8200
rect 150 8150 400 9550
rect -1800 7650 -1750 8150
rect -650 7800 400 8150
rect -650 7650 -600 7800
rect -1800 7600 -600 7650
rect -100 7740 400 7800
rect -100 7600 200 7740
rect 1540 7640 1900 9100
rect 1500 7600 1900 7640
rect 6200 8400 10700 11600
rect 11100 8400 11200 11600
rect 6200 8300 11200 8400
rect 0 7580 200 7600
rect -6800 6400 -200 7200
rect 0 7120 20 7580
rect 180 7120 200 7580
rect 0 7100 200 7120
rect 6200 6800 9000 8300
rect 10200 7580 11200 7600
rect 10200 7420 10220 7580
rect 10380 7420 11200 7580
rect 10200 7400 11200 7420
rect 5400 6700 9500 6800
rect -100 6480 200 6500
rect -100 6400 20 6480
rect -6800 6120 20 6400
rect 180 6120 200 6480
rect -6800 6000 200 6120
rect -9600 5800 200 6000
rect -1600 2400 200 5800
rect 5500 939 9000 1100
rect 5800 -400 9000 939
rect 11000 400 11200 7400
rect 10200 380 11200 400
rect 10200 220 10220 380
rect 10380 220 11200 380
rect 10200 200 11200 220
rect 11000 0 11200 200
rect 11000 -200 11600 0
rect 5800 -500 10800 -400
rect 5800 -3700 10300 -500
rect 10700 -3700 10800 -500
rect 5800 -3800 10800 -3700
rect 11400 -4000 11600 -200
<< via3 >>
rect -5150 12050 -650 12550
rect -300 9950 800 11550
rect -9400 6000 -6800 8400
rect -5150 7850 -2650 8350
rect -1750 7650 -650 8150
rect 10700 8400 11100 11600
rect 10300 -3700 10700 -500
<< mimcap >>
rect -5150 11700 -650 11750
rect -5150 8700 -5100 11700
rect -700 8700 -650 11700
rect -5150 8650 -650 8700
rect 6300 11500 10100 11600
rect 6300 8500 6400 11500
rect 10000 8500 10100 11500
rect 6300 8400 10100 8500
rect 5900 -600 9700 -500
rect 5900 -3600 6000 -600
rect 9600 -3600 9700 -600
rect 5900 -3700 9700 -3600
<< mimcapcontact >>
rect -5100 8700 -700 11700
rect 6400 8500 10000 11500
rect 6000 -3600 9600 -600
<< metal4 >>
rect -5200 12550 -600 12600
rect -5200 12050 -5150 12550
rect -650 12050 -600 12550
rect -5200 12000 -600 12050
rect -5200 11700 -450 11800
rect -5200 8700 -5100 11700
rect -700 11600 -450 11700
rect -700 11550 850 11600
rect -700 9950 -300 11550
rect 800 9950 850 11550
rect 6200 11500 10200 11700
rect 6200 11400 6400 11500
rect -700 9900 850 9950
rect 1900 11200 6400 11400
rect 1900 9900 2000 11200
rect -700 8700 -600 9900
rect -5200 8600 -600 8700
rect -9600 8400 -6600 8600
rect -9600 6000 -9400 8400
rect -6800 6000 -6600 8400
rect -5200 8350 -2550 8400
rect -5200 7850 -5150 8350
rect -2650 7850 -2550 8350
rect 1800 8200 2000 9900
rect 4200 8500 6400 11200
rect 10000 8500 10200 11500
rect 4200 8300 10200 8500
rect 10600 11600 11200 11700
rect 10600 8400 10700 11600
rect 11100 8400 11200 11600
rect 10600 8300 11200 8400
rect 4200 8200 4439 8300
rect -5200 7800 -2550 7850
rect -1800 8150 -600 8200
rect -1800 7650 -1750 8150
rect -650 7650 -600 8150
rect 1800 8001 4439 8200
rect 1800 8000 4400 8001
rect -1800 7600 -600 7650
rect -9600 5800 -6600 6000
rect 10200 1800 17800 6000
rect 3700 -400 4400 400
rect 3700 -600 9800 -400
rect 3700 -3600 6000 -600
rect 9600 -3600 9800 -600
rect 3700 -3800 9800 -3600
rect 10200 -500 10800 -400
rect 10200 -3700 10300 -500
rect 10700 -3700 10800 -500
rect 10200 -3800 10800 -3700
rect 11800 -4000 16400 1800
<< via4 >>
rect -5150 12050 -650 12550
rect -9400 6000 -6800 8400
rect -5150 7850 -2650 8350
rect 2000 8200 4200 11200
rect 10700 8400 11100 11600
rect -1750 7650 -650 8150
rect 10300 -3700 10700 -500
<< mimcap2 >>
rect -5150 11700 -650 11750
rect -5150 8700 -5100 11700
rect -700 8700 -650 11700
rect -5150 8650 -650 8700
rect 6300 11500 10100 11600
rect 6300 8500 6400 11500
rect 10000 8500 10100 11500
rect 6300 8400 10100 8500
rect 5900 -600 9700 -500
rect 5900 -3600 6000 -600
rect 9600 -3600 9700 -600
rect 5900 -3700 9700 -3600
<< mimcap2contact >>
rect -5100 8700 -700 11700
rect 6400 8500 10000 11500
rect 6000 -3600 9600 -600
<< metal5 >>
rect -5200 12550 -600 12600
rect -5200 12050 -5150 12550
rect -650 12050 -600 12550
rect -5200 11700 -600 12050
rect -9600 8400 -6600 10600
rect -9600 6000 -9400 8400
rect -6800 6000 -6600 8400
rect -5200 8700 -5100 11700
rect -700 8700 -600 11700
rect 6200 11600 11200 11700
rect 6200 11500 10700 11600
rect -5200 8350 -600 8700
rect -5200 7850 -5150 8350
rect -2650 8150 -600 8350
rect -2650 7850 -1750 8150
rect -5200 7800 -1750 7850
rect -1800 7650 -1750 7800
rect -650 7650 -600 8150
rect -1800 7600 -600 7650
rect 1800 11200 4400 11400
rect 1800 8200 2000 11200
rect 4200 8200 4400 11200
rect 6200 8500 6400 11500
rect 10000 8500 10700 11500
rect 6200 8400 10700 8500
rect 11100 8400 11200 11600
rect 6200 8300 11200 8400
rect 1800 8100 4400 8200
rect 1800 7600 5900 8100
rect -9600 5800 -6600 6000
rect 5800 -500 10800 -400
rect 5800 -600 10300 -500
rect 5800 -3600 6000 -600
rect 9600 -3600 10300 -600
rect 5800 -3700 10300 -3600
rect 10700 -3700 10800 -500
rect 5800 -3800 10800 -3700
use PA_core_1  PA_core_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/PA/./
timestamp 1660789662
transform 0 -1 10000 1 0 700
box -700 -500 7196 10000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1662263286
transform 1 0 1900 0 1 7640
box 0 0 4000 4000
use nfet_diode_1  nfet_diode_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660705385
transform 1 0 40 0 1 0
box 340 7600 1560 9660
use sky130_fd_pr__res_high_po_0p35_ZE2H5K  sky130_fd_pr__res_high_po_0p35_ZE2H5K_0
timestamp 1660277336
transform 1 0 101 0 1 6798
box -201 -898 201 898
<< labels >>
rlabel metal4 16400 1800 17800 6000 1 OUTPUT
rlabel metal5 1800 10000 4400 11400 1 GND
rlabel metal5 9800 -2400 10800 -400 1 VGATE_CAS
rlabel metal5 10200 9700 11200 11700 1 VGATE_CAS
rlabel metal5 -9600 8700 -6600 10600 1 INPUT
rlabel metal3 -5174 8426 -2634 8636 1 IREF_L
<< end >>
