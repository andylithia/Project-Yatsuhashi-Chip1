magic
tech sky130B
magscale 1 2
timestamp 1666841414
<< pwell >>
rect -5370 19520 -5330 19530
<< locali >>
rect -5380 20650 -4270 20660
rect -5380 20640 -5290 20650
rect -5380 19530 -5370 20640
rect -5336 20610 -5290 20640
rect -4360 20640 -4270 20650
rect -4360 20610 -4310 20640
rect -5336 20600 -4310 20610
rect -5336 19570 -5330 20600
rect -4320 19570 -4310 20600
rect -5336 19560 -4310 19570
rect -5336 19530 -5290 19560
rect -5380 19520 -5290 19530
rect -4360 19530 -4310 19560
rect -4276 19530 -4270 20640
rect -4360 19520 -4270 19530
rect -5380 19510 -4270 19520
<< viali >>
rect -5370 19530 -5336 20640
rect -5290 20610 -4360 20650
rect -5290 19520 -4360 19560
rect -4310 19530 -4276 20640
<< metal1 >>
rect -5500 21100 -2500 21200
rect -5500 21080 -5380 21100
rect -5120 21080 -4880 21100
rect -4620 21080 -4380 21100
rect -4120 21080 -3880 21100
rect -3620 21080 -3380 21100
rect -3120 21080 -2880 21100
rect -2620 21080 -2500 21100
rect -5500 20820 -5400 21080
rect -5100 20820 -4900 21080
rect -4600 20820 -4400 21080
rect -4100 20820 -3900 21080
rect -3600 20820 -3400 21080
rect -3100 20820 -2900 21080
rect -2600 20820 -2500 21080
rect -5500 20800 -5380 20820
rect -5120 20800 -4880 20820
rect -4620 20800 -4380 20820
rect -4120 20800 -3880 20820
rect -3620 20800 -3380 20820
rect -3120 20800 -2880 20820
rect -2620 20800 -2500 20820
rect -5500 20700 -2500 20800
rect 5500 21100 11500 21200
rect 5500 21080 5620 21100
rect 5880 21080 6120 21100
rect 6380 21080 6620 21100
rect 6880 21080 7120 21100
rect 7380 21080 7620 21100
rect 7880 21080 8120 21100
rect 8380 21080 8620 21100
rect 8880 21080 9120 21100
rect 9380 21080 9620 21100
rect 9880 21080 10120 21100
rect 10380 21080 10620 21100
rect 10880 21080 11120 21100
rect 11380 21080 11500 21100
rect 5500 20820 5600 21080
rect 5900 20820 6100 21080
rect 6400 20820 6600 21080
rect 6900 20820 7100 21080
rect 7400 20820 7600 21080
rect 7900 20820 8100 21080
rect 8400 20820 8600 21080
rect 8900 20820 9100 21080
rect 9400 20820 9600 21080
rect 9900 20820 10100 21080
rect 10400 20820 10600 21080
rect 10900 20820 11100 21080
rect 11400 20820 11500 21080
rect 5500 20800 5620 20820
rect 5880 20800 6120 20820
rect 6380 20800 6620 20820
rect 6880 20800 7120 20820
rect 7380 20800 7620 20820
rect 7880 20800 8120 20820
rect 8380 20800 8620 20820
rect 8880 20800 9120 20820
rect 9380 20800 9620 20820
rect 9880 20800 10120 20820
rect 10380 20800 10620 20820
rect 10880 20800 11120 20820
rect 11380 20800 11500 20820
rect -4276 20660 -4100 20700
rect -5380 20650 -4100 20660
rect -5380 20640 -5290 20650
rect -21500 20100 -13000 20200
rect -21500 20080 -21380 20100
rect -21120 20080 -20880 20100
rect -20620 20080 -20380 20100
rect -20120 20080 -19880 20100
rect -19620 20080 -19380 20100
rect -19120 20080 -18880 20100
rect -18620 20080 -18380 20100
rect -18120 20080 -17880 20100
rect -17620 20080 -17380 20100
rect -17120 20080 -16880 20100
rect -16620 20080 -16380 20100
rect -16120 20080 -15880 20100
rect -15620 20080 -15380 20100
rect -15120 20080 -14880 20100
rect -14620 20080 -14380 20100
rect -14120 20080 -13880 20100
rect -13620 20080 -13380 20100
rect -13120 20080 -13000 20100
rect -21500 19820 -21400 20080
rect -21100 19820 -20900 20080
rect -20600 19820 -20400 20080
rect -20100 19820 -19900 20080
rect -19600 19820 -19400 20080
rect -19100 19820 -18900 20080
rect -18600 19820 -18400 20080
rect -18100 19820 -17900 20080
rect -17600 19820 -17400 20080
rect -17100 19820 -16900 20080
rect -16600 19820 -16400 20080
rect -16100 19820 -15900 20080
rect -15600 19820 -15400 20080
rect -15100 19820 -14900 20080
rect -14600 19820 -14400 20080
rect -14100 19820 -13900 20080
rect -13600 19820 -13400 20080
rect -13100 19820 -13000 20080
rect -21500 19800 -21380 19820
rect -21120 19800 -20880 19820
rect -20620 19800 -20380 19820
rect -20120 19800 -19880 19820
rect -19620 19800 -19380 19820
rect -19120 19800 -18880 19820
rect -18620 19800 -18380 19820
rect -18120 19800 -17880 19820
rect -17620 19800 -17380 19820
rect -17120 19800 -16880 19820
rect -16620 19800 -16380 19820
rect -16120 19800 -15880 19820
rect -15620 19800 -15380 19820
rect -15120 19800 -14880 19820
rect -14620 19800 -14380 19820
rect -14120 19800 -13880 19820
rect -13620 19800 -13380 19820
rect -13120 19800 -13000 19820
rect -21500 19600 -13000 19800
rect -21500 19580 -21380 19600
rect -21120 19580 -20880 19600
rect -20620 19580 -20380 19600
rect -20120 19580 -19880 19600
rect -19620 19580 -19380 19600
rect -19120 19580 -18880 19600
rect -18620 19580 -18380 19600
rect -18120 19580 -17880 19600
rect -17620 19580 -17380 19600
rect -17120 19580 -16880 19600
rect -16620 19580 -16380 19600
rect -16120 19580 -15880 19600
rect -15620 19580 -15380 19600
rect -15120 19580 -14880 19600
rect -14620 19580 -14380 19600
rect -14120 19580 -13880 19600
rect -13620 19580 -13380 19600
rect -13120 19580 -13000 19600
rect -21500 19320 -21400 19580
rect -21100 19320 -20900 19580
rect -20600 19320 -20400 19580
rect -20100 19320 -19900 19580
rect -19600 19320 -19400 19580
rect -19100 19320 -18900 19580
rect -18600 19320 -18400 19580
rect -18100 19320 -17900 19580
rect -17600 19320 -17400 19580
rect -17100 19320 -16900 19580
rect -16600 19320 -16400 19580
rect -16100 19320 -15900 19580
rect -15600 19320 -15400 19580
rect -15100 19320 -14900 19580
rect -14600 19320 -14400 19580
rect -14100 19320 -13900 19580
rect -13600 19320 -13400 19580
rect -13100 19320 -13000 19580
rect -5380 19530 -5370 20640
rect -5336 20610 -5290 20640
rect -4360 20640 -4100 20650
rect -4360 20610 -4310 20640
rect -5336 20600 -4310 20610
rect -5336 20510 -5330 20600
rect -5140 20550 -5050 20560
rect -5336 20430 -5170 20510
rect -5140 20440 -5130 20550
rect -5060 20440 -5050 20550
rect -4600 20550 -4510 20560
rect -5140 20430 -5050 20440
rect -5021 20437 -4847 20509
rect -4805 20437 -4631 20509
rect -4600 20440 -4590 20550
rect -4520 20440 -4510 20550
rect -4320 20510 -4310 20600
rect -4600 20430 -4510 20440
rect -4480 20430 -4310 20510
rect -5336 19740 -5330 20430
rect -5336 19660 -5170 19740
rect -5129 19663 -4955 19735
rect -5336 19570 -5330 19660
rect -4920 19570 -4730 19750
rect -4320 19740 -4310 20430
rect -4700 19730 -4520 19740
rect -4700 19630 -4690 19730
rect -4530 19630 -4520 19730
rect -4490 19660 -4310 19740
rect -4320 19570 -4310 19660
rect -5336 19560 -4310 19570
rect -5336 19530 -5290 19560
rect -5380 19520 -5290 19530
rect -4360 19530 -4310 19560
rect -4276 20600 -4100 20640
rect 5500 20600 11500 20800
rect -4276 20200 -4000 20600
rect 5500 20580 5620 20600
rect 5880 20580 6120 20600
rect 6380 20580 6620 20600
rect 6880 20580 7120 20600
rect 7380 20580 7620 20600
rect 7880 20580 8120 20600
rect 8380 20580 8620 20600
rect 8880 20580 9120 20600
rect 9380 20580 9620 20600
rect 9880 20580 10120 20600
rect 10380 20580 10620 20600
rect 10880 20580 11120 20600
rect 11380 20580 11500 20600
rect 5500 20320 5600 20580
rect 5900 20320 6100 20580
rect 6400 20320 6600 20580
rect 6900 20320 7100 20580
rect 7400 20320 7600 20580
rect 7900 20320 8100 20580
rect 8400 20320 8600 20580
rect 8900 20320 9100 20580
rect 9400 20320 9600 20580
rect 9900 20320 10100 20580
rect 10400 20320 10600 20580
rect 10900 20320 11100 20580
rect 11400 20320 11500 20580
rect 5500 20300 5620 20320
rect 5880 20300 6120 20320
rect 6380 20300 6620 20320
rect 6880 20300 7120 20320
rect 7380 20300 7620 20320
rect 7880 20300 8120 20320
rect 8380 20300 8620 20320
rect 8880 20300 9120 20320
rect 9380 20300 9620 20320
rect 9880 20300 10120 20320
rect 10380 20300 10620 20320
rect 10880 20300 11120 20320
rect 11380 20300 11500 20320
rect -4276 20100 -4100 20200
rect 5500 20100 11500 20300
rect -4276 19700 -4000 20100
rect 5500 20080 5620 20100
rect 5880 20080 6120 20100
rect 6380 20080 6620 20100
rect 6880 20080 7120 20100
rect 7380 20080 7620 20100
rect 7880 20080 8120 20100
rect 8380 20080 8620 20100
rect 8880 20080 9120 20100
rect 9380 20080 9620 20100
rect 9880 20080 10120 20100
rect 10380 20080 10620 20100
rect 10880 20080 11120 20100
rect 11380 20080 11500 20100
rect 5500 19820 5600 20080
rect 5900 19820 6100 20080
rect 6400 19820 6600 20080
rect 6900 19820 7100 20080
rect 7400 19820 7600 20080
rect 7900 19820 8100 20080
rect 8400 19820 8600 20080
rect 8900 19820 9100 20080
rect 9400 19820 9600 20080
rect 9900 19820 10100 20080
rect 10400 19820 10600 20080
rect 10900 19820 11100 20080
rect 11400 19820 11500 20080
rect 5500 19800 5620 19820
rect 5880 19800 6120 19820
rect 6380 19800 6620 19820
rect 6880 19800 7120 19820
rect 7380 19800 7620 19820
rect 7880 19800 8120 19820
rect 8380 19800 8620 19820
rect 8880 19800 9120 19820
rect 9380 19800 9620 19820
rect 9880 19800 10120 19820
rect 10380 19800 10620 19820
rect 10880 19800 11120 19820
rect 11380 19800 11500 19820
rect 5500 19700 11500 19800
rect -4276 19600 -4100 19700
rect -4000 19600 500 19700
rect -4276 19530 -4270 19600
rect -4360 19520 -4270 19530
rect -5380 19510 -4270 19520
rect -4000 19580 -3880 19600
rect -3620 19580 -3380 19600
rect -3120 19580 -2880 19600
rect -2620 19580 -2380 19600
rect -2120 19580 -1880 19600
rect -1620 19580 -1380 19600
rect -1120 19580 -880 19600
rect -620 19580 -380 19600
rect -120 19580 120 19600
rect 380 19580 500 19600
rect -21500 19300 -21380 19320
rect -21120 19300 -20880 19320
rect -20620 19300 -20380 19320
rect -20120 19300 -19880 19320
rect -19620 19300 -19380 19320
rect -19120 19300 -18880 19320
rect -18620 19300 -18380 19320
rect -18120 19300 -17880 19320
rect -17620 19300 -17380 19320
rect -17120 19300 -16880 19320
rect -16620 19300 -16380 19320
rect -16120 19300 -15880 19320
rect -15620 19300 -15380 19320
rect -15120 19300 -14880 19320
rect -14620 19300 -14380 19320
rect -14120 19300 -13880 19320
rect -13620 19300 -13380 19320
rect -13120 19300 -13000 19320
rect -21500 19100 -13000 19300
rect -4000 19320 -3900 19580
rect -3600 19320 -3400 19580
rect -3100 19320 -2900 19580
rect -2600 19320 -2400 19580
rect -2100 19320 -1900 19580
rect -1600 19320 -1400 19580
rect -1100 19320 -900 19580
rect -600 19320 -400 19580
rect -100 19320 100 19580
rect 400 19320 500 19580
rect -4000 19300 -3880 19320
rect -3620 19300 -3380 19320
rect -3120 19300 -2880 19320
rect -2620 19300 -2380 19320
rect -2120 19300 -1880 19320
rect -1620 19300 -1380 19320
rect -1120 19300 -880 19320
rect -620 19300 -380 19320
rect -120 19300 120 19320
rect 380 19300 500 19320
rect 3700 19600 11500 19700
rect 3700 19580 4120 19600
rect 4380 19580 4620 19600
rect 4880 19580 5120 19600
rect 5380 19580 5620 19600
rect 5880 19580 6120 19600
rect 6380 19580 6620 19600
rect 6880 19580 7120 19600
rect 7380 19580 7620 19600
rect 7880 19580 8120 19600
rect 8380 19580 8620 19600
rect 8880 19580 9120 19600
rect 9380 19580 9620 19600
rect 9880 19580 10120 19600
rect 10380 19580 10620 19600
rect 10880 19580 11120 19600
rect 11380 19580 11500 19600
rect 3700 19320 4100 19580
rect 4400 19320 4600 19580
rect 4900 19320 5100 19580
rect 5400 19320 5600 19580
rect 5900 19320 6100 19580
rect 6400 19320 6600 19580
rect 6900 19320 7100 19580
rect 7400 19320 7600 19580
rect 7900 19320 8100 19580
rect 8400 19320 8600 19580
rect 8900 19320 9100 19580
rect 9400 19320 9600 19580
rect 9900 19320 10100 19580
rect 10400 19320 10600 19580
rect 10900 19320 11100 19580
rect 11400 19320 11500 19580
rect 3700 19300 4120 19320
rect 4380 19300 4620 19320
rect 4880 19300 5120 19320
rect 5380 19300 5620 19320
rect 5880 19300 6120 19320
rect 6380 19300 6620 19320
rect 6880 19300 7120 19320
rect 7380 19300 7620 19320
rect 7880 19300 8120 19320
rect 8380 19300 8620 19320
rect 8880 19300 9120 19320
rect 9380 19300 9620 19320
rect 9880 19300 10120 19320
rect 10380 19300 10620 19320
rect 10880 19300 11120 19320
rect 11380 19300 11500 19320
rect -4000 19200 500 19300
rect -21500 19080 -21380 19100
rect -21120 19080 -20880 19100
rect -20620 19080 -20380 19100
rect -20120 19080 -19880 19100
rect -19620 19080 -19380 19100
rect -19120 19080 -18880 19100
rect -18620 19080 -18380 19100
rect -18120 19080 -17880 19100
rect -17620 19080 -17380 19100
rect -17120 19080 -16880 19100
rect -16620 19080 -16380 19100
rect -16120 19080 -15880 19100
rect -15620 19080 -15380 19100
rect -15120 19080 -14880 19100
rect -14620 19080 -14380 19100
rect -14120 19080 -13880 19100
rect -13620 19080 -13380 19100
rect -13120 19080 -13000 19100
rect -21500 18820 -21400 19080
rect -21100 18820 -20900 19080
rect -20600 18820 -20400 19080
rect -20100 18820 -19900 19080
rect -19600 18820 -19400 19080
rect -19100 18820 -18900 19080
rect -18600 18820 -18400 19080
rect -18100 18820 -17900 19080
rect -17600 18820 -17400 19080
rect -17100 18820 -16900 19080
rect -16600 18820 -16400 19080
rect -16100 18820 -15900 19080
rect -15600 18820 -15400 19080
rect -15100 18820 -14900 19080
rect -14600 18820 -14400 19080
rect -14100 18820 -13900 19080
rect -13600 18820 -13400 19080
rect -13100 18820 -13000 19080
rect -21500 18800 -21380 18820
rect -21120 18800 -20880 18820
rect -20620 18800 -20380 18820
rect -20120 18800 -19880 18820
rect -19620 18800 -19380 18820
rect -19120 18800 -18880 18820
rect -18620 18800 -18380 18820
rect -18120 18800 -17880 18820
rect -17620 18800 -17380 18820
rect -17120 18800 -16880 18820
rect -16620 18800 -16380 18820
rect -16120 18800 -15880 18820
rect -15620 18800 -15380 18820
rect -15120 18800 -14880 18820
rect -14620 18800 -14380 18820
rect -14120 18800 -13880 18820
rect -13620 18800 -13380 18820
rect -13120 18800 -13000 18820
rect -21500 18600 -13000 18800
rect -21500 18580 -21380 18600
rect -21120 18580 -20880 18600
rect -20620 18580 -20380 18600
rect -20120 18580 -19880 18600
rect -19620 18580 -19380 18600
rect -19120 18580 -18880 18600
rect -18620 18580 -18380 18600
rect -18120 18580 -17880 18600
rect -17620 18580 -17380 18600
rect -17120 18580 -16880 18600
rect -16620 18580 -16380 18600
rect -16120 18580 -15880 18600
rect -15620 18580 -15380 18600
rect -15120 18580 -14880 18600
rect -14620 18580 -14380 18600
rect -14120 18580 -13880 18600
rect -13620 18580 -13380 18600
rect -13120 18580 -13000 18600
rect -21500 18320 -21400 18580
rect -21100 18320 -20900 18580
rect -20600 18320 -20400 18580
rect -20100 18320 -19900 18580
rect -19600 18320 -19400 18580
rect -19100 18320 -18900 18580
rect -18600 18320 -18400 18580
rect -18100 18320 -17900 18580
rect -17600 18320 -17400 18580
rect -17100 18320 -16900 18580
rect -16600 18320 -16400 18580
rect -16100 18320 -15900 18580
rect -15600 18320 -15400 18580
rect -15100 18320 -14900 18580
rect -14600 18320 -14400 18580
rect -14100 18320 -13900 18580
rect -13600 18320 -13400 18580
rect -13100 18320 -13000 18580
rect -21500 18300 -21380 18320
rect -21120 18300 -20880 18320
rect -20620 18300 -20380 18320
rect -20120 18300 -19880 18320
rect -19620 18300 -19380 18320
rect -19120 18300 -18880 18320
rect -18620 18300 -18380 18320
rect -18120 18300 -17880 18320
rect -17620 18300 -17380 18320
rect -17120 18300 -16880 18320
rect -16620 18300 -16380 18320
rect -16120 18300 -15880 18320
rect -15620 18300 -15380 18320
rect -15120 18300 -14880 18320
rect -14620 18300 -14380 18320
rect -14120 18300 -13880 18320
rect -13620 18300 -13380 18320
rect -13120 18300 -13000 18320
rect -21500 18100 -13000 18300
rect -5500 19100 500 19200
rect -5500 19080 -5380 19100
rect -5120 19080 -4880 19100
rect -4620 19080 -4380 19100
rect -4120 19080 -3880 19100
rect -3620 19080 -3380 19100
rect -3120 19080 -2880 19100
rect -2620 19080 -2380 19100
rect -2120 19080 -1880 19100
rect -1620 19080 -1380 19100
rect -1120 19080 -880 19100
rect -620 19080 -380 19100
rect -120 19080 120 19100
rect 380 19080 500 19100
rect -5500 18820 -5400 19080
rect -5100 18820 -4900 19080
rect -4600 18820 -4400 19080
rect -4100 18820 -3900 19080
rect -3600 18820 -3400 19080
rect -3100 18820 -2900 19080
rect -2600 18820 -2400 19080
rect -2100 18820 -1900 19080
rect -1600 18820 -1400 19080
rect -1100 18820 -900 19080
rect -600 18820 -400 19080
rect -100 18820 100 19080
rect 400 18820 500 19080
rect -5500 18800 -5380 18820
rect -5120 18800 -4880 18820
rect -4620 18800 -4380 18820
rect -4120 18800 -3880 18820
rect -3620 18800 -3380 18820
rect -3120 18800 -2880 18820
rect -2620 18800 -2380 18820
rect -2120 18800 -1880 18820
rect -1620 18800 -1380 18820
rect -1120 18800 -880 18820
rect -620 18800 -380 18820
rect -120 18800 120 18820
rect 380 18800 500 18820
rect -5500 18600 500 18800
rect -5500 18580 -5380 18600
rect -5120 18580 -4880 18600
rect -4620 18580 -4380 18600
rect -4120 18580 -3880 18600
rect -3620 18580 -3380 18600
rect -3120 18580 -2880 18600
rect -2620 18580 -2380 18600
rect -2120 18580 -1880 18600
rect -1620 18580 -1380 18600
rect -1120 18580 -880 18600
rect -620 18580 -380 18600
rect -120 18580 120 18600
rect 380 18580 500 18600
rect -5500 18320 -5400 18580
rect -5100 18320 -4900 18580
rect -4600 18320 -4400 18580
rect -4100 18320 -3900 18580
rect -3600 18320 -3400 18580
rect -3100 18320 -2900 18580
rect -2600 18320 -2400 18580
rect -2100 18320 -1900 18580
rect -1600 18320 -1400 18580
rect -1100 18320 -900 18580
rect -600 18320 -400 18580
rect -100 18320 100 18580
rect 400 18320 500 18580
rect -5500 18300 -5380 18320
rect -5120 18300 -4880 18320
rect -4620 18300 -4380 18320
rect -4120 18300 -3880 18320
rect -3620 18300 -3380 18320
rect -3120 18300 -2880 18320
rect -2620 18300 -2380 18320
rect -2120 18300 -1880 18320
rect -1620 18300 -1380 18320
rect -1120 18300 -880 18320
rect -620 18300 -380 18320
rect -120 18300 120 18320
rect 380 18300 500 18320
rect -5500 18200 500 18300
rect -21500 18080 -21380 18100
rect -21120 18080 -20880 18100
rect -20620 18080 -20380 18100
rect -20120 18080 -19880 18100
rect -19620 18080 -19380 18100
rect -19120 18080 -18880 18100
rect -18620 18080 -18380 18100
rect -18120 18080 -17880 18100
rect -17620 18080 -17380 18100
rect -17120 18080 -16880 18100
rect -16620 18080 -16380 18100
rect -16120 18080 -15880 18100
rect -15620 18080 -15380 18100
rect -15120 18080 -14880 18100
rect -14620 18080 -14380 18100
rect -14120 18080 -13880 18100
rect -13620 18080 -13380 18100
rect -13120 18080 -13000 18100
rect -21500 17820 -21400 18080
rect -21100 17820 -20900 18080
rect -20600 17820 -20400 18080
rect -20100 17820 -19900 18080
rect -19600 17820 -19400 18080
rect -19100 17820 -18900 18080
rect -18600 17820 -18400 18080
rect -18100 17820 -17900 18080
rect -17600 17820 -17400 18080
rect -17100 17820 -16900 18080
rect -16600 17820 -16400 18080
rect -16100 17820 -15900 18080
rect -15600 17820 -15400 18080
rect -15100 17820 -14900 18080
rect -14600 17820 -14400 18080
rect -14100 17820 -13900 18080
rect -13600 17820 -13400 18080
rect -13100 17820 -13000 18080
rect -21500 17800 -21380 17820
rect -21120 17800 -20880 17820
rect -20620 17800 -20380 17820
rect -20120 17800 -19880 17820
rect -19620 17800 -19380 17820
rect -19120 17800 -18880 17820
rect -18620 17800 -18380 17820
rect -18120 17800 -17880 17820
rect -17620 17800 -17380 17820
rect -17120 17800 -16880 17820
rect -16620 17800 -16380 17820
rect -16120 17800 -15880 17820
rect -15620 17800 -15380 17820
rect -15120 17800 -14880 17820
rect -14620 17800 -14380 17820
rect -14120 17800 -13880 17820
rect -13620 17800 -13380 17820
rect -13120 17800 -13000 17820
rect -21500 17600 -13000 17800
rect -21500 17580 -21380 17600
rect -21120 17580 -20880 17600
rect -20620 17580 -20380 17600
rect -20120 17580 -19880 17600
rect -19620 17580 -19380 17600
rect -19120 17580 -18880 17600
rect -18620 17580 -18380 17600
rect -18120 17580 -17880 17600
rect -17620 17580 -17380 17600
rect -17120 17580 -16880 17600
rect -16620 17580 -16380 17600
rect -16120 17580 -15880 17600
rect -15620 17580 -15380 17600
rect -15120 17580 -14880 17600
rect -14620 17580 -14380 17600
rect -14120 17580 -13880 17600
rect -13620 17580 -13380 17600
rect -13120 17580 -13000 17600
rect -21500 17320 -21400 17580
rect -21100 17320 -20900 17580
rect -20600 17320 -20400 17580
rect -20100 17320 -19900 17580
rect -19600 17320 -19400 17580
rect -19100 17320 -18900 17580
rect -18600 17320 -18400 17580
rect -18100 17320 -17900 17580
rect -17600 17320 -17400 17580
rect -17100 17320 -16900 17580
rect -16600 17320 -16400 17580
rect -16100 17320 -15900 17580
rect -15600 17320 -15400 17580
rect -15100 17320 -14900 17580
rect -14600 17320 -14400 17580
rect -14100 17320 -13900 17580
rect -13600 17320 -13400 17580
rect -13100 17320 -13000 17580
rect -21500 17300 -21380 17320
rect -21120 17300 -20880 17320
rect -20620 17300 -20380 17320
rect -20120 17300 -19880 17320
rect -19620 17300 -19380 17320
rect -19120 17300 -18880 17320
rect -18620 17300 -18380 17320
rect -18120 17300 -17880 17320
rect -17620 17300 -17380 17320
rect -17120 17300 -16880 17320
rect -16620 17300 -16380 17320
rect -16120 17300 -15880 17320
rect -15620 17300 -15380 17320
rect -15120 17300 -14880 17320
rect -14620 17300 -14380 17320
rect -14120 17300 -13880 17320
rect -13620 17300 -13380 17320
rect -13120 17300 -13000 17320
rect -21500 17100 -13000 17300
rect -2500 18100 500 18200
rect -2500 18080 -2380 18100
rect -2120 18080 -1880 18100
rect -1620 18080 -1380 18100
rect -1120 18080 -880 18100
rect -620 18080 -380 18100
rect -120 18080 120 18100
rect 380 18080 500 18100
rect -2500 17820 -2400 18080
rect -2100 17820 -1900 18080
rect -1600 17820 -1400 18080
rect -1100 17820 -900 18080
rect -600 17820 -400 18080
rect -100 17820 100 18080
rect 400 18000 500 18080
rect 3650 19100 11500 19300
rect 3650 19080 4120 19100
rect 4380 19080 4620 19100
rect 4880 19080 5120 19100
rect 5380 19080 5620 19100
rect 5880 19080 6120 19100
rect 6380 19080 6620 19100
rect 6880 19080 7120 19100
rect 7380 19080 7620 19100
rect 7880 19080 8120 19100
rect 8380 19080 8620 19100
rect 8880 19080 9120 19100
rect 9380 19080 9620 19100
rect 9880 19080 10120 19100
rect 10380 19080 10620 19100
rect 10880 19080 11120 19100
rect 11380 19080 11500 19100
rect 3650 18820 4100 19080
rect 4400 18820 4600 19080
rect 4900 18820 5100 19080
rect 5400 18820 5600 19080
rect 5900 18820 6100 19080
rect 6400 18820 6600 19080
rect 6900 18820 7100 19080
rect 7400 18820 7600 19080
rect 7900 18820 8100 19080
rect 8400 18820 8600 19080
rect 8900 18820 9100 19080
rect 9400 18820 9600 19080
rect 9900 18820 10100 19080
rect 10400 18820 10600 19080
rect 10900 18820 11100 19080
rect 11400 18820 11500 19080
rect 3650 18800 4120 18820
rect 4380 18800 4620 18820
rect 4880 18800 5120 18820
rect 5380 18800 5620 18820
rect 5880 18800 6120 18820
rect 6380 18800 6620 18820
rect 6880 18800 7120 18820
rect 7380 18800 7620 18820
rect 7880 18800 8120 18820
rect 8380 18800 8620 18820
rect 8880 18800 9120 18820
rect 9380 18800 9620 18820
rect 9880 18800 10120 18820
rect 10380 18800 10620 18820
rect 10880 18800 11120 18820
rect 11380 18800 11500 18820
rect 3650 18600 11500 18800
rect 3650 18580 4120 18600
rect 4380 18580 4620 18600
rect 4880 18580 5120 18600
rect 5380 18580 5620 18600
rect 5880 18580 6120 18600
rect 6380 18580 6620 18600
rect 6880 18580 7120 18600
rect 7380 18580 7620 18600
rect 7880 18580 8120 18600
rect 8380 18580 8620 18600
rect 8880 18580 9120 18600
rect 9380 18580 9620 18600
rect 9880 18580 10120 18600
rect 10380 18580 10620 18600
rect 10880 18580 11120 18600
rect 11380 18580 11500 18600
rect 3650 18320 4100 18580
rect 4400 18320 4600 18580
rect 4900 18320 5100 18580
rect 5400 18320 5600 18580
rect 5900 18320 6100 18580
rect 6400 18320 6600 18580
rect 6900 18320 7100 18580
rect 7400 18320 7600 18580
rect 7900 18320 8100 18580
rect 8400 18320 8600 18580
rect 8900 18320 9100 18580
rect 9400 18320 9600 18580
rect 9900 18320 10100 18580
rect 10400 18320 10600 18580
rect 10900 18320 11100 18580
rect 11400 18320 11500 18580
rect 3650 18300 4120 18320
rect 4380 18300 4620 18320
rect 4880 18300 5120 18320
rect 5380 18300 5620 18320
rect 5880 18300 6120 18320
rect 6380 18300 6620 18320
rect 6880 18300 7120 18320
rect 7380 18300 7620 18320
rect 7880 18300 8120 18320
rect 8380 18300 8620 18320
rect 8880 18300 9120 18320
rect 9380 18300 9620 18320
rect 9880 18300 10120 18320
rect 10380 18300 10620 18320
rect 10880 18300 11120 18320
rect 11380 18300 11500 18320
rect 3650 18100 11500 18300
rect 3650 18080 4120 18100
rect 4380 18080 4620 18100
rect 4880 18080 5120 18100
rect 5380 18080 5620 18100
rect 5880 18080 6120 18100
rect 6380 18080 6620 18100
rect 6880 18080 7120 18100
rect 7380 18080 7620 18100
rect 7880 18080 8120 18100
rect 8380 18080 8620 18100
rect 8880 18080 9120 18100
rect 9380 18080 9620 18100
rect 9880 18080 10120 18100
rect 10380 18080 10620 18100
rect 10880 18080 11120 18100
rect 11380 18080 11500 18100
rect 3650 18000 4100 18080
rect 400 17820 4100 18000
rect 4400 17820 4600 18080
rect 4900 17820 5100 18080
rect 5400 17820 5600 18080
rect 5900 17820 6100 18080
rect 6400 17820 6600 18080
rect 6900 17820 7100 18080
rect 7400 17820 7600 18080
rect 7900 17820 8100 18080
rect 8400 17820 8600 18080
rect 8900 17820 9100 18080
rect 9400 17820 9600 18080
rect 9900 17820 10100 18080
rect 10400 17820 10600 18080
rect 10900 17820 11100 18080
rect 11400 17820 11500 18080
rect -2500 17800 -2380 17820
rect -2120 17800 -1880 17820
rect -1620 17800 -1380 17820
rect -1120 17800 -880 17820
rect -620 17800 -380 17820
rect -120 17800 120 17820
rect 380 17800 4120 17820
rect 4380 17800 4620 17820
rect 4880 17800 5120 17820
rect 5380 17800 5620 17820
rect 5880 17800 6120 17820
rect 6380 17800 6620 17820
rect 6880 17800 7120 17820
rect 7380 17800 7620 17820
rect 7880 17800 8120 17820
rect 8380 17800 8620 17820
rect 8880 17800 9120 17820
rect 9380 17800 9620 17820
rect 9880 17800 10120 17820
rect 10380 17800 10620 17820
rect 10880 17800 11120 17820
rect 11380 17800 11500 17820
rect -2500 17600 11500 17800
rect -2500 17580 -2380 17600
rect -2120 17580 -1880 17600
rect -1620 17580 -1380 17600
rect -1120 17580 -880 17600
rect -620 17580 -380 17600
rect -120 17580 120 17600
rect 380 17580 620 17600
rect 880 17580 1120 17600
rect 1380 17580 1620 17600
rect 1880 17580 2120 17600
rect 2380 17580 2620 17600
rect 2880 17580 3120 17600
rect 3380 17580 3620 17600
rect 3880 17580 4120 17600
rect 4380 17580 4620 17600
rect 4880 17580 5120 17600
rect 5380 17580 5620 17600
rect 5880 17580 6120 17600
rect 6380 17580 6620 17600
rect 6880 17580 7120 17600
rect 7380 17580 7620 17600
rect 7880 17580 8120 17600
rect 8380 17580 8620 17600
rect 8880 17580 9120 17600
rect 9380 17580 9620 17600
rect 9880 17580 10120 17600
rect 10380 17580 10620 17600
rect 10880 17580 11120 17600
rect 11380 17580 11500 17600
rect -2500 17320 -2400 17580
rect -2100 17320 -1900 17580
rect -1600 17320 -1400 17580
rect -1100 17320 -900 17580
rect -600 17320 -400 17580
rect -100 17320 100 17580
rect 400 17320 600 17580
rect 900 17320 1100 17580
rect 1400 17320 1600 17580
rect 1900 17320 2100 17580
rect 2400 17320 2600 17580
rect 2900 17320 3100 17580
rect 3400 17320 3600 17580
rect 3900 17320 4100 17580
rect 4400 17320 4600 17580
rect 4900 17320 5100 17580
rect 5400 17320 5600 17580
rect 5900 17320 6100 17580
rect 6400 17320 6600 17580
rect 6900 17320 7100 17580
rect 7400 17320 7600 17580
rect 7900 17320 8100 17580
rect 8400 17320 8600 17580
rect 8900 17320 9100 17580
rect 9400 17320 9600 17580
rect 9900 17320 10100 17580
rect 10400 17320 10600 17580
rect 10900 17320 11100 17580
rect 11400 17320 11500 17580
rect -2500 17300 -2380 17320
rect -2120 17300 -1880 17320
rect -1620 17300 -1380 17320
rect -1120 17300 -880 17320
rect -620 17300 -380 17320
rect -120 17300 120 17320
rect 380 17300 620 17320
rect 880 17300 1120 17320
rect 1380 17300 1620 17320
rect 1880 17300 2120 17320
rect 2380 17300 2620 17320
rect 2880 17300 3120 17320
rect 3380 17300 3620 17320
rect 3880 17300 4120 17320
rect 4380 17300 4620 17320
rect 4880 17300 5120 17320
rect 5380 17300 5620 17320
rect 5880 17300 6120 17320
rect 6380 17300 6620 17320
rect 6880 17300 7120 17320
rect 7380 17300 7620 17320
rect 7880 17300 8120 17320
rect 8380 17300 8620 17320
rect 8880 17300 9120 17320
rect 9380 17300 9620 17320
rect 9880 17300 10120 17320
rect 10380 17300 10620 17320
rect 10880 17300 11120 17320
rect 11380 17300 11500 17320
rect -2500 17200 11500 17300
rect -21500 17080 -21380 17100
rect -21120 17080 -20880 17100
rect -20620 17080 -20380 17100
rect -20120 17080 -19880 17100
rect -19620 17080 -19380 17100
rect -19120 17080 -18880 17100
rect -18620 17080 -18380 17100
rect -18120 17080 -17880 17100
rect -17620 17080 -17380 17100
rect -17120 17080 -16880 17100
rect -16620 17080 -16380 17100
rect -16120 17080 -15880 17100
rect -15620 17080 -15380 17100
rect -15120 17080 -14880 17100
rect -14620 17080 -14380 17100
rect -14120 17080 -13880 17100
rect -13620 17080 -13380 17100
rect -13120 17080 -13000 17100
rect -21500 16820 -21400 17080
rect -21100 16820 -20900 17080
rect -20600 16820 -20400 17080
rect -20100 16820 -19900 17080
rect -19600 16820 -19400 17080
rect -19100 16820 -18900 17080
rect -18600 16820 -18400 17080
rect -18100 16820 -17900 17080
rect -17600 16820 -17400 17080
rect -17100 16820 -16900 17080
rect -16600 16820 -16400 17080
rect -16100 16820 -15900 17080
rect -15600 16820 -15400 17080
rect -15100 16820 -14900 17080
rect -14600 16820 -14400 17080
rect -14100 16820 -13900 17080
rect -13600 16820 -13400 17080
rect -13100 16820 -13000 17080
rect -21500 16800 -21380 16820
rect -21120 16800 -20880 16820
rect -20620 16800 -20380 16820
rect -20120 16800 -19880 16820
rect -19620 16800 -19380 16820
rect -19120 16800 -18880 16820
rect -18620 16800 -18380 16820
rect -18120 16800 -17880 16820
rect -17620 16800 -17380 16820
rect -17120 16800 -16880 16820
rect -16620 16800 -16380 16820
rect -16120 16800 -15880 16820
rect -15620 16800 -15380 16820
rect -15120 16800 -14880 16820
rect -14620 16800 -14380 16820
rect -14120 16800 -13880 16820
rect -13620 16800 -13380 16820
rect -13120 16800 -13000 16820
rect -21500 16600 -13000 16800
rect -21500 16580 -21380 16600
rect -21120 16580 -20880 16600
rect -20620 16580 -20380 16600
rect -20120 16580 -19880 16600
rect -19620 16580 -19380 16600
rect -19120 16580 -18880 16600
rect -18620 16580 -18380 16600
rect -18120 16580 -17880 16600
rect -17620 16580 -17380 16600
rect -17120 16580 -16880 16600
rect -16620 16580 -16380 16600
rect -16120 16580 -15880 16600
rect -15620 16580 -15380 16600
rect -15120 16580 -14880 16600
rect -14620 16580 -14380 16600
rect -14120 16580 -13880 16600
rect -13620 16580 -13380 16600
rect -13120 16580 -13000 16600
rect -21500 16320 -21400 16580
rect -21100 16320 -20900 16580
rect -20600 16320 -20400 16580
rect -20100 16320 -19900 16580
rect -19600 16320 -19400 16580
rect -19100 16320 -18900 16580
rect -18600 16320 -18400 16580
rect -18100 16320 -17900 16580
rect -17600 16320 -17400 16580
rect -17100 16320 -16900 16580
rect -16600 16320 -16400 16580
rect -16100 16320 -15900 16580
rect -15600 16320 -15400 16580
rect -15100 16320 -14900 16580
rect -14600 16320 -14400 16580
rect -14100 16320 -13900 16580
rect -13600 16320 -13400 16580
rect -13100 16320 -13000 16580
rect -21500 16300 -21380 16320
rect -21120 16300 -20880 16320
rect -20620 16300 -20380 16320
rect -20120 16300 -19880 16320
rect -19620 16300 -19380 16320
rect -19120 16300 -18880 16320
rect -18620 16300 -18380 16320
rect -18120 16300 -17880 16320
rect -17620 16300 -17380 16320
rect -17120 16300 -16880 16320
rect -16620 16300 -16380 16320
rect -16120 16300 -15880 16320
rect -15620 16300 -15380 16320
rect -15120 16300 -14880 16320
rect -14620 16300 -14380 16320
rect -14120 16300 -13880 16320
rect -13620 16300 -13380 16320
rect -13120 16300 -13000 16320
rect -21500 16100 -13000 16300
rect -21500 16080 -21380 16100
rect -21120 16080 -20880 16100
rect -20620 16080 -20380 16100
rect -20120 16080 -19880 16100
rect -19620 16080 -19380 16100
rect -19120 16080 -18880 16100
rect -18620 16080 -18380 16100
rect -18120 16080 -17880 16100
rect -17620 16080 -17380 16100
rect -17120 16080 -16880 16100
rect -16620 16080 -16380 16100
rect -16120 16080 -15880 16100
rect -15620 16080 -15380 16100
rect -15120 16080 -14880 16100
rect -14620 16080 -14380 16100
rect -14120 16080 -13880 16100
rect -13620 16080 -13380 16100
rect -13120 16080 -13000 16100
rect -21500 15820 -21400 16080
rect -21100 15820 -20900 16080
rect -20600 15820 -20400 16080
rect -20100 15820 -19900 16080
rect -19600 15820 -19400 16080
rect -19100 15820 -18900 16080
rect -18600 15820 -18400 16080
rect -18100 15820 -17900 16080
rect -17600 15820 -17400 16080
rect -17100 15820 -16900 16080
rect -16600 15820 -16400 16080
rect -16100 15820 -15900 16080
rect -15600 15820 -15400 16080
rect -15100 15820 -14900 16080
rect -14600 15820 -14400 16080
rect -14100 15820 -13900 16080
rect -13600 15820 -13400 16080
rect -13100 15820 -13000 16080
rect -21500 15800 -21380 15820
rect -21120 15800 -20880 15820
rect -20620 15800 -20380 15820
rect -20120 15800 -19880 15820
rect -19620 15800 -19380 15820
rect -19120 15800 -18880 15820
rect -18620 15800 -18380 15820
rect -18120 15800 -17880 15820
rect -17620 15800 -17380 15820
rect -17120 15800 -16880 15820
rect -16620 15800 -16380 15820
rect -16120 15800 -15880 15820
rect -15620 15800 -15380 15820
rect -15120 15800 -14880 15820
rect -14620 15800 -14380 15820
rect -14120 15800 -13880 15820
rect -13620 15800 -13380 15820
rect -13120 15800 -13000 15820
rect -21500 15600 -13000 15800
rect 5500 17100 11500 17200
rect 5500 17080 5620 17100
rect 5880 17080 6120 17100
rect 6380 17080 6620 17100
rect 6880 17080 7120 17100
rect 7380 17080 7620 17100
rect 7880 17080 8120 17100
rect 8380 17080 8620 17100
rect 8880 17080 9120 17100
rect 9380 17080 9620 17100
rect 9880 17080 10120 17100
rect 10380 17080 10620 17100
rect 10880 17080 11120 17100
rect 11380 17080 11500 17100
rect 5500 16820 5600 17080
rect 5900 16820 6100 17080
rect 6400 16820 6600 17080
rect 6900 16820 7100 17080
rect 7400 16820 7600 17080
rect 7900 16820 8100 17080
rect 8400 16820 8600 17080
rect 8900 16820 9100 17080
rect 9400 16820 9600 17080
rect 9900 16820 10100 17080
rect 10400 16820 10600 17080
rect 10900 16820 11100 17080
rect 11400 16820 11500 17080
rect 5500 16800 5620 16820
rect 5880 16800 6120 16820
rect 6380 16800 6620 16820
rect 6880 16800 7120 16820
rect 7380 16800 7620 16820
rect 7880 16800 8120 16820
rect 8380 16800 8620 16820
rect 8880 16800 9120 16820
rect 9380 16800 9620 16820
rect 9880 16800 10120 16820
rect 10380 16800 10620 16820
rect 10880 16800 11120 16820
rect 11380 16800 11500 16820
rect 5500 16600 11500 16800
rect 5500 16580 5620 16600
rect 5880 16580 6120 16600
rect 6380 16580 6620 16600
rect 6880 16580 7120 16600
rect 7380 16580 7620 16600
rect 7880 16580 8120 16600
rect 8380 16580 8620 16600
rect 8880 16580 9120 16600
rect 9380 16580 9620 16600
rect 9880 16580 10120 16600
rect 10380 16580 10620 16600
rect 10880 16580 11120 16600
rect 11380 16580 11500 16600
rect 5500 16320 5600 16580
rect 5900 16320 6100 16580
rect 6400 16320 6600 16580
rect 6900 16320 7100 16580
rect 7400 16320 7600 16580
rect 7900 16320 8100 16580
rect 8400 16320 8600 16580
rect 8900 16320 9100 16580
rect 9400 16320 9600 16580
rect 9900 16320 10100 16580
rect 10400 16320 10600 16580
rect 10900 16320 11100 16580
rect 11400 16320 11500 16580
rect 5500 16300 5620 16320
rect 5880 16300 6120 16320
rect 6380 16300 6620 16320
rect 6880 16300 7120 16320
rect 7380 16300 7620 16320
rect 7880 16300 8120 16320
rect 8380 16300 8620 16320
rect 8880 16300 9120 16320
rect 9380 16300 9620 16320
rect 9880 16300 10120 16320
rect 10380 16300 10620 16320
rect 10880 16300 11120 16320
rect 11380 16300 11500 16320
rect 5500 16100 11500 16300
rect 5500 16080 5620 16100
rect 5880 16080 6120 16100
rect 6380 16080 6620 16100
rect 6880 16080 7120 16100
rect 7380 16080 7620 16100
rect 7880 16080 8120 16100
rect 8380 16080 8620 16100
rect 8880 16080 9120 16100
rect 9380 16080 9620 16100
rect 9880 16080 10120 16100
rect 10380 16080 10620 16100
rect 10880 16080 11120 16100
rect 11380 16080 11500 16100
rect 5500 15820 5600 16080
rect 5900 15820 6100 16080
rect 6400 15820 6600 16080
rect 6900 15820 7100 16080
rect 7400 15820 7600 16080
rect 7900 15820 8100 16080
rect 8400 15820 8600 16080
rect 8900 15820 9100 16080
rect 9400 15820 9600 16080
rect 9900 15820 10100 16080
rect 10400 15820 10600 16080
rect 10900 15820 11100 16080
rect 11400 15820 11500 16080
rect 5500 15800 5620 15820
rect 5880 15800 6120 15820
rect 6380 15800 6620 15820
rect 6880 15800 7120 15820
rect 7380 15800 7620 15820
rect 7880 15800 8120 15820
rect 8380 15800 8620 15820
rect 8880 15800 9120 15820
rect 9380 15800 9620 15820
rect 9880 15800 10120 15820
rect 10380 15800 10620 15820
rect 10880 15800 11120 15820
rect 11380 15800 11500 15820
rect 5500 15700 11500 15800
rect -21500 15580 -21380 15600
rect -21120 15580 -20880 15600
rect -20620 15580 -20380 15600
rect -20120 15580 -19880 15600
rect -19620 15580 -19380 15600
rect -19120 15580 -18880 15600
rect -18620 15580 -18380 15600
rect -18120 15580 -17880 15600
rect -17620 15580 -17380 15600
rect -17120 15580 -16880 15600
rect -16620 15580 -16380 15600
rect -16120 15580 -15880 15600
rect -15620 15580 -15380 15600
rect -15120 15580 -14880 15600
rect -14620 15580 -14380 15600
rect -14120 15580 -13880 15600
rect -13620 15580 -13380 15600
rect -13120 15580 -13000 15600
rect -21500 15320 -21400 15580
rect -21100 15320 -20900 15580
rect -20600 15320 -20400 15580
rect -20100 15320 -19900 15580
rect -19600 15320 -19400 15580
rect -19100 15320 -18900 15580
rect -18600 15320 -18400 15580
rect -18100 15320 -17900 15580
rect -17600 15320 -17400 15580
rect -17100 15320 -16900 15580
rect -16600 15320 -16400 15580
rect -16100 15320 -15900 15580
rect -15600 15320 -15400 15580
rect -15100 15320 -14900 15580
rect -14600 15320 -14400 15580
rect -14100 15320 -13900 15580
rect -13600 15320 -13400 15580
rect -13100 15320 -13000 15580
rect -21500 15300 -21380 15320
rect -21120 15300 -20880 15320
rect -20620 15300 -20380 15320
rect -20120 15300 -19880 15320
rect -19620 15300 -19380 15320
rect -19120 15300 -18880 15320
rect -18620 15300 -18380 15320
rect -18120 15300 -17880 15320
rect -17620 15300 -17380 15320
rect -17120 15300 -16880 15320
rect -16620 15300 -16380 15320
rect -16120 15300 -15880 15320
rect -15620 15300 -15380 15320
rect -15120 15300 -14880 15320
rect -14620 15300 -14380 15320
rect -14120 15300 -13880 15320
rect -13620 15300 -13380 15320
rect -13120 15300 -13000 15320
rect -21500 15100 -13000 15300
rect 7500 15600 11500 15700
rect 7500 15580 7620 15600
rect 7880 15580 8120 15600
rect 8380 15580 8620 15600
rect 8880 15580 9120 15600
rect 9380 15580 9620 15600
rect 9880 15580 10120 15600
rect 10380 15580 10620 15600
rect 10880 15580 11120 15600
rect 11380 15580 11500 15600
rect 7500 15320 7600 15580
rect 7900 15320 8100 15580
rect 8400 15320 8600 15580
rect 8900 15320 9100 15580
rect 9400 15320 9600 15580
rect 9900 15320 10100 15580
rect 10400 15320 10600 15580
rect 10900 15320 11100 15580
rect 11400 15320 11500 15580
rect 7500 15300 7620 15320
rect 7880 15300 8120 15320
rect 8380 15300 8620 15320
rect 8880 15300 9120 15320
rect 9380 15300 9620 15320
rect 9880 15300 10120 15320
rect 10380 15300 10620 15320
rect 10880 15300 11120 15320
rect 11380 15300 11500 15320
rect 7500 15200 11500 15300
rect -21500 15080 -21380 15100
rect -21120 15080 -20880 15100
rect -20620 15080 -20380 15100
rect -20120 15080 -19880 15100
rect -19620 15080 -19380 15100
rect -19120 15080 -18880 15100
rect -18620 15080 -18380 15100
rect -18120 15080 -17880 15100
rect -17620 15080 -17380 15100
rect -17120 15080 -16880 15100
rect -16620 15080 -16380 15100
rect -16120 15080 -15880 15100
rect -15620 15080 -15380 15100
rect -15120 15080 -14880 15100
rect -14620 15080 -14380 15100
rect -14120 15080 -13880 15100
rect -13620 15080 -13380 15100
rect -13120 15080 -13000 15100
rect -21500 14820 -21400 15080
rect -21100 14820 -20900 15080
rect -20600 14820 -20400 15080
rect -20100 14820 -19900 15080
rect -19600 14820 -19400 15080
rect -19100 14820 -18900 15080
rect -18600 14820 -18400 15080
rect -18100 14820 -17900 15080
rect -17600 14820 -17400 15080
rect -17100 14820 -16900 15080
rect -16600 14820 -16400 15080
rect -16100 14820 -15900 15080
rect -15600 14820 -15400 15080
rect -15100 14820 -14900 15080
rect -14600 14820 -14400 15080
rect -14100 14820 -13900 15080
rect -13600 14820 -13400 15080
rect -13100 14820 -13000 15080
rect -21500 14800 -21380 14820
rect -21120 14800 -20880 14820
rect -20620 14800 -20380 14820
rect -20120 14800 -19880 14820
rect -19620 14800 -19380 14820
rect -19120 14800 -18880 14820
rect -18620 14800 -18380 14820
rect -18120 14800 -17880 14820
rect -17620 14800 -17380 14820
rect -17120 14800 -16880 14820
rect -16620 14800 -16380 14820
rect -16120 14800 -15880 14820
rect -15620 14800 -15380 14820
rect -15120 14800 -14880 14820
rect -14620 14800 -14380 14820
rect -14120 14800 -13880 14820
rect -13620 14800 -13380 14820
rect -13120 14800 -13000 14820
rect -21500 14600 -13000 14800
rect 8000 15100 11500 15200
rect 8000 15080 8120 15100
rect 8380 15080 8620 15100
rect 8880 15080 9120 15100
rect 9380 15080 9620 15100
rect 9880 15080 10120 15100
rect 10380 15080 10620 15100
rect 10880 15080 11120 15100
rect 11380 15080 11500 15100
rect 8000 14820 8100 15080
rect 8400 14820 8600 15080
rect 8900 14820 9100 15080
rect 9400 14820 9600 15080
rect 9900 14820 10100 15080
rect 10400 14820 10600 15080
rect 10900 14820 11100 15080
rect 11400 14820 11500 15080
rect 8000 14800 8120 14820
rect 8380 14800 8620 14820
rect 8880 14800 9120 14820
rect 9380 14800 9620 14820
rect 9880 14800 10120 14820
rect 10380 14800 10620 14820
rect 10880 14800 11120 14820
rect 11380 14800 11500 14820
rect 8000 14700 11500 14800
rect -21500 14580 -21380 14600
rect -21120 14580 -20880 14600
rect -20620 14580 -20380 14600
rect -20120 14580 -19880 14600
rect -19620 14580 -19380 14600
rect -19120 14580 -18880 14600
rect -18620 14580 -18380 14600
rect -18120 14580 -17880 14600
rect -17620 14580 -17380 14600
rect -17120 14580 -16880 14600
rect -16620 14580 -16380 14600
rect -16120 14580 -15880 14600
rect -15620 14580 -15380 14600
rect -15120 14580 -14880 14600
rect -14620 14580 -14380 14600
rect -14120 14580 -13880 14600
rect -13620 14580 -13380 14600
rect -13120 14580 -13000 14600
rect -21500 14320 -21400 14580
rect -21100 14320 -20900 14580
rect -20600 14320 -20400 14580
rect -20100 14320 -19900 14580
rect -19600 14320 -19400 14580
rect -19100 14320 -18900 14580
rect -18600 14320 -18400 14580
rect -18100 14320 -17900 14580
rect -17600 14320 -17400 14580
rect -17100 14320 -16900 14580
rect -16600 14320 -16400 14580
rect -16100 14320 -15900 14580
rect -15600 14320 -15400 14580
rect -15100 14320 -14900 14580
rect -14600 14320 -14400 14580
rect -14100 14320 -13900 14580
rect -13600 14320 -13400 14580
rect -13100 14320 -13000 14580
rect -21500 14300 -21380 14320
rect -21120 14300 -20880 14320
rect -20620 14300 -20380 14320
rect -20120 14300 -19880 14320
rect -19620 14300 -19380 14320
rect -19120 14300 -18880 14320
rect -18620 14300 -18380 14320
rect -18120 14300 -17880 14320
rect -17620 14300 -17380 14320
rect -17120 14300 -16880 14320
rect -16620 14300 -16380 14320
rect -16120 14300 -15880 14320
rect -15620 14300 -15380 14320
rect -15120 14300 -14880 14320
rect -14620 14300 -14380 14320
rect -14120 14300 -13880 14320
rect -13620 14300 -13380 14320
rect -13120 14300 -13000 14320
rect -21500 14100 -13000 14300
rect 8500 14600 11500 14700
rect 8500 14580 8620 14600
rect 8880 14580 9120 14600
rect 9380 14580 9620 14600
rect 9880 14580 10120 14600
rect 10380 14580 10620 14600
rect 10880 14580 11120 14600
rect 11380 14580 11500 14600
rect 8500 14320 8600 14580
rect 8900 14320 9100 14580
rect 9400 14320 9600 14580
rect 9900 14320 10100 14580
rect 10400 14320 10600 14580
rect 10900 14320 11100 14580
rect 11400 14320 11500 14580
rect 8500 14300 8620 14320
rect 8880 14300 9120 14320
rect 9380 14300 9620 14320
rect 9880 14300 10120 14320
rect 10380 14300 10620 14320
rect 10880 14300 11120 14320
rect 11380 14300 11500 14320
rect 8500 14200 11500 14300
rect -21500 14080 -21380 14100
rect -21120 14080 -20880 14100
rect -20620 14080 -20380 14100
rect -20120 14080 -19880 14100
rect -19620 14080 -19380 14100
rect -19120 14080 -18880 14100
rect -18620 14080 -18380 14100
rect -18120 14080 -17880 14100
rect -17620 14080 -17380 14100
rect -17120 14080 -16880 14100
rect -16620 14080 -16380 14100
rect -16120 14080 -15880 14100
rect -15620 14080 -15380 14100
rect -15120 14080 -14880 14100
rect -14620 14080 -14380 14100
rect -14120 14080 -13880 14100
rect -13620 14080 -13380 14100
rect -13120 14080 -13000 14100
rect -21500 13820 -21400 14080
rect -21100 13820 -20900 14080
rect -20600 13820 -20400 14080
rect -20100 13820 -19900 14080
rect -19600 13820 -19400 14080
rect -19100 13820 -18900 14080
rect -18600 13820 -18400 14080
rect -18100 13820 -17900 14080
rect -17600 13820 -17400 14080
rect -17100 13820 -16900 14080
rect -16600 13820 -16400 14080
rect -16100 13820 -15900 14080
rect -15600 13820 -15400 14080
rect -15100 13820 -14900 14080
rect -14600 13820 -14400 14080
rect -14100 13820 -13900 14080
rect -13600 13820 -13400 14080
rect -13100 13820 -13000 14080
rect -21500 13800 -21380 13820
rect -21120 13800 -20880 13820
rect -20620 13800 -20380 13820
rect -20120 13800 -19880 13820
rect -19620 13800 -19380 13820
rect -19120 13800 -18880 13820
rect -18620 13800 -18380 13820
rect -18120 13800 -17880 13820
rect -17620 13800 -17380 13820
rect -17120 13800 -16880 13820
rect -16620 13800 -16380 13820
rect -16120 13800 -15880 13820
rect -15620 13800 -15380 13820
rect -15120 13800 -14880 13820
rect -14620 13800 -14380 13820
rect -14120 13800 -13880 13820
rect -13620 13800 -13380 13820
rect -13120 13800 -13000 13820
rect -21500 13700 -13000 13800
rect 9000 14100 11500 14200
rect 9000 14080 9120 14100
rect 9380 14080 9620 14100
rect 9880 14080 10120 14100
rect 10380 14080 10620 14100
rect 10880 14080 11120 14100
rect 11380 14080 11500 14100
rect 9000 13820 9100 14080
rect 9400 13820 9600 14080
rect 9900 13820 10100 14080
rect 10400 13820 10600 14080
rect 10900 13820 11100 14080
rect 11400 13820 11500 14080
rect 9000 13800 9120 13820
rect 9380 13800 9620 13820
rect 9880 13800 10120 13820
rect 10380 13800 10620 13820
rect 10880 13800 11120 13820
rect 11380 13800 11500 13820
rect 9000 13700 11500 13800
rect -21500 13600 -13500 13700
rect -21500 13580 -21380 13600
rect -21120 13580 -20880 13600
rect -20620 13580 -20380 13600
rect -20120 13580 -19880 13600
rect -19620 13580 -19380 13600
rect -19120 13580 -18880 13600
rect -18620 13580 -18380 13600
rect -18120 13580 -17880 13600
rect -17620 13580 -17380 13600
rect -17120 13580 -16880 13600
rect -16620 13580 -16380 13600
rect -16120 13580 -15880 13600
rect -15620 13580 -15380 13600
rect -15120 13580 -14880 13600
rect -14620 13580 -14380 13600
rect -14120 13580 -13880 13600
rect -13620 13580 -13500 13600
rect -21500 13320 -21400 13580
rect -21100 13320 -20900 13580
rect -20600 13320 -20400 13580
rect -20100 13320 -19900 13580
rect -19600 13320 -19400 13580
rect -19100 13320 -18900 13580
rect -18600 13320 -18400 13580
rect -18100 13320 -17900 13580
rect -17600 13320 -17400 13580
rect -17100 13320 -16900 13580
rect -16600 13320 -16400 13580
rect -16100 13320 -15900 13580
rect -15600 13320 -15400 13580
rect -15100 13320 -14900 13580
rect -14600 13320 -14400 13580
rect -14100 13320 -13900 13580
rect -13600 13320 -13500 13580
rect -21500 13300 -21380 13320
rect -21120 13300 -20880 13320
rect -20620 13300 -20380 13320
rect -20120 13300 -19880 13320
rect -19620 13300 -19380 13320
rect -19120 13300 -18880 13320
rect -18620 13300 -18380 13320
rect -18120 13300 -17880 13320
rect -17620 13300 -17380 13320
rect -17120 13300 -16880 13320
rect -16620 13300 -16380 13320
rect -16120 13300 -15880 13320
rect -15620 13300 -15380 13320
rect -15120 13300 -14880 13320
rect -14620 13300 -14380 13320
rect -14120 13300 -13880 13320
rect -13620 13300 -13500 13320
rect -21500 13200 -13500 13300
rect 9500 13600 11500 13700
rect 9500 13580 9620 13600
rect 9880 13580 10120 13600
rect 10380 13580 10620 13600
rect 10880 13580 11120 13600
rect 11380 13580 11500 13600
rect 9500 13320 9600 13580
rect 9900 13320 10100 13580
rect 10400 13320 10600 13580
rect 10900 13320 11100 13580
rect 11400 13320 11500 13580
rect 9500 13300 9620 13320
rect 9880 13300 10120 13320
rect 10380 13300 10620 13320
rect 10880 13300 11120 13320
rect 11380 13300 11500 13320
rect 9500 13200 11500 13300
rect -21500 13100 -14000 13200
rect -21500 13080 -21380 13100
rect -21120 13080 -20880 13100
rect -20620 13080 -20380 13100
rect -20120 13080 -19880 13100
rect -19620 13080 -19380 13100
rect -19120 13080 -18880 13100
rect -18620 13080 -18380 13100
rect -18120 13080 -17880 13100
rect -17620 13080 -17380 13100
rect -17120 13080 -16880 13100
rect -16620 13080 -16380 13100
rect -16120 13080 -15880 13100
rect -15620 13080 -15380 13100
rect -15120 13080 -14880 13100
rect -14620 13080 -14380 13100
rect -14120 13080 -14000 13100
rect -21500 12820 -21400 13080
rect -21100 12820 -20900 13080
rect -20600 12820 -20400 13080
rect -20100 12820 -19900 13080
rect -19600 12820 -19400 13080
rect -19100 12820 -18900 13080
rect -18600 12820 -18400 13080
rect -18100 12820 -17900 13080
rect -17600 12820 -17400 13080
rect -17100 12820 -16900 13080
rect -16600 12820 -16400 13080
rect -16100 12820 -15900 13080
rect -15600 12820 -15400 13080
rect -15100 12820 -14900 13080
rect -14600 12820 -14400 13080
rect -14100 12820 -14000 13080
rect -21500 12800 -21380 12820
rect -21120 12800 -20880 12820
rect -20620 12800 -20380 12820
rect -20120 12800 -19880 12820
rect -19620 12800 -19380 12820
rect -19120 12800 -18880 12820
rect -18620 12800 -18380 12820
rect -18120 12800 -17880 12820
rect -17620 12800 -17380 12820
rect -17120 12800 -16880 12820
rect -16620 12800 -16380 12820
rect -16120 12800 -15880 12820
rect -15620 12800 -15380 12820
rect -15120 12800 -14880 12820
rect -14620 12800 -14380 12820
rect -14120 12800 -14000 12820
rect -21500 12700 -14000 12800
rect 10000 13100 11500 13200
rect 10000 13080 10120 13100
rect 10380 13080 10620 13100
rect 10880 13080 11120 13100
rect 11380 13080 11500 13100
rect 10000 12820 10100 13080
rect 10400 12820 10600 13080
rect 10900 12820 11100 13080
rect 11400 12820 11500 13080
rect 10000 12800 10120 12820
rect 10380 12800 10620 12820
rect 10880 12800 11120 12820
rect 11380 12800 11500 12820
rect 10000 12700 11500 12800
rect -21500 12600 -14500 12700
rect -21500 12580 -21380 12600
rect -21120 12580 -20880 12600
rect -20620 12580 -20380 12600
rect -20120 12580 -19880 12600
rect -19620 12580 -19380 12600
rect -19120 12580 -18880 12600
rect -18620 12580 -18380 12600
rect -18120 12580 -17880 12600
rect -17620 12580 -17380 12600
rect -17120 12580 -16880 12600
rect -16620 12580 -16380 12600
rect -16120 12580 -15880 12600
rect -15620 12580 -15380 12600
rect -15120 12580 -14880 12600
rect -14620 12580 -14500 12600
rect -21500 12320 -21400 12580
rect -21100 12320 -20900 12580
rect -20600 12320 -20400 12580
rect -20100 12320 -19900 12580
rect -19600 12320 -19400 12580
rect -19100 12320 -18900 12580
rect -18600 12320 -18400 12580
rect -18100 12320 -17900 12580
rect -17600 12320 -17400 12580
rect -17100 12320 -16900 12580
rect -16600 12320 -16400 12580
rect -16100 12320 -15900 12580
rect -15600 12320 -15400 12580
rect -15100 12320 -14900 12580
rect -14600 12320 -14500 12580
rect -21500 12300 -21380 12320
rect -21120 12300 -20880 12320
rect -20620 12300 -20380 12320
rect -20120 12300 -19880 12320
rect -19620 12300 -19380 12320
rect -19120 12300 -18880 12320
rect -18620 12300 -18380 12320
rect -18120 12300 -17880 12320
rect -17620 12300 -17380 12320
rect -17120 12300 -16880 12320
rect -16620 12300 -16380 12320
rect -16120 12300 -15880 12320
rect -15620 12300 -15380 12320
rect -15120 12300 -14880 12320
rect -14620 12300 -14500 12320
rect -21500 12200 -14500 12300
rect 10500 12600 11500 12700
rect 10500 12580 10620 12600
rect 10880 12580 11120 12600
rect 11380 12580 11500 12600
rect 10500 12320 10600 12580
rect 10900 12320 11100 12580
rect 11400 12320 11500 12580
rect 10500 12300 10620 12320
rect 10880 12300 11120 12320
rect 11380 12300 11500 12320
rect 10500 12200 11500 12300
rect 11000 12100 11500 12200
rect 11000 12080 11120 12100
rect 11380 12080 11500 12100
rect 11000 11820 11100 12080
rect 11400 11820 11500 12080
rect 11000 11800 11120 11820
rect 11380 11800 11500 11820
rect 11000 11700 11500 11800
<< via1 >>
rect -5130 20440 -5060 20550
rect -4590 20440 -4520 20550
rect -4690 19630 -4530 19730
<< metal2 >>
rect -5210 20840 -5010 20860
rect -5210 20580 -5190 20840
rect -5030 20580 -5010 20840
rect -5210 20560 -5010 20580
rect -4650 20840 -4450 20860
rect -4650 20580 -4630 20840
rect -4470 20580 -4450 20840
rect -4650 20560 -4450 20580
rect -5140 20550 -5050 20560
rect -5140 20440 -5130 20550
rect -5060 20440 -5050 20550
rect -5140 20430 -5050 20440
rect -4600 20550 -4510 20560
rect -4600 20440 -4590 20550
rect -4520 20440 -4510 20550
rect -4600 20430 -4510 20440
rect -14800 19800 -14000 19850
rect -14800 15500 -14750 19800
rect -14050 19600 -12700 19800
rect -4700 19730 -4520 19740
rect -9500 19600 -9050 19650
rect -14050 19400 -14000 19600
rect -14050 19200 -12700 19400
rect -14050 19000 -14000 19200
rect -14050 18800 -12700 19000
rect -14050 18600 -14000 18800
rect -14050 18400 -12700 18600
rect -14050 18200 -14000 18400
rect -14050 18000 -12700 18200
rect -9500 18000 -9450 19600
rect -9100 18000 -9050 19600
rect -4700 19540 -4690 19730
rect -4530 19540 -4520 19730
rect -4700 19530 -4520 19540
rect -14050 17800 -14000 18000
rect -9500 17950 -9050 18000
rect -14050 17600 -12700 17800
rect -14050 17400 -14000 17600
rect -14050 17200 -12700 17400
rect -14050 17000 -14000 17200
rect -14050 16800 -12700 17000
rect -14050 16600 -14000 16800
rect -14050 16400 -12700 16600
rect -14050 16200 -14000 16400
rect -14050 16000 -12700 16200
rect -14050 15500 -14000 16000
rect -14800 15450 -14000 15500
<< via2 >>
rect -5190 20580 -5030 20840
rect -4630 20580 -4470 20840
rect -14750 15500 -14050 19800
rect -9450 18000 -9100 19600
rect -4690 19630 -4530 19730
rect -4690 19540 -4530 19630
<< metal3 >>
rect -5300 20900 -5000 21400
rect -5210 20860 -5000 20900
rect -4700 20900 -4400 21400
rect -4700 20860 -4450 20900
rect -5210 20840 -5010 20860
rect -5210 20580 -5190 20840
rect -5030 20580 -5010 20840
rect -5210 20560 -5010 20580
rect -4650 20840 -4450 20860
rect -4650 20580 -4630 20840
rect -4470 20580 -4450 20840
rect -4650 20560 -4450 20580
rect 5950 20500 11100 20600
rect -20400 19800 -15000 19900
rect -9500 19850 -8900 19900
rect -20400 15500 -20300 19800
rect -19700 15500 -15000 19800
rect -20400 15400 -15000 15500
rect -14800 19800 -14000 19850
rect -14800 15500 -14750 19800
rect -14050 15500 -14000 19800
rect -9500 17750 -9450 19850
rect -8900 17800 -8850 19800
rect -4700 19790 -4520 19800
rect -4700 19540 -4690 19790
rect -4530 19540 -4520 19790
rect -4700 19530 -4520 19540
rect -4900 19000 0 19450
rect -4900 18600 300 19000
rect -4900 18350 0 18600
rect -9500 17700 -8900 17750
rect -13600 17200 -12400 17400
rect -11350 17230 -11160 17240
rect -13600 15500 -13500 17200
rect -11350 17110 -11330 17230
rect -11170 17110 -11160 17230
rect -11350 17100 -11160 17110
rect -13400 16900 -12400 17100
rect -13400 15500 -13300 16900
rect -13200 16600 -12400 16800
rect -13200 15500 -13100 16600
rect -13000 16300 -12400 16500
rect -13000 15500 -12900 16300
rect -12800 16000 -12400 16200
rect 5950 16100 10350 20500
rect 10850 16100 11100 20500
rect 5950 16000 11100 16100
rect -12800 15500 -12700 16000
rect -14800 15450 -14000 15500
<< via3 >>
rect -20300 15500 -19700 19800
rect -14750 15500 -14050 19800
rect -9450 19600 -8900 19850
rect -9450 18000 -9100 19600
rect -9100 18000 -8900 19600
rect -9450 17750 -8900 18000
rect -4690 19730 -4530 19790
rect -4690 19540 -4530 19730
rect -11330 17110 -11170 17230
rect 10350 16100 10850 20500
<< mimcap >>
rect 6050 20400 10050 20500
rect -19200 19700 -15100 19800
rect -19200 15600 -19100 19700
rect -15200 15600 -15100 19700
rect -4850 19350 -50 19400
rect -4850 18450 -4800 19350
rect -100 18450 -50 19350
rect -4850 18400 -50 18450
rect 6050 16200 6150 20400
rect 9950 16200 10050 20400
rect 6050 16100 10050 16200
rect -19200 15500 -15100 15600
<< mimcapcontact >>
rect -19100 15600 -15200 19700
rect -4800 18450 -100 19350
rect 6150 16200 9950 20400
<< metal4 >>
rect 5950 20400 10150 20600
rect -20400 19800 -19600 19900
rect -20400 15500 -20300 19800
rect -19700 15500 -19600 19800
rect -20400 15400 -19600 15500
rect -19400 19850 -14800 19900
rect -9500 19850 -6500 19900
rect -19400 19800 -13900 19850
rect -19400 19700 -14750 19800
rect -19400 15600 -19100 19700
rect -15200 15600 -14750 19700
rect -19400 15500 -14750 15600
rect -14050 15500 -13900 19800
rect -9500 17750 -9450 19850
rect -8900 19800 -6500 19850
rect -8900 17750 -8700 19800
rect -9500 17700 -8700 17750
rect -11370 17230 -11130 17240
rect -11134 16990 -11130 17230
rect -11370 16980 -11130 16990
rect -8800 15600 -8700 17700
rect -6600 15600 -6500 19800
rect -4700 19790 -4520 19800
rect -4700 19540 -4690 19790
rect -4530 19540 -4520 19790
rect -4700 19400 -4520 19540
rect -4850 19350 -50 19400
rect -4850 18450 -4800 19350
rect -100 18450 -50 19350
rect -4850 18400 -50 18450
rect 5950 18200 6150 20400
rect 4150 17400 6150 18200
rect 1150 16300 2650 17400
rect 1100 15800 3100 16300
rect 5950 16200 6150 17400
rect 9950 16200 10150 20400
rect 5950 16000 10150 16200
rect 10250 20500 10950 20600
rect 10250 16100 10350 20500
rect 10850 16100 10950 20500
rect 10250 16000 10950 16100
rect -8800 15500 -6500 15600
rect -19400 15400 -13900 15500
<< via4 >>
rect -20300 15500 -19700 19800
rect -11370 17110 -11330 17230
rect -11330 17110 -11170 17230
rect -11170 17110 -11134 17230
rect -11370 16990 -11134 17110
rect -8700 15600 -6600 19800
rect 10350 16100 10850 20500
<< mimcap2 >>
rect 6050 20400 10050 20500
rect -19200 19700 -15100 19800
rect -19200 15600 -19100 19700
rect -15200 15600 -15100 19700
rect 6050 16200 6150 20400
rect 9950 16200 10050 20400
rect 6050 16100 10050 16200
rect -19200 15500 -15100 15600
<< mimcap2contact >>
rect -19100 15600 -15200 19700
rect 6150 16200 9950 20400
<< metal5 >>
rect 5950 20500 10950 20600
rect 5950 20400 10350 20500
rect -20400 19800 -15000 19900
rect -20400 15500 -20300 19800
rect -19700 19700 -15000 19800
rect -19700 15600 -19100 19700
rect -15200 15600 -15000 19700
rect -8900 19800 -6500 19900
rect -11700 17230 -10900 17350
rect -11700 16990 -11370 17230
rect -11134 16990 -10900 17230
rect -11700 16750 -10900 16990
rect -19700 15500 -15000 15600
rect -20400 15400 -15000 15500
rect -8900 15600 -8700 19800
rect -6600 18000 -6500 19800
rect -6600 16000 -5200 18000
rect 5950 16200 6150 20400
rect 9950 16200 10350 20400
rect 5950 16100 10350 16200
rect 10850 16100 10950 20500
rect 5950 16000 10950 16100
rect -8900 14500 -6900 15600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660275339
transform 1 0 -1100 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_1
timestamp 1660275339
transform 1 0 -1600 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_2
timestamp 1660275339
transform 1 0 -2100 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_3
timestamp 1660275339
transform 1 0 -2600 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_4
timestamp 1660275339
transform 1 0 -3100 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_5
timestamp 1660275339
transform 1 0 -3600 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_6
timestamp 1660275339
transform 1 0 -600 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_7
timestamp 1660275339
transform 1 0 -4100 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_8
timestamp 1660275339
transform 1 0 -4100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_9
timestamp 1660275339
transform 1 0 -3600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_10
timestamp 1660275339
transform 1 0 -3100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_11
timestamp 1660275339
transform 1 0 3400 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_12
timestamp 1660275339
transform 1 0 3900 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_13
timestamp 1660275339
transform 1 0 4400 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_14
timestamp 1660275339
transform 1 0 4900 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_15
timestamp 1660275339
transform 1 0 3900 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_16
timestamp 1660275339
transform 1 0 -100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_17
timestamp 1660275339
transform 1 0 400 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_18
timestamp 1660275339
transform 1 0 900 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_19
timestamp 1660275339
transform 1 0 1400 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_20
timestamp 1660275339
transform 1 0 1900 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_21
timestamp 1660275339
transform 1 0 2400 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_22
timestamp 1660275339
transform 1 0 2900 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_23
timestamp 1660275339
transform 1 0 4400 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_24
timestamp 1660275339
transform 1 0 3400 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_25
timestamp 1660275339
transform 1 0 4900 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_26
timestamp 1660275339
transform 1 0 3900 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_27
timestamp 1660275339
transform 1 0 4400 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_28
timestamp 1660275339
transform 1 0 3900 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_29
timestamp 1660275339
transform 1 0 4400 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_30
timestamp 1660275339
transform 1 0 4900 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_31
timestamp 1660275339
transform 1 0 3900 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_32
timestamp 1660275339
transform 1 0 4400 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_33
timestamp 1660275339
transform 1 0 4900 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_34
timestamp 1660275339
transform 1 0 3900 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_35
timestamp 1660275339
transform 1 0 4400 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_36
timestamp 1660275339
transform 1 0 4900 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_37
timestamp 1660275339
transform 1 0 4900 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_38
timestamp 1660275339
transform 1 0 -6100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_39
timestamp 1660275339
transform 1 0 -6100 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_40
timestamp 1660275339
transform 1 0 -6100 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_41
timestamp 1660275339
transform 1 0 -6100 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_42
timestamp 1660275339
transform 1 0 -6100 0 1 19300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_43
timestamp 1660275339
transform 1 0 -9100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_44
timestamp 1660275339
transform 1 0 -10600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_45
timestamp 1660275339
transform 1 0 -10100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_46
timestamp 1660275339
transform 1 0 -9600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_47
timestamp 1660275339
transform 1 0 -11100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_48
timestamp 1660275339
transform 1 0 -11600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_49
timestamp 1660275339
transform 1 0 -12100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_50
timestamp 1660275339
transform 1 0 -12600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_51
timestamp 1660275339
transform 1 0 -13600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_52
timestamp 1660275339
transform 1 0 -13100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_53
timestamp 1660275339
transform 1 0 -14100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_54
timestamp 1660275339
transform 1 0 -14600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_55
timestamp 1660275339
transform 1 0 -12100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_56
timestamp 1660275339
transform 1 0 -7100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_57
timestamp 1660275339
transform 1 0 -6600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_58
timestamp 1660275339
transform 1 0 -6100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_59
timestamp 1660275339
transform 1 0 -12600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_60
timestamp 1660275339
transform 1 0 -13600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_61
timestamp 1660275339
transform 1 0 -13100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_62
timestamp 1660275339
transform 1 0 -8600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_63
timestamp 1660275339
transform 1 0 -8100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_64
timestamp 1660275339
transform 1 0 -7600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_65
timestamp 1660275339
transform 1 0 -14100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_66
timestamp 1660275339
transform 1 0 -14600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_67
timestamp 1660275339
transform 1 0 -9100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_68
timestamp 1660275339
transform 1 0 -9600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_69
timestamp 1660275339
transform 1 0 -10600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_70
timestamp 1660275339
transform 1 0 -10100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_71
timestamp 1660275339
transform 1 0 -11100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_72
timestamp 1660275339
transform 1 0 -11600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_73
timestamp 1660275339
transform 1 0 -15600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_74
timestamp 1660275339
transform 1 0 -15100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_75
timestamp 1660275339
transform 1 0 -15100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_76
timestamp 1660275339
transform 1 0 -15600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_77
timestamp 1660275339
transform 1 0 -16600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_78
timestamp 1660275339
transform 1 0 -16100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_79
timestamp 1660275339
transform 1 0 -16100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_80
timestamp 1660275339
transform 1 0 -16600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_81
timestamp 1660275339
transform 1 0 -17600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_82
timestamp 1660275339
transform 1 0 -17100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_83
timestamp 1660275339
transform 1 0 -17100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_84
timestamp 1660275339
transform 1 0 -17600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_85
timestamp 1660275339
transform 1 0 -18600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_86
timestamp 1660275339
transform 1 0 -18100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_87
timestamp 1660275339
transform 1 0 -18100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_88
timestamp 1660275339
transform 1 0 -18600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_89
timestamp 1660275339
transform 1 0 -19600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_90
timestamp 1660275339
transform 1 0 -19100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_91
timestamp 1660275339
transform 1 0 -19100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_92
timestamp 1660275339
transform 1 0 -19600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_93
timestamp 1660275339
transform 1 0 -20600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_94
timestamp 1660275339
transform 1 0 -20100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_95
timestamp 1660275339
transform 1 0 -20100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_96
timestamp 1660275339
transform 1 0 -20600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_97
timestamp 1660275339
transform 1 0 -21600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_98
timestamp 1660275339
transform 1 0 -21100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_99
timestamp 1660275339
transform 1 0 -21100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_100
timestamp 1660275339
transform 1 0 -21600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_101
timestamp 1660275339
transform 1 0 -8100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_102
timestamp 1660275339
transform 1 0 -8600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_103
timestamp 1660275339
transform 1 0 -7600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_104
timestamp 1660275339
transform 1 0 -7100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_105
timestamp 1660275339
transform 1 0 -6600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_106
timestamp 1660275339
transform 1 0 -1600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_107
timestamp 1660275339
transform 1 0 -2600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_108
timestamp 1660275339
transform 1 0 -2100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_109
timestamp 1660275339
transform 1 0 -1100 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_110
timestamp 1660275339
transform 1 0 -600 0 1 21300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_111
timestamp 1660275339
transform 1 0 -3100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_112
timestamp 1660275339
transform 1 0 -4100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_113
timestamp 1660275339
transform 1 0 -3600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_114
timestamp 1660275339
transform 1 0 -1600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_115
timestamp 1660275339
transform 1 0 -2600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_116
timestamp 1660275339
transform 1 0 -2100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_117
timestamp 1660275339
transform 1 0 -100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_118
timestamp 1660275339
transform 1 0 -1100 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_119
timestamp 1660275339
transform 1 0 -600 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_120
timestamp 1660275339
transform 1 0 1400 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_121
timestamp 1660275339
transform 1 0 400 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_122
timestamp 1660275339
transform 1 0 900 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_123
timestamp 1660275339
transform 1 0 2900 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_124
timestamp 1660275339
transform 1 0 1900 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_125
timestamp 1660275339
transform 1 0 2400 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_126
timestamp 1660275339
transform 1 0 4400 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_127
timestamp 1660275339
transform 1 0 3900 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_128
timestamp 1660275339
transform 1 0 3400 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_129
timestamp 1660275339
transform 1 0 4900 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_130
timestamp 1660275339
transform 1 0 -600 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_131
timestamp 1660275339
transform 1 0 -1100 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_132
timestamp 1660275339
transform 1 0 -1600 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_133
timestamp 1660275339
transform 1 0 -600 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_134
timestamp 1660275339
transform 1 0 -1100 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_135
timestamp 1660275339
transform 1 0 -1600 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_136
timestamp 1660275339
transform 1 0 -21100 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_137
timestamp 1660275339
transform 1 0 -21600 0 1 20300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_138
timestamp 1660275339
transform 1 0 -21600 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_139
timestamp 1660275339
transform 1 0 -21100 0 1 20800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_140
timestamp 1660275339
transform 1 0 -21100 0 1 19300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_141
timestamp 1660275339
transform 1 0 -21600 0 1 19300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_142
timestamp 1660275339
transform 1 0 -21600 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_143
timestamp 1660275339
transform 1 0 -21100 0 1 19800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_144
timestamp 1660275339
transform 1 0 -21100 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_145
timestamp 1660275339
transform 1 0 -21600 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_146
timestamp 1660275339
transform 1 0 -21600 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_147
timestamp 1660275339
transform 1 0 -21100 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_148
timestamp 1660275339
transform 1 0 -21100 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_149
timestamp 1660275339
transform 1 0 -21600 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_150
timestamp 1660275339
transform 1 0 -21600 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_151
timestamp 1660275339
transform 1 0 -21100 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_152
timestamp 1660275339
transform 1 0 -21100 0 1 16300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_153
timestamp 1660275339
transform 1 0 -21600 0 1 16300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_154
timestamp 1660275339
transform 1 0 -21600 0 1 16800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_155
timestamp 1660275339
transform 1 0 -21100 0 1 16800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_156
timestamp 1660275339
transform 1 0 -21100 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_157
timestamp 1660275339
transform 1 0 -21600 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_158
timestamp 1660275339
transform 1 0 -21600 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_159
timestamp 1660275339
transform 1 0 -21100 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_160
timestamp 1660275339
transform 1 0 -20100 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_161
timestamp 1660275339
transform 1 0 -20600 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_162
timestamp 1660275339
transform 1 0 -20600 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_163
timestamp 1660275339
transform 1 0 -20100 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_164
timestamp 1660275339
transform 1 0 -19100 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_165
timestamp 1660275339
transform 1 0 -19600 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_166
timestamp 1660275339
transform 1 0 -19600 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_167
timestamp 1660275339
transform 1 0 -19100 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_168
timestamp 1660275339
transform 1 0 -18100 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_169
timestamp 1660275339
transform 1 0 -18600 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_170
timestamp 1660275339
transform 1 0 -18600 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_171
timestamp 1660275339
transform 1 0 -18100 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_172
timestamp 1660275339
transform 1 0 -17100 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_173
timestamp 1660275339
transform 1 0 -17600 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_174
timestamp 1660275339
transform 1 0 -17600 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_175
timestamp 1660275339
transform 1 0 -17100 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_176
timestamp 1660275339
transform 1 0 -16100 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_177
timestamp 1660275339
transform 1 0 -16600 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_178
timestamp 1660275339
transform 1 0 -16600 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_179
timestamp 1660275339
transform 1 0 -16100 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_180
timestamp 1660275339
transform 1 0 -15100 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_181
timestamp 1660275339
transform 1 0 -15600 0 1 15300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_182
timestamp 1660275339
transform 1 0 -15600 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_183
timestamp 1660275339
transform 1 0 -15100 0 1 15800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_184
timestamp 1660275339
transform 1 0 -1600 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_185
timestamp 1660275339
transform 1 0 -1100 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_186
timestamp 1660275339
transform 1 0 -600 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_187
timestamp 1660275339
transform 1 0 -600 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_188
timestamp 1660275339
transform 1 0 -1100 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_189
timestamp 1660275339
transform 1 0 -1600 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_190
timestamp 1660275339
transform 1 0 -3100 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_191
timestamp 1660275339
transform 1 0 -2600 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_192
timestamp 1660275339
transform 1 0 -2100 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_193
timestamp 1660275339
transform 1 0 -2100 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_194
timestamp 1660275339
transform 1 0 -2600 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_195
timestamp 1660275339
transform 1 0 -3100 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_196
timestamp 1660275339
transform 1 0 -3100 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_197
timestamp 1660275339
transform 1 0 -2600 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_198
timestamp 1660275339
transform 1 0 -2100 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_199
timestamp 1660275339
transform 1 0 -2100 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_200
timestamp 1660275339
transform 1 0 -2600 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_201
timestamp 1660275339
transform 1 0 -3100 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_202
timestamp 1660275339
transform 1 0 -3600 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_203
timestamp 1660275339
transform 1 0 -3600 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_204
timestamp 1660275339
transform 1 0 -3600 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_205
timestamp 1660275339
transform 1 0 -3600 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_206
timestamp 1660275339
transform 1 0 -4100 0 1 18800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_207
timestamp 1660275339
transform 1 0 -4100 0 1 18300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_208
timestamp 1660275339
transform 1 0 -4100 0 1 17800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_209
timestamp 1660275339
transform 1 0 -4100 0 1 17300
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_210
timestamp 1660275339
transform 1 0 5400 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_211
timestamp 1660275339
transform 1 0 5900 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_212
timestamp 1660275339
transform 1 0 6400 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_213
timestamp 1660275339
transform 1 0 6900 0 1 21800
box 100 -1100 600 -600
use hash_m1m2m3_W2p5L2p5  hash_m1m2m3_W2p5L2p5_214
timestamp 1660275339
transform 1 0 7400 0 1 21800
box 100 -1100 600 -600
use octal_ind_0p700n_5GHz  octal_ind_0p700n_5GHz_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1660787815
transform 0 -1 -20900 -1 0 -15900
box -33800 -32500 -8800 -7500
use pmirror_pfet_64x_complete  pmirror_pfet_64x_complete_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660185098
transform 0 1 -12800 -1 0 20150
box 0 0 4280 3344
use rfbcsa_1  rfbcsa_1_0
timestamp 1662654558
transform 1 0 600 0 1 18200
box -650 -800 3840 2000
use sky130_fd_pr__res_generic_po_3TQ83P  sky130_fd_pr__res_generic_po_3TQ83P_0
timestamp 1659923628
transform 1 0 -4826 0 1 20086
box -577 -589 577 589
<< labels >>
rlabel metal4 4150 17550 4450 18150 1 D
rlabel metal5 -11700 16750 -10900 17350 3 IREF
rlabel metal3 10900 16000 11100 20600 1 OUT
rlabel metal3 -5300 21200 -5000 21400 1 IN_DUMMY
rlabel metal3 -4700 21200 -4400 21400 1 IN
rlabel metal5 -20400 15400 -19600 19900 1 VLO
rlabel metal3 -12800 15500 -12700 15700 1 G8
rlabel metal3 -13000 15500 -12900 15700 1 G4
rlabel metal3 -13200 15500 -13100 15700 1 G2
rlabel metal3 -13400 15500 -13300 15700 1 G16
rlabel metal3 -13600 15500 -13500 15700 1 G32
rlabel metal4 -15000 15400 -13900 15500 1 VHI
<< end >>
