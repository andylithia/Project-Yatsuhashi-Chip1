magic
tech sky130B
magscale 1 2
timestamp 1659929390
<< pwell >>
rect -500 3412 714 3420
rect -500 3390 860 3412
rect -506 2319 870 3390
rect -506 2270 832 2319
rect 845 2270 870 2319
rect -506 2244 870 2270
rect -506 2230 -430 2244
rect -420 2230 870 2244
rect -500 2220 860 2230
<< psubdiff >>
rect -500 3354 -430 3390
rect -500 3320 -480 3354
rect -446 3320 -430 3354
rect -500 3284 -430 3320
rect -500 3250 -480 3284
rect -446 3250 -430 3284
rect -500 3214 -430 3250
rect -500 3180 -480 3214
rect -446 3180 -430 3214
rect -500 3144 -430 3180
rect -500 3110 -480 3144
rect -446 3110 -430 3144
rect -500 3074 -430 3110
rect -500 3040 -480 3074
rect -446 3040 -430 3074
rect -500 3004 -430 3040
rect -500 2970 -480 3004
rect -446 2970 -430 3004
rect -500 2934 -430 2970
rect -500 2900 -480 2934
rect -446 2900 -430 2934
rect -500 2864 -430 2900
rect -500 2830 -480 2864
rect -446 2830 -430 2864
rect -500 2794 -430 2830
rect -500 2760 -480 2794
rect -446 2760 -430 2794
rect -500 2724 -430 2760
rect -500 2690 -480 2724
rect -446 2690 -430 2724
rect -500 2654 -430 2690
rect -500 2620 -480 2654
rect -446 2620 -430 2654
rect -500 2584 -430 2620
rect -500 2550 -480 2584
rect -446 2550 -430 2584
rect -500 2514 -430 2550
rect -500 2480 -480 2514
rect -446 2480 -430 2514
rect -500 2444 -430 2480
rect -500 2410 -480 2444
rect -446 2410 -430 2444
rect -500 2374 -430 2410
rect -500 2340 -480 2374
rect -446 2340 -430 2374
rect -500 2310 -430 2340
rect 790 3354 870 3390
rect 790 3320 810 3354
rect 844 3320 870 3354
rect 790 3284 870 3320
rect 790 3250 810 3284
rect 844 3250 870 3284
rect 790 3214 870 3250
rect 790 3180 810 3214
rect 844 3180 870 3214
rect 790 3144 870 3180
rect 790 3110 810 3144
rect 844 3110 870 3144
rect 790 3074 870 3110
rect 790 3040 810 3074
rect 844 3040 870 3074
rect 790 3004 870 3040
rect 790 2970 810 3004
rect 844 2970 870 3004
rect 790 2934 870 2970
rect 790 2900 810 2934
rect 844 2900 870 2934
rect 790 2864 870 2900
rect 790 2830 810 2864
rect 844 2830 870 2864
rect 790 2794 870 2830
rect 790 2760 810 2794
rect 844 2760 870 2794
rect 790 2724 870 2760
rect 790 2690 810 2724
rect 844 2690 870 2724
rect 790 2654 870 2690
rect 790 2620 810 2654
rect 844 2620 870 2654
rect 790 2584 870 2620
rect 790 2550 810 2584
rect 844 2550 870 2584
rect 790 2514 870 2550
rect 790 2480 810 2514
rect 844 2480 870 2514
rect 790 2444 870 2480
rect 790 2410 810 2444
rect 844 2410 870 2444
rect 790 2374 870 2410
rect 790 2340 810 2374
rect 844 2340 870 2374
rect 790 2310 870 2340
rect -500 2284 870 2310
rect -500 2250 -400 2284
rect -366 2250 -330 2284
rect -296 2250 -260 2284
rect -226 2250 -190 2284
rect -156 2250 -120 2284
rect -86 2250 -50 2284
rect -16 2250 20 2284
rect 54 2250 90 2284
rect 124 2250 160 2284
rect 194 2250 230 2284
rect 264 2250 300 2284
rect 334 2250 370 2284
rect 404 2250 440 2284
rect 474 2250 510 2284
rect 544 2250 580 2284
rect 614 2250 650 2284
rect 684 2250 720 2284
rect 754 2250 870 2284
rect -500 2230 870 2250
<< psubdiffcont >>
rect -480 3320 -446 3354
rect -480 3250 -446 3284
rect -480 3180 -446 3214
rect -480 3110 -446 3144
rect -480 3040 -446 3074
rect -480 2970 -446 3004
rect -480 2900 -446 2934
rect -480 2830 -446 2864
rect -480 2760 -446 2794
rect -480 2690 -446 2724
rect -480 2620 -446 2654
rect -480 2550 -446 2584
rect -480 2480 -446 2514
rect -480 2410 -446 2444
rect -480 2340 -446 2374
rect 810 3320 844 3354
rect 810 3250 844 3284
rect 810 3180 844 3214
rect 810 3110 844 3144
rect 810 3040 844 3074
rect 810 2970 844 3004
rect 810 2900 844 2934
rect 810 2830 844 2864
rect 810 2760 844 2794
rect 810 2690 844 2724
rect 810 2620 844 2654
rect 810 2550 844 2584
rect 810 2480 844 2514
rect 810 2410 844 2444
rect 810 2340 844 2374
rect -400 2250 -366 2284
rect -330 2250 -296 2284
rect -260 2250 -226 2284
rect -190 2250 -156 2284
rect -120 2250 -86 2284
rect -50 2250 -16 2284
rect 20 2250 54 2284
rect 90 2250 124 2284
rect 160 2250 194 2284
rect 230 2250 264 2284
rect 300 2250 334 2284
rect 370 2250 404 2284
rect 440 2250 474 2284
rect 510 2250 544 2284
rect 580 2250 614 2284
rect 650 2250 684 2284
rect 720 2250 754 2284
<< poly >>
rect -5 3479 17 3483
rect -5 3417 24 3479
rect 2 3413 24 3417
<< polycont >>
rect -316 3429 -282 3463
rect -44 3429 -10 3463
rect 24 3429 58 3463
rect 300 3429 334 3463
rect 368 3429 402 3463
<< locali >>
rect -332 3429 -316 3463
rect -282 3429 -44 3463
rect -10 3429 24 3463
rect 58 3429 300 3463
rect 334 3429 368 3463
rect 402 3429 714 3463
rect -490 3354 -440 3370
rect -490 3320 -480 3354
rect -446 3320 -440 3354
rect -490 3284 -440 3320
rect -490 3240 -480 3284
rect -446 3240 -440 3284
rect -490 3214 -440 3240
rect -490 3160 -480 3214
rect -446 3160 -440 3214
rect -490 3144 -440 3160
rect -490 3080 -480 3144
rect -446 3080 -440 3144
rect -490 3074 -440 3080
rect -490 3040 -480 3074
rect -446 3040 -440 3074
rect -490 3034 -440 3040
rect -490 2970 -480 3034
rect -446 2970 -440 3034
rect -490 2954 -440 2970
rect -490 2900 -480 2954
rect -446 2900 -440 2954
rect -490 2874 -440 2900
rect -490 2830 -480 2874
rect -446 2830 -440 2874
rect -490 2794 -440 2830
rect -490 2760 -480 2794
rect -446 2760 -440 2794
rect -490 2724 -440 2760
rect -490 2680 -480 2724
rect -446 2680 -440 2724
rect -490 2654 -440 2680
rect -490 2600 -480 2654
rect -446 2600 -440 2654
rect -490 2584 -440 2600
rect -490 2520 -480 2584
rect -446 2520 -440 2584
rect -490 2514 -440 2520
rect -490 2480 -480 2514
rect -446 2480 -440 2514
rect -490 2474 -440 2480
rect -490 2410 -480 2474
rect -446 2410 -440 2474
rect -490 2394 -440 2410
rect -490 2340 -480 2394
rect -446 2340 -440 2394
rect -490 2300 -440 2340
rect 800 3354 860 3370
rect 800 3320 810 3354
rect 844 3320 860 3354
rect 800 3284 860 3320
rect 800 3240 810 3284
rect 844 3240 860 3284
rect 800 3214 860 3240
rect 800 3160 810 3214
rect 844 3160 860 3214
rect 800 3144 860 3160
rect 800 3080 810 3144
rect 844 3080 860 3144
rect 800 3074 860 3080
rect 800 3040 810 3074
rect 844 3040 860 3074
rect 800 3034 860 3040
rect 800 2970 810 3034
rect 844 2970 860 3034
rect 800 2954 860 2970
rect 800 2900 810 2954
rect 844 2900 860 2954
rect 800 2874 860 2900
rect 800 2830 810 2874
rect 844 2830 860 2874
rect 800 2794 860 2830
rect 800 2760 810 2794
rect 844 2760 860 2794
rect 800 2724 860 2760
rect 800 2680 810 2724
rect 844 2680 860 2724
rect 800 2654 860 2680
rect 800 2600 810 2654
rect 844 2600 860 2654
rect 800 2584 860 2600
rect 800 2520 810 2584
rect 844 2520 860 2584
rect 800 2514 860 2520
rect 800 2480 810 2514
rect 844 2480 860 2514
rect 800 2474 860 2480
rect 800 2410 810 2474
rect 844 2410 860 2474
rect 800 2394 860 2410
rect 800 2340 810 2394
rect 844 2340 860 2394
rect 800 2300 860 2340
rect -490 2284 860 2300
rect -490 2250 -400 2284
rect -356 2250 -330 2284
rect -276 2250 -260 2284
rect -196 2250 -190 2284
rect -156 2250 -150 2284
rect -86 2250 -70 2284
rect -16 2250 10 2284
rect 54 2250 90 2284
rect 124 2250 160 2284
rect 204 2250 230 2284
rect 284 2250 300 2284
rect 364 2250 370 2284
rect 404 2250 410 2284
rect 474 2250 490 2284
rect 544 2250 570 2284
rect 614 2250 650 2284
rect 684 2250 720 2284
rect 754 2250 860 2284
rect -490 2240 860 2250
<< viali >>
rect -480 3320 -446 3354
rect -480 3250 -446 3274
rect -480 3240 -446 3250
rect -480 3180 -446 3194
rect -480 3160 -446 3180
rect -480 3110 -446 3114
rect -480 3080 -446 3110
rect -480 3004 -446 3034
rect -480 3000 -446 3004
rect -480 2934 -446 2954
rect -480 2920 -446 2934
rect -480 2864 -446 2874
rect -480 2840 -446 2864
rect -480 2760 -446 2794
rect -480 2690 -446 2714
rect -480 2680 -446 2690
rect -480 2620 -446 2634
rect -480 2600 -446 2620
rect -480 2550 -446 2554
rect -480 2520 -446 2550
rect -480 2444 -446 2474
rect -480 2440 -446 2444
rect -480 2374 -446 2394
rect -480 2360 -446 2374
rect 810 3320 844 3354
rect 810 3250 844 3274
rect 810 3240 844 3250
rect 810 3180 844 3194
rect 810 3160 844 3180
rect 810 3110 844 3114
rect 810 3080 844 3110
rect 810 3004 844 3034
rect 810 3000 844 3004
rect 810 2934 844 2954
rect 810 2920 844 2934
rect 810 2864 844 2874
rect 810 2840 844 2864
rect 810 2760 844 2794
rect 810 2690 844 2714
rect 810 2680 844 2690
rect 810 2620 844 2634
rect 810 2600 844 2620
rect 810 2550 844 2554
rect 810 2520 844 2550
rect 810 2444 844 2474
rect 810 2440 844 2444
rect 810 2374 844 2394
rect 810 2360 844 2374
rect -390 2250 -366 2284
rect -366 2250 -356 2284
rect -310 2250 -296 2284
rect -296 2250 -276 2284
rect -230 2250 -226 2284
rect -226 2250 -196 2284
rect -150 2250 -120 2284
rect -120 2250 -116 2284
rect -70 2250 -50 2284
rect -50 2250 -36 2284
rect 10 2250 20 2284
rect 20 2250 44 2284
rect 90 2250 124 2284
rect 170 2250 194 2284
rect 194 2250 204 2284
rect 250 2250 264 2284
rect 264 2250 284 2284
rect 330 2250 334 2284
rect 334 2250 364 2284
rect 410 2250 440 2284
rect 440 2250 444 2284
rect 490 2250 510 2284
rect 510 2250 524 2284
rect 570 2250 580 2284
rect 580 2250 604 2284
rect 650 2250 684 2284
<< metal1 >>
rect -340 3520 710 3580
rect -5 3417 17 3483
rect -500 3380 -430 3390
rect 790 3380 860 3390
rect -500 3354 -310 3380
rect -500 3320 -480 3354
rect -446 3320 -310 3354
rect -500 3274 -310 3320
rect -500 3240 -480 3274
rect -446 3240 -310 3274
rect -500 3194 -310 3240
rect -500 3160 -480 3194
rect -446 3160 -310 3194
rect -500 3114 -310 3160
rect -500 3080 -480 3114
rect -446 3080 -310 3114
rect -500 3034 -310 3080
rect -500 3000 -480 3034
rect -446 3000 -310 3034
rect -500 2954 -310 3000
rect -500 2920 -480 2954
rect -446 2920 -310 2954
rect -500 2874 -310 2920
rect -500 2840 -480 2874
rect -446 2840 -310 2874
rect -500 2794 -310 2840
rect -500 2760 -480 2794
rect -446 2760 -310 2794
rect -500 2714 -310 2760
rect -500 2680 -480 2714
rect -446 2680 -310 2714
rect -500 2634 -310 2680
rect -500 2600 -480 2634
rect -446 2600 -310 2634
rect -500 2554 -310 2600
rect -500 2520 -480 2554
rect -446 2520 -310 2554
rect -500 2474 -310 2520
rect -500 2440 -480 2474
rect -446 2440 -310 2474
rect -500 2394 -310 2440
rect -500 2360 -480 2394
rect -446 2360 -310 2394
rect -500 2284 -310 2360
rect 680 3354 860 3380
rect 680 3320 810 3354
rect 844 3320 860 3354
rect 680 3274 860 3320
rect 680 3240 810 3274
rect 844 3240 860 3274
rect 680 3194 860 3240
rect 680 3160 810 3194
rect 844 3160 860 3194
rect 680 3114 860 3160
rect 680 3080 810 3114
rect 844 3080 860 3114
rect 680 3034 860 3080
rect 680 3000 810 3034
rect 844 3000 860 3034
rect 680 2954 860 3000
rect 680 2920 810 2954
rect 844 2920 860 2954
rect 680 2874 860 2920
rect 680 2840 810 2874
rect 844 2840 860 2874
rect 680 2794 860 2840
rect 680 2760 810 2794
rect 844 2760 860 2794
rect 680 2714 860 2760
rect 680 2680 810 2714
rect 844 2680 860 2714
rect 680 2634 860 2680
rect 680 2600 810 2634
rect 844 2600 860 2634
rect 680 2554 860 2600
rect 680 2520 810 2554
rect 844 2520 860 2554
rect 680 2474 860 2520
rect 680 2440 810 2474
rect 844 2440 860 2474
rect 680 2394 860 2440
rect 680 2360 810 2394
rect 844 2360 860 2394
rect 680 2284 860 2360
rect -500 2250 -390 2284
rect -356 2250 -310 2284
rect 684 2250 860 2284
rect -500 2230 860 2250
rect -490 2210 -370 2230
<< metal2 >>
rect -340 3420 730 3500
use sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap  sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_0
timestamp 1659107442
transform 1 0 -501 0 1 2289
box 100 -41 576 1290
use sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap  sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_1
timestamp 1659107442
transform 1 0 -157 0 1 2289
box 100 -41 576 1290
use sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap  sky130_fd_pr__rf_nfet_01v8_aM04_W5p00L0p15_notap_2
timestamp 1659107442
transform 1 0 187 0 1 2289
box 100 -41 576 1290
<< labels >>
rlabel metal1 -490 2210 -370 2230 1 S
rlabel metal1 -340 3520 -310 3580 1 G
rlabel metal2 -340 3420 -300 3500 1 SD
<< end >>
