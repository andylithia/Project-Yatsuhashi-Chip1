magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< locali >>
rect 70 282 136 316
rect 549 314 970 348
rect 70 174 136 208
rect 936 170 970 314
rect 1505 103 3722 137
<< metal1 >>
rect 246 -30 294 402
rect 670 -32 720 402
rect 1524 0 1552 395
rect 2972 0 3000 395
use sky130_fd_bd_sram__openram_dp_nand2_dec  sky130_fd_bd_sram__openram_dp_nand2_dec_0
timestamp 1661296025
transform 1 0 0 0 1 0
box 70 -56 888 476
use sky130_sram_1r1w_24x128_8_pinv_dec_0  sky130_sram_1r1w_24x128_8_pinv_dec_0_0
timestamp 1661296025
transform 1 0 876 0 1 0
box 44 0 2864 490
<< labels >>
rlabel locali s 2613 120 2613 120 4 Z
port 1 nsew
rlabel locali s 103 299 103 299 4 A
port 2 nsew
rlabel locali s 103 191 103 191 4 B
port 3 nsew
rlabel metal1 s 670 -32 720 402 4 vdd
port 4 nsew
rlabel metal1 s 2972 0 3000 395 4 vdd
port 4 nsew
rlabel metal1 s 1524 0 1552 395 4 gnd
port 5 nsew
rlabel metal1 s 246 -30 294 402 4 gnd
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 3722 395
<< end >>
