* SPICE3 file created from ./COMMON/mimcap_W1L5.ext - technology: sky130A

X0 top bot sky130_fd_pr__cap_mim_m3_1 l=1e+06u w=5e+06u
