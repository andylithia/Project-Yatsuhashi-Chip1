** sch_path: /home/andylithia/openmpw/Project-Yatsuhashi-Chip1/xschem/untitled-4.sch
**.subckt untitled-4
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1.26 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
V1 net1 GND 1.2
V2 net2 GND 1.2
**** begin user architecture code
.lib /home/andylithia/openmpw/pdk_1/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/andylithia/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.control
ac dec 10 1 10K
plot V(vmid) V(vin)

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
