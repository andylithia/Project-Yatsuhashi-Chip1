magic
tech sky130B
magscale 1 2
timestamp 1662185799
<< locali >>
rect 9740 103740 9860 103760
rect 9740 101420 9760 103740
rect 9840 101420 9860 103740
rect 9740 101400 9860 101420
<< viali >>
rect 9760 101420 9840 103740
<< metal1 >>
rect 14000 121900 58000 122000
rect 14000 121880 14120 121900
rect 14380 121880 14620 121900
rect 14880 121880 15120 121900
rect 15380 121880 15620 121900
rect 15880 121880 16120 121900
rect 16380 121880 16620 121900
rect 16880 121880 17120 121900
rect 17380 121880 17620 121900
rect 17880 121880 18120 121900
rect 18380 121880 18620 121900
rect 18880 121880 19120 121900
rect 19380 121880 19620 121900
rect 19880 121880 20120 121900
rect 20380 121880 20620 121900
rect 20880 121880 21120 121900
rect 21380 121880 21620 121900
rect 21880 121880 22120 121900
rect 22380 121880 22620 121900
rect 22880 121880 23120 121900
rect 23380 121880 23620 121900
rect 23880 121880 24120 121900
rect 24380 121880 24620 121900
rect 24880 121880 25120 121900
rect 25380 121880 25620 121900
rect 25880 121880 26120 121900
rect 26380 121880 26620 121900
rect 26880 121880 27120 121900
rect 27380 121880 27620 121900
rect 27880 121880 28120 121900
rect 28380 121880 28620 121900
rect 28880 121880 29120 121900
rect 29380 121880 29620 121900
rect 29880 121880 30120 121900
rect 30380 121880 30620 121900
rect 30880 121880 31120 121900
rect 31380 121880 31620 121900
rect 31880 121880 32120 121900
rect 32380 121880 32620 121900
rect 32880 121880 33120 121900
rect 33380 121880 33620 121900
rect 33880 121880 34120 121900
rect 34380 121880 34620 121900
rect 34880 121880 35120 121900
rect 35380 121880 35620 121900
rect 35880 121880 36120 121900
rect 36380 121880 36620 121900
rect 36880 121880 37120 121900
rect 37380 121880 37620 121900
rect 37880 121880 38120 121900
rect 38380 121880 38620 121900
rect 38880 121880 39120 121900
rect 39380 121880 39620 121900
rect 39880 121880 40120 121900
rect 40380 121880 40620 121900
rect 40880 121880 41120 121900
rect 41380 121880 41620 121900
rect 41880 121880 42120 121900
rect 42380 121880 42620 121900
rect 42880 121880 43120 121900
rect 43380 121880 43620 121900
rect 43880 121880 44120 121900
rect 44380 121880 44620 121900
rect 44880 121880 45120 121900
rect 45380 121880 45620 121900
rect 45880 121880 46120 121900
rect 46380 121880 46620 121900
rect 46880 121880 47120 121900
rect 47380 121880 47620 121900
rect 47880 121880 48120 121900
rect 48380 121880 48620 121900
rect 48880 121880 49120 121900
rect 49380 121880 49620 121900
rect 49880 121880 50120 121900
rect 50380 121880 50620 121900
rect 50880 121880 51120 121900
rect 51380 121880 51620 121900
rect 51880 121880 52120 121900
rect 52380 121880 52620 121900
rect 52880 121880 53120 121900
rect 53380 121880 53620 121900
rect 53880 121880 54120 121900
rect 54380 121880 54620 121900
rect 54880 121880 55120 121900
rect 55380 121880 55620 121900
rect 55880 121880 56120 121900
rect 56380 121880 56620 121900
rect 56880 121880 57120 121900
rect 57380 121880 57620 121900
rect 57880 121880 58000 121900
rect 14000 121620 14100 121880
rect 14400 121620 14600 121880
rect 14900 121620 15100 121880
rect 15400 121620 15600 121880
rect 15900 121620 16100 121880
rect 16400 121620 16600 121880
rect 16900 121620 17100 121880
rect 17400 121620 17600 121880
rect 17900 121620 18100 121880
rect 18400 121620 18600 121880
rect 18900 121620 19100 121880
rect 19400 121620 19600 121880
rect 19900 121620 20100 121880
rect 20400 121620 20600 121880
rect 20900 121620 21100 121880
rect 21400 121620 21600 121880
rect 21900 121620 22100 121880
rect 22400 121620 22600 121880
rect 22900 121620 23100 121880
rect 23400 121620 23600 121880
rect 23900 121620 24100 121880
rect 24400 121620 24600 121880
rect 24900 121620 25100 121880
rect 25400 121620 25600 121880
rect 25900 121620 26100 121880
rect 26400 121620 26600 121880
rect 26900 121620 27100 121880
rect 27400 121620 27600 121880
rect 27900 121620 28100 121880
rect 28400 121620 28600 121880
rect 28900 121620 29100 121880
rect 29400 121620 29600 121880
rect 29900 121620 30100 121880
rect 30400 121620 30600 121880
rect 30900 121620 31100 121880
rect 31400 121620 31600 121880
rect 31900 121620 32100 121880
rect 32400 121620 32600 121880
rect 32900 121620 33100 121880
rect 33400 121620 33600 121880
rect 33900 121620 34100 121880
rect 34400 121620 34600 121880
rect 34900 121620 35100 121880
rect 35400 121620 35600 121880
rect 35900 121620 36100 121880
rect 36400 121620 36600 121880
rect 36900 121620 37100 121880
rect 37400 121620 37600 121880
rect 37900 121620 38100 121880
rect 38400 121620 38600 121880
rect 38900 121620 39100 121880
rect 39400 121620 39600 121880
rect 39900 121620 40100 121880
rect 40400 121620 40600 121880
rect 40900 121620 41100 121880
rect 41400 121620 41600 121880
rect 41900 121620 42100 121880
rect 42400 121620 42600 121880
rect 42900 121620 43100 121880
rect 43400 121620 43600 121880
rect 43900 121620 44100 121880
rect 44400 121620 44600 121880
rect 44900 121620 45100 121880
rect 45400 121620 45600 121880
rect 45900 121620 46100 121880
rect 46400 121620 46600 121880
rect 46900 121620 47100 121880
rect 47400 121620 47600 121880
rect 47900 121620 48100 121880
rect 48400 121620 48600 121880
rect 48900 121620 49100 121880
rect 49400 121620 49600 121880
rect 49900 121620 50100 121880
rect 50400 121620 50600 121880
rect 50900 121620 51100 121880
rect 51400 121620 51600 121880
rect 51900 121620 52100 121880
rect 52400 121620 52600 121880
rect 52900 121620 53100 121880
rect 53400 121620 53600 121880
rect 53900 121620 54100 121880
rect 54400 121620 54600 121880
rect 54900 121620 55100 121880
rect 55400 121620 55600 121880
rect 55900 121620 56100 121880
rect 56400 121620 56600 121880
rect 56900 121620 57100 121880
rect 57400 121620 57600 121880
rect 57900 121620 58000 121880
rect 14000 121600 14120 121620
rect 14380 121600 14620 121620
rect 14880 121600 15120 121620
rect 15380 121600 15620 121620
rect 15880 121600 16120 121620
rect 16380 121600 16620 121620
rect 16880 121600 17120 121620
rect 17380 121600 17620 121620
rect 17880 121600 18120 121620
rect 18380 121600 18620 121620
rect 18880 121600 19120 121620
rect 19380 121600 19620 121620
rect 19880 121600 20120 121620
rect 20380 121600 20620 121620
rect 20880 121600 21120 121620
rect 21380 121600 21620 121620
rect 21880 121600 22120 121620
rect 22380 121600 22620 121620
rect 22880 121600 23120 121620
rect 23380 121600 23620 121620
rect 23880 121600 24120 121620
rect 24380 121600 24620 121620
rect 24880 121600 25120 121620
rect 25380 121600 25620 121620
rect 25880 121600 26120 121620
rect 26380 121600 26620 121620
rect 26880 121600 27120 121620
rect 27380 121600 27620 121620
rect 27880 121600 28120 121620
rect 28380 121600 28620 121620
rect 28880 121600 29120 121620
rect 29380 121600 29620 121620
rect 29880 121600 30120 121620
rect 30380 121600 30620 121620
rect 30880 121600 31120 121620
rect 31380 121600 31620 121620
rect 31880 121600 32120 121620
rect 32380 121600 32620 121620
rect 32880 121600 33120 121620
rect 33380 121600 33620 121620
rect 33880 121600 34120 121620
rect 34380 121600 34620 121620
rect 34880 121600 35120 121620
rect 35380 121600 35620 121620
rect 35880 121600 36120 121620
rect 36380 121600 36620 121620
rect 36880 121600 37120 121620
rect 37380 121600 37620 121620
rect 37880 121600 38120 121620
rect 38380 121600 38620 121620
rect 38880 121600 39120 121620
rect 39380 121600 39620 121620
rect 39880 121600 40120 121620
rect 40380 121600 40620 121620
rect 40880 121600 41120 121620
rect 41380 121600 41620 121620
rect 41880 121600 42120 121620
rect 42380 121600 42620 121620
rect 42880 121600 43120 121620
rect 43380 121600 43620 121620
rect 43880 121600 44120 121620
rect 44380 121600 44620 121620
rect 44880 121600 45120 121620
rect 45380 121600 45620 121620
rect 45880 121600 46120 121620
rect 46380 121600 46620 121620
rect 46880 121600 47120 121620
rect 47380 121600 47620 121620
rect 47880 121600 48120 121620
rect 48380 121600 48620 121620
rect 48880 121600 49120 121620
rect 49380 121600 49620 121620
rect 49880 121600 50120 121620
rect 50380 121600 50620 121620
rect 50880 121600 51120 121620
rect 51380 121600 51620 121620
rect 51880 121600 52120 121620
rect 52380 121600 52620 121620
rect 52880 121600 53120 121620
rect 53380 121600 53620 121620
rect 53880 121600 54120 121620
rect 54380 121600 54620 121620
rect 54880 121600 55120 121620
rect 55380 121600 55620 121620
rect 55880 121600 56120 121620
rect 56380 121600 56620 121620
rect 56880 121600 57120 121620
rect 57380 121600 57620 121620
rect 57880 121600 58000 121620
rect 14000 121400 58000 121600
rect 14000 121380 14120 121400
rect 14380 121380 14620 121400
rect 14880 121380 15120 121400
rect 15380 121380 15620 121400
rect 15880 121380 16120 121400
rect 16380 121380 16620 121400
rect 16880 121380 17120 121400
rect 17380 121380 17620 121400
rect 17880 121380 18120 121400
rect 18380 121380 18620 121400
rect 18880 121380 19120 121400
rect 19380 121380 19620 121400
rect 19880 121380 20120 121400
rect 20380 121380 20620 121400
rect 20880 121380 21120 121400
rect 21380 121380 21620 121400
rect 21880 121380 22120 121400
rect 22380 121380 22620 121400
rect 22880 121380 23120 121400
rect 23380 121380 23620 121400
rect 23880 121380 24120 121400
rect 24380 121380 24620 121400
rect 24880 121380 25120 121400
rect 25380 121380 25620 121400
rect 25880 121380 26120 121400
rect 26380 121380 26620 121400
rect 26880 121380 27120 121400
rect 27380 121380 27620 121400
rect 27880 121380 28120 121400
rect 28380 121380 28620 121400
rect 28880 121380 29120 121400
rect 29380 121380 29620 121400
rect 29880 121380 30120 121400
rect 30380 121380 30620 121400
rect 30880 121380 31120 121400
rect 31380 121380 31620 121400
rect 31880 121380 32120 121400
rect 32380 121380 32620 121400
rect 32880 121380 33120 121400
rect 33380 121380 33620 121400
rect 33880 121380 34120 121400
rect 34380 121380 34620 121400
rect 34880 121380 35120 121400
rect 35380 121380 35620 121400
rect 35880 121380 36120 121400
rect 36380 121380 36620 121400
rect 36880 121380 37120 121400
rect 37380 121380 37620 121400
rect 37880 121380 38120 121400
rect 38380 121380 38620 121400
rect 38880 121380 39120 121400
rect 39380 121380 39620 121400
rect 39880 121380 40120 121400
rect 40380 121380 40620 121400
rect 40880 121380 41120 121400
rect 41380 121380 41620 121400
rect 41880 121380 42120 121400
rect 42380 121380 42620 121400
rect 42880 121380 43120 121400
rect 43380 121380 43620 121400
rect 43880 121380 44120 121400
rect 44380 121380 44620 121400
rect 44880 121380 45120 121400
rect 45380 121380 45620 121400
rect 45880 121380 46120 121400
rect 46380 121380 46620 121400
rect 46880 121380 47120 121400
rect 47380 121380 47620 121400
rect 47880 121380 48120 121400
rect 48380 121380 48620 121400
rect 48880 121380 49120 121400
rect 49380 121380 49620 121400
rect 49880 121380 50120 121400
rect 50380 121380 50620 121400
rect 50880 121380 51120 121400
rect 51380 121380 51620 121400
rect 51880 121380 52120 121400
rect 52380 121380 52620 121400
rect 52880 121380 53120 121400
rect 53380 121380 53620 121400
rect 53880 121380 54120 121400
rect 54380 121380 54620 121400
rect 54880 121380 55120 121400
rect 55380 121380 55620 121400
rect 55880 121380 56120 121400
rect 56380 121380 56620 121400
rect 56880 121380 57120 121400
rect 57380 121380 57620 121400
rect 57880 121380 58000 121400
rect 14000 121120 14100 121380
rect 14400 121120 14600 121380
rect 14900 121120 15100 121380
rect 15400 121120 15600 121380
rect 15900 121120 16100 121380
rect 16400 121120 16600 121380
rect 16900 121120 17100 121380
rect 17400 121120 17600 121380
rect 17900 121120 18100 121380
rect 18400 121120 18600 121380
rect 18900 121120 19100 121380
rect 19400 121120 19600 121380
rect 19900 121120 20100 121380
rect 20400 121120 20600 121380
rect 20900 121120 21100 121380
rect 21400 121120 21600 121380
rect 21900 121120 22100 121380
rect 22400 121120 22600 121380
rect 22900 121120 23100 121380
rect 23400 121120 23600 121380
rect 23900 121120 24100 121380
rect 24400 121120 24600 121380
rect 24900 121120 25100 121380
rect 25400 121120 25600 121380
rect 25900 121120 26100 121380
rect 26400 121120 26600 121380
rect 26900 121120 27100 121380
rect 27400 121120 27600 121380
rect 27900 121120 28100 121380
rect 28400 121120 28600 121380
rect 28900 121120 29100 121380
rect 29400 121120 29600 121380
rect 29900 121120 30100 121380
rect 30400 121120 30600 121380
rect 30900 121120 31100 121380
rect 31400 121120 31600 121380
rect 31900 121120 32100 121380
rect 32400 121120 32600 121380
rect 32900 121120 33100 121380
rect 33400 121120 33600 121380
rect 33900 121120 34100 121380
rect 34400 121120 34600 121380
rect 34900 121120 35100 121380
rect 35400 121120 35600 121380
rect 35900 121120 36100 121380
rect 36400 121120 36600 121380
rect 36900 121120 37100 121380
rect 37400 121120 37600 121380
rect 37900 121120 38100 121380
rect 38400 121120 38600 121380
rect 38900 121120 39100 121380
rect 39400 121120 39600 121380
rect 39900 121120 40100 121380
rect 40400 121120 40600 121380
rect 40900 121120 41100 121380
rect 41400 121120 41600 121380
rect 41900 121120 42100 121380
rect 42400 121120 42600 121380
rect 42900 121120 43100 121380
rect 43400 121120 43600 121380
rect 43900 121120 44100 121380
rect 44400 121120 44600 121380
rect 44900 121120 45100 121380
rect 45400 121120 45600 121380
rect 45900 121120 46100 121380
rect 46400 121120 46600 121380
rect 46900 121120 47100 121380
rect 47400 121120 47600 121380
rect 47900 121120 48100 121380
rect 48400 121120 48600 121380
rect 48900 121120 49100 121380
rect 49400 121120 49600 121380
rect 49900 121120 50100 121380
rect 50400 121120 50600 121380
rect 50900 121120 51100 121380
rect 51400 121120 51600 121380
rect 51900 121120 52100 121380
rect 52400 121120 52600 121380
rect 52900 121120 53100 121380
rect 53400 121120 53600 121380
rect 53900 121120 54100 121380
rect 54400 121120 54600 121380
rect 54900 121120 55100 121380
rect 55400 121120 55600 121380
rect 55900 121120 56100 121380
rect 56400 121120 56600 121380
rect 56900 121120 57100 121380
rect 57400 121120 57600 121380
rect 57900 121120 58000 121380
rect 14000 121100 14120 121120
rect 14380 121100 14620 121120
rect 14880 121100 15120 121120
rect 15380 121100 15620 121120
rect 15880 121100 16120 121120
rect 16380 121100 16620 121120
rect 16880 121100 17120 121120
rect 17380 121100 17620 121120
rect 17880 121100 18120 121120
rect 18380 121100 18620 121120
rect 18880 121100 19120 121120
rect 19380 121100 19620 121120
rect 19880 121100 20120 121120
rect 20380 121100 20620 121120
rect 20880 121100 21120 121120
rect 21380 121100 21620 121120
rect 21880 121100 22120 121120
rect 22380 121100 22620 121120
rect 22880 121100 23120 121120
rect 23380 121100 23620 121120
rect 23880 121100 24120 121120
rect 24380 121100 24620 121120
rect 24880 121100 25120 121120
rect 25380 121100 25620 121120
rect 25880 121100 26120 121120
rect 26380 121100 26620 121120
rect 26880 121100 27120 121120
rect 27380 121100 27620 121120
rect 27880 121100 28120 121120
rect 28380 121100 28620 121120
rect 28880 121100 29120 121120
rect 29380 121100 29620 121120
rect 29880 121100 30120 121120
rect 30380 121100 30620 121120
rect 30880 121100 31120 121120
rect 31380 121100 31620 121120
rect 31880 121100 32120 121120
rect 32380 121100 32620 121120
rect 32880 121100 33120 121120
rect 33380 121100 33620 121120
rect 33880 121100 34120 121120
rect 34380 121100 34620 121120
rect 34880 121100 35120 121120
rect 35380 121100 35620 121120
rect 35880 121100 36120 121120
rect 36380 121100 36620 121120
rect 36880 121100 37120 121120
rect 37380 121100 37620 121120
rect 37880 121100 38120 121120
rect 38380 121100 38620 121120
rect 38880 121100 39120 121120
rect 39380 121100 39620 121120
rect 39880 121100 40120 121120
rect 40380 121100 40620 121120
rect 40880 121100 41120 121120
rect 41380 121100 41620 121120
rect 41880 121100 42120 121120
rect 42380 121100 42620 121120
rect 42880 121100 43120 121120
rect 43380 121100 43620 121120
rect 43880 121100 44120 121120
rect 44380 121100 44620 121120
rect 44880 121100 45120 121120
rect 45380 121100 45620 121120
rect 45880 121100 46120 121120
rect 46380 121100 46620 121120
rect 46880 121100 47120 121120
rect 47380 121100 47620 121120
rect 47880 121100 48120 121120
rect 48380 121100 48620 121120
rect 48880 121100 49120 121120
rect 49380 121100 49620 121120
rect 49880 121100 50120 121120
rect 50380 121100 50620 121120
rect 50880 121100 51120 121120
rect 51380 121100 51620 121120
rect 51880 121100 52120 121120
rect 52380 121100 52620 121120
rect 52880 121100 53120 121120
rect 53380 121100 53620 121120
rect 53880 121100 54120 121120
rect 54380 121100 54620 121120
rect 54880 121100 55120 121120
rect 55380 121100 55620 121120
rect 55880 121100 56120 121120
rect 56380 121100 56620 121120
rect 56880 121100 57120 121120
rect 57380 121100 57620 121120
rect 57880 121100 58000 121120
rect 14000 120900 58000 121100
rect 14000 120880 14120 120900
rect 14380 120880 14620 120900
rect 14880 120880 15120 120900
rect 15380 120880 15620 120900
rect 15880 120880 16120 120900
rect 16380 120880 16620 120900
rect 16880 120880 17120 120900
rect 17380 120880 17620 120900
rect 17880 120880 18120 120900
rect 18380 120880 18620 120900
rect 18880 120880 19120 120900
rect 19380 120880 19620 120900
rect 19880 120880 20120 120900
rect 20380 120880 20620 120900
rect 20880 120880 21120 120900
rect 21380 120880 21620 120900
rect 21880 120880 22120 120900
rect 22380 120880 22620 120900
rect 22880 120880 23120 120900
rect 23380 120880 23620 120900
rect 23880 120880 24120 120900
rect 24380 120880 24620 120900
rect 24880 120880 25120 120900
rect 25380 120880 25620 120900
rect 25880 120880 26120 120900
rect 26380 120880 26620 120900
rect 26880 120880 27120 120900
rect 27380 120880 27620 120900
rect 27880 120880 28120 120900
rect 28380 120880 28620 120900
rect 28880 120880 29120 120900
rect 29380 120880 29620 120900
rect 29880 120880 30120 120900
rect 30380 120880 30620 120900
rect 30880 120880 31120 120900
rect 31380 120880 31620 120900
rect 31880 120880 32120 120900
rect 32380 120880 32620 120900
rect 32880 120880 33120 120900
rect 33380 120880 33620 120900
rect 33880 120880 34120 120900
rect 34380 120880 34620 120900
rect 34880 120880 35120 120900
rect 35380 120880 35620 120900
rect 35880 120880 36120 120900
rect 36380 120880 36620 120900
rect 36880 120880 37120 120900
rect 37380 120880 37620 120900
rect 37880 120880 38120 120900
rect 38380 120880 38620 120900
rect 38880 120880 39120 120900
rect 39380 120880 39620 120900
rect 39880 120880 40120 120900
rect 40380 120880 40620 120900
rect 40880 120880 41120 120900
rect 41380 120880 41620 120900
rect 41880 120880 42120 120900
rect 42380 120880 42620 120900
rect 42880 120880 43120 120900
rect 43380 120880 43620 120900
rect 43880 120880 44120 120900
rect 44380 120880 44620 120900
rect 44880 120880 45120 120900
rect 45380 120880 45620 120900
rect 45880 120880 46120 120900
rect 46380 120880 46620 120900
rect 46880 120880 47120 120900
rect 47380 120880 47620 120900
rect 47880 120880 48120 120900
rect 48380 120880 48620 120900
rect 48880 120880 49120 120900
rect 49380 120880 49620 120900
rect 49880 120880 50120 120900
rect 50380 120880 50620 120900
rect 50880 120880 51120 120900
rect 51380 120880 51620 120900
rect 51880 120880 52120 120900
rect 52380 120880 52620 120900
rect 52880 120880 53120 120900
rect 53380 120880 53620 120900
rect 53880 120880 54120 120900
rect 54380 120880 54620 120900
rect 54880 120880 55120 120900
rect 55380 120880 55620 120900
rect 55880 120880 56120 120900
rect 56380 120880 56620 120900
rect 56880 120880 57120 120900
rect 57380 120880 57620 120900
rect 57880 120880 58000 120900
rect 14000 120620 14100 120880
rect 14400 120620 14600 120880
rect 14900 120620 15100 120880
rect 15400 120620 15600 120880
rect 15900 120620 16100 120880
rect 16400 120620 16600 120880
rect 16900 120620 17100 120880
rect 17400 120620 17600 120880
rect 17900 120620 18100 120880
rect 18400 120620 18600 120880
rect 18900 120620 19100 120880
rect 19400 120620 19600 120880
rect 19900 120620 20100 120880
rect 20400 120620 20600 120880
rect 20900 120620 21100 120880
rect 21400 120620 21600 120880
rect 21900 120620 22100 120880
rect 22400 120620 22600 120880
rect 22900 120620 23100 120880
rect 23400 120620 23600 120880
rect 23900 120620 24100 120880
rect 24400 120620 24600 120880
rect 24900 120620 25100 120880
rect 25400 120620 25600 120880
rect 25900 120620 26100 120880
rect 26400 120620 26600 120880
rect 26900 120620 27100 120880
rect 27400 120620 27600 120880
rect 27900 120620 28100 120880
rect 28400 120620 28600 120880
rect 28900 120620 29100 120880
rect 29400 120620 29600 120880
rect 29900 120620 30100 120880
rect 30400 120620 30600 120880
rect 30900 120620 31100 120880
rect 31400 120620 31600 120880
rect 31900 120620 32100 120880
rect 32400 120620 32600 120880
rect 32900 120620 33100 120880
rect 33400 120620 33600 120880
rect 33900 120620 34100 120880
rect 34400 120620 34600 120880
rect 34900 120620 35100 120880
rect 35400 120620 35600 120880
rect 35900 120620 36100 120880
rect 36400 120620 36600 120880
rect 36900 120620 37100 120880
rect 37400 120620 37600 120880
rect 37900 120620 38100 120880
rect 38400 120620 38600 120880
rect 38900 120620 39100 120880
rect 39400 120620 39600 120880
rect 39900 120620 40100 120880
rect 40400 120620 40600 120880
rect 40900 120620 41100 120880
rect 41400 120620 41600 120880
rect 41900 120620 42100 120880
rect 42400 120620 42600 120880
rect 42900 120620 43100 120880
rect 43400 120620 43600 120880
rect 43900 120620 44100 120880
rect 44400 120620 44600 120880
rect 44900 120620 45100 120880
rect 45400 120620 45600 120880
rect 45900 120620 46100 120880
rect 46400 120620 46600 120880
rect 46900 120620 47100 120880
rect 47400 120620 47600 120880
rect 47900 120620 48100 120880
rect 48400 120620 48600 120880
rect 48900 120620 49100 120880
rect 49400 120620 49600 120880
rect 49900 120620 50100 120880
rect 50400 120620 50600 120880
rect 50900 120620 51100 120880
rect 51400 120620 51600 120880
rect 51900 120620 52100 120880
rect 52400 120620 52600 120880
rect 52900 120620 53100 120880
rect 53400 120620 53600 120880
rect 53900 120620 54100 120880
rect 54400 120620 54600 120880
rect 54900 120620 55100 120880
rect 55400 120620 55600 120880
rect 55900 120620 56100 120880
rect 56400 120620 56600 120880
rect 56900 120620 57100 120880
rect 57400 120620 57600 120880
rect 57900 120620 58000 120880
rect 14000 120600 14120 120620
rect 14380 120600 14620 120620
rect 14880 120600 15120 120620
rect 15380 120600 15620 120620
rect 15880 120600 16120 120620
rect 16380 120600 16620 120620
rect 16880 120600 17120 120620
rect 17380 120600 17620 120620
rect 17880 120600 18120 120620
rect 18380 120600 18620 120620
rect 18880 120600 19120 120620
rect 19380 120600 19620 120620
rect 19880 120600 20120 120620
rect 20380 120600 20620 120620
rect 20880 120600 21120 120620
rect 21380 120600 21620 120620
rect 21880 120600 22120 120620
rect 22380 120600 22620 120620
rect 22880 120600 23120 120620
rect 23380 120600 23620 120620
rect 23880 120600 24120 120620
rect 24380 120600 24620 120620
rect 24880 120600 25120 120620
rect 25380 120600 25620 120620
rect 25880 120600 26120 120620
rect 26380 120600 26620 120620
rect 26880 120600 27120 120620
rect 27380 120600 27620 120620
rect 27880 120600 28120 120620
rect 28380 120600 28620 120620
rect 28880 120600 29120 120620
rect 29380 120600 29620 120620
rect 29880 120600 30120 120620
rect 30380 120600 30620 120620
rect 30880 120600 31120 120620
rect 31380 120600 31620 120620
rect 31880 120600 32120 120620
rect 32380 120600 32620 120620
rect 32880 120600 33120 120620
rect 33380 120600 33620 120620
rect 33880 120600 34120 120620
rect 34380 120600 34620 120620
rect 34880 120600 35120 120620
rect 35380 120600 35620 120620
rect 35880 120600 36120 120620
rect 36380 120600 36620 120620
rect 36880 120600 37120 120620
rect 37380 120600 37620 120620
rect 37880 120600 38120 120620
rect 38380 120600 38620 120620
rect 38880 120600 39120 120620
rect 39380 120600 39620 120620
rect 39880 120600 40120 120620
rect 40380 120600 40620 120620
rect 40880 120600 41120 120620
rect 41380 120600 41620 120620
rect 41880 120600 42120 120620
rect 42380 120600 42620 120620
rect 42880 120600 43120 120620
rect 43380 120600 43620 120620
rect 43880 120600 44120 120620
rect 44380 120600 44620 120620
rect 44880 120600 45120 120620
rect 45380 120600 45620 120620
rect 45880 120600 46120 120620
rect 46380 120600 46620 120620
rect 46880 120600 47120 120620
rect 47380 120600 47620 120620
rect 47880 120600 48120 120620
rect 48380 120600 48620 120620
rect 48880 120600 49120 120620
rect 49380 120600 49620 120620
rect 49880 120600 50120 120620
rect 50380 120600 50620 120620
rect 50880 120600 51120 120620
rect 51380 120600 51620 120620
rect 51880 120600 52120 120620
rect 52380 120600 52620 120620
rect 52880 120600 53120 120620
rect 53380 120600 53620 120620
rect 53880 120600 54120 120620
rect 54380 120600 54620 120620
rect 54880 120600 55120 120620
rect 55380 120600 55620 120620
rect 55880 120600 56120 120620
rect 56380 120600 56620 120620
rect 56880 120600 57120 120620
rect 57380 120600 57620 120620
rect 57880 120600 58000 120620
rect 14000 120400 58000 120600
rect 14000 120380 14120 120400
rect 14380 120380 14620 120400
rect 14880 120380 15120 120400
rect 15380 120380 15620 120400
rect 15880 120380 16120 120400
rect 16380 120380 16620 120400
rect 16880 120380 17120 120400
rect 17380 120380 17620 120400
rect 17880 120380 18120 120400
rect 18380 120380 18620 120400
rect 18880 120380 19120 120400
rect 19380 120380 19620 120400
rect 19880 120380 20120 120400
rect 20380 120380 20620 120400
rect 20880 120380 21120 120400
rect 21380 120380 21620 120400
rect 21880 120380 22120 120400
rect 22380 120380 22620 120400
rect 22880 120380 23120 120400
rect 23380 120380 23620 120400
rect 23880 120380 24120 120400
rect 24380 120380 24620 120400
rect 24880 120380 25120 120400
rect 25380 120380 25620 120400
rect 25880 120380 26120 120400
rect 26380 120380 26620 120400
rect 26880 120380 27120 120400
rect 27380 120380 27620 120400
rect 27880 120380 28120 120400
rect 28380 120380 28620 120400
rect 28880 120380 29120 120400
rect 29380 120380 29620 120400
rect 29880 120380 30120 120400
rect 30380 120380 30620 120400
rect 30880 120380 31120 120400
rect 31380 120380 31620 120400
rect 31880 120380 32120 120400
rect 32380 120380 32620 120400
rect 32880 120380 33120 120400
rect 33380 120380 33620 120400
rect 33880 120380 34120 120400
rect 34380 120380 34620 120400
rect 34880 120380 35120 120400
rect 35380 120380 35620 120400
rect 35880 120380 36120 120400
rect 36380 120380 36620 120400
rect 36880 120380 37120 120400
rect 37380 120380 37620 120400
rect 37880 120380 38120 120400
rect 38380 120380 38620 120400
rect 38880 120380 39120 120400
rect 39380 120380 39620 120400
rect 39880 120380 40120 120400
rect 40380 120380 40620 120400
rect 40880 120380 41120 120400
rect 41380 120380 41620 120400
rect 41880 120380 42120 120400
rect 42380 120380 42620 120400
rect 42880 120380 43120 120400
rect 43380 120380 43620 120400
rect 43880 120380 44120 120400
rect 44380 120380 44620 120400
rect 44880 120380 45120 120400
rect 45380 120380 45620 120400
rect 45880 120380 46120 120400
rect 46380 120380 46620 120400
rect 46880 120380 47120 120400
rect 47380 120380 47620 120400
rect 47880 120380 48120 120400
rect 48380 120380 48620 120400
rect 48880 120380 49120 120400
rect 49380 120380 49620 120400
rect 49880 120380 50120 120400
rect 50380 120380 50620 120400
rect 50880 120380 51120 120400
rect 51380 120380 51620 120400
rect 51880 120380 52120 120400
rect 52380 120380 52620 120400
rect 52880 120380 53120 120400
rect 53380 120380 53620 120400
rect 53880 120380 54120 120400
rect 54380 120380 54620 120400
rect 54880 120380 55120 120400
rect 55380 120380 55620 120400
rect 55880 120380 56120 120400
rect 56380 120380 56620 120400
rect 56880 120380 57120 120400
rect 57380 120380 57620 120400
rect 57880 120380 58000 120400
rect 14000 120120 14100 120380
rect 14400 120120 14600 120380
rect 14900 120120 15100 120380
rect 15400 120120 15600 120380
rect 15900 120120 16100 120380
rect 16400 120120 16600 120380
rect 16900 120120 17100 120380
rect 17400 120120 17600 120380
rect 17900 120120 18100 120380
rect 18400 120120 18600 120380
rect 18900 120120 19100 120380
rect 19400 120120 19600 120380
rect 19900 120120 20100 120380
rect 20400 120120 20600 120380
rect 20900 120120 21100 120380
rect 21400 120120 21600 120380
rect 21900 120120 22100 120380
rect 22400 120120 22600 120380
rect 22900 120120 23100 120380
rect 23400 120120 23600 120380
rect 23900 120120 24100 120380
rect 24400 120120 24600 120380
rect 24900 120120 25100 120380
rect 25400 120120 25600 120380
rect 25900 120120 26100 120380
rect 26400 120120 26600 120380
rect 26900 120120 27100 120380
rect 27400 120120 27600 120380
rect 27900 120120 28100 120380
rect 28400 120120 28600 120380
rect 28900 120120 29100 120380
rect 29400 120120 29600 120380
rect 29900 120120 30100 120380
rect 30400 120120 30600 120380
rect 30900 120120 31100 120380
rect 31400 120120 31600 120380
rect 31900 120120 32100 120380
rect 32400 120120 32600 120380
rect 32900 120120 33100 120380
rect 33400 120120 33600 120380
rect 33900 120120 34100 120380
rect 34400 120120 34600 120380
rect 34900 120120 35100 120380
rect 35400 120120 35600 120380
rect 35900 120120 36100 120380
rect 36400 120120 36600 120380
rect 36900 120120 37100 120380
rect 37400 120120 37600 120380
rect 37900 120120 38100 120380
rect 38400 120120 38600 120380
rect 38900 120120 39100 120380
rect 39400 120120 39600 120380
rect 39900 120120 40100 120380
rect 40400 120120 40600 120380
rect 40900 120120 41100 120380
rect 41400 120120 41600 120380
rect 41900 120120 42100 120380
rect 42400 120120 42600 120380
rect 42900 120120 43100 120380
rect 43400 120120 43600 120380
rect 43900 120120 44100 120380
rect 44400 120120 44600 120380
rect 44900 120120 45100 120380
rect 45400 120120 45600 120380
rect 45900 120120 46100 120380
rect 46400 120120 46600 120380
rect 46900 120120 47100 120380
rect 47400 120120 47600 120380
rect 47900 120120 48100 120380
rect 48400 120120 48600 120380
rect 48900 120120 49100 120380
rect 49400 120120 49600 120380
rect 49900 120120 50100 120380
rect 50400 120120 50600 120380
rect 50900 120120 51100 120380
rect 51400 120120 51600 120380
rect 51900 120120 52100 120380
rect 52400 120120 52600 120380
rect 52900 120120 53100 120380
rect 53400 120120 53600 120380
rect 53900 120120 54100 120380
rect 54400 120120 54600 120380
rect 54900 120120 55100 120380
rect 55400 120120 55600 120380
rect 55900 120120 56100 120380
rect 56400 120120 56600 120380
rect 56900 120120 57100 120380
rect 57400 120120 57600 120380
rect 57900 120120 58000 120380
rect 14000 120100 14120 120120
rect 14380 120100 14620 120120
rect 14880 120100 15120 120120
rect 15380 120100 15620 120120
rect 15880 120100 16120 120120
rect 16380 120100 16620 120120
rect 16880 120100 17120 120120
rect 17380 120100 17620 120120
rect 17880 120100 18120 120120
rect 18380 120100 18620 120120
rect 18880 120100 19120 120120
rect 19380 120100 19620 120120
rect 19880 120100 20120 120120
rect 20380 120100 20620 120120
rect 20880 120100 21120 120120
rect 21380 120100 21620 120120
rect 21880 120100 22120 120120
rect 22380 120100 22620 120120
rect 22880 120100 23120 120120
rect 23380 120100 23620 120120
rect 23880 120100 24120 120120
rect 24380 120100 24620 120120
rect 24880 120100 25120 120120
rect 25380 120100 25620 120120
rect 25880 120100 26120 120120
rect 26380 120100 26620 120120
rect 26880 120100 27120 120120
rect 27380 120100 27620 120120
rect 27880 120100 28120 120120
rect 28380 120100 28620 120120
rect 28880 120100 29120 120120
rect 29380 120100 29620 120120
rect 29880 120100 30120 120120
rect 30380 120100 30620 120120
rect 30880 120100 31120 120120
rect 31380 120100 31620 120120
rect 31880 120100 32120 120120
rect 32380 120100 32620 120120
rect 32880 120100 33120 120120
rect 33380 120100 33620 120120
rect 33880 120100 34120 120120
rect 34380 120100 34620 120120
rect 34880 120100 35120 120120
rect 35380 120100 35620 120120
rect 35880 120100 36120 120120
rect 36380 120100 36620 120120
rect 36880 120100 37120 120120
rect 37380 120100 37620 120120
rect 37880 120100 38120 120120
rect 38380 120100 38620 120120
rect 38880 120100 39120 120120
rect 39380 120100 39620 120120
rect 39880 120100 40120 120120
rect 40380 120100 40620 120120
rect 40880 120100 41120 120120
rect 41380 120100 41620 120120
rect 41880 120100 42120 120120
rect 42380 120100 42620 120120
rect 42880 120100 43120 120120
rect 43380 120100 43620 120120
rect 43880 120100 44120 120120
rect 44380 120100 44620 120120
rect 44880 120100 45120 120120
rect 45380 120100 45620 120120
rect 45880 120100 46120 120120
rect 46380 120100 46620 120120
rect 46880 120100 47120 120120
rect 47380 120100 47620 120120
rect 47880 120100 48120 120120
rect 48380 120100 48620 120120
rect 48880 120100 49120 120120
rect 49380 120100 49620 120120
rect 49880 120100 50120 120120
rect 50380 120100 50620 120120
rect 50880 120100 51120 120120
rect 51380 120100 51620 120120
rect 51880 120100 52120 120120
rect 52380 120100 52620 120120
rect 52880 120100 53120 120120
rect 53380 120100 53620 120120
rect 53880 120100 54120 120120
rect 54380 120100 54620 120120
rect 54880 120100 55120 120120
rect 55380 120100 55620 120120
rect 55880 120100 56120 120120
rect 56380 120100 56620 120120
rect 56880 120100 57120 120120
rect 57380 120100 57620 120120
rect 57880 120100 58000 120120
rect 14000 119900 58000 120100
rect 14000 119880 14120 119900
rect 14380 119880 14620 119900
rect 14880 119880 15120 119900
rect 15380 119880 15620 119900
rect 15880 119880 16120 119900
rect 16380 119880 16620 119900
rect 16880 119880 17120 119900
rect 17380 119880 17620 119900
rect 17880 119880 18120 119900
rect 18380 119880 18620 119900
rect 18880 119880 19120 119900
rect 19380 119880 19620 119900
rect 19880 119880 20120 119900
rect 20380 119880 20620 119900
rect 20880 119880 21120 119900
rect 21380 119880 21620 119900
rect 21880 119880 22120 119900
rect 22380 119880 22620 119900
rect 22880 119880 23120 119900
rect 23380 119880 23620 119900
rect 23880 119880 24120 119900
rect 24380 119880 24620 119900
rect 24880 119880 25120 119900
rect 25380 119880 25620 119900
rect 25880 119880 26120 119900
rect 26380 119880 26620 119900
rect 26880 119880 27120 119900
rect 27380 119880 27620 119900
rect 27880 119880 28120 119900
rect 28380 119880 28620 119900
rect 28880 119880 29120 119900
rect 29380 119880 29620 119900
rect 29880 119880 30120 119900
rect 30380 119880 30620 119900
rect 30880 119880 31120 119900
rect 31380 119880 31620 119900
rect 31880 119880 32120 119900
rect 32380 119880 32620 119900
rect 32880 119880 33120 119900
rect 33380 119880 33620 119900
rect 33880 119880 34120 119900
rect 34380 119880 34620 119900
rect 34880 119880 35120 119900
rect 35380 119880 35620 119900
rect 35880 119880 36120 119900
rect 36380 119880 36620 119900
rect 36880 119880 37120 119900
rect 37380 119880 37620 119900
rect 37880 119880 38120 119900
rect 38380 119880 38620 119900
rect 38880 119880 39120 119900
rect 39380 119880 39620 119900
rect 39880 119880 40120 119900
rect 40380 119880 40620 119900
rect 40880 119880 41120 119900
rect 41380 119880 41620 119900
rect 41880 119880 42120 119900
rect 42380 119880 42620 119900
rect 42880 119880 43120 119900
rect 43380 119880 43620 119900
rect 43880 119880 44120 119900
rect 44380 119880 44620 119900
rect 44880 119880 45120 119900
rect 45380 119880 45620 119900
rect 45880 119880 46120 119900
rect 46380 119880 46620 119900
rect 46880 119880 47120 119900
rect 47380 119880 47620 119900
rect 47880 119880 48120 119900
rect 48380 119880 48620 119900
rect 48880 119880 49120 119900
rect 49380 119880 49620 119900
rect 49880 119880 50120 119900
rect 50380 119880 50620 119900
rect 50880 119880 51120 119900
rect 51380 119880 51620 119900
rect 51880 119880 52120 119900
rect 52380 119880 52620 119900
rect 52880 119880 53120 119900
rect 53380 119880 53620 119900
rect 53880 119880 54120 119900
rect 54380 119880 54620 119900
rect 54880 119880 55120 119900
rect 55380 119880 55620 119900
rect 55880 119880 56120 119900
rect 56380 119880 56620 119900
rect 56880 119880 57120 119900
rect 57380 119880 57620 119900
rect 57880 119880 58000 119900
rect 14000 119620 14100 119880
rect 14400 119620 14600 119880
rect 14900 119620 15100 119880
rect 15400 119620 15600 119880
rect 15900 119620 16100 119880
rect 16400 119620 16600 119880
rect 16900 119620 17100 119880
rect 17400 119620 17600 119880
rect 17900 119620 18100 119880
rect 18400 119620 18600 119880
rect 18900 119620 19100 119880
rect 19400 119620 19600 119880
rect 19900 119620 20100 119880
rect 20400 119620 20600 119880
rect 20900 119620 21100 119880
rect 21400 119620 21600 119880
rect 21900 119620 22100 119880
rect 22400 119620 22600 119880
rect 22900 119620 23100 119880
rect 23400 119620 23600 119880
rect 23900 119620 24100 119880
rect 24400 119620 24600 119880
rect 24900 119620 25100 119880
rect 25400 119620 25600 119880
rect 25900 119620 26100 119880
rect 26400 119620 26600 119880
rect 26900 119620 27100 119880
rect 27400 119620 27600 119880
rect 27900 119620 28100 119880
rect 28400 119620 28600 119880
rect 28900 119620 29100 119880
rect 29400 119620 29600 119880
rect 29900 119620 30100 119880
rect 30400 119620 30600 119880
rect 30900 119620 31100 119880
rect 31400 119620 31600 119880
rect 31900 119620 32100 119880
rect 32400 119620 32600 119880
rect 32900 119620 33100 119880
rect 33400 119620 33600 119880
rect 33900 119620 34100 119880
rect 34400 119620 34600 119880
rect 34900 119620 35100 119880
rect 35400 119620 35600 119880
rect 35900 119620 36100 119880
rect 36400 119620 36600 119880
rect 36900 119620 37100 119880
rect 37400 119620 37600 119880
rect 37900 119620 38100 119880
rect 38400 119620 38600 119880
rect 38900 119620 39100 119880
rect 39400 119620 39600 119880
rect 39900 119620 40100 119880
rect 40400 119620 40600 119880
rect 40900 119620 41100 119880
rect 41400 119620 41600 119880
rect 41900 119620 42100 119880
rect 42400 119620 42600 119880
rect 42900 119620 43100 119880
rect 43400 119620 43600 119880
rect 43900 119620 44100 119880
rect 44400 119620 44600 119880
rect 44900 119620 45100 119880
rect 45400 119620 45600 119880
rect 45900 119620 46100 119880
rect 46400 119620 46600 119880
rect 46900 119620 47100 119880
rect 47400 119620 47600 119880
rect 47900 119620 48100 119880
rect 48400 119620 48600 119880
rect 48900 119620 49100 119880
rect 49400 119620 49600 119880
rect 49900 119620 50100 119880
rect 50400 119620 50600 119880
rect 50900 119620 51100 119880
rect 51400 119620 51600 119880
rect 51900 119620 52100 119880
rect 52400 119620 52600 119880
rect 52900 119620 53100 119880
rect 53400 119620 53600 119880
rect 53900 119620 54100 119880
rect 54400 119620 54600 119880
rect 54900 119620 55100 119880
rect 55400 119620 55600 119880
rect 55900 119620 56100 119880
rect 56400 119620 56600 119880
rect 56900 119620 57100 119880
rect 57400 119620 57600 119880
rect 57900 119620 58000 119880
rect 14000 119600 14120 119620
rect 14380 119600 14620 119620
rect 14880 119600 15120 119620
rect 15380 119600 15620 119620
rect 15880 119600 16120 119620
rect 16380 119600 16620 119620
rect 16880 119600 17120 119620
rect 17380 119600 17620 119620
rect 17880 119600 18120 119620
rect 18380 119600 18620 119620
rect 18880 119600 19120 119620
rect 19380 119600 19620 119620
rect 19880 119600 20120 119620
rect 20380 119600 20620 119620
rect 20880 119600 21120 119620
rect 21380 119600 21620 119620
rect 21880 119600 22120 119620
rect 22380 119600 22620 119620
rect 22880 119600 23120 119620
rect 23380 119600 23620 119620
rect 23880 119600 24120 119620
rect 24380 119600 24620 119620
rect 24880 119600 25120 119620
rect 25380 119600 25620 119620
rect 25880 119600 26120 119620
rect 26380 119600 26620 119620
rect 26880 119600 27120 119620
rect 27380 119600 27620 119620
rect 27880 119600 28120 119620
rect 28380 119600 28620 119620
rect 28880 119600 29120 119620
rect 29380 119600 29620 119620
rect 29880 119600 30120 119620
rect 30380 119600 30620 119620
rect 30880 119600 31120 119620
rect 31380 119600 31620 119620
rect 31880 119600 32120 119620
rect 32380 119600 32620 119620
rect 32880 119600 33120 119620
rect 33380 119600 33620 119620
rect 33880 119600 34120 119620
rect 34380 119600 34620 119620
rect 34880 119600 35120 119620
rect 35380 119600 35620 119620
rect 35880 119600 36120 119620
rect 36380 119600 36620 119620
rect 36880 119600 37120 119620
rect 37380 119600 37620 119620
rect 37880 119600 38120 119620
rect 38380 119600 38620 119620
rect 38880 119600 39120 119620
rect 39380 119600 39620 119620
rect 39880 119600 40120 119620
rect 40380 119600 40620 119620
rect 40880 119600 41120 119620
rect 41380 119600 41620 119620
rect 41880 119600 42120 119620
rect 42380 119600 42620 119620
rect 42880 119600 43120 119620
rect 43380 119600 43620 119620
rect 43880 119600 44120 119620
rect 44380 119600 44620 119620
rect 44880 119600 45120 119620
rect 45380 119600 45620 119620
rect 45880 119600 46120 119620
rect 46380 119600 46620 119620
rect 46880 119600 47120 119620
rect 47380 119600 47620 119620
rect 47880 119600 48120 119620
rect 48380 119600 48620 119620
rect 48880 119600 49120 119620
rect 49380 119600 49620 119620
rect 49880 119600 50120 119620
rect 50380 119600 50620 119620
rect 50880 119600 51120 119620
rect 51380 119600 51620 119620
rect 51880 119600 52120 119620
rect 52380 119600 52620 119620
rect 52880 119600 53120 119620
rect 53380 119600 53620 119620
rect 53880 119600 54120 119620
rect 54380 119600 54620 119620
rect 54880 119600 55120 119620
rect 55380 119600 55620 119620
rect 55880 119600 56120 119620
rect 56380 119600 56620 119620
rect 56880 119600 57120 119620
rect 57380 119600 57620 119620
rect 57880 119600 58000 119620
rect 14000 119400 58000 119600
rect 14000 119380 14120 119400
rect 14380 119380 14620 119400
rect 14880 119380 15120 119400
rect 15380 119380 15620 119400
rect 15880 119380 16120 119400
rect 16380 119380 16620 119400
rect 16880 119380 17120 119400
rect 17380 119380 17620 119400
rect 17880 119380 18120 119400
rect 18380 119380 18620 119400
rect 18880 119380 19120 119400
rect 19380 119380 19620 119400
rect 19880 119380 20120 119400
rect 20380 119380 20620 119400
rect 20880 119380 21120 119400
rect 21380 119380 21620 119400
rect 21880 119380 22120 119400
rect 22380 119380 22620 119400
rect 22880 119380 23120 119400
rect 23380 119380 23620 119400
rect 23880 119380 24120 119400
rect 24380 119380 24620 119400
rect 24880 119380 25120 119400
rect 25380 119380 25620 119400
rect 25880 119380 26120 119400
rect 26380 119380 26620 119400
rect 26880 119380 27120 119400
rect 27380 119380 27620 119400
rect 27880 119380 28120 119400
rect 28380 119380 28620 119400
rect 28880 119380 29120 119400
rect 29380 119380 29620 119400
rect 29880 119380 30120 119400
rect 30380 119380 30620 119400
rect 30880 119380 31120 119400
rect 31380 119380 31620 119400
rect 31880 119380 32120 119400
rect 32380 119380 32620 119400
rect 32880 119380 33120 119400
rect 33380 119380 33620 119400
rect 33880 119380 34120 119400
rect 34380 119380 34620 119400
rect 34880 119380 35120 119400
rect 35380 119380 35620 119400
rect 35880 119380 36120 119400
rect 36380 119380 36620 119400
rect 36880 119380 37120 119400
rect 37380 119380 37620 119400
rect 37880 119380 38120 119400
rect 38380 119380 38620 119400
rect 38880 119380 39120 119400
rect 39380 119380 39620 119400
rect 39880 119380 40120 119400
rect 40380 119380 40620 119400
rect 40880 119380 41120 119400
rect 41380 119380 41620 119400
rect 41880 119380 42120 119400
rect 42380 119380 42620 119400
rect 42880 119380 43120 119400
rect 43380 119380 43620 119400
rect 43880 119380 44120 119400
rect 44380 119380 44620 119400
rect 44880 119380 45120 119400
rect 45380 119380 45620 119400
rect 45880 119380 46120 119400
rect 46380 119380 46620 119400
rect 46880 119380 47120 119400
rect 47380 119380 47620 119400
rect 47880 119380 48120 119400
rect 48380 119380 48620 119400
rect 48880 119380 49120 119400
rect 49380 119380 49620 119400
rect 49880 119380 50120 119400
rect 50380 119380 50620 119400
rect 50880 119380 51120 119400
rect 51380 119380 51620 119400
rect 51880 119380 52120 119400
rect 52380 119380 52620 119400
rect 52880 119380 53120 119400
rect 53380 119380 53620 119400
rect 53880 119380 54120 119400
rect 54380 119380 54620 119400
rect 54880 119380 55120 119400
rect 55380 119380 55620 119400
rect 55880 119380 56120 119400
rect 56380 119380 56620 119400
rect 56880 119380 57120 119400
rect 57380 119380 57620 119400
rect 57880 119380 58000 119400
rect 14000 119120 14100 119380
rect 14400 119120 14600 119380
rect 14900 119120 15100 119380
rect 15400 119120 15600 119380
rect 15900 119120 16100 119380
rect 16400 119120 16600 119380
rect 16900 119120 17100 119380
rect 17400 119120 17600 119380
rect 17900 119120 18100 119380
rect 18400 119120 18600 119380
rect 18900 119120 19100 119380
rect 19400 119120 19600 119380
rect 19900 119120 20100 119380
rect 20400 119120 20600 119380
rect 20900 119120 21100 119380
rect 21400 119120 21600 119380
rect 21900 119120 22100 119380
rect 22400 119120 22600 119380
rect 22900 119120 23100 119380
rect 23400 119120 23600 119380
rect 23900 119120 24100 119380
rect 24400 119120 24600 119380
rect 24900 119120 25100 119380
rect 25400 119120 25600 119380
rect 25900 119120 26100 119380
rect 26400 119120 26600 119380
rect 26900 119120 27100 119380
rect 27400 119120 27600 119380
rect 27900 119120 28100 119380
rect 28400 119120 28600 119380
rect 28900 119120 29100 119380
rect 29400 119120 29600 119380
rect 29900 119120 30100 119380
rect 30400 119120 30600 119380
rect 30900 119120 31100 119380
rect 31400 119120 31600 119380
rect 31900 119120 32100 119380
rect 32400 119120 32600 119380
rect 32900 119120 33100 119380
rect 33400 119120 33600 119380
rect 33900 119120 34100 119380
rect 34400 119120 34600 119380
rect 34900 119120 35100 119380
rect 35400 119120 35600 119380
rect 35900 119120 36100 119380
rect 36400 119120 36600 119380
rect 36900 119120 37100 119380
rect 37400 119120 37600 119380
rect 37900 119120 38100 119380
rect 38400 119120 38600 119380
rect 38900 119120 39100 119380
rect 39400 119120 39600 119380
rect 39900 119120 40100 119380
rect 40400 119120 40600 119380
rect 40900 119120 41100 119380
rect 41400 119120 41600 119380
rect 41900 119120 42100 119380
rect 42400 119120 42600 119380
rect 42900 119120 43100 119380
rect 43400 119120 43600 119380
rect 43900 119120 44100 119380
rect 44400 119120 44600 119380
rect 44900 119120 45100 119380
rect 45400 119120 45600 119380
rect 45900 119120 46100 119380
rect 46400 119120 46600 119380
rect 46900 119120 47100 119380
rect 47400 119120 47600 119380
rect 47900 119120 48100 119380
rect 48400 119120 48600 119380
rect 48900 119120 49100 119380
rect 49400 119120 49600 119380
rect 49900 119120 50100 119380
rect 50400 119120 50600 119380
rect 50900 119120 51100 119380
rect 51400 119120 51600 119380
rect 51900 119120 52100 119380
rect 52400 119120 52600 119380
rect 52900 119120 53100 119380
rect 53400 119120 53600 119380
rect 53900 119120 54100 119380
rect 54400 119120 54600 119380
rect 54900 119120 55100 119380
rect 55400 119120 55600 119380
rect 55900 119120 56100 119380
rect 56400 119120 56600 119380
rect 56900 119120 57100 119380
rect 57400 119120 57600 119380
rect 57900 119120 58000 119380
rect 14000 119100 14120 119120
rect 14380 119100 14620 119120
rect 14880 119100 15120 119120
rect 15380 119100 15620 119120
rect 15880 119100 16120 119120
rect 16380 119100 16620 119120
rect 16880 119100 17120 119120
rect 17380 119100 17620 119120
rect 17880 119100 18120 119120
rect 18380 119100 18620 119120
rect 18880 119100 19120 119120
rect 19380 119100 19620 119120
rect 19880 119100 20120 119120
rect 20380 119100 20620 119120
rect 20880 119100 21120 119120
rect 21380 119100 21620 119120
rect 21880 119100 22120 119120
rect 22380 119100 22620 119120
rect 22880 119100 23120 119120
rect 23380 119100 23620 119120
rect 23880 119100 24120 119120
rect 24380 119100 24620 119120
rect 24880 119100 25120 119120
rect 25380 119100 25620 119120
rect 25880 119100 26120 119120
rect 26380 119100 26620 119120
rect 26880 119100 27120 119120
rect 27380 119100 27620 119120
rect 27880 119100 28120 119120
rect 28380 119100 28620 119120
rect 28880 119100 29120 119120
rect 29380 119100 29620 119120
rect 29880 119100 30120 119120
rect 30380 119100 30620 119120
rect 30880 119100 31120 119120
rect 31380 119100 31620 119120
rect 31880 119100 32120 119120
rect 32380 119100 32620 119120
rect 32880 119100 33120 119120
rect 33380 119100 33620 119120
rect 33880 119100 34120 119120
rect 34380 119100 34620 119120
rect 34880 119100 35120 119120
rect 35380 119100 35620 119120
rect 35880 119100 36120 119120
rect 36380 119100 36620 119120
rect 36880 119100 37120 119120
rect 37380 119100 37620 119120
rect 37880 119100 38120 119120
rect 38380 119100 38620 119120
rect 38880 119100 39120 119120
rect 39380 119100 39620 119120
rect 39880 119100 40120 119120
rect 40380 119100 40620 119120
rect 40880 119100 41120 119120
rect 41380 119100 41620 119120
rect 41880 119100 42120 119120
rect 42380 119100 42620 119120
rect 42880 119100 43120 119120
rect 43380 119100 43620 119120
rect 43880 119100 44120 119120
rect 44380 119100 44620 119120
rect 44880 119100 45120 119120
rect 45380 119100 45620 119120
rect 45880 119100 46120 119120
rect 46380 119100 46620 119120
rect 46880 119100 47120 119120
rect 47380 119100 47620 119120
rect 47880 119100 48120 119120
rect 48380 119100 48620 119120
rect 48880 119100 49120 119120
rect 49380 119100 49620 119120
rect 49880 119100 50120 119120
rect 50380 119100 50620 119120
rect 50880 119100 51120 119120
rect 51380 119100 51620 119120
rect 51880 119100 52120 119120
rect 52380 119100 52620 119120
rect 52880 119100 53120 119120
rect 53380 119100 53620 119120
rect 53880 119100 54120 119120
rect 54380 119100 54620 119120
rect 54880 119100 55120 119120
rect 55380 119100 55620 119120
rect 55880 119100 56120 119120
rect 56380 119100 56620 119120
rect 56880 119100 57120 119120
rect 57380 119100 57620 119120
rect 57880 119100 58000 119120
rect 14000 118900 58000 119100
rect 14000 118880 14120 118900
rect 14380 118880 14620 118900
rect 14880 118880 15120 118900
rect 15380 118880 15620 118900
rect 15880 118880 16120 118900
rect 16380 118880 16620 118900
rect 16880 118880 17120 118900
rect 17380 118880 17620 118900
rect 17880 118880 18120 118900
rect 18380 118880 18620 118900
rect 18880 118880 19120 118900
rect 19380 118880 19620 118900
rect 19880 118880 20120 118900
rect 20380 118880 20620 118900
rect 20880 118880 21120 118900
rect 21380 118880 21620 118900
rect 21880 118880 22120 118900
rect 22380 118880 22620 118900
rect 22880 118880 23120 118900
rect 23380 118880 23620 118900
rect 23880 118880 24120 118900
rect 24380 118880 24620 118900
rect 24880 118880 25120 118900
rect 25380 118880 25620 118900
rect 25880 118880 26120 118900
rect 26380 118880 26620 118900
rect 26880 118880 27120 118900
rect 27380 118880 27620 118900
rect 27880 118880 28120 118900
rect 28380 118880 28620 118900
rect 28880 118880 29120 118900
rect 29380 118880 29620 118900
rect 29880 118880 30120 118900
rect 30380 118880 30620 118900
rect 30880 118880 31120 118900
rect 31380 118880 31620 118900
rect 31880 118880 32120 118900
rect 32380 118880 32620 118900
rect 32880 118880 33120 118900
rect 33380 118880 33620 118900
rect 33880 118880 34120 118900
rect 34380 118880 34620 118900
rect 34880 118880 35120 118900
rect 35380 118880 35620 118900
rect 35880 118880 36120 118900
rect 36380 118880 36620 118900
rect 36880 118880 37120 118900
rect 37380 118880 37620 118900
rect 37880 118880 38120 118900
rect 38380 118880 38620 118900
rect 38880 118880 39120 118900
rect 39380 118880 39620 118900
rect 39880 118880 40120 118900
rect 40380 118880 40620 118900
rect 40880 118880 41120 118900
rect 41380 118880 41620 118900
rect 41880 118880 42120 118900
rect 42380 118880 42620 118900
rect 42880 118880 43120 118900
rect 43380 118880 43620 118900
rect 43880 118880 44120 118900
rect 44380 118880 44620 118900
rect 44880 118880 45120 118900
rect 45380 118880 45620 118900
rect 45880 118880 46120 118900
rect 46380 118880 46620 118900
rect 46880 118880 47120 118900
rect 47380 118880 47620 118900
rect 47880 118880 48120 118900
rect 48380 118880 48620 118900
rect 48880 118880 49120 118900
rect 49380 118880 49620 118900
rect 49880 118880 50120 118900
rect 50380 118880 50620 118900
rect 50880 118880 51120 118900
rect 51380 118880 51620 118900
rect 51880 118880 52120 118900
rect 52380 118880 52620 118900
rect 52880 118880 53120 118900
rect 53380 118880 53620 118900
rect 53880 118880 54120 118900
rect 54380 118880 54620 118900
rect 54880 118880 55120 118900
rect 55380 118880 55620 118900
rect 55880 118880 56120 118900
rect 56380 118880 56620 118900
rect 56880 118880 57120 118900
rect 57380 118880 57620 118900
rect 57880 118880 58000 118900
rect 14000 118620 14100 118880
rect 14400 118620 14600 118880
rect 14900 118620 15100 118880
rect 15400 118620 15600 118880
rect 15900 118620 16100 118880
rect 16400 118620 16600 118880
rect 16900 118620 17100 118880
rect 17400 118620 17600 118880
rect 17900 118620 18100 118880
rect 18400 118620 18600 118880
rect 18900 118620 19100 118880
rect 19400 118620 19600 118880
rect 19900 118620 20100 118880
rect 20400 118620 20600 118880
rect 20900 118620 21100 118880
rect 21400 118620 21600 118880
rect 21900 118620 22100 118880
rect 22400 118620 22600 118880
rect 22900 118620 23100 118880
rect 23400 118620 23600 118880
rect 23900 118620 24100 118880
rect 24400 118620 24600 118880
rect 24900 118620 25100 118880
rect 25400 118620 25600 118880
rect 25900 118620 26100 118880
rect 26400 118620 26600 118880
rect 26900 118620 27100 118880
rect 27400 118620 27600 118880
rect 27900 118620 28100 118880
rect 28400 118620 28600 118880
rect 28900 118620 29100 118880
rect 29400 118620 29600 118880
rect 29900 118620 30100 118880
rect 30400 118620 30600 118880
rect 30900 118620 31100 118880
rect 31400 118620 31600 118880
rect 31900 118620 32100 118880
rect 32400 118620 32600 118880
rect 32900 118620 33100 118880
rect 33400 118620 33600 118880
rect 33900 118620 34100 118880
rect 34400 118620 34600 118880
rect 34900 118620 35100 118880
rect 35400 118620 35600 118880
rect 35900 118620 36100 118880
rect 36400 118620 36600 118880
rect 36900 118620 37100 118880
rect 37400 118620 37600 118880
rect 37900 118620 38100 118880
rect 38400 118620 38600 118880
rect 38900 118620 39100 118880
rect 39400 118620 39600 118880
rect 39900 118620 40100 118880
rect 40400 118620 40600 118880
rect 40900 118620 41100 118880
rect 41400 118620 41600 118880
rect 41900 118620 42100 118880
rect 42400 118620 42600 118880
rect 42900 118620 43100 118880
rect 43400 118620 43600 118880
rect 43900 118620 44100 118880
rect 44400 118620 44600 118880
rect 44900 118620 45100 118880
rect 45400 118620 45600 118880
rect 45900 118620 46100 118880
rect 46400 118620 46600 118880
rect 46900 118620 47100 118880
rect 47400 118620 47600 118880
rect 47900 118620 48100 118880
rect 48400 118620 48600 118880
rect 48900 118620 49100 118880
rect 49400 118620 49600 118880
rect 49900 118620 50100 118880
rect 50400 118620 50600 118880
rect 50900 118620 51100 118880
rect 51400 118620 51600 118880
rect 51900 118620 52100 118880
rect 52400 118620 52600 118880
rect 52900 118620 53100 118880
rect 53400 118620 53600 118880
rect 53900 118620 54100 118880
rect 54400 118620 54600 118880
rect 54900 118620 55100 118880
rect 55400 118620 55600 118880
rect 55900 118620 56100 118880
rect 56400 118620 56600 118880
rect 56900 118620 57100 118880
rect 57400 118620 57600 118880
rect 57900 118620 58000 118880
rect 14000 118600 14120 118620
rect 14380 118600 14620 118620
rect 14880 118600 15120 118620
rect 15380 118600 15620 118620
rect 15880 118600 16120 118620
rect 16380 118600 16620 118620
rect 16880 118600 17120 118620
rect 17380 118600 17620 118620
rect 17880 118600 18120 118620
rect 18380 118600 18620 118620
rect 18880 118600 19120 118620
rect 19380 118600 19620 118620
rect 19880 118600 20120 118620
rect 20380 118600 20620 118620
rect 20880 118600 21120 118620
rect 21380 118600 21620 118620
rect 21880 118600 22120 118620
rect 22380 118600 22620 118620
rect 22880 118600 23120 118620
rect 23380 118600 23620 118620
rect 23880 118600 24120 118620
rect 24380 118600 24620 118620
rect 24880 118600 25120 118620
rect 25380 118600 25620 118620
rect 25880 118600 26120 118620
rect 26380 118600 26620 118620
rect 26880 118600 27120 118620
rect 27380 118600 27620 118620
rect 27880 118600 28120 118620
rect 28380 118600 28620 118620
rect 28880 118600 29120 118620
rect 29380 118600 29620 118620
rect 29880 118600 30120 118620
rect 30380 118600 30620 118620
rect 30880 118600 31120 118620
rect 31380 118600 31620 118620
rect 31880 118600 32120 118620
rect 32380 118600 32620 118620
rect 32880 118600 33120 118620
rect 33380 118600 33620 118620
rect 33880 118600 34120 118620
rect 34380 118600 34620 118620
rect 34880 118600 35120 118620
rect 35380 118600 35620 118620
rect 35880 118600 36120 118620
rect 36380 118600 36620 118620
rect 36880 118600 37120 118620
rect 37380 118600 37620 118620
rect 37880 118600 38120 118620
rect 38380 118600 38620 118620
rect 38880 118600 39120 118620
rect 39380 118600 39620 118620
rect 39880 118600 40120 118620
rect 40380 118600 40620 118620
rect 40880 118600 41120 118620
rect 41380 118600 41620 118620
rect 41880 118600 42120 118620
rect 42380 118600 42620 118620
rect 42880 118600 43120 118620
rect 43380 118600 43620 118620
rect 43880 118600 44120 118620
rect 44380 118600 44620 118620
rect 44880 118600 45120 118620
rect 45380 118600 45620 118620
rect 45880 118600 46120 118620
rect 46380 118600 46620 118620
rect 46880 118600 47120 118620
rect 47380 118600 47620 118620
rect 47880 118600 48120 118620
rect 48380 118600 48620 118620
rect 48880 118600 49120 118620
rect 49380 118600 49620 118620
rect 49880 118600 50120 118620
rect 50380 118600 50620 118620
rect 50880 118600 51120 118620
rect 51380 118600 51620 118620
rect 51880 118600 52120 118620
rect 52380 118600 52620 118620
rect 52880 118600 53120 118620
rect 53380 118600 53620 118620
rect 53880 118600 54120 118620
rect 54380 118600 54620 118620
rect 54880 118600 55120 118620
rect 55380 118600 55620 118620
rect 55880 118600 56120 118620
rect 56380 118600 56620 118620
rect 56880 118600 57120 118620
rect 57380 118600 57620 118620
rect 57880 118600 58000 118620
rect 14000 118400 58000 118600
rect 14000 118380 14120 118400
rect 14380 118380 14620 118400
rect 14880 118380 15120 118400
rect 15380 118380 15620 118400
rect 15880 118380 16120 118400
rect 16380 118380 16620 118400
rect 16880 118380 17120 118400
rect 17380 118380 17620 118400
rect 17880 118380 18120 118400
rect 18380 118380 18620 118400
rect 18880 118380 19120 118400
rect 19380 118380 19620 118400
rect 19880 118380 20120 118400
rect 20380 118380 20620 118400
rect 20880 118380 21120 118400
rect 21380 118380 21620 118400
rect 21880 118380 22120 118400
rect 22380 118380 22620 118400
rect 22880 118380 23120 118400
rect 23380 118380 23620 118400
rect 23880 118380 24120 118400
rect 24380 118380 24620 118400
rect 24880 118380 25120 118400
rect 25380 118380 25620 118400
rect 25880 118380 26120 118400
rect 26380 118380 26620 118400
rect 26880 118380 27120 118400
rect 27380 118380 27620 118400
rect 27880 118380 28120 118400
rect 28380 118380 28620 118400
rect 28880 118380 29120 118400
rect 29380 118380 29620 118400
rect 29880 118380 30120 118400
rect 30380 118380 30620 118400
rect 30880 118380 31120 118400
rect 31380 118380 31620 118400
rect 31880 118380 32120 118400
rect 32380 118380 32620 118400
rect 32880 118380 33120 118400
rect 33380 118380 33620 118400
rect 33880 118380 34120 118400
rect 34380 118380 34620 118400
rect 34880 118380 35120 118400
rect 35380 118380 35620 118400
rect 35880 118380 36120 118400
rect 36380 118380 36620 118400
rect 36880 118380 37120 118400
rect 37380 118380 37620 118400
rect 37880 118380 38120 118400
rect 38380 118380 38620 118400
rect 38880 118380 39120 118400
rect 39380 118380 39620 118400
rect 39880 118380 40120 118400
rect 40380 118380 40620 118400
rect 40880 118380 41120 118400
rect 41380 118380 41620 118400
rect 41880 118380 42120 118400
rect 42380 118380 42620 118400
rect 42880 118380 43120 118400
rect 43380 118380 43620 118400
rect 43880 118380 44120 118400
rect 44380 118380 44620 118400
rect 44880 118380 45120 118400
rect 45380 118380 45620 118400
rect 45880 118380 46120 118400
rect 46380 118380 46620 118400
rect 46880 118380 47120 118400
rect 47380 118380 47620 118400
rect 47880 118380 48120 118400
rect 48380 118380 48620 118400
rect 48880 118380 49120 118400
rect 49380 118380 49620 118400
rect 49880 118380 50120 118400
rect 50380 118380 50620 118400
rect 50880 118380 51120 118400
rect 51380 118380 51620 118400
rect 51880 118380 52120 118400
rect 52380 118380 52620 118400
rect 52880 118380 53120 118400
rect 53380 118380 53620 118400
rect 53880 118380 54120 118400
rect 54380 118380 54620 118400
rect 54880 118380 55120 118400
rect 55380 118380 55620 118400
rect 55880 118380 56120 118400
rect 56380 118380 56620 118400
rect 56880 118380 57120 118400
rect 57380 118380 57620 118400
rect 57880 118380 58000 118400
rect 14000 118120 14100 118380
rect 14400 118120 14600 118380
rect 14900 118120 15100 118380
rect 15400 118120 15600 118380
rect 15900 118120 16100 118380
rect 16400 118120 16600 118380
rect 16900 118120 17100 118380
rect 17400 118120 17600 118380
rect 17900 118120 18100 118380
rect 18400 118120 18600 118380
rect 18900 118120 19100 118380
rect 19400 118120 19600 118380
rect 19900 118120 20100 118380
rect 20400 118120 20600 118380
rect 20900 118120 21100 118380
rect 21400 118120 21600 118380
rect 21900 118120 22100 118380
rect 22400 118120 22600 118380
rect 22900 118120 23100 118380
rect 23400 118120 23600 118380
rect 23900 118120 24100 118380
rect 24400 118120 24600 118380
rect 24900 118120 25100 118380
rect 25400 118120 25600 118380
rect 25900 118120 26100 118380
rect 26400 118120 26600 118380
rect 26900 118120 27100 118380
rect 27400 118120 27600 118380
rect 27900 118120 28100 118380
rect 28400 118120 28600 118380
rect 28900 118120 29100 118380
rect 29400 118120 29600 118380
rect 29900 118120 30100 118380
rect 30400 118120 30600 118380
rect 30900 118120 31100 118380
rect 31400 118120 31600 118380
rect 31900 118120 32100 118380
rect 32400 118120 32600 118380
rect 32900 118120 33100 118380
rect 33400 118120 33600 118380
rect 33900 118120 34100 118380
rect 34400 118120 34600 118380
rect 34900 118120 35100 118380
rect 35400 118120 35600 118380
rect 35900 118120 36100 118380
rect 36400 118120 36600 118380
rect 36900 118120 37100 118380
rect 37400 118120 37600 118380
rect 37900 118120 38100 118380
rect 38400 118120 38600 118380
rect 38900 118120 39100 118380
rect 39400 118120 39600 118380
rect 39900 118120 40100 118380
rect 40400 118120 40600 118380
rect 40900 118120 41100 118380
rect 41400 118120 41600 118380
rect 41900 118120 42100 118380
rect 42400 118120 42600 118380
rect 42900 118120 43100 118380
rect 43400 118120 43600 118380
rect 43900 118120 44100 118380
rect 44400 118120 44600 118380
rect 44900 118120 45100 118380
rect 45400 118120 45600 118380
rect 45900 118120 46100 118380
rect 46400 118120 46600 118380
rect 46900 118120 47100 118380
rect 47400 118120 47600 118380
rect 47900 118120 48100 118380
rect 48400 118120 48600 118380
rect 48900 118120 49100 118380
rect 49400 118120 49600 118380
rect 49900 118120 50100 118380
rect 50400 118120 50600 118380
rect 50900 118120 51100 118380
rect 51400 118120 51600 118380
rect 51900 118120 52100 118380
rect 52400 118120 52600 118380
rect 52900 118120 53100 118380
rect 53400 118120 53600 118380
rect 53900 118120 54100 118380
rect 54400 118120 54600 118380
rect 54900 118120 55100 118380
rect 55400 118120 55600 118380
rect 55900 118120 56100 118380
rect 56400 118120 56600 118380
rect 56900 118120 57100 118380
rect 57400 118120 57600 118380
rect 57900 118120 58000 118380
rect 14000 118100 14120 118120
rect 14380 118100 14620 118120
rect 14880 118100 15120 118120
rect 15380 118100 15620 118120
rect 15880 118100 16120 118120
rect 16380 118100 16620 118120
rect 16880 118100 17120 118120
rect 17380 118100 17620 118120
rect 17880 118100 18120 118120
rect 18380 118100 18620 118120
rect 18880 118100 19120 118120
rect 19380 118100 19620 118120
rect 19880 118100 20120 118120
rect 20380 118100 20620 118120
rect 20880 118100 21120 118120
rect 21380 118100 21620 118120
rect 21880 118100 22120 118120
rect 22380 118100 22620 118120
rect 22880 118100 23120 118120
rect 23380 118100 23620 118120
rect 23880 118100 24120 118120
rect 24380 118100 24620 118120
rect 24880 118100 25120 118120
rect 25380 118100 25620 118120
rect 25880 118100 26120 118120
rect 26380 118100 26620 118120
rect 26880 118100 27120 118120
rect 27380 118100 27620 118120
rect 27880 118100 28120 118120
rect 28380 118100 28620 118120
rect 28880 118100 29120 118120
rect 29380 118100 29620 118120
rect 29880 118100 30120 118120
rect 30380 118100 30620 118120
rect 30880 118100 31120 118120
rect 31380 118100 31620 118120
rect 31880 118100 32120 118120
rect 32380 118100 32620 118120
rect 32880 118100 33120 118120
rect 33380 118100 33620 118120
rect 33880 118100 34120 118120
rect 34380 118100 34620 118120
rect 34880 118100 35120 118120
rect 35380 118100 35620 118120
rect 35880 118100 36120 118120
rect 36380 118100 36620 118120
rect 36880 118100 37120 118120
rect 37380 118100 37620 118120
rect 37880 118100 38120 118120
rect 38380 118100 38620 118120
rect 38880 118100 39120 118120
rect 39380 118100 39620 118120
rect 39880 118100 40120 118120
rect 40380 118100 40620 118120
rect 40880 118100 41120 118120
rect 41380 118100 41620 118120
rect 41880 118100 42120 118120
rect 42380 118100 42620 118120
rect 42880 118100 43120 118120
rect 43380 118100 43620 118120
rect 43880 118100 44120 118120
rect 44380 118100 44620 118120
rect 44880 118100 45120 118120
rect 45380 118100 45620 118120
rect 45880 118100 46120 118120
rect 46380 118100 46620 118120
rect 46880 118100 47120 118120
rect 47380 118100 47620 118120
rect 47880 118100 48120 118120
rect 48380 118100 48620 118120
rect 48880 118100 49120 118120
rect 49380 118100 49620 118120
rect 49880 118100 50120 118120
rect 50380 118100 50620 118120
rect 50880 118100 51120 118120
rect 51380 118100 51620 118120
rect 51880 118100 52120 118120
rect 52380 118100 52620 118120
rect 52880 118100 53120 118120
rect 53380 118100 53620 118120
rect 53880 118100 54120 118120
rect 54380 118100 54620 118120
rect 54880 118100 55120 118120
rect 55380 118100 55620 118120
rect 55880 118100 56120 118120
rect 56380 118100 56620 118120
rect 56880 118100 57120 118120
rect 57380 118100 57620 118120
rect 57880 118100 58000 118120
rect 14000 117900 58000 118100
rect 14000 117880 14120 117900
rect 14380 117880 14620 117900
rect 14880 117880 15120 117900
rect 15380 117880 15620 117900
rect 15880 117880 16120 117900
rect 16380 117880 16620 117900
rect 16880 117880 17120 117900
rect 17380 117880 17620 117900
rect 17880 117880 18120 117900
rect 18380 117880 18620 117900
rect 18880 117880 19120 117900
rect 19380 117880 19620 117900
rect 19880 117880 20120 117900
rect 20380 117880 20620 117900
rect 20880 117880 21120 117900
rect 21380 117880 21620 117900
rect 21880 117880 22120 117900
rect 22380 117880 22620 117900
rect 22880 117880 23120 117900
rect 23380 117880 23620 117900
rect 23880 117880 24120 117900
rect 24380 117880 24620 117900
rect 24880 117880 25120 117900
rect 25380 117880 25620 117900
rect 25880 117880 26120 117900
rect 26380 117880 26620 117900
rect 26880 117880 27120 117900
rect 27380 117880 27620 117900
rect 27880 117880 28120 117900
rect 28380 117880 28620 117900
rect 28880 117880 29120 117900
rect 29380 117880 29620 117900
rect 29880 117880 30120 117900
rect 30380 117880 30620 117900
rect 30880 117880 31120 117900
rect 31380 117880 31620 117900
rect 31880 117880 32120 117900
rect 32380 117880 32620 117900
rect 32880 117880 33120 117900
rect 33380 117880 33620 117900
rect 33880 117880 34120 117900
rect 34380 117880 34620 117900
rect 34880 117880 35120 117900
rect 35380 117880 35620 117900
rect 35880 117880 36120 117900
rect 36380 117880 36620 117900
rect 36880 117880 37120 117900
rect 37380 117880 37620 117900
rect 37880 117880 38120 117900
rect 38380 117880 38620 117900
rect 38880 117880 39120 117900
rect 39380 117880 39620 117900
rect 39880 117880 40120 117900
rect 40380 117880 40620 117900
rect 40880 117880 41120 117900
rect 41380 117880 41620 117900
rect 41880 117880 42120 117900
rect 42380 117880 42620 117900
rect 42880 117880 43120 117900
rect 43380 117880 43620 117900
rect 43880 117880 44120 117900
rect 44380 117880 44620 117900
rect 44880 117880 45120 117900
rect 45380 117880 45620 117900
rect 45880 117880 46120 117900
rect 46380 117880 46620 117900
rect 46880 117880 47120 117900
rect 47380 117880 47620 117900
rect 47880 117880 48120 117900
rect 48380 117880 48620 117900
rect 48880 117880 49120 117900
rect 49380 117880 49620 117900
rect 49880 117880 50120 117900
rect 50380 117880 50620 117900
rect 50880 117880 51120 117900
rect 51380 117880 51620 117900
rect 51880 117880 52120 117900
rect 52380 117880 52620 117900
rect 52880 117880 53120 117900
rect 53380 117880 53620 117900
rect 53880 117880 54120 117900
rect 54380 117880 54620 117900
rect 54880 117880 55120 117900
rect 55380 117880 55620 117900
rect 55880 117880 56120 117900
rect 56380 117880 56620 117900
rect 56880 117880 57120 117900
rect 57380 117880 57620 117900
rect 57880 117880 58000 117900
rect 14000 117620 14100 117880
rect 14400 117620 14600 117880
rect 14900 117620 15100 117880
rect 15400 117620 15600 117880
rect 15900 117620 16100 117880
rect 16400 117620 16600 117880
rect 16900 117620 17100 117880
rect 17400 117620 17600 117880
rect 17900 117620 18100 117880
rect 18400 117620 18600 117880
rect 18900 117620 19100 117880
rect 19400 117620 19600 117880
rect 19900 117620 20100 117880
rect 20400 117620 20600 117880
rect 20900 117620 21100 117880
rect 21400 117620 21600 117880
rect 21900 117620 22100 117880
rect 22400 117620 22600 117880
rect 22900 117620 23100 117880
rect 23400 117620 23600 117880
rect 23900 117620 24100 117880
rect 24400 117620 24600 117880
rect 24900 117620 25100 117880
rect 25400 117620 25600 117880
rect 25900 117620 26100 117880
rect 26400 117620 26600 117880
rect 26900 117620 27100 117880
rect 27400 117620 27600 117880
rect 27900 117620 28100 117880
rect 28400 117620 28600 117880
rect 28900 117620 29100 117880
rect 29400 117620 29600 117880
rect 29900 117620 30100 117880
rect 30400 117620 30600 117880
rect 30900 117620 31100 117880
rect 31400 117620 31600 117880
rect 31900 117620 32100 117880
rect 32400 117620 32600 117880
rect 32900 117620 33100 117880
rect 33400 117620 33600 117880
rect 33900 117620 34100 117880
rect 34400 117620 34600 117880
rect 34900 117620 35100 117880
rect 35400 117620 35600 117880
rect 35900 117620 36100 117880
rect 36400 117620 36600 117880
rect 36900 117620 37100 117880
rect 37400 117620 37600 117880
rect 37900 117620 38100 117880
rect 38400 117620 38600 117880
rect 38900 117620 39100 117880
rect 39400 117620 39600 117880
rect 39900 117620 40100 117880
rect 40400 117620 40600 117880
rect 40900 117620 41100 117880
rect 41400 117620 41600 117880
rect 41900 117620 42100 117880
rect 42400 117620 42600 117880
rect 42900 117620 43100 117880
rect 43400 117620 43600 117880
rect 43900 117620 44100 117880
rect 44400 117620 44600 117880
rect 44900 117620 45100 117880
rect 45400 117620 45600 117880
rect 45900 117620 46100 117880
rect 46400 117620 46600 117880
rect 46900 117620 47100 117880
rect 47400 117620 47600 117880
rect 47900 117620 48100 117880
rect 48400 117620 48600 117880
rect 48900 117620 49100 117880
rect 49400 117620 49600 117880
rect 49900 117620 50100 117880
rect 50400 117620 50600 117880
rect 50900 117620 51100 117880
rect 51400 117620 51600 117880
rect 51900 117620 52100 117880
rect 52400 117620 52600 117880
rect 52900 117620 53100 117880
rect 53400 117620 53600 117880
rect 53900 117620 54100 117880
rect 54400 117620 54600 117880
rect 54900 117620 55100 117880
rect 55400 117620 55600 117880
rect 55900 117620 56100 117880
rect 56400 117620 56600 117880
rect 56900 117620 57100 117880
rect 57400 117620 57600 117880
rect 57900 117620 58000 117880
rect 14000 117600 14120 117620
rect 14380 117600 14620 117620
rect 14880 117600 15120 117620
rect 15380 117600 15620 117620
rect 15880 117600 16120 117620
rect 16380 117600 16620 117620
rect 16880 117600 17120 117620
rect 17380 117600 17620 117620
rect 17880 117600 18120 117620
rect 18380 117600 18620 117620
rect 18880 117600 19120 117620
rect 19380 117600 19620 117620
rect 19880 117600 20120 117620
rect 20380 117600 20620 117620
rect 20880 117600 21120 117620
rect 21380 117600 21620 117620
rect 21880 117600 22120 117620
rect 22380 117600 22620 117620
rect 22880 117600 23120 117620
rect 23380 117600 23620 117620
rect 23880 117600 24120 117620
rect 24380 117600 24620 117620
rect 24880 117600 25120 117620
rect 25380 117600 25620 117620
rect 25880 117600 26120 117620
rect 26380 117600 26620 117620
rect 26880 117600 27120 117620
rect 27380 117600 27620 117620
rect 27880 117600 28120 117620
rect 28380 117600 28620 117620
rect 28880 117600 29120 117620
rect 29380 117600 29620 117620
rect 29880 117600 30120 117620
rect 30380 117600 30620 117620
rect 30880 117600 31120 117620
rect 31380 117600 31620 117620
rect 31880 117600 32120 117620
rect 32380 117600 32620 117620
rect 32880 117600 33120 117620
rect 33380 117600 33620 117620
rect 33880 117600 34120 117620
rect 34380 117600 34620 117620
rect 34880 117600 35120 117620
rect 35380 117600 35620 117620
rect 35880 117600 36120 117620
rect 36380 117600 36620 117620
rect 36880 117600 37120 117620
rect 37380 117600 37620 117620
rect 37880 117600 38120 117620
rect 38380 117600 38620 117620
rect 38880 117600 39120 117620
rect 39380 117600 39620 117620
rect 39880 117600 40120 117620
rect 40380 117600 40620 117620
rect 40880 117600 41120 117620
rect 41380 117600 41620 117620
rect 41880 117600 42120 117620
rect 42380 117600 42620 117620
rect 42880 117600 43120 117620
rect 43380 117600 43620 117620
rect 43880 117600 44120 117620
rect 44380 117600 44620 117620
rect 44880 117600 45120 117620
rect 45380 117600 45620 117620
rect 45880 117600 46120 117620
rect 46380 117600 46620 117620
rect 46880 117600 47120 117620
rect 47380 117600 47620 117620
rect 47880 117600 48120 117620
rect 48380 117600 48620 117620
rect 48880 117600 49120 117620
rect 49380 117600 49620 117620
rect 49880 117600 50120 117620
rect 50380 117600 50620 117620
rect 50880 117600 51120 117620
rect 51380 117600 51620 117620
rect 51880 117600 52120 117620
rect 52380 117600 52620 117620
rect 52880 117600 53120 117620
rect 53380 117600 53620 117620
rect 53880 117600 54120 117620
rect 54380 117600 54620 117620
rect 54880 117600 55120 117620
rect 55380 117600 55620 117620
rect 55880 117600 56120 117620
rect 56380 117600 56620 117620
rect 56880 117600 57120 117620
rect 57380 117600 57620 117620
rect 57880 117600 58000 117620
rect 14000 117400 58000 117600
rect 14000 117380 14120 117400
rect 14380 117380 14620 117400
rect 14880 117380 15120 117400
rect 15380 117380 15620 117400
rect 15880 117380 16120 117400
rect 16380 117380 16620 117400
rect 16880 117380 17120 117400
rect 17380 117380 17620 117400
rect 17880 117380 18120 117400
rect 18380 117380 18620 117400
rect 18880 117380 19120 117400
rect 19380 117380 19620 117400
rect 19880 117380 20120 117400
rect 20380 117380 20620 117400
rect 20880 117380 21120 117400
rect 21380 117380 21620 117400
rect 21880 117380 22120 117400
rect 22380 117380 22620 117400
rect 22880 117380 23120 117400
rect 23380 117380 23620 117400
rect 23880 117380 24120 117400
rect 24380 117380 24620 117400
rect 24880 117380 25120 117400
rect 25380 117380 25620 117400
rect 25880 117380 26120 117400
rect 26380 117380 26620 117400
rect 26880 117380 27120 117400
rect 27380 117380 27620 117400
rect 27880 117380 28120 117400
rect 28380 117380 28620 117400
rect 28880 117380 29120 117400
rect 29380 117380 29620 117400
rect 29880 117380 30120 117400
rect 30380 117380 30620 117400
rect 30880 117380 31120 117400
rect 31380 117380 31620 117400
rect 31880 117380 32120 117400
rect 32380 117380 32620 117400
rect 32880 117380 33120 117400
rect 33380 117380 33620 117400
rect 33880 117380 34120 117400
rect 34380 117380 34620 117400
rect 34880 117380 35120 117400
rect 35380 117380 35620 117400
rect 35880 117380 36120 117400
rect 36380 117380 36620 117400
rect 36880 117380 37120 117400
rect 37380 117380 37620 117400
rect 37880 117380 38120 117400
rect 38380 117380 38620 117400
rect 38880 117380 39120 117400
rect 39380 117380 39620 117400
rect 39880 117380 40120 117400
rect 40380 117380 40620 117400
rect 40880 117380 41120 117400
rect 41380 117380 41620 117400
rect 41880 117380 42120 117400
rect 42380 117380 42620 117400
rect 42880 117380 43120 117400
rect 43380 117380 43620 117400
rect 43880 117380 44120 117400
rect 44380 117380 44620 117400
rect 44880 117380 45120 117400
rect 45380 117380 45620 117400
rect 45880 117380 46120 117400
rect 46380 117380 46620 117400
rect 46880 117380 47120 117400
rect 47380 117380 47620 117400
rect 47880 117380 48120 117400
rect 48380 117380 48620 117400
rect 48880 117380 49120 117400
rect 49380 117380 49620 117400
rect 49880 117380 50120 117400
rect 50380 117380 50620 117400
rect 50880 117380 51120 117400
rect 51380 117380 51620 117400
rect 51880 117380 52120 117400
rect 52380 117380 52620 117400
rect 52880 117380 53120 117400
rect 53380 117380 53620 117400
rect 53880 117380 54120 117400
rect 54380 117380 54620 117400
rect 54880 117380 55120 117400
rect 55380 117380 55620 117400
rect 55880 117380 56120 117400
rect 56380 117380 56620 117400
rect 56880 117380 57120 117400
rect 57380 117380 57620 117400
rect 57880 117380 58000 117400
rect 14000 117120 14100 117380
rect 14400 117120 14600 117380
rect 14900 117120 15100 117380
rect 15400 117120 15600 117380
rect 15900 117120 16100 117380
rect 16400 117120 16600 117380
rect 16900 117120 17100 117380
rect 17400 117120 17600 117380
rect 17900 117120 18100 117380
rect 18400 117120 18600 117380
rect 18900 117120 19100 117380
rect 19400 117120 19600 117380
rect 19900 117120 20100 117380
rect 20400 117120 20600 117380
rect 20900 117120 21100 117380
rect 21400 117120 21600 117380
rect 21900 117120 22100 117380
rect 22400 117120 22600 117380
rect 22900 117120 23100 117380
rect 23400 117120 23600 117380
rect 23900 117120 24100 117380
rect 24400 117120 24600 117380
rect 24900 117120 25100 117380
rect 25400 117120 25600 117380
rect 25900 117120 26100 117380
rect 26400 117120 26600 117380
rect 26900 117120 27100 117380
rect 27400 117120 27600 117380
rect 27900 117120 28100 117380
rect 28400 117120 28600 117380
rect 28900 117120 29100 117380
rect 29400 117120 29600 117380
rect 29900 117120 30100 117380
rect 30400 117120 30600 117380
rect 30900 117120 31100 117380
rect 31400 117120 31600 117380
rect 31900 117120 32100 117380
rect 32400 117120 32600 117380
rect 32900 117120 33100 117380
rect 33400 117120 33600 117380
rect 33900 117120 34100 117380
rect 34400 117120 34600 117380
rect 34900 117120 35100 117380
rect 35400 117120 35600 117380
rect 35900 117120 36100 117380
rect 36400 117120 36600 117380
rect 36900 117120 37100 117380
rect 37400 117120 37600 117380
rect 37900 117120 38100 117380
rect 38400 117120 38600 117380
rect 38900 117120 39100 117380
rect 39400 117120 39600 117380
rect 39900 117120 40100 117380
rect 40400 117120 40600 117380
rect 40900 117120 41100 117380
rect 41400 117120 41600 117380
rect 41900 117120 42100 117380
rect 42400 117120 42600 117380
rect 42900 117120 43100 117380
rect 43400 117120 43600 117380
rect 43900 117120 44100 117380
rect 44400 117120 44600 117380
rect 44900 117120 45100 117380
rect 45400 117120 45600 117380
rect 45900 117120 46100 117380
rect 46400 117120 46600 117380
rect 46900 117120 47100 117380
rect 47400 117120 47600 117380
rect 47900 117120 48100 117380
rect 48400 117120 48600 117380
rect 48900 117120 49100 117380
rect 49400 117120 49600 117380
rect 49900 117120 50100 117380
rect 50400 117120 50600 117380
rect 50900 117120 51100 117380
rect 51400 117120 51600 117380
rect 51900 117120 52100 117380
rect 52400 117120 52600 117380
rect 52900 117120 53100 117380
rect 53400 117120 53600 117380
rect 53900 117120 54100 117380
rect 54400 117120 54600 117380
rect 54900 117120 55100 117380
rect 55400 117120 55600 117380
rect 55900 117120 56100 117380
rect 56400 117120 56600 117380
rect 56900 117120 57100 117380
rect 57400 117120 57600 117380
rect 57900 117120 58000 117380
rect 14000 117100 14120 117120
rect 14380 117100 14620 117120
rect 14880 117100 15120 117120
rect 15380 117100 15620 117120
rect 15880 117100 16120 117120
rect 16380 117100 16620 117120
rect 16880 117100 17120 117120
rect 17380 117100 17620 117120
rect 17880 117100 18120 117120
rect 18380 117100 18620 117120
rect 18880 117100 19120 117120
rect 19380 117100 19620 117120
rect 19880 117100 20120 117120
rect 20380 117100 20620 117120
rect 20880 117100 21120 117120
rect 21380 117100 21620 117120
rect 21880 117100 22120 117120
rect 22380 117100 22620 117120
rect 22880 117100 23120 117120
rect 23380 117100 23620 117120
rect 23880 117100 24120 117120
rect 24380 117100 24620 117120
rect 24880 117100 25120 117120
rect 25380 117100 25620 117120
rect 25880 117100 26120 117120
rect 26380 117100 26620 117120
rect 26880 117100 27120 117120
rect 27380 117100 27620 117120
rect 27880 117100 28120 117120
rect 28380 117100 28620 117120
rect 28880 117100 29120 117120
rect 29380 117100 29620 117120
rect 29880 117100 30120 117120
rect 30380 117100 30620 117120
rect 30880 117100 31120 117120
rect 31380 117100 31620 117120
rect 31880 117100 32120 117120
rect 32380 117100 32620 117120
rect 32880 117100 33120 117120
rect 33380 117100 33620 117120
rect 33880 117100 34120 117120
rect 34380 117100 34620 117120
rect 34880 117100 35120 117120
rect 35380 117100 35620 117120
rect 35880 117100 36120 117120
rect 36380 117100 36620 117120
rect 36880 117100 37120 117120
rect 37380 117100 37620 117120
rect 37880 117100 38120 117120
rect 38380 117100 38620 117120
rect 38880 117100 39120 117120
rect 39380 117100 39620 117120
rect 39880 117100 40120 117120
rect 40380 117100 40620 117120
rect 40880 117100 41120 117120
rect 41380 117100 41620 117120
rect 41880 117100 42120 117120
rect 42380 117100 42620 117120
rect 42880 117100 43120 117120
rect 43380 117100 43620 117120
rect 43880 117100 44120 117120
rect 44380 117100 44620 117120
rect 44880 117100 45120 117120
rect 45380 117100 45620 117120
rect 45880 117100 46120 117120
rect 46380 117100 46620 117120
rect 46880 117100 47120 117120
rect 47380 117100 47620 117120
rect 47880 117100 48120 117120
rect 48380 117100 48620 117120
rect 48880 117100 49120 117120
rect 49380 117100 49620 117120
rect 49880 117100 50120 117120
rect 50380 117100 50620 117120
rect 50880 117100 51120 117120
rect 51380 117100 51620 117120
rect 51880 117100 52120 117120
rect 52380 117100 52620 117120
rect 52880 117100 53120 117120
rect 53380 117100 53620 117120
rect 53880 117100 54120 117120
rect 54380 117100 54620 117120
rect 54880 117100 55120 117120
rect 55380 117100 55620 117120
rect 55880 117100 56120 117120
rect 56380 117100 56620 117120
rect 56880 117100 57120 117120
rect 57380 117100 57620 117120
rect 57880 117100 58000 117120
rect 14000 116900 58000 117100
rect 14000 116880 14120 116900
rect 14380 116880 14620 116900
rect 14880 116880 15120 116900
rect 15380 116880 15620 116900
rect 15880 116880 16120 116900
rect 16380 116880 16620 116900
rect 16880 116880 17120 116900
rect 17380 116880 17620 116900
rect 17880 116880 18120 116900
rect 18380 116880 18620 116900
rect 18880 116880 19120 116900
rect 19380 116880 19620 116900
rect 19880 116880 20120 116900
rect 20380 116880 20620 116900
rect 20880 116880 21120 116900
rect 21380 116880 21620 116900
rect 21880 116880 22120 116900
rect 22380 116880 22620 116900
rect 22880 116880 23120 116900
rect 23380 116880 23620 116900
rect 23880 116880 24120 116900
rect 24380 116880 24620 116900
rect 24880 116880 25120 116900
rect 25380 116880 25620 116900
rect 25880 116880 26120 116900
rect 26380 116880 26620 116900
rect 26880 116880 27120 116900
rect 27380 116880 27620 116900
rect 27880 116880 28120 116900
rect 28380 116880 28620 116900
rect 28880 116880 29120 116900
rect 29380 116880 29620 116900
rect 29880 116880 30120 116900
rect 30380 116880 30620 116900
rect 30880 116880 31120 116900
rect 31380 116880 31620 116900
rect 31880 116880 32120 116900
rect 32380 116880 32620 116900
rect 32880 116880 33120 116900
rect 33380 116880 33620 116900
rect 33880 116880 34120 116900
rect 34380 116880 34620 116900
rect 34880 116880 35120 116900
rect 35380 116880 35620 116900
rect 35880 116880 36120 116900
rect 36380 116880 36620 116900
rect 36880 116880 37120 116900
rect 37380 116880 37620 116900
rect 37880 116880 38120 116900
rect 38380 116880 38620 116900
rect 38880 116880 39120 116900
rect 39380 116880 39620 116900
rect 39880 116880 40120 116900
rect 40380 116880 40620 116900
rect 40880 116880 41120 116900
rect 41380 116880 41620 116900
rect 41880 116880 42120 116900
rect 42380 116880 42620 116900
rect 42880 116880 43120 116900
rect 43380 116880 43620 116900
rect 43880 116880 44120 116900
rect 44380 116880 44620 116900
rect 44880 116880 45120 116900
rect 45380 116880 45620 116900
rect 45880 116880 46120 116900
rect 46380 116880 46620 116900
rect 46880 116880 47120 116900
rect 47380 116880 47620 116900
rect 47880 116880 48120 116900
rect 48380 116880 48620 116900
rect 48880 116880 49120 116900
rect 49380 116880 49620 116900
rect 49880 116880 50120 116900
rect 50380 116880 50620 116900
rect 50880 116880 51120 116900
rect 51380 116880 51620 116900
rect 51880 116880 52120 116900
rect 52380 116880 52620 116900
rect 52880 116880 53120 116900
rect 53380 116880 53620 116900
rect 53880 116880 54120 116900
rect 54380 116880 54620 116900
rect 54880 116880 55120 116900
rect 55380 116880 55620 116900
rect 55880 116880 56120 116900
rect 56380 116880 56620 116900
rect 56880 116880 57120 116900
rect 57380 116880 57620 116900
rect 57880 116880 58000 116900
rect 14000 116620 14100 116880
rect 14400 116620 14600 116880
rect 14900 116620 15100 116880
rect 15400 116620 15600 116880
rect 15900 116620 16100 116880
rect 16400 116620 16600 116880
rect 16900 116620 17100 116880
rect 17400 116620 17600 116880
rect 17900 116620 18100 116880
rect 18400 116620 18600 116880
rect 18900 116620 19100 116880
rect 19400 116620 19600 116880
rect 19900 116620 20100 116880
rect 20400 116620 20600 116880
rect 20900 116620 21100 116880
rect 21400 116620 21600 116880
rect 21900 116620 22100 116880
rect 22400 116620 22600 116880
rect 22900 116620 23100 116880
rect 23400 116620 23600 116880
rect 23900 116620 24100 116880
rect 24400 116620 24600 116880
rect 24900 116620 25100 116880
rect 25400 116620 25600 116880
rect 25900 116620 26100 116880
rect 26400 116620 26600 116880
rect 26900 116620 27100 116880
rect 27400 116620 27600 116880
rect 27900 116620 28100 116880
rect 28400 116620 28600 116880
rect 28900 116620 29100 116880
rect 29400 116620 29600 116880
rect 29900 116620 30100 116880
rect 30400 116620 30600 116880
rect 30900 116620 31100 116880
rect 31400 116620 31600 116880
rect 31900 116620 32100 116880
rect 32400 116620 32600 116880
rect 32900 116620 33100 116880
rect 33400 116620 33600 116880
rect 33900 116620 34100 116880
rect 34400 116620 34600 116880
rect 34900 116620 35100 116880
rect 35400 116620 35600 116880
rect 35900 116620 36100 116880
rect 36400 116620 36600 116880
rect 36900 116620 37100 116880
rect 37400 116620 37600 116880
rect 37900 116620 38100 116880
rect 38400 116620 38600 116880
rect 38900 116620 39100 116880
rect 39400 116620 39600 116880
rect 39900 116620 40100 116880
rect 40400 116620 40600 116880
rect 40900 116620 41100 116880
rect 41400 116620 41600 116880
rect 41900 116620 42100 116880
rect 42400 116620 42600 116880
rect 42900 116620 43100 116880
rect 43400 116620 43600 116880
rect 43900 116620 44100 116880
rect 44400 116620 44600 116880
rect 44900 116620 45100 116880
rect 45400 116620 45600 116880
rect 45900 116620 46100 116880
rect 46400 116620 46600 116880
rect 46900 116620 47100 116880
rect 47400 116620 47600 116880
rect 47900 116620 48100 116880
rect 48400 116620 48600 116880
rect 48900 116620 49100 116880
rect 49400 116620 49600 116880
rect 49900 116620 50100 116880
rect 50400 116620 50600 116880
rect 50900 116620 51100 116880
rect 51400 116620 51600 116880
rect 51900 116620 52100 116880
rect 52400 116620 52600 116880
rect 52900 116620 53100 116880
rect 53400 116620 53600 116880
rect 53900 116620 54100 116880
rect 54400 116620 54600 116880
rect 54900 116620 55100 116880
rect 55400 116620 55600 116880
rect 55900 116620 56100 116880
rect 56400 116620 56600 116880
rect 56900 116620 57100 116880
rect 57400 116620 57600 116880
rect 57900 116620 58000 116880
rect 14000 116600 14120 116620
rect 14380 116600 14620 116620
rect 14880 116600 15120 116620
rect 15380 116600 15620 116620
rect 15880 116600 16120 116620
rect 16380 116600 16620 116620
rect 16880 116600 17120 116620
rect 17380 116600 17620 116620
rect 17880 116600 18120 116620
rect 18380 116600 18620 116620
rect 18880 116600 19120 116620
rect 19380 116600 19620 116620
rect 19880 116600 20120 116620
rect 20380 116600 20620 116620
rect 20880 116600 21120 116620
rect 21380 116600 21620 116620
rect 21880 116600 22120 116620
rect 22380 116600 22620 116620
rect 22880 116600 23120 116620
rect 23380 116600 23620 116620
rect 23880 116600 24120 116620
rect 24380 116600 24620 116620
rect 24880 116600 25120 116620
rect 25380 116600 25620 116620
rect 25880 116600 26120 116620
rect 26380 116600 26620 116620
rect 26880 116600 27120 116620
rect 27380 116600 27620 116620
rect 27880 116600 28120 116620
rect 28380 116600 28620 116620
rect 28880 116600 29120 116620
rect 29380 116600 29620 116620
rect 29880 116600 30120 116620
rect 30380 116600 30620 116620
rect 30880 116600 31120 116620
rect 31380 116600 31620 116620
rect 31880 116600 32120 116620
rect 32380 116600 32620 116620
rect 32880 116600 33120 116620
rect 33380 116600 33620 116620
rect 33880 116600 34120 116620
rect 34380 116600 34620 116620
rect 34880 116600 35120 116620
rect 35380 116600 35620 116620
rect 35880 116600 36120 116620
rect 36380 116600 36620 116620
rect 36880 116600 37120 116620
rect 37380 116600 37620 116620
rect 37880 116600 38120 116620
rect 38380 116600 38620 116620
rect 38880 116600 39120 116620
rect 39380 116600 39620 116620
rect 39880 116600 40120 116620
rect 40380 116600 40620 116620
rect 40880 116600 41120 116620
rect 41380 116600 41620 116620
rect 41880 116600 42120 116620
rect 42380 116600 42620 116620
rect 42880 116600 43120 116620
rect 43380 116600 43620 116620
rect 43880 116600 44120 116620
rect 44380 116600 44620 116620
rect 44880 116600 45120 116620
rect 45380 116600 45620 116620
rect 45880 116600 46120 116620
rect 46380 116600 46620 116620
rect 46880 116600 47120 116620
rect 47380 116600 47620 116620
rect 47880 116600 48120 116620
rect 48380 116600 48620 116620
rect 48880 116600 49120 116620
rect 49380 116600 49620 116620
rect 49880 116600 50120 116620
rect 50380 116600 50620 116620
rect 50880 116600 51120 116620
rect 51380 116600 51620 116620
rect 51880 116600 52120 116620
rect 52380 116600 52620 116620
rect 52880 116600 53120 116620
rect 53380 116600 53620 116620
rect 53880 116600 54120 116620
rect 54380 116600 54620 116620
rect 54880 116600 55120 116620
rect 55380 116600 55620 116620
rect 55880 116600 56120 116620
rect 56380 116600 56620 116620
rect 56880 116600 57120 116620
rect 57380 116600 57620 116620
rect 57880 116600 58000 116620
rect 14000 116400 58000 116600
rect 14000 116380 14120 116400
rect 14380 116380 14620 116400
rect 14880 116380 15120 116400
rect 15380 116380 15620 116400
rect 15880 116380 16120 116400
rect 16380 116380 16620 116400
rect 16880 116380 17120 116400
rect 17380 116380 17620 116400
rect 17880 116380 18120 116400
rect 18380 116380 18620 116400
rect 18880 116380 19120 116400
rect 19380 116380 19620 116400
rect 19880 116380 20120 116400
rect 20380 116380 20620 116400
rect 20880 116380 21120 116400
rect 21380 116380 21620 116400
rect 21880 116380 22120 116400
rect 22380 116380 22620 116400
rect 22880 116380 23120 116400
rect 23380 116380 23620 116400
rect 23880 116380 24120 116400
rect 24380 116380 24620 116400
rect 24880 116380 25120 116400
rect 25380 116380 25620 116400
rect 25880 116380 26120 116400
rect 26380 116380 26620 116400
rect 26880 116380 27120 116400
rect 27380 116380 27620 116400
rect 27880 116380 28120 116400
rect 28380 116380 28620 116400
rect 28880 116380 29120 116400
rect 29380 116380 29620 116400
rect 29880 116380 30120 116400
rect 30380 116380 30620 116400
rect 30880 116380 31120 116400
rect 31380 116380 31620 116400
rect 31880 116380 32120 116400
rect 32380 116380 32620 116400
rect 32880 116380 33120 116400
rect 33380 116380 33620 116400
rect 33880 116380 34120 116400
rect 34380 116380 34620 116400
rect 34880 116380 35120 116400
rect 35380 116380 35620 116400
rect 35880 116380 36120 116400
rect 36380 116380 36620 116400
rect 36880 116380 37120 116400
rect 37380 116380 37620 116400
rect 37880 116380 38120 116400
rect 38380 116380 38620 116400
rect 38880 116380 39120 116400
rect 39380 116380 39620 116400
rect 39880 116380 40120 116400
rect 40380 116380 40620 116400
rect 40880 116380 41120 116400
rect 41380 116380 41620 116400
rect 41880 116380 42120 116400
rect 42380 116380 42620 116400
rect 42880 116380 43120 116400
rect 43380 116380 43620 116400
rect 43880 116380 44120 116400
rect 44380 116380 44620 116400
rect 44880 116380 45120 116400
rect 45380 116380 45620 116400
rect 45880 116380 46120 116400
rect 46380 116380 46620 116400
rect 46880 116380 47120 116400
rect 47380 116380 47620 116400
rect 47880 116380 48120 116400
rect 48380 116380 48620 116400
rect 48880 116380 49120 116400
rect 49380 116380 49620 116400
rect 49880 116380 50120 116400
rect 50380 116380 50620 116400
rect 50880 116380 51120 116400
rect 51380 116380 51620 116400
rect 51880 116380 52120 116400
rect 52380 116380 52620 116400
rect 52880 116380 53120 116400
rect 53380 116380 53620 116400
rect 53880 116380 54120 116400
rect 54380 116380 54620 116400
rect 54880 116380 55120 116400
rect 55380 116380 55620 116400
rect 55880 116380 56120 116400
rect 56380 116380 56620 116400
rect 56880 116380 57120 116400
rect 57380 116380 57620 116400
rect 57880 116380 58000 116400
rect 14000 116120 14100 116380
rect 14400 116120 14600 116380
rect 14900 116120 15100 116380
rect 15400 116120 15600 116380
rect 15900 116120 16100 116380
rect 16400 116120 16600 116380
rect 16900 116120 17100 116380
rect 17400 116120 17600 116380
rect 17900 116120 18100 116380
rect 18400 116120 18600 116380
rect 18900 116120 19100 116380
rect 19400 116120 19600 116380
rect 19900 116120 20100 116380
rect 20400 116120 20600 116380
rect 20900 116120 21100 116380
rect 21400 116120 21600 116380
rect 21900 116120 22100 116380
rect 22400 116120 22600 116380
rect 22900 116120 23100 116380
rect 23400 116120 23600 116380
rect 23900 116120 24100 116380
rect 24400 116120 24600 116380
rect 24900 116120 25100 116380
rect 25400 116120 25600 116380
rect 25900 116120 26100 116380
rect 26400 116120 26600 116380
rect 26900 116120 27100 116380
rect 27400 116120 27600 116380
rect 27900 116120 28100 116380
rect 28400 116120 28600 116380
rect 28900 116120 29100 116380
rect 29400 116120 29600 116380
rect 29900 116120 30100 116380
rect 30400 116120 30600 116380
rect 30900 116120 31100 116380
rect 31400 116120 31600 116380
rect 31900 116120 32100 116380
rect 32400 116120 32600 116380
rect 32900 116120 33100 116380
rect 33400 116120 33600 116380
rect 33900 116120 34100 116380
rect 34400 116120 34600 116380
rect 34900 116120 35100 116380
rect 35400 116120 35600 116380
rect 35900 116120 36100 116380
rect 36400 116120 36600 116380
rect 36900 116120 37100 116380
rect 37400 116120 37600 116380
rect 37900 116120 38100 116380
rect 38400 116120 38600 116380
rect 38900 116120 39100 116380
rect 39400 116120 39600 116380
rect 39900 116120 40100 116380
rect 40400 116120 40600 116380
rect 40900 116120 41100 116380
rect 41400 116120 41600 116380
rect 41900 116120 42100 116380
rect 42400 116120 42600 116380
rect 42900 116120 43100 116380
rect 43400 116120 43600 116380
rect 43900 116120 44100 116380
rect 44400 116120 44600 116380
rect 44900 116120 45100 116380
rect 45400 116120 45600 116380
rect 45900 116120 46100 116380
rect 46400 116120 46600 116380
rect 46900 116120 47100 116380
rect 47400 116120 47600 116380
rect 47900 116120 48100 116380
rect 48400 116120 48600 116380
rect 48900 116120 49100 116380
rect 49400 116120 49600 116380
rect 49900 116120 50100 116380
rect 50400 116120 50600 116380
rect 50900 116120 51100 116380
rect 51400 116120 51600 116380
rect 51900 116120 52100 116380
rect 52400 116120 52600 116380
rect 52900 116120 53100 116380
rect 53400 116120 53600 116380
rect 53900 116120 54100 116380
rect 54400 116120 54600 116380
rect 54900 116120 55100 116380
rect 55400 116120 55600 116380
rect 55900 116120 56100 116380
rect 56400 116120 56600 116380
rect 56900 116120 57100 116380
rect 57400 116120 57600 116380
rect 57900 116120 58000 116380
rect 14000 116100 14120 116120
rect 14380 116100 14620 116120
rect 14880 116100 15120 116120
rect 15380 116100 15620 116120
rect 15880 116100 16120 116120
rect 16380 116100 16620 116120
rect 16880 116100 17120 116120
rect 17380 116100 17620 116120
rect 17880 116100 18120 116120
rect 18380 116100 18620 116120
rect 18880 116100 19120 116120
rect 19380 116100 19620 116120
rect 19880 116100 20120 116120
rect 20380 116100 20620 116120
rect 20880 116100 21120 116120
rect 21380 116100 21620 116120
rect 21880 116100 22120 116120
rect 22380 116100 22620 116120
rect 22880 116100 23120 116120
rect 23380 116100 23620 116120
rect 23880 116100 24120 116120
rect 24380 116100 24620 116120
rect 24880 116100 25120 116120
rect 25380 116100 25620 116120
rect 25880 116100 26120 116120
rect 26380 116100 26620 116120
rect 26880 116100 27120 116120
rect 27380 116100 27620 116120
rect 27880 116100 28120 116120
rect 28380 116100 28620 116120
rect 28880 116100 29120 116120
rect 29380 116100 29620 116120
rect 29880 116100 30120 116120
rect 30380 116100 30620 116120
rect 30880 116100 31120 116120
rect 31380 116100 31620 116120
rect 31880 116100 32120 116120
rect 32380 116100 32620 116120
rect 32880 116100 33120 116120
rect 33380 116100 33620 116120
rect 33880 116100 34120 116120
rect 34380 116100 34620 116120
rect 34880 116100 35120 116120
rect 35380 116100 35620 116120
rect 35880 116100 36120 116120
rect 36380 116100 36620 116120
rect 36880 116100 37120 116120
rect 37380 116100 37620 116120
rect 37880 116100 38120 116120
rect 38380 116100 38620 116120
rect 38880 116100 39120 116120
rect 39380 116100 39620 116120
rect 39880 116100 40120 116120
rect 40380 116100 40620 116120
rect 40880 116100 41120 116120
rect 41380 116100 41620 116120
rect 41880 116100 42120 116120
rect 42380 116100 42620 116120
rect 42880 116100 43120 116120
rect 43380 116100 43620 116120
rect 43880 116100 44120 116120
rect 44380 116100 44620 116120
rect 44880 116100 45120 116120
rect 45380 116100 45620 116120
rect 45880 116100 46120 116120
rect 46380 116100 46620 116120
rect 46880 116100 47120 116120
rect 47380 116100 47620 116120
rect 47880 116100 48120 116120
rect 48380 116100 48620 116120
rect 48880 116100 49120 116120
rect 49380 116100 49620 116120
rect 49880 116100 50120 116120
rect 50380 116100 50620 116120
rect 50880 116100 51120 116120
rect 51380 116100 51620 116120
rect 51880 116100 52120 116120
rect 52380 116100 52620 116120
rect 52880 116100 53120 116120
rect 53380 116100 53620 116120
rect 53880 116100 54120 116120
rect 54380 116100 54620 116120
rect 54880 116100 55120 116120
rect 55380 116100 55620 116120
rect 55880 116100 56120 116120
rect 56380 116100 56620 116120
rect 56880 116100 57120 116120
rect 57380 116100 57620 116120
rect 57880 116100 58000 116120
rect 14000 115900 58000 116100
rect 14000 115880 14120 115900
rect 14380 115880 14620 115900
rect 14880 115880 15120 115900
rect 15380 115880 15620 115900
rect 15880 115880 16120 115900
rect 16380 115880 16620 115900
rect 16880 115880 17120 115900
rect 17380 115880 17620 115900
rect 17880 115880 18120 115900
rect 18380 115880 18620 115900
rect 18880 115880 19120 115900
rect 19380 115880 19620 115900
rect 19880 115880 20120 115900
rect 20380 115880 20620 115900
rect 20880 115880 21120 115900
rect 21380 115880 21620 115900
rect 21880 115880 22120 115900
rect 22380 115880 22620 115900
rect 22880 115880 23120 115900
rect 23380 115880 23620 115900
rect 23880 115880 24120 115900
rect 24380 115880 24620 115900
rect 24880 115880 25120 115900
rect 25380 115880 25620 115900
rect 25880 115880 26120 115900
rect 26380 115880 26620 115900
rect 26880 115880 27120 115900
rect 27380 115880 27620 115900
rect 27880 115880 28120 115900
rect 28380 115880 28620 115900
rect 28880 115880 29120 115900
rect 29380 115880 29620 115900
rect 29880 115880 30120 115900
rect 30380 115880 30620 115900
rect 30880 115880 31120 115900
rect 31380 115880 31620 115900
rect 31880 115880 32120 115900
rect 32380 115880 32620 115900
rect 32880 115880 33120 115900
rect 33380 115880 33620 115900
rect 33880 115880 34120 115900
rect 34380 115880 34620 115900
rect 34880 115880 35120 115900
rect 35380 115880 35620 115900
rect 35880 115880 36120 115900
rect 36380 115880 36620 115900
rect 36880 115880 37120 115900
rect 37380 115880 37620 115900
rect 37880 115880 38120 115900
rect 38380 115880 38620 115900
rect 38880 115880 39120 115900
rect 39380 115880 39620 115900
rect 39880 115880 40120 115900
rect 40380 115880 40620 115900
rect 40880 115880 41120 115900
rect 41380 115880 41620 115900
rect 41880 115880 42120 115900
rect 42380 115880 42620 115900
rect 42880 115880 43120 115900
rect 43380 115880 43620 115900
rect 43880 115880 44120 115900
rect 44380 115880 44620 115900
rect 44880 115880 45120 115900
rect 45380 115880 45620 115900
rect 45880 115880 46120 115900
rect 46380 115880 46620 115900
rect 46880 115880 47120 115900
rect 47380 115880 47620 115900
rect 47880 115880 48120 115900
rect 48380 115880 48620 115900
rect 48880 115880 49120 115900
rect 49380 115880 49620 115900
rect 49880 115880 50120 115900
rect 50380 115880 50620 115900
rect 50880 115880 51120 115900
rect 51380 115880 51620 115900
rect 51880 115880 52120 115900
rect 52380 115880 52620 115900
rect 52880 115880 53120 115900
rect 53380 115880 53620 115900
rect 53880 115880 54120 115900
rect 54380 115880 54620 115900
rect 54880 115880 55120 115900
rect 55380 115880 55620 115900
rect 55880 115880 56120 115900
rect 56380 115880 56620 115900
rect 56880 115880 57120 115900
rect 57380 115880 57620 115900
rect 57880 115880 58000 115900
rect 14000 115620 14100 115880
rect 14400 115620 14600 115880
rect 14900 115620 15100 115880
rect 15400 115620 15600 115880
rect 15900 115620 16100 115880
rect 16400 115620 16600 115880
rect 16900 115620 17100 115880
rect 17400 115620 17600 115880
rect 17900 115620 18100 115880
rect 18400 115620 18600 115880
rect 18900 115620 19100 115880
rect 19400 115620 19600 115880
rect 19900 115620 20100 115880
rect 20400 115620 20600 115880
rect 20900 115620 21100 115880
rect 21400 115620 21600 115880
rect 21900 115620 22100 115880
rect 22400 115620 22600 115880
rect 22900 115620 23100 115880
rect 23400 115620 23600 115880
rect 23900 115620 24100 115880
rect 24400 115620 24600 115880
rect 24900 115620 25100 115880
rect 25400 115620 25600 115880
rect 25900 115620 26100 115880
rect 26400 115620 26600 115880
rect 26900 115620 27100 115880
rect 27400 115620 27600 115880
rect 27900 115620 28100 115880
rect 28400 115620 28600 115880
rect 28900 115620 29100 115880
rect 29400 115620 29600 115880
rect 29900 115620 30100 115880
rect 30400 115620 30600 115880
rect 30900 115620 31100 115880
rect 31400 115620 31600 115880
rect 31900 115620 32100 115880
rect 32400 115620 32600 115880
rect 32900 115620 33100 115880
rect 33400 115620 33600 115880
rect 33900 115620 34100 115880
rect 34400 115620 34600 115880
rect 34900 115620 35100 115880
rect 35400 115620 35600 115880
rect 35900 115620 36100 115880
rect 36400 115620 36600 115880
rect 36900 115620 37100 115880
rect 37400 115620 37600 115880
rect 37900 115620 38100 115880
rect 38400 115620 38600 115880
rect 38900 115620 39100 115880
rect 39400 115620 39600 115880
rect 39900 115620 40100 115880
rect 40400 115620 40600 115880
rect 40900 115620 41100 115880
rect 41400 115620 41600 115880
rect 41900 115620 42100 115880
rect 42400 115620 42600 115880
rect 42900 115620 43100 115880
rect 43400 115620 43600 115880
rect 43900 115620 44100 115880
rect 44400 115620 44600 115880
rect 44900 115620 45100 115880
rect 45400 115620 45600 115880
rect 45900 115620 46100 115880
rect 46400 115620 46600 115880
rect 46900 115620 47100 115880
rect 47400 115620 47600 115880
rect 47900 115620 48100 115880
rect 48400 115620 48600 115880
rect 48900 115620 49100 115880
rect 49400 115620 49600 115880
rect 49900 115620 50100 115880
rect 50400 115620 50600 115880
rect 50900 115620 51100 115880
rect 51400 115620 51600 115880
rect 51900 115620 52100 115880
rect 52400 115620 52600 115880
rect 52900 115620 53100 115880
rect 53400 115620 53600 115880
rect 53900 115620 54100 115880
rect 54400 115620 54600 115880
rect 54900 115620 55100 115880
rect 55400 115620 55600 115880
rect 55900 115620 56100 115880
rect 56400 115620 56600 115880
rect 56900 115620 57100 115880
rect 57400 115620 57600 115880
rect 57900 115620 58000 115880
rect 14000 115600 14120 115620
rect 14380 115600 14620 115620
rect 14880 115600 15120 115620
rect 15380 115600 15620 115620
rect 15880 115600 16120 115620
rect 16380 115600 16620 115620
rect 16880 115600 17120 115620
rect 17380 115600 17620 115620
rect 17880 115600 18120 115620
rect 18380 115600 18620 115620
rect 18880 115600 19120 115620
rect 19380 115600 19620 115620
rect 19880 115600 20120 115620
rect 20380 115600 20620 115620
rect 20880 115600 21120 115620
rect 21380 115600 21620 115620
rect 21880 115600 22120 115620
rect 22380 115600 22620 115620
rect 22880 115600 23120 115620
rect 23380 115600 23620 115620
rect 23880 115600 24120 115620
rect 24380 115600 24620 115620
rect 24880 115600 25120 115620
rect 25380 115600 25620 115620
rect 25880 115600 26120 115620
rect 26380 115600 26620 115620
rect 26880 115600 27120 115620
rect 27380 115600 27620 115620
rect 27880 115600 28120 115620
rect 28380 115600 28620 115620
rect 28880 115600 29120 115620
rect 29380 115600 29620 115620
rect 29880 115600 30120 115620
rect 30380 115600 30620 115620
rect 30880 115600 31120 115620
rect 31380 115600 31620 115620
rect 31880 115600 32120 115620
rect 32380 115600 32620 115620
rect 32880 115600 33120 115620
rect 33380 115600 33620 115620
rect 33880 115600 34120 115620
rect 34380 115600 34620 115620
rect 34880 115600 35120 115620
rect 35380 115600 35620 115620
rect 35880 115600 36120 115620
rect 36380 115600 36620 115620
rect 36880 115600 37120 115620
rect 37380 115600 37620 115620
rect 37880 115600 38120 115620
rect 38380 115600 38620 115620
rect 38880 115600 39120 115620
rect 39380 115600 39620 115620
rect 39880 115600 40120 115620
rect 40380 115600 40620 115620
rect 40880 115600 41120 115620
rect 41380 115600 41620 115620
rect 41880 115600 42120 115620
rect 42380 115600 42620 115620
rect 42880 115600 43120 115620
rect 43380 115600 43620 115620
rect 43880 115600 44120 115620
rect 44380 115600 44620 115620
rect 44880 115600 45120 115620
rect 45380 115600 45620 115620
rect 45880 115600 46120 115620
rect 46380 115600 46620 115620
rect 46880 115600 47120 115620
rect 47380 115600 47620 115620
rect 47880 115600 48120 115620
rect 48380 115600 48620 115620
rect 48880 115600 49120 115620
rect 49380 115600 49620 115620
rect 49880 115600 50120 115620
rect 50380 115600 50620 115620
rect 50880 115600 51120 115620
rect 51380 115600 51620 115620
rect 51880 115600 52120 115620
rect 52380 115600 52620 115620
rect 52880 115600 53120 115620
rect 53380 115600 53620 115620
rect 53880 115600 54120 115620
rect 54380 115600 54620 115620
rect 54880 115600 55120 115620
rect 55380 115600 55620 115620
rect 55880 115600 56120 115620
rect 56380 115600 56620 115620
rect 56880 115600 57120 115620
rect 57380 115600 57620 115620
rect 57880 115600 58000 115620
rect 14000 115400 58000 115600
rect 14000 115380 14120 115400
rect 14380 115380 14620 115400
rect 14880 115380 15120 115400
rect 15380 115380 15620 115400
rect 15880 115380 16120 115400
rect 16380 115380 16620 115400
rect 16880 115380 17120 115400
rect 17380 115380 17620 115400
rect 17880 115380 18120 115400
rect 18380 115380 18620 115400
rect 18880 115380 19120 115400
rect 19380 115380 19620 115400
rect 19880 115380 20120 115400
rect 20380 115380 20620 115400
rect 20880 115380 21120 115400
rect 21380 115380 21620 115400
rect 21880 115380 22120 115400
rect 22380 115380 22620 115400
rect 22880 115380 23120 115400
rect 23380 115380 23620 115400
rect 23880 115380 24120 115400
rect 24380 115380 24620 115400
rect 24880 115380 25120 115400
rect 25380 115380 25620 115400
rect 25880 115380 26120 115400
rect 26380 115380 26620 115400
rect 26880 115380 27120 115400
rect 27380 115380 27620 115400
rect 27880 115380 28120 115400
rect 28380 115380 28620 115400
rect 28880 115380 29120 115400
rect 29380 115380 29620 115400
rect 29880 115380 30120 115400
rect 30380 115380 30620 115400
rect 30880 115380 31120 115400
rect 31380 115380 31620 115400
rect 31880 115380 32120 115400
rect 32380 115380 32620 115400
rect 32880 115380 33120 115400
rect 33380 115380 33620 115400
rect 33880 115380 34120 115400
rect 34380 115380 34620 115400
rect 34880 115380 35120 115400
rect 35380 115380 35620 115400
rect 35880 115380 36120 115400
rect 36380 115380 36620 115400
rect 36880 115380 37120 115400
rect 37380 115380 37620 115400
rect 37880 115380 38120 115400
rect 38380 115380 38620 115400
rect 38880 115380 39120 115400
rect 39380 115380 39620 115400
rect 39880 115380 40120 115400
rect 40380 115380 40620 115400
rect 40880 115380 41120 115400
rect 41380 115380 41620 115400
rect 41880 115380 42120 115400
rect 42380 115380 42620 115400
rect 42880 115380 43120 115400
rect 43380 115380 43620 115400
rect 43880 115380 44120 115400
rect 44380 115380 44620 115400
rect 44880 115380 45120 115400
rect 45380 115380 45620 115400
rect 45880 115380 46120 115400
rect 46380 115380 46620 115400
rect 46880 115380 47120 115400
rect 47380 115380 47620 115400
rect 47880 115380 48120 115400
rect 48380 115380 48620 115400
rect 48880 115380 49120 115400
rect 49380 115380 49620 115400
rect 49880 115380 50120 115400
rect 50380 115380 50620 115400
rect 50880 115380 51120 115400
rect 51380 115380 51620 115400
rect 51880 115380 52120 115400
rect 52380 115380 52620 115400
rect 52880 115380 53120 115400
rect 53380 115380 53620 115400
rect 53880 115380 54120 115400
rect 54380 115380 54620 115400
rect 54880 115380 55120 115400
rect 55380 115380 55620 115400
rect 55880 115380 56120 115400
rect 56380 115380 56620 115400
rect 56880 115380 57120 115400
rect 57380 115380 57620 115400
rect 57880 115380 58000 115400
rect 14000 115120 14100 115380
rect 14400 115120 14600 115380
rect 14900 115120 15100 115380
rect 15400 115120 15600 115380
rect 15900 115120 16100 115380
rect 16400 115120 16600 115380
rect 16900 115120 17100 115380
rect 17400 115120 17600 115380
rect 17900 115120 18100 115380
rect 18400 115120 18600 115380
rect 18900 115120 19100 115380
rect 19400 115120 19600 115380
rect 19900 115120 20100 115380
rect 20400 115120 20600 115380
rect 20900 115120 21100 115380
rect 21400 115120 21600 115380
rect 21900 115120 22100 115380
rect 22400 115120 22600 115380
rect 22900 115120 23100 115380
rect 23400 115120 23600 115380
rect 23900 115120 24100 115380
rect 24400 115120 24600 115380
rect 24900 115120 25100 115380
rect 25400 115120 25600 115380
rect 25900 115120 26100 115380
rect 26400 115120 26600 115380
rect 26900 115120 27100 115380
rect 27400 115120 27600 115380
rect 27900 115120 28100 115380
rect 28400 115120 28600 115380
rect 28900 115120 29100 115380
rect 29400 115120 29600 115380
rect 29900 115120 30100 115380
rect 30400 115120 30600 115380
rect 30900 115120 31100 115380
rect 31400 115120 31600 115380
rect 31900 115120 32100 115380
rect 32400 115120 32600 115380
rect 32900 115120 33100 115380
rect 33400 115120 33600 115380
rect 33900 115120 34100 115380
rect 34400 115120 34600 115380
rect 34900 115120 35100 115380
rect 35400 115120 35600 115380
rect 35900 115120 36100 115380
rect 36400 115120 36600 115380
rect 36900 115120 37100 115380
rect 37400 115120 37600 115380
rect 37900 115120 38100 115380
rect 38400 115120 38600 115380
rect 38900 115120 39100 115380
rect 39400 115120 39600 115380
rect 39900 115120 40100 115380
rect 40400 115120 40600 115380
rect 40900 115120 41100 115380
rect 41400 115120 41600 115380
rect 41900 115120 42100 115380
rect 42400 115120 42600 115380
rect 42900 115120 43100 115380
rect 43400 115120 43600 115380
rect 43900 115120 44100 115380
rect 44400 115120 44600 115380
rect 44900 115120 45100 115380
rect 45400 115120 45600 115380
rect 45900 115120 46100 115380
rect 46400 115120 46600 115380
rect 46900 115120 47100 115380
rect 47400 115120 47600 115380
rect 47900 115120 48100 115380
rect 48400 115120 48600 115380
rect 48900 115120 49100 115380
rect 49400 115120 49600 115380
rect 49900 115120 50100 115380
rect 50400 115120 50600 115380
rect 50900 115120 51100 115380
rect 51400 115120 51600 115380
rect 51900 115120 52100 115380
rect 52400 115120 52600 115380
rect 52900 115120 53100 115380
rect 53400 115120 53600 115380
rect 53900 115120 54100 115380
rect 54400 115120 54600 115380
rect 54900 115120 55100 115380
rect 55400 115120 55600 115380
rect 55900 115120 56100 115380
rect 56400 115120 56600 115380
rect 56900 115120 57100 115380
rect 57400 115120 57600 115380
rect 57900 115120 58000 115380
rect 14000 115100 14120 115120
rect 14380 115100 14620 115120
rect 14880 115100 15120 115120
rect 15380 115100 15620 115120
rect 15880 115100 16120 115120
rect 16380 115100 16620 115120
rect 16880 115100 17120 115120
rect 17380 115100 17620 115120
rect 17880 115100 18120 115120
rect 18380 115100 18620 115120
rect 18880 115100 19120 115120
rect 19380 115100 19620 115120
rect 19880 115100 20120 115120
rect 20380 115100 20620 115120
rect 20880 115100 21120 115120
rect 21380 115100 21620 115120
rect 21880 115100 22120 115120
rect 22380 115100 22620 115120
rect 22880 115100 23120 115120
rect 23380 115100 23620 115120
rect 23880 115100 24120 115120
rect 24380 115100 24620 115120
rect 24880 115100 25120 115120
rect 25380 115100 25620 115120
rect 25880 115100 26120 115120
rect 26380 115100 26620 115120
rect 26880 115100 27120 115120
rect 27380 115100 27620 115120
rect 27880 115100 28120 115120
rect 28380 115100 28620 115120
rect 28880 115100 29120 115120
rect 29380 115100 29620 115120
rect 29880 115100 30120 115120
rect 30380 115100 30620 115120
rect 30880 115100 31120 115120
rect 31380 115100 31620 115120
rect 31880 115100 32120 115120
rect 32380 115100 32620 115120
rect 32880 115100 33120 115120
rect 33380 115100 33620 115120
rect 33880 115100 34120 115120
rect 34380 115100 34620 115120
rect 34880 115100 35120 115120
rect 35380 115100 35620 115120
rect 35880 115100 36120 115120
rect 36380 115100 36620 115120
rect 36880 115100 37120 115120
rect 37380 115100 37620 115120
rect 37880 115100 38120 115120
rect 38380 115100 38620 115120
rect 38880 115100 39120 115120
rect 39380 115100 39620 115120
rect 39880 115100 40120 115120
rect 40380 115100 40620 115120
rect 40880 115100 41120 115120
rect 41380 115100 41620 115120
rect 41880 115100 42120 115120
rect 42380 115100 42620 115120
rect 42880 115100 43120 115120
rect 43380 115100 43620 115120
rect 43880 115100 44120 115120
rect 44380 115100 44620 115120
rect 44880 115100 45120 115120
rect 45380 115100 45620 115120
rect 45880 115100 46120 115120
rect 46380 115100 46620 115120
rect 46880 115100 47120 115120
rect 47380 115100 47620 115120
rect 47880 115100 48120 115120
rect 48380 115100 48620 115120
rect 48880 115100 49120 115120
rect 49380 115100 49620 115120
rect 49880 115100 50120 115120
rect 50380 115100 50620 115120
rect 50880 115100 51120 115120
rect 51380 115100 51620 115120
rect 51880 115100 52120 115120
rect 52380 115100 52620 115120
rect 52880 115100 53120 115120
rect 53380 115100 53620 115120
rect 53880 115100 54120 115120
rect 54380 115100 54620 115120
rect 54880 115100 55120 115120
rect 55380 115100 55620 115120
rect 55880 115100 56120 115120
rect 56380 115100 56620 115120
rect 56880 115100 57120 115120
rect 57380 115100 57620 115120
rect 57880 115100 58000 115120
rect 14000 114900 58000 115100
rect 14000 114880 14120 114900
rect 14380 114880 14620 114900
rect 14880 114880 15120 114900
rect 15380 114880 15620 114900
rect 15880 114880 16120 114900
rect 16380 114880 16620 114900
rect 16880 114880 17120 114900
rect 17380 114880 17620 114900
rect 17880 114880 18120 114900
rect 18380 114880 18620 114900
rect 18880 114880 19120 114900
rect 19380 114880 19620 114900
rect 19880 114880 20120 114900
rect 20380 114880 20620 114900
rect 20880 114880 21120 114900
rect 21380 114880 21620 114900
rect 21880 114880 22120 114900
rect 22380 114880 22620 114900
rect 22880 114880 23120 114900
rect 23380 114880 23620 114900
rect 23880 114880 24120 114900
rect 24380 114880 24620 114900
rect 24880 114880 25120 114900
rect 25380 114880 25620 114900
rect 25880 114880 26120 114900
rect 26380 114880 26620 114900
rect 26880 114880 27120 114900
rect 27380 114880 27620 114900
rect 27880 114880 28120 114900
rect 28380 114880 28620 114900
rect 28880 114880 29120 114900
rect 29380 114880 29620 114900
rect 29880 114880 30120 114900
rect 30380 114880 30620 114900
rect 30880 114880 31120 114900
rect 31380 114880 31620 114900
rect 31880 114880 32120 114900
rect 32380 114880 32620 114900
rect 32880 114880 33120 114900
rect 33380 114880 33620 114900
rect 33880 114880 34120 114900
rect 34380 114880 34620 114900
rect 34880 114880 35120 114900
rect 35380 114880 35620 114900
rect 35880 114880 36120 114900
rect 36380 114880 36620 114900
rect 36880 114880 37120 114900
rect 37380 114880 37620 114900
rect 37880 114880 38120 114900
rect 38380 114880 38620 114900
rect 38880 114880 39120 114900
rect 39380 114880 39620 114900
rect 39880 114880 40120 114900
rect 40380 114880 40620 114900
rect 40880 114880 41120 114900
rect 41380 114880 41620 114900
rect 41880 114880 42120 114900
rect 42380 114880 42620 114900
rect 42880 114880 43120 114900
rect 43380 114880 43620 114900
rect 43880 114880 44120 114900
rect 44380 114880 44620 114900
rect 44880 114880 45120 114900
rect 45380 114880 45620 114900
rect 45880 114880 46120 114900
rect 46380 114880 46620 114900
rect 46880 114880 47120 114900
rect 47380 114880 47620 114900
rect 47880 114880 48120 114900
rect 48380 114880 48620 114900
rect 48880 114880 49120 114900
rect 49380 114880 49620 114900
rect 49880 114880 50120 114900
rect 50380 114880 50620 114900
rect 50880 114880 51120 114900
rect 51380 114880 51620 114900
rect 51880 114880 52120 114900
rect 52380 114880 52620 114900
rect 52880 114880 53120 114900
rect 53380 114880 53620 114900
rect 53880 114880 54120 114900
rect 54380 114880 54620 114900
rect 54880 114880 55120 114900
rect 55380 114880 55620 114900
rect 55880 114880 56120 114900
rect 56380 114880 56620 114900
rect 56880 114880 57120 114900
rect 57380 114880 57620 114900
rect 57880 114880 58000 114900
rect 14000 114620 14100 114880
rect 14400 114620 14600 114880
rect 14900 114620 15100 114880
rect 15400 114620 15600 114880
rect 15900 114620 16100 114880
rect 16400 114620 16600 114880
rect 16900 114620 17100 114880
rect 17400 114620 17600 114880
rect 17900 114620 18100 114880
rect 18400 114620 18600 114880
rect 18900 114620 19100 114880
rect 19400 114620 19600 114880
rect 19900 114620 20100 114880
rect 20400 114620 20600 114880
rect 20900 114620 21100 114880
rect 21400 114620 21600 114880
rect 21900 114620 22100 114880
rect 22400 114620 22600 114880
rect 22900 114620 23100 114880
rect 23400 114620 23600 114880
rect 23900 114620 24100 114880
rect 24400 114620 24600 114880
rect 24900 114620 25100 114880
rect 25400 114620 25600 114880
rect 25900 114620 26100 114880
rect 26400 114620 26600 114880
rect 26900 114620 27100 114880
rect 27400 114620 27600 114880
rect 27900 114620 28100 114880
rect 28400 114620 28600 114880
rect 28900 114620 29100 114880
rect 29400 114620 29600 114880
rect 29900 114620 30100 114880
rect 30400 114620 30600 114880
rect 30900 114620 31100 114880
rect 31400 114620 31600 114880
rect 31900 114620 32100 114880
rect 32400 114620 32600 114880
rect 32900 114620 33100 114880
rect 33400 114620 33600 114880
rect 33900 114620 34100 114880
rect 34400 114620 34600 114880
rect 34900 114620 35100 114880
rect 35400 114620 35600 114880
rect 35900 114620 36100 114880
rect 36400 114620 36600 114880
rect 36900 114620 37100 114880
rect 37400 114620 37600 114880
rect 37900 114620 38100 114880
rect 38400 114620 38600 114880
rect 38900 114620 39100 114880
rect 39400 114620 39600 114880
rect 39900 114620 40100 114880
rect 40400 114620 40600 114880
rect 40900 114620 41100 114880
rect 41400 114620 41600 114880
rect 41900 114620 42100 114880
rect 42400 114620 42600 114880
rect 42900 114620 43100 114880
rect 43400 114620 43600 114880
rect 43900 114620 44100 114880
rect 44400 114620 44600 114880
rect 44900 114620 45100 114880
rect 45400 114620 45600 114880
rect 45900 114620 46100 114880
rect 46400 114620 46600 114880
rect 46900 114620 47100 114880
rect 47400 114620 47600 114880
rect 47900 114620 48100 114880
rect 48400 114620 48600 114880
rect 48900 114620 49100 114880
rect 49400 114620 49600 114880
rect 49900 114620 50100 114880
rect 50400 114620 50600 114880
rect 50900 114620 51100 114880
rect 51400 114620 51600 114880
rect 51900 114620 52100 114880
rect 52400 114620 52600 114880
rect 52900 114620 53100 114880
rect 53400 114620 53600 114880
rect 53900 114620 54100 114880
rect 54400 114620 54600 114880
rect 54900 114620 55100 114880
rect 55400 114620 55600 114880
rect 55900 114620 56100 114880
rect 56400 114620 56600 114880
rect 56900 114620 57100 114880
rect 57400 114620 57600 114880
rect 57900 114620 58000 114880
rect 14000 114600 14120 114620
rect 14380 114600 14620 114620
rect 14880 114600 15120 114620
rect 15380 114600 15620 114620
rect 15880 114600 16120 114620
rect 16380 114600 16620 114620
rect 16880 114600 17120 114620
rect 17380 114600 17620 114620
rect 17880 114600 18120 114620
rect 18380 114600 18620 114620
rect 18880 114600 19120 114620
rect 19380 114600 19620 114620
rect 19880 114600 20120 114620
rect 20380 114600 20620 114620
rect 20880 114600 21120 114620
rect 21380 114600 21620 114620
rect 21880 114600 22120 114620
rect 22380 114600 22620 114620
rect 22880 114600 23120 114620
rect 23380 114600 23620 114620
rect 23880 114600 24120 114620
rect 24380 114600 24620 114620
rect 24880 114600 25120 114620
rect 25380 114600 25620 114620
rect 25880 114600 26120 114620
rect 26380 114600 26620 114620
rect 26880 114600 27120 114620
rect 27380 114600 27620 114620
rect 27880 114600 28120 114620
rect 28380 114600 28620 114620
rect 28880 114600 29120 114620
rect 29380 114600 29620 114620
rect 29880 114600 30120 114620
rect 30380 114600 30620 114620
rect 30880 114600 31120 114620
rect 31380 114600 31620 114620
rect 31880 114600 32120 114620
rect 32380 114600 32620 114620
rect 32880 114600 33120 114620
rect 33380 114600 33620 114620
rect 33880 114600 34120 114620
rect 34380 114600 34620 114620
rect 34880 114600 35120 114620
rect 35380 114600 35620 114620
rect 35880 114600 36120 114620
rect 36380 114600 36620 114620
rect 36880 114600 37120 114620
rect 37380 114600 37620 114620
rect 37880 114600 38120 114620
rect 38380 114600 38620 114620
rect 38880 114600 39120 114620
rect 39380 114600 39620 114620
rect 39880 114600 40120 114620
rect 40380 114600 40620 114620
rect 40880 114600 41120 114620
rect 41380 114600 41620 114620
rect 41880 114600 42120 114620
rect 42380 114600 42620 114620
rect 42880 114600 43120 114620
rect 43380 114600 43620 114620
rect 43880 114600 44120 114620
rect 44380 114600 44620 114620
rect 44880 114600 45120 114620
rect 45380 114600 45620 114620
rect 45880 114600 46120 114620
rect 46380 114600 46620 114620
rect 46880 114600 47120 114620
rect 47380 114600 47620 114620
rect 47880 114600 48120 114620
rect 48380 114600 48620 114620
rect 48880 114600 49120 114620
rect 49380 114600 49620 114620
rect 49880 114600 50120 114620
rect 50380 114600 50620 114620
rect 50880 114600 51120 114620
rect 51380 114600 51620 114620
rect 51880 114600 52120 114620
rect 52380 114600 52620 114620
rect 52880 114600 53120 114620
rect 53380 114600 53620 114620
rect 53880 114600 54120 114620
rect 54380 114600 54620 114620
rect 54880 114600 55120 114620
rect 55380 114600 55620 114620
rect 55880 114600 56120 114620
rect 56380 114600 56620 114620
rect 56880 114600 57120 114620
rect 57380 114600 57620 114620
rect 57880 114600 58000 114620
rect 14000 114400 58000 114600
rect 14000 114380 14120 114400
rect 14380 114380 14620 114400
rect 14880 114380 15120 114400
rect 15380 114380 15620 114400
rect 15880 114380 16120 114400
rect 16380 114380 16620 114400
rect 16880 114380 17120 114400
rect 17380 114380 17620 114400
rect 17880 114380 18120 114400
rect 18380 114380 18620 114400
rect 18880 114380 19120 114400
rect 19380 114380 19620 114400
rect 19880 114380 20120 114400
rect 20380 114380 20620 114400
rect 20880 114380 21120 114400
rect 21380 114380 21620 114400
rect 21880 114380 22120 114400
rect 22380 114380 22620 114400
rect 22880 114380 23120 114400
rect 23380 114380 23620 114400
rect 23880 114380 24120 114400
rect 24380 114380 24620 114400
rect 24880 114380 25120 114400
rect 25380 114380 25620 114400
rect 25880 114380 26120 114400
rect 26380 114380 26620 114400
rect 26880 114380 27120 114400
rect 27380 114380 27620 114400
rect 27880 114380 28120 114400
rect 28380 114380 28620 114400
rect 28880 114380 29120 114400
rect 29380 114380 29620 114400
rect 29880 114380 30120 114400
rect 30380 114380 30620 114400
rect 30880 114380 31120 114400
rect 31380 114380 31620 114400
rect 31880 114380 32120 114400
rect 32380 114380 32620 114400
rect 32880 114380 33120 114400
rect 33380 114380 33620 114400
rect 33880 114380 34120 114400
rect 34380 114380 34620 114400
rect 34880 114380 35120 114400
rect 35380 114380 35620 114400
rect 35880 114380 36120 114400
rect 36380 114380 36620 114400
rect 36880 114380 37120 114400
rect 37380 114380 37620 114400
rect 37880 114380 38120 114400
rect 38380 114380 38620 114400
rect 38880 114380 39120 114400
rect 39380 114380 39620 114400
rect 39880 114380 40120 114400
rect 40380 114380 40620 114400
rect 40880 114380 41120 114400
rect 41380 114380 41620 114400
rect 41880 114380 42120 114400
rect 42380 114380 42620 114400
rect 42880 114380 43120 114400
rect 43380 114380 43620 114400
rect 43880 114380 44120 114400
rect 44380 114380 44620 114400
rect 44880 114380 45120 114400
rect 45380 114380 45620 114400
rect 45880 114380 46120 114400
rect 46380 114380 46620 114400
rect 46880 114380 47120 114400
rect 47380 114380 47620 114400
rect 47880 114380 48120 114400
rect 48380 114380 48620 114400
rect 48880 114380 49120 114400
rect 49380 114380 49620 114400
rect 49880 114380 50120 114400
rect 50380 114380 50620 114400
rect 50880 114380 51120 114400
rect 51380 114380 51620 114400
rect 51880 114380 52120 114400
rect 52380 114380 52620 114400
rect 52880 114380 53120 114400
rect 53380 114380 53620 114400
rect 53880 114380 54120 114400
rect 54380 114380 54620 114400
rect 54880 114380 55120 114400
rect 55380 114380 55620 114400
rect 55880 114380 56120 114400
rect 56380 114380 56620 114400
rect 56880 114380 57120 114400
rect 57380 114380 57620 114400
rect 57880 114380 58000 114400
rect 14000 114120 14100 114380
rect 14400 114120 14600 114380
rect 14900 114120 15100 114380
rect 15400 114120 15600 114380
rect 15900 114120 16100 114380
rect 16400 114120 16600 114380
rect 16900 114120 17100 114380
rect 17400 114120 17600 114380
rect 17900 114120 18100 114380
rect 18400 114120 18600 114380
rect 18900 114120 19100 114380
rect 19400 114120 19600 114380
rect 19900 114120 20100 114380
rect 20400 114120 20600 114380
rect 20900 114120 21100 114380
rect 21400 114120 21600 114380
rect 21900 114120 22100 114380
rect 22400 114120 22600 114380
rect 22900 114120 23100 114380
rect 23400 114120 23600 114380
rect 23900 114120 24100 114380
rect 24400 114120 24600 114380
rect 24900 114120 25100 114380
rect 25400 114120 25600 114380
rect 25900 114120 26100 114380
rect 26400 114120 26600 114380
rect 26900 114120 27100 114380
rect 27400 114120 27600 114380
rect 27900 114120 28100 114380
rect 28400 114120 28600 114380
rect 28900 114120 29100 114380
rect 29400 114120 29600 114380
rect 29900 114120 30100 114380
rect 30400 114120 30600 114380
rect 30900 114120 31100 114380
rect 31400 114120 31600 114380
rect 31900 114120 32100 114380
rect 32400 114120 32600 114380
rect 32900 114120 33100 114380
rect 33400 114120 33600 114380
rect 33900 114120 34100 114380
rect 34400 114120 34600 114380
rect 34900 114120 35100 114380
rect 35400 114120 35600 114380
rect 35900 114120 36100 114380
rect 36400 114120 36600 114380
rect 36900 114120 37100 114380
rect 37400 114120 37600 114380
rect 37900 114120 38100 114380
rect 38400 114120 38600 114380
rect 38900 114120 39100 114380
rect 39400 114120 39600 114380
rect 39900 114120 40100 114380
rect 40400 114120 40600 114380
rect 40900 114120 41100 114380
rect 41400 114120 41600 114380
rect 41900 114120 42100 114380
rect 42400 114120 42600 114380
rect 42900 114120 43100 114380
rect 43400 114120 43600 114380
rect 43900 114120 44100 114380
rect 44400 114120 44600 114380
rect 44900 114120 45100 114380
rect 45400 114120 45600 114380
rect 45900 114120 46100 114380
rect 46400 114120 46600 114380
rect 46900 114120 47100 114380
rect 47400 114120 47600 114380
rect 47900 114120 48100 114380
rect 48400 114120 48600 114380
rect 48900 114120 49100 114380
rect 49400 114120 49600 114380
rect 49900 114120 50100 114380
rect 50400 114120 50600 114380
rect 50900 114120 51100 114380
rect 51400 114120 51600 114380
rect 51900 114120 52100 114380
rect 52400 114120 52600 114380
rect 52900 114120 53100 114380
rect 53400 114120 53600 114380
rect 53900 114120 54100 114380
rect 54400 114120 54600 114380
rect 54900 114120 55100 114380
rect 55400 114120 55600 114380
rect 55900 114120 56100 114380
rect 56400 114120 56600 114380
rect 56900 114120 57100 114380
rect 57400 114120 57600 114380
rect 57900 114120 58000 114380
rect 14000 114100 14120 114120
rect 14380 114100 14620 114120
rect 14880 114100 15120 114120
rect 15380 114100 15620 114120
rect 15880 114100 16120 114120
rect 16380 114100 16620 114120
rect 16880 114100 17120 114120
rect 17380 114100 17620 114120
rect 17880 114100 18120 114120
rect 18380 114100 18620 114120
rect 18880 114100 19120 114120
rect 19380 114100 19620 114120
rect 19880 114100 20120 114120
rect 20380 114100 20620 114120
rect 20880 114100 21120 114120
rect 21380 114100 21620 114120
rect 21880 114100 22120 114120
rect 22380 114100 22620 114120
rect 22880 114100 23120 114120
rect 23380 114100 23620 114120
rect 23880 114100 24120 114120
rect 24380 114100 24620 114120
rect 24880 114100 25120 114120
rect 25380 114100 25620 114120
rect 25880 114100 26120 114120
rect 26380 114100 26620 114120
rect 26880 114100 27120 114120
rect 27380 114100 27620 114120
rect 27880 114100 28120 114120
rect 28380 114100 28620 114120
rect 28880 114100 29120 114120
rect 29380 114100 29620 114120
rect 29880 114100 30120 114120
rect 30380 114100 30620 114120
rect 30880 114100 31120 114120
rect 31380 114100 31620 114120
rect 31880 114100 32120 114120
rect 32380 114100 32620 114120
rect 32880 114100 33120 114120
rect 33380 114100 33620 114120
rect 33880 114100 34120 114120
rect 34380 114100 34620 114120
rect 34880 114100 35120 114120
rect 35380 114100 35620 114120
rect 35880 114100 36120 114120
rect 36380 114100 36620 114120
rect 36880 114100 37120 114120
rect 37380 114100 37620 114120
rect 37880 114100 38120 114120
rect 38380 114100 38620 114120
rect 38880 114100 39120 114120
rect 39380 114100 39620 114120
rect 39880 114100 40120 114120
rect 40380 114100 40620 114120
rect 40880 114100 41120 114120
rect 41380 114100 41620 114120
rect 41880 114100 42120 114120
rect 42380 114100 42620 114120
rect 42880 114100 43120 114120
rect 43380 114100 43620 114120
rect 43880 114100 44120 114120
rect 44380 114100 44620 114120
rect 44880 114100 45120 114120
rect 45380 114100 45620 114120
rect 45880 114100 46120 114120
rect 46380 114100 46620 114120
rect 46880 114100 47120 114120
rect 47380 114100 47620 114120
rect 47880 114100 48120 114120
rect 48380 114100 48620 114120
rect 48880 114100 49120 114120
rect 49380 114100 49620 114120
rect 49880 114100 50120 114120
rect 50380 114100 50620 114120
rect 50880 114100 51120 114120
rect 51380 114100 51620 114120
rect 51880 114100 52120 114120
rect 52380 114100 52620 114120
rect 52880 114100 53120 114120
rect 53380 114100 53620 114120
rect 53880 114100 54120 114120
rect 54380 114100 54620 114120
rect 54880 114100 55120 114120
rect 55380 114100 55620 114120
rect 55880 114100 56120 114120
rect 56380 114100 56620 114120
rect 56880 114100 57120 114120
rect 57380 114100 57620 114120
rect 57880 114100 58000 114120
rect 14000 114000 58000 114100
rect 118000 121900 142000 122000
rect 118000 121880 118120 121900
rect 118380 121880 118620 121900
rect 118880 121880 119120 121900
rect 119380 121880 119620 121900
rect 119880 121880 120120 121900
rect 120380 121880 120620 121900
rect 120880 121880 121120 121900
rect 121380 121880 121620 121900
rect 121880 121880 122120 121900
rect 122380 121880 122620 121900
rect 122880 121880 123120 121900
rect 123380 121880 123620 121900
rect 123880 121880 124120 121900
rect 124380 121880 124620 121900
rect 124880 121880 125120 121900
rect 125380 121880 125620 121900
rect 125880 121880 126120 121900
rect 126380 121880 126620 121900
rect 126880 121880 127120 121900
rect 127380 121880 127620 121900
rect 127880 121880 128120 121900
rect 128380 121880 128620 121900
rect 128880 121880 129120 121900
rect 129380 121880 129620 121900
rect 129880 121880 130120 121900
rect 130380 121880 130620 121900
rect 130880 121880 131120 121900
rect 131380 121880 131620 121900
rect 131880 121880 132120 121900
rect 132380 121880 132620 121900
rect 132880 121880 133120 121900
rect 133380 121880 133620 121900
rect 133880 121880 134120 121900
rect 134380 121880 134620 121900
rect 134880 121880 135120 121900
rect 135380 121880 135620 121900
rect 135880 121880 136120 121900
rect 136380 121880 136620 121900
rect 136880 121880 137120 121900
rect 137380 121880 137620 121900
rect 137880 121880 138120 121900
rect 138380 121880 138620 121900
rect 138880 121880 139120 121900
rect 139380 121880 139620 121900
rect 139880 121880 140120 121900
rect 140380 121880 140620 121900
rect 140880 121880 141120 121900
rect 141380 121880 141620 121900
rect 141880 121880 142000 121900
rect 118000 121620 118100 121880
rect 118400 121620 118600 121880
rect 118900 121620 119100 121880
rect 119400 121620 119600 121880
rect 119900 121620 120100 121880
rect 120400 121620 120600 121880
rect 120900 121620 121100 121880
rect 121400 121620 121600 121880
rect 121900 121620 122100 121880
rect 122400 121620 122600 121880
rect 122900 121620 123100 121880
rect 123400 121620 123600 121880
rect 123900 121620 124100 121880
rect 124400 121620 124600 121880
rect 124900 121620 125100 121880
rect 125400 121620 125600 121880
rect 125900 121620 126100 121880
rect 126400 121620 126600 121880
rect 126900 121620 127100 121880
rect 127400 121620 127600 121880
rect 127900 121620 128100 121880
rect 128400 121620 128600 121880
rect 128900 121620 129100 121880
rect 129400 121620 129600 121880
rect 129900 121620 130100 121880
rect 130400 121620 130600 121880
rect 130900 121620 131100 121880
rect 131400 121620 131600 121880
rect 131900 121620 132100 121880
rect 132400 121620 132600 121880
rect 132900 121620 133100 121880
rect 133400 121620 133600 121880
rect 133900 121620 134100 121880
rect 134400 121620 134600 121880
rect 134900 121620 135100 121880
rect 135400 121620 135600 121880
rect 135900 121620 136100 121880
rect 136400 121620 136600 121880
rect 136900 121620 137100 121880
rect 137400 121620 137600 121880
rect 137900 121620 138100 121880
rect 138400 121620 138600 121880
rect 138900 121620 139100 121880
rect 139400 121620 139600 121880
rect 139900 121620 140100 121880
rect 140400 121620 140600 121880
rect 140900 121620 141100 121880
rect 141400 121620 141600 121880
rect 141900 121620 142000 121880
rect 118000 121600 118120 121620
rect 118380 121600 118620 121620
rect 118880 121600 119120 121620
rect 119380 121600 119620 121620
rect 119880 121600 120120 121620
rect 120380 121600 120620 121620
rect 120880 121600 121120 121620
rect 121380 121600 121620 121620
rect 121880 121600 122120 121620
rect 122380 121600 122620 121620
rect 122880 121600 123120 121620
rect 123380 121600 123620 121620
rect 123880 121600 124120 121620
rect 124380 121600 124620 121620
rect 124880 121600 125120 121620
rect 125380 121600 125620 121620
rect 125880 121600 126120 121620
rect 126380 121600 126620 121620
rect 126880 121600 127120 121620
rect 127380 121600 127620 121620
rect 127880 121600 128120 121620
rect 128380 121600 128620 121620
rect 128880 121600 129120 121620
rect 129380 121600 129620 121620
rect 129880 121600 130120 121620
rect 130380 121600 130620 121620
rect 130880 121600 131120 121620
rect 131380 121600 131620 121620
rect 131880 121600 132120 121620
rect 132380 121600 132620 121620
rect 132880 121600 133120 121620
rect 133380 121600 133620 121620
rect 133880 121600 134120 121620
rect 134380 121600 134620 121620
rect 134880 121600 135120 121620
rect 135380 121600 135620 121620
rect 135880 121600 136120 121620
rect 136380 121600 136620 121620
rect 136880 121600 137120 121620
rect 137380 121600 137620 121620
rect 137880 121600 138120 121620
rect 138380 121600 138620 121620
rect 138880 121600 139120 121620
rect 139380 121600 139620 121620
rect 139880 121600 140120 121620
rect 140380 121600 140620 121620
rect 140880 121600 141120 121620
rect 141380 121600 141620 121620
rect 141880 121600 142000 121620
rect 118000 121400 142000 121600
rect 118000 121380 118120 121400
rect 118380 121380 118620 121400
rect 118880 121380 119120 121400
rect 119380 121380 119620 121400
rect 119880 121380 120120 121400
rect 120380 121380 120620 121400
rect 120880 121380 121120 121400
rect 121380 121380 121620 121400
rect 121880 121380 122120 121400
rect 122380 121380 122620 121400
rect 122880 121380 123120 121400
rect 123380 121380 123620 121400
rect 123880 121380 124120 121400
rect 124380 121380 124620 121400
rect 124880 121380 125120 121400
rect 125380 121380 125620 121400
rect 125880 121380 126120 121400
rect 126380 121380 126620 121400
rect 126880 121380 127120 121400
rect 127380 121380 127620 121400
rect 127880 121380 128120 121400
rect 128380 121380 128620 121400
rect 128880 121380 129120 121400
rect 129380 121380 129620 121400
rect 129880 121380 130120 121400
rect 130380 121380 130620 121400
rect 130880 121380 131120 121400
rect 131380 121380 131620 121400
rect 131880 121380 132120 121400
rect 132380 121380 132620 121400
rect 132880 121380 133120 121400
rect 133380 121380 133620 121400
rect 133880 121380 134120 121400
rect 134380 121380 134620 121400
rect 134880 121380 135120 121400
rect 135380 121380 135620 121400
rect 135880 121380 136120 121400
rect 136380 121380 136620 121400
rect 136880 121380 137120 121400
rect 137380 121380 137620 121400
rect 137880 121380 138120 121400
rect 138380 121380 138620 121400
rect 138880 121380 139120 121400
rect 139380 121380 139620 121400
rect 139880 121380 140120 121400
rect 140380 121380 140620 121400
rect 140880 121380 141120 121400
rect 141380 121380 141620 121400
rect 141880 121380 142000 121400
rect 118000 121120 118100 121380
rect 118400 121120 118600 121380
rect 118900 121120 119100 121380
rect 119400 121120 119600 121380
rect 119900 121120 120100 121380
rect 120400 121120 120600 121380
rect 120900 121120 121100 121380
rect 121400 121120 121600 121380
rect 121900 121120 122100 121380
rect 122400 121120 122600 121380
rect 122900 121120 123100 121380
rect 123400 121120 123600 121380
rect 123900 121120 124100 121380
rect 124400 121120 124600 121380
rect 124900 121120 125100 121380
rect 125400 121120 125600 121380
rect 125900 121120 126100 121380
rect 126400 121120 126600 121380
rect 126900 121120 127100 121380
rect 127400 121120 127600 121380
rect 127900 121120 128100 121380
rect 128400 121120 128600 121380
rect 128900 121120 129100 121380
rect 129400 121120 129600 121380
rect 129900 121120 130100 121380
rect 130400 121120 130600 121380
rect 130900 121120 131100 121380
rect 131400 121120 131600 121380
rect 131900 121120 132100 121380
rect 132400 121120 132600 121380
rect 132900 121120 133100 121380
rect 133400 121120 133600 121380
rect 133900 121120 134100 121380
rect 134400 121120 134600 121380
rect 134900 121120 135100 121380
rect 135400 121120 135600 121380
rect 135900 121120 136100 121380
rect 136400 121120 136600 121380
rect 136900 121120 137100 121380
rect 137400 121120 137600 121380
rect 137900 121120 138100 121380
rect 138400 121120 138600 121380
rect 138900 121120 139100 121380
rect 139400 121120 139600 121380
rect 139900 121120 140100 121380
rect 140400 121120 140600 121380
rect 140900 121120 141100 121380
rect 141400 121120 141600 121380
rect 141900 121120 142000 121380
rect 118000 121100 118120 121120
rect 118380 121100 118620 121120
rect 118880 121100 119120 121120
rect 119380 121100 119620 121120
rect 119880 121100 120120 121120
rect 120380 121100 120620 121120
rect 120880 121100 121120 121120
rect 121380 121100 121620 121120
rect 121880 121100 122120 121120
rect 122380 121100 122620 121120
rect 122880 121100 123120 121120
rect 123380 121100 123620 121120
rect 123880 121100 124120 121120
rect 124380 121100 124620 121120
rect 124880 121100 125120 121120
rect 125380 121100 125620 121120
rect 125880 121100 126120 121120
rect 126380 121100 126620 121120
rect 126880 121100 127120 121120
rect 127380 121100 127620 121120
rect 127880 121100 128120 121120
rect 128380 121100 128620 121120
rect 128880 121100 129120 121120
rect 129380 121100 129620 121120
rect 129880 121100 130120 121120
rect 130380 121100 130620 121120
rect 130880 121100 131120 121120
rect 131380 121100 131620 121120
rect 131880 121100 132120 121120
rect 132380 121100 132620 121120
rect 132880 121100 133120 121120
rect 133380 121100 133620 121120
rect 133880 121100 134120 121120
rect 134380 121100 134620 121120
rect 134880 121100 135120 121120
rect 135380 121100 135620 121120
rect 135880 121100 136120 121120
rect 136380 121100 136620 121120
rect 136880 121100 137120 121120
rect 137380 121100 137620 121120
rect 137880 121100 138120 121120
rect 138380 121100 138620 121120
rect 138880 121100 139120 121120
rect 139380 121100 139620 121120
rect 139880 121100 140120 121120
rect 140380 121100 140620 121120
rect 140880 121100 141120 121120
rect 141380 121100 141620 121120
rect 141880 121100 142000 121120
rect 118000 120900 142000 121100
rect 118000 120880 118120 120900
rect 118380 120880 118620 120900
rect 118880 120880 119120 120900
rect 119380 120880 119620 120900
rect 119880 120880 120120 120900
rect 120380 120880 120620 120900
rect 120880 120880 121120 120900
rect 121380 120880 121620 120900
rect 121880 120880 122120 120900
rect 122380 120880 122620 120900
rect 122880 120880 123120 120900
rect 123380 120880 123620 120900
rect 123880 120880 124120 120900
rect 124380 120880 124620 120900
rect 124880 120880 125120 120900
rect 125380 120880 125620 120900
rect 125880 120880 126120 120900
rect 126380 120880 126620 120900
rect 126880 120880 127120 120900
rect 127380 120880 127620 120900
rect 127880 120880 128120 120900
rect 128380 120880 128620 120900
rect 128880 120880 129120 120900
rect 129380 120880 129620 120900
rect 129880 120880 130120 120900
rect 130380 120880 130620 120900
rect 130880 120880 131120 120900
rect 131380 120880 131620 120900
rect 131880 120880 132120 120900
rect 132380 120880 132620 120900
rect 132880 120880 133120 120900
rect 133380 120880 133620 120900
rect 133880 120880 134120 120900
rect 134380 120880 134620 120900
rect 134880 120880 135120 120900
rect 135380 120880 135620 120900
rect 135880 120880 136120 120900
rect 136380 120880 136620 120900
rect 136880 120880 137120 120900
rect 137380 120880 137620 120900
rect 137880 120880 138120 120900
rect 138380 120880 138620 120900
rect 138880 120880 139120 120900
rect 139380 120880 139620 120900
rect 139880 120880 140120 120900
rect 140380 120880 140620 120900
rect 140880 120880 141120 120900
rect 141380 120880 141620 120900
rect 141880 120880 142000 120900
rect 118000 120620 118100 120880
rect 118400 120620 118600 120880
rect 118900 120620 119100 120880
rect 119400 120620 119600 120880
rect 119900 120620 120100 120880
rect 120400 120620 120600 120880
rect 120900 120620 121100 120880
rect 121400 120620 121600 120880
rect 121900 120620 122100 120880
rect 122400 120620 122600 120880
rect 122900 120620 123100 120880
rect 123400 120620 123600 120880
rect 123900 120620 124100 120880
rect 124400 120620 124600 120880
rect 124900 120620 125100 120880
rect 125400 120620 125600 120880
rect 125900 120620 126100 120880
rect 126400 120620 126600 120880
rect 126900 120620 127100 120880
rect 127400 120620 127600 120880
rect 127900 120620 128100 120880
rect 128400 120620 128600 120880
rect 128900 120620 129100 120880
rect 129400 120620 129600 120880
rect 129900 120620 130100 120880
rect 130400 120620 130600 120880
rect 130900 120620 131100 120880
rect 131400 120620 131600 120880
rect 131900 120620 132100 120880
rect 132400 120620 132600 120880
rect 132900 120620 133100 120880
rect 133400 120620 133600 120880
rect 133900 120620 134100 120880
rect 134400 120620 134600 120880
rect 134900 120620 135100 120880
rect 135400 120620 135600 120880
rect 135900 120620 136100 120880
rect 136400 120620 136600 120880
rect 136900 120620 137100 120880
rect 137400 120620 137600 120880
rect 137900 120620 138100 120880
rect 138400 120620 138600 120880
rect 138900 120620 139100 120880
rect 139400 120620 139600 120880
rect 139900 120620 140100 120880
rect 140400 120620 140600 120880
rect 140900 120620 141100 120880
rect 141400 120620 141600 120880
rect 141900 120620 142000 120880
rect 118000 120600 118120 120620
rect 118380 120600 118620 120620
rect 118880 120600 119120 120620
rect 119380 120600 119620 120620
rect 119880 120600 120120 120620
rect 120380 120600 120620 120620
rect 120880 120600 121120 120620
rect 121380 120600 121620 120620
rect 121880 120600 122120 120620
rect 122380 120600 122620 120620
rect 122880 120600 123120 120620
rect 123380 120600 123620 120620
rect 123880 120600 124120 120620
rect 124380 120600 124620 120620
rect 124880 120600 125120 120620
rect 125380 120600 125620 120620
rect 125880 120600 126120 120620
rect 126380 120600 126620 120620
rect 126880 120600 127120 120620
rect 127380 120600 127620 120620
rect 127880 120600 128120 120620
rect 128380 120600 128620 120620
rect 128880 120600 129120 120620
rect 129380 120600 129620 120620
rect 129880 120600 130120 120620
rect 130380 120600 130620 120620
rect 130880 120600 131120 120620
rect 131380 120600 131620 120620
rect 131880 120600 132120 120620
rect 132380 120600 132620 120620
rect 132880 120600 133120 120620
rect 133380 120600 133620 120620
rect 133880 120600 134120 120620
rect 134380 120600 134620 120620
rect 134880 120600 135120 120620
rect 135380 120600 135620 120620
rect 135880 120600 136120 120620
rect 136380 120600 136620 120620
rect 136880 120600 137120 120620
rect 137380 120600 137620 120620
rect 137880 120600 138120 120620
rect 138380 120600 138620 120620
rect 138880 120600 139120 120620
rect 139380 120600 139620 120620
rect 139880 120600 140120 120620
rect 140380 120600 140620 120620
rect 140880 120600 141120 120620
rect 141380 120600 141620 120620
rect 141880 120600 142000 120620
rect 118000 120400 142000 120600
rect 118000 120380 118120 120400
rect 118380 120380 118620 120400
rect 118880 120380 119120 120400
rect 119380 120380 119620 120400
rect 119880 120380 120120 120400
rect 120380 120380 120620 120400
rect 120880 120380 121120 120400
rect 121380 120380 121620 120400
rect 121880 120380 122120 120400
rect 122380 120380 122620 120400
rect 122880 120380 123120 120400
rect 123380 120380 123620 120400
rect 123880 120380 124120 120400
rect 124380 120380 124620 120400
rect 124880 120380 125120 120400
rect 125380 120380 125620 120400
rect 125880 120380 126120 120400
rect 126380 120380 126620 120400
rect 126880 120380 127120 120400
rect 127380 120380 127620 120400
rect 127880 120380 128120 120400
rect 128380 120380 128620 120400
rect 128880 120380 129120 120400
rect 129380 120380 129620 120400
rect 129880 120380 130120 120400
rect 130380 120380 130620 120400
rect 130880 120380 131120 120400
rect 131380 120380 131620 120400
rect 131880 120380 132120 120400
rect 132380 120380 132620 120400
rect 132880 120380 133120 120400
rect 133380 120380 133620 120400
rect 133880 120380 134120 120400
rect 134380 120380 134620 120400
rect 134880 120380 135120 120400
rect 135380 120380 135620 120400
rect 135880 120380 136120 120400
rect 136380 120380 136620 120400
rect 136880 120380 137120 120400
rect 137380 120380 137620 120400
rect 137880 120380 138120 120400
rect 138380 120380 138620 120400
rect 138880 120380 139120 120400
rect 139380 120380 139620 120400
rect 139880 120380 140120 120400
rect 140380 120380 140620 120400
rect 140880 120380 141120 120400
rect 141380 120380 141620 120400
rect 141880 120380 142000 120400
rect 118000 120120 118100 120380
rect 118400 120120 118600 120380
rect 118900 120120 119100 120380
rect 119400 120120 119600 120380
rect 119900 120120 120100 120380
rect 120400 120120 120600 120380
rect 120900 120120 121100 120380
rect 121400 120120 121600 120380
rect 121900 120120 122100 120380
rect 122400 120120 122600 120380
rect 122900 120120 123100 120380
rect 123400 120120 123600 120380
rect 123900 120120 124100 120380
rect 124400 120120 124600 120380
rect 124900 120120 125100 120380
rect 125400 120120 125600 120380
rect 125900 120120 126100 120380
rect 126400 120120 126600 120380
rect 126900 120120 127100 120380
rect 127400 120120 127600 120380
rect 127900 120120 128100 120380
rect 128400 120120 128600 120380
rect 128900 120120 129100 120380
rect 129400 120120 129600 120380
rect 129900 120120 130100 120380
rect 130400 120120 130600 120380
rect 130900 120120 131100 120380
rect 131400 120120 131600 120380
rect 131900 120120 132100 120380
rect 132400 120120 132600 120380
rect 132900 120120 133100 120380
rect 133400 120120 133600 120380
rect 133900 120120 134100 120380
rect 134400 120120 134600 120380
rect 134900 120120 135100 120380
rect 135400 120120 135600 120380
rect 135900 120120 136100 120380
rect 136400 120120 136600 120380
rect 136900 120120 137100 120380
rect 137400 120120 137600 120380
rect 137900 120120 138100 120380
rect 138400 120120 138600 120380
rect 138900 120120 139100 120380
rect 139400 120120 139600 120380
rect 139900 120120 140100 120380
rect 140400 120120 140600 120380
rect 140900 120120 141100 120380
rect 141400 120120 141600 120380
rect 141900 120120 142000 120380
rect 118000 120100 118120 120120
rect 118380 120100 118620 120120
rect 118880 120100 119120 120120
rect 119380 120100 119620 120120
rect 119880 120100 120120 120120
rect 120380 120100 120620 120120
rect 120880 120100 121120 120120
rect 121380 120100 121620 120120
rect 121880 120100 122120 120120
rect 122380 120100 122620 120120
rect 122880 120100 123120 120120
rect 123380 120100 123620 120120
rect 123880 120100 124120 120120
rect 124380 120100 124620 120120
rect 124880 120100 125120 120120
rect 125380 120100 125620 120120
rect 125880 120100 126120 120120
rect 126380 120100 126620 120120
rect 126880 120100 127120 120120
rect 127380 120100 127620 120120
rect 127880 120100 128120 120120
rect 128380 120100 128620 120120
rect 128880 120100 129120 120120
rect 129380 120100 129620 120120
rect 129880 120100 130120 120120
rect 130380 120100 130620 120120
rect 130880 120100 131120 120120
rect 131380 120100 131620 120120
rect 131880 120100 132120 120120
rect 132380 120100 132620 120120
rect 132880 120100 133120 120120
rect 133380 120100 133620 120120
rect 133880 120100 134120 120120
rect 134380 120100 134620 120120
rect 134880 120100 135120 120120
rect 135380 120100 135620 120120
rect 135880 120100 136120 120120
rect 136380 120100 136620 120120
rect 136880 120100 137120 120120
rect 137380 120100 137620 120120
rect 137880 120100 138120 120120
rect 138380 120100 138620 120120
rect 138880 120100 139120 120120
rect 139380 120100 139620 120120
rect 139880 120100 140120 120120
rect 140380 120100 140620 120120
rect 140880 120100 141120 120120
rect 141380 120100 141620 120120
rect 141880 120100 142000 120120
rect 118000 119900 142000 120100
rect 118000 119880 118120 119900
rect 118380 119880 118620 119900
rect 118880 119880 119120 119900
rect 119380 119880 119620 119900
rect 119880 119880 120120 119900
rect 120380 119880 120620 119900
rect 120880 119880 121120 119900
rect 121380 119880 121620 119900
rect 121880 119880 122120 119900
rect 122380 119880 122620 119900
rect 122880 119880 123120 119900
rect 123380 119880 123620 119900
rect 123880 119880 124120 119900
rect 124380 119880 124620 119900
rect 124880 119880 125120 119900
rect 125380 119880 125620 119900
rect 125880 119880 126120 119900
rect 126380 119880 126620 119900
rect 126880 119880 127120 119900
rect 127380 119880 127620 119900
rect 127880 119880 128120 119900
rect 128380 119880 128620 119900
rect 128880 119880 129120 119900
rect 129380 119880 129620 119900
rect 129880 119880 130120 119900
rect 130380 119880 130620 119900
rect 130880 119880 131120 119900
rect 131380 119880 131620 119900
rect 131880 119880 132120 119900
rect 132380 119880 132620 119900
rect 132880 119880 133120 119900
rect 133380 119880 133620 119900
rect 133880 119880 134120 119900
rect 134380 119880 134620 119900
rect 134880 119880 135120 119900
rect 135380 119880 135620 119900
rect 135880 119880 136120 119900
rect 136380 119880 136620 119900
rect 136880 119880 137120 119900
rect 137380 119880 137620 119900
rect 137880 119880 138120 119900
rect 138380 119880 138620 119900
rect 138880 119880 139120 119900
rect 139380 119880 139620 119900
rect 139880 119880 140120 119900
rect 140380 119880 140620 119900
rect 140880 119880 141120 119900
rect 141380 119880 141620 119900
rect 141880 119880 142000 119900
rect 118000 119620 118100 119880
rect 118400 119620 118600 119880
rect 118900 119620 119100 119880
rect 119400 119620 119600 119880
rect 119900 119620 120100 119880
rect 120400 119620 120600 119880
rect 120900 119620 121100 119880
rect 121400 119620 121600 119880
rect 121900 119620 122100 119880
rect 122400 119620 122600 119880
rect 122900 119620 123100 119880
rect 123400 119620 123600 119880
rect 123900 119620 124100 119880
rect 124400 119620 124600 119880
rect 124900 119620 125100 119880
rect 125400 119620 125600 119880
rect 125900 119620 126100 119880
rect 126400 119620 126600 119880
rect 126900 119620 127100 119880
rect 127400 119620 127600 119880
rect 127900 119620 128100 119880
rect 128400 119620 128600 119880
rect 128900 119620 129100 119880
rect 129400 119620 129600 119880
rect 129900 119620 130100 119880
rect 130400 119620 130600 119880
rect 130900 119620 131100 119880
rect 131400 119620 131600 119880
rect 131900 119620 132100 119880
rect 132400 119620 132600 119880
rect 132900 119620 133100 119880
rect 133400 119620 133600 119880
rect 133900 119620 134100 119880
rect 134400 119620 134600 119880
rect 134900 119620 135100 119880
rect 135400 119620 135600 119880
rect 135900 119620 136100 119880
rect 136400 119620 136600 119880
rect 136900 119620 137100 119880
rect 137400 119620 137600 119880
rect 137900 119620 138100 119880
rect 138400 119620 138600 119880
rect 138900 119620 139100 119880
rect 139400 119620 139600 119880
rect 139900 119620 140100 119880
rect 140400 119620 140600 119880
rect 140900 119620 141100 119880
rect 141400 119620 141600 119880
rect 141900 119620 142000 119880
rect 118000 119600 118120 119620
rect 118380 119600 118620 119620
rect 118880 119600 119120 119620
rect 119380 119600 119620 119620
rect 119880 119600 120120 119620
rect 120380 119600 120620 119620
rect 120880 119600 121120 119620
rect 121380 119600 121620 119620
rect 121880 119600 122120 119620
rect 122380 119600 122620 119620
rect 122880 119600 123120 119620
rect 123380 119600 123620 119620
rect 123880 119600 124120 119620
rect 124380 119600 124620 119620
rect 124880 119600 125120 119620
rect 125380 119600 125620 119620
rect 125880 119600 126120 119620
rect 126380 119600 126620 119620
rect 126880 119600 127120 119620
rect 127380 119600 127620 119620
rect 127880 119600 128120 119620
rect 128380 119600 128620 119620
rect 128880 119600 129120 119620
rect 129380 119600 129620 119620
rect 129880 119600 130120 119620
rect 130380 119600 130620 119620
rect 130880 119600 131120 119620
rect 131380 119600 131620 119620
rect 131880 119600 132120 119620
rect 132380 119600 132620 119620
rect 132880 119600 133120 119620
rect 133380 119600 133620 119620
rect 133880 119600 134120 119620
rect 134380 119600 134620 119620
rect 134880 119600 135120 119620
rect 135380 119600 135620 119620
rect 135880 119600 136120 119620
rect 136380 119600 136620 119620
rect 136880 119600 137120 119620
rect 137380 119600 137620 119620
rect 137880 119600 138120 119620
rect 138380 119600 138620 119620
rect 138880 119600 139120 119620
rect 139380 119600 139620 119620
rect 139880 119600 140120 119620
rect 140380 119600 140620 119620
rect 140880 119600 141120 119620
rect 141380 119600 141620 119620
rect 141880 119600 142000 119620
rect 118000 119400 142000 119600
rect 118000 119380 118120 119400
rect 118380 119380 118620 119400
rect 118880 119380 119120 119400
rect 119380 119380 119620 119400
rect 119880 119380 120120 119400
rect 120380 119380 120620 119400
rect 120880 119380 121120 119400
rect 121380 119380 121620 119400
rect 121880 119380 122120 119400
rect 122380 119380 122620 119400
rect 122880 119380 123120 119400
rect 123380 119380 123620 119400
rect 123880 119380 124120 119400
rect 124380 119380 124620 119400
rect 124880 119380 125120 119400
rect 125380 119380 125620 119400
rect 125880 119380 126120 119400
rect 126380 119380 126620 119400
rect 126880 119380 127120 119400
rect 127380 119380 127620 119400
rect 127880 119380 128120 119400
rect 128380 119380 128620 119400
rect 128880 119380 129120 119400
rect 129380 119380 129620 119400
rect 129880 119380 130120 119400
rect 130380 119380 130620 119400
rect 130880 119380 131120 119400
rect 131380 119380 131620 119400
rect 131880 119380 132120 119400
rect 132380 119380 132620 119400
rect 132880 119380 133120 119400
rect 133380 119380 133620 119400
rect 133880 119380 134120 119400
rect 134380 119380 134620 119400
rect 134880 119380 135120 119400
rect 135380 119380 135620 119400
rect 135880 119380 136120 119400
rect 136380 119380 136620 119400
rect 136880 119380 137120 119400
rect 137380 119380 137620 119400
rect 137880 119380 138120 119400
rect 138380 119380 138620 119400
rect 138880 119380 139120 119400
rect 139380 119380 139620 119400
rect 139880 119380 140120 119400
rect 140380 119380 140620 119400
rect 140880 119380 141120 119400
rect 141380 119380 141620 119400
rect 141880 119380 142000 119400
rect 118000 119120 118100 119380
rect 118400 119120 118600 119380
rect 118900 119120 119100 119380
rect 119400 119120 119600 119380
rect 119900 119120 120100 119380
rect 120400 119120 120600 119380
rect 120900 119120 121100 119380
rect 121400 119120 121600 119380
rect 121900 119120 122100 119380
rect 122400 119120 122600 119380
rect 122900 119120 123100 119380
rect 123400 119120 123600 119380
rect 123900 119120 124100 119380
rect 124400 119120 124600 119380
rect 124900 119120 125100 119380
rect 125400 119120 125600 119380
rect 125900 119120 126100 119380
rect 126400 119120 126600 119380
rect 126900 119120 127100 119380
rect 127400 119120 127600 119380
rect 127900 119120 128100 119380
rect 128400 119120 128600 119380
rect 128900 119120 129100 119380
rect 129400 119120 129600 119380
rect 129900 119120 130100 119380
rect 130400 119120 130600 119380
rect 130900 119120 131100 119380
rect 131400 119120 131600 119380
rect 131900 119120 132100 119380
rect 132400 119120 132600 119380
rect 132900 119120 133100 119380
rect 133400 119120 133600 119380
rect 133900 119120 134100 119380
rect 134400 119120 134600 119380
rect 134900 119120 135100 119380
rect 135400 119120 135600 119380
rect 135900 119120 136100 119380
rect 136400 119120 136600 119380
rect 136900 119120 137100 119380
rect 137400 119120 137600 119380
rect 137900 119120 138100 119380
rect 138400 119120 138600 119380
rect 138900 119120 139100 119380
rect 139400 119120 139600 119380
rect 139900 119120 140100 119380
rect 140400 119120 140600 119380
rect 140900 119120 141100 119380
rect 141400 119120 141600 119380
rect 141900 119120 142000 119380
rect 118000 119100 118120 119120
rect 118380 119100 118620 119120
rect 118880 119100 119120 119120
rect 119380 119100 119620 119120
rect 119880 119100 120120 119120
rect 120380 119100 120620 119120
rect 120880 119100 121120 119120
rect 121380 119100 121620 119120
rect 121880 119100 122120 119120
rect 122380 119100 122620 119120
rect 122880 119100 123120 119120
rect 123380 119100 123620 119120
rect 123880 119100 124120 119120
rect 124380 119100 124620 119120
rect 124880 119100 125120 119120
rect 125380 119100 125620 119120
rect 125880 119100 126120 119120
rect 126380 119100 126620 119120
rect 126880 119100 127120 119120
rect 127380 119100 127620 119120
rect 127880 119100 128120 119120
rect 128380 119100 128620 119120
rect 128880 119100 129120 119120
rect 129380 119100 129620 119120
rect 129880 119100 130120 119120
rect 130380 119100 130620 119120
rect 130880 119100 131120 119120
rect 131380 119100 131620 119120
rect 131880 119100 132120 119120
rect 132380 119100 132620 119120
rect 132880 119100 133120 119120
rect 133380 119100 133620 119120
rect 133880 119100 134120 119120
rect 134380 119100 134620 119120
rect 134880 119100 135120 119120
rect 135380 119100 135620 119120
rect 135880 119100 136120 119120
rect 136380 119100 136620 119120
rect 136880 119100 137120 119120
rect 137380 119100 137620 119120
rect 137880 119100 138120 119120
rect 138380 119100 138620 119120
rect 138880 119100 139120 119120
rect 139380 119100 139620 119120
rect 139880 119100 140120 119120
rect 140380 119100 140620 119120
rect 140880 119100 141120 119120
rect 141380 119100 141620 119120
rect 141880 119100 142000 119120
rect 118000 118900 142000 119100
rect 118000 118880 118120 118900
rect 118380 118880 118620 118900
rect 118880 118880 119120 118900
rect 119380 118880 119620 118900
rect 119880 118880 120120 118900
rect 120380 118880 120620 118900
rect 120880 118880 121120 118900
rect 121380 118880 121620 118900
rect 121880 118880 122120 118900
rect 122380 118880 122620 118900
rect 122880 118880 123120 118900
rect 123380 118880 123620 118900
rect 123880 118880 124120 118900
rect 124380 118880 124620 118900
rect 124880 118880 125120 118900
rect 125380 118880 125620 118900
rect 125880 118880 126120 118900
rect 126380 118880 126620 118900
rect 126880 118880 127120 118900
rect 127380 118880 127620 118900
rect 127880 118880 128120 118900
rect 128380 118880 128620 118900
rect 128880 118880 129120 118900
rect 129380 118880 129620 118900
rect 129880 118880 130120 118900
rect 130380 118880 130620 118900
rect 130880 118880 131120 118900
rect 131380 118880 131620 118900
rect 131880 118880 132120 118900
rect 132380 118880 132620 118900
rect 132880 118880 133120 118900
rect 133380 118880 133620 118900
rect 133880 118880 134120 118900
rect 134380 118880 134620 118900
rect 134880 118880 135120 118900
rect 135380 118880 135620 118900
rect 135880 118880 136120 118900
rect 136380 118880 136620 118900
rect 136880 118880 137120 118900
rect 137380 118880 137620 118900
rect 137880 118880 138120 118900
rect 138380 118880 138620 118900
rect 138880 118880 139120 118900
rect 139380 118880 139620 118900
rect 139880 118880 140120 118900
rect 140380 118880 140620 118900
rect 140880 118880 141120 118900
rect 141380 118880 141620 118900
rect 141880 118880 142000 118900
rect 118000 118620 118100 118880
rect 118400 118620 118600 118880
rect 118900 118620 119100 118880
rect 119400 118620 119600 118880
rect 119900 118620 120100 118880
rect 120400 118620 120600 118880
rect 120900 118620 121100 118880
rect 121400 118620 121600 118880
rect 121900 118620 122100 118880
rect 122400 118620 122600 118880
rect 122900 118620 123100 118880
rect 123400 118620 123600 118880
rect 123900 118620 124100 118880
rect 124400 118620 124600 118880
rect 124900 118620 125100 118880
rect 125400 118620 125600 118880
rect 125900 118620 126100 118880
rect 126400 118620 126600 118880
rect 126900 118620 127100 118880
rect 127400 118620 127600 118880
rect 127900 118620 128100 118880
rect 128400 118620 128600 118880
rect 128900 118620 129100 118880
rect 129400 118620 129600 118880
rect 129900 118620 130100 118880
rect 130400 118620 130600 118880
rect 130900 118620 131100 118880
rect 131400 118620 131600 118880
rect 131900 118620 132100 118880
rect 132400 118620 132600 118880
rect 132900 118620 133100 118880
rect 133400 118620 133600 118880
rect 133900 118620 134100 118880
rect 134400 118620 134600 118880
rect 134900 118620 135100 118880
rect 135400 118620 135600 118880
rect 135900 118620 136100 118880
rect 136400 118620 136600 118880
rect 136900 118620 137100 118880
rect 137400 118620 137600 118880
rect 137900 118620 138100 118880
rect 138400 118620 138600 118880
rect 138900 118620 139100 118880
rect 139400 118620 139600 118880
rect 139900 118620 140100 118880
rect 140400 118620 140600 118880
rect 140900 118620 141100 118880
rect 141400 118620 141600 118880
rect 141900 118620 142000 118880
rect 118000 118600 118120 118620
rect 118380 118600 118620 118620
rect 118880 118600 119120 118620
rect 119380 118600 119620 118620
rect 119880 118600 120120 118620
rect 120380 118600 120620 118620
rect 120880 118600 121120 118620
rect 121380 118600 121620 118620
rect 121880 118600 122120 118620
rect 122380 118600 122620 118620
rect 122880 118600 123120 118620
rect 123380 118600 123620 118620
rect 123880 118600 124120 118620
rect 124380 118600 124620 118620
rect 124880 118600 125120 118620
rect 125380 118600 125620 118620
rect 125880 118600 126120 118620
rect 126380 118600 126620 118620
rect 126880 118600 127120 118620
rect 127380 118600 127620 118620
rect 127880 118600 128120 118620
rect 128380 118600 128620 118620
rect 128880 118600 129120 118620
rect 129380 118600 129620 118620
rect 129880 118600 130120 118620
rect 130380 118600 130620 118620
rect 130880 118600 131120 118620
rect 131380 118600 131620 118620
rect 131880 118600 132120 118620
rect 132380 118600 132620 118620
rect 132880 118600 133120 118620
rect 133380 118600 133620 118620
rect 133880 118600 134120 118620
rect 134380 118600 134620 118620
rect 134880 118600 135120 118620
rect 135380 118600 135620 118620
rect 135880 118600 136120 118620
rect 136380 118600 136620 118620
rect 136880 118600 137120 118620
rect 137380 118600 137620 118620
rect 137880 118600 138120 118620
rect 138380 118600 138620 118620
rect 138880 118600 139120 118620
rect 139380 118600 139620 118620
rect 139880 118600 140120 118620
rect 140380 118600 140620 118620
rect 140880 118600 141120 118620
rect 141380 118600 141620 118620
rect 141880 118600 142000 118620
rect 118000 118400 142000 118600
rect 118000 118380 118120 118400
rect 118380 118380 118620 118400
rect 118880 118380 119120 118400
rect 119380 118380 119620 118400
rect 119880 118380 120120 118400
rect 120380 118380 120620 118400
rect 120880 118380 121120 118400
rect 121380 118380 121620 118400
rect 121880 118380 122120 118400
rect 122380 118380 122620 118400
rect 122880 118380 123120 118400
rect 123380 118380 123620 118400
rect 123880 118380 124120 118400
rect 124380 118380 124620 118400
rect 124880 118380 125120 118400
rect 125380 118380 125620 118400
rect 125880 118380 126120 118400
rect 126380 118380 126620 118400
rect 126880 118380 127120 118400
rect 127380 118380 127620 118400
rect 127880 118380 128120 118400
rect 128380 118380 128620 118400
rect 128880 118380 129120 118400
rect 129380 118380 129620 118400
rect 129880 118380 130120 118400
rect 130380 118380 130620 118400
rect 130880 118380 131120 118400
rect 131380 118380 131620 118400
rect 131880 118380 132120 118400
rect 132380 118380 132620 118400
rect 132880 118380 133120 118400
rect 133380 118380 133620 118400
rect 133880 118380 134120 118400
rect 134380 118380 134620 118400
rect 134880 118380 135120 118400
rect 135380 118380 135620 118400
rect 135880 118380 136120 118400
rect 136380 118380 136620 118400
rect 136880 118380 137120 118400
rect 137380 118380 137620 118400
rect 137880 118380 138120 118400
rect 138380 118380 138620 118400
rect 138880 118380 139120 118400
rect 139380 118380 139620 118400
rect 139880 118380 140120 118400
rect 140380 118380 140620 118400
rect 140880 118380 141120 118400
rect 141380 118380 141620 118400
rect 141880 118380 142000 118400
rect 118000 118120 118100 118380
rect 118400 118120 118600 118380
rect 118900 118120 119100 118380
rect 119400 118120 119600 118380
rect 119900 118120 120100 118380
rect 120400 118120 120600 118380
rect 120900 118120 121100 118380
rect 121400 118120 121600 118380
rect 121900 118120 122100 118380
rect 122400 118120 122600 118380
rect 122900 118120 123100 118380
rect 123400 118120 123600 118380
rect 123900 118120 124100 118380
rect 124400 118120 124600 118380
rect 124900 118120 125100 118380
rect 125400 118120 125600 118380
rect 125900 118120 126100 118380
rect 126400 118120 126600 118380
rect 126900 118120 127100 118380
rect 127400 118120 127600 118380
rect 127900 118120 128100 118380
rect 128400 118120 128600 118380
rect 128900 118120 129100 118380
rect 129400 118120 129600 118380
rect 129900 118120 130100 118380
rect 130400 118120 130600 118380
rect 130900 118120 131100 118380
rect 131400 118120 131600 118380
rect 131900 118120 132100 118380
rect 132400 118120 132600 118380
rect 132900 118120 133100 118380
rect 133400 118120 133600 118380
rect 133900 118120 134100 118380
rect 134400 118120 134600 118380
rect 134900 118120 135100 118380
rect 135400 118120 135600 118380
rect 135900 118120 136100 118380
rect 136400 118120 136600 118380
rect 136900 118120 137100 118380
rect 137400 118120 137600 118380
rect 137900 118120 138100 118380
rect 138400 118120 138600 118380
rect 138900 118120 139100 118380
rect 139400 118120 139600 118380
rect 139900 118120 140100 118380
rect 140400 118120 140600 118380
rect 140900 118120 141100 118380
rect 141400 118120 141600 118380
rect 141900 118120 142000 118380
rect 118000 118100 118120 118120
rect 118380 118100 118620 118120
rect 118880 118100 119120 118120
rect 119380 118100 119620 118120
rect 119880 118100 120120 118120
rect 120380 118100 120620 118120
rect 120880 118100 121120 118120
rect 121380 118100 121620 118120
rect 121880 118100 122120 118120
rect 122380 118100 122620 118120
rect 122880 118100 123120 118120
rect 123380 118100 123620 118120
rect 123880 118100 124120 118120
rect 124380 118100 124620 118120
rect 124880 118100 125120 118120
rect 125380 118100 125620 118120
rect 125880 118100 126120 118120
rect 126380 118100 126620 118120
rect 126880 118100 127120 118120
rect 127380 118100 127620 118120
rect 127880 118100 128120 118120
rect 128380 118100 128620 118120
rect 128880 118100 129120 118120
rect 129380 118100 129620 118120
rect 129880 118100 130120 118120
rect 130380 118100 130620 118120
rect 130880 118100 131120 118120
rect 131380 118100 131620 118120
rect 131880 118100 132120 118120
rect 132380 118100 132620 118120
rect 132880 118100 133120 118120
rect 133380 118100 133620 118120
rect 133880 118100 134120 118120
rect 134380 118100 134620 118120
rect 134880 118100 135120 118120
rect 135380 118100 135620 118120
rect 135880 118100 136120 118120
rect 136380 118100 136620 118120
rect 136880 118100 137120 118120
rect 137380 118100 137620 118120
rect 137880 118100 138120 118120
rect 138380 118100 138620 118120
rect 138880 118100 139120 118120
rect 139380 118100 139620 118120
rect 139880 118100 140120 118120
rect 140380 118100 140620 118120
rect 140880 118100 141120 118120
rect 141380 118100 141620 118120
rect 141880 118100 142000 118120
rect 118000 117900 142000 118100
rect 118000 117880 118120 117900
rect 118380 117880 118620 117900
rect 118880 117880 119120 117900
rect 119380 117880 119620 117900
rect 119880 117880 120120 117900
rect 120380 117880 120620 117900
rect 120880 117880 121120 117900
rect 121380 117880 121620 117900
rect 121880 117880 122120 117900
rect 122380 117880 122620 117900
rect 122880 117880 123120 117900
rect 123380 117880 123620 117900
rect 123880 117880 124120 117900
rect 124380 117880 124620 117900
rect 124880 117880 125120 117900
rect 125380 117880 125620 117900
rect 125880 117880 126120 117900
rect 126380 117880 126620 117900
rect 126880 117880 127120 117900
rect 127380 117880 127620 117900
rect 127880 117880 128120 117900
rect 128380 117880 128620 117900
rect 128880 117880 129120 117900
rect 129380 117880 129620 117900
rect 129880 117880 130120 117900
rect 130380 117880 130620 117900
rect 130880 117880 131120 117900
rect 131380 117880 131620 117900
rect 131880 117880 132120 117900
rect 132380 117880 132620 117900
rect 132880 117880 133120 117900
rect 133380 117880 133620 117900
rect 133880 117880 134120 117900
rect 134380 117880 134620 117900
rect 134880 117880 135120 117900
rect 135380 117880 135620 117900
rect 135880 117880 136120 117900
rect 136380 117880 136620 117900
rect 136880 117880 137120 117900
rect 137380 117880 137620 117900
rect 137880 117880 138120 117900
rect 138380 117880 138620 117900
rect 138880 117880 139120 117900
rect 139380 117880 139620 117900
rect 139880 117880 140120 117900
rect 140380 117880 140620 117900
rect 140880 117880 141120 117900
rect 141380 117880 141620 117900
rect 141880 117880 142000 117900
rect 118000 117620 118100 117880
rect 118400 117620 118600 117880
rect 118900 117620 119100 117880
rect 119400 117620 119600 117880
rect 119900 117620 120100 117880
rect 120400 117620 120600 117880
rect 120900 117620 121100 117880
rect 121400 117620 121600 117880
rect 121900 117620 122100 117880
rect 122400 117620 122600 117880
rect 122900 117620 123100 117880
rect 123400 117620 123600 117880
rect 123900 117620 124100 117880
rect 124400 117620 124600 117880
rect 124900 117620 125100 117880
rect 125400 117620 125600 117880
rect 125900 117620 126100 117880
rect 126400 117620 126600 117880
rect 126900 117620 127100 117880
rect 127400 117620 127600 117880
rect 127900 117620 128100 117880
rect 128400 117620 128600 117880
rect 128900 117620 129100 117880
rect 129400 117620 129600 117880
rect 129900 117620 130100 117880
rect 130400 117620 130600 117880
rect 130900 117620 131100 117880
rect 131400 117620 131600 117880
rect 131900 117620 132100 117880
rect 132400 117620 132600 117880
rect 132900 117620 133100 117880
rect 133400 117620 133600 117880
rect 133900 117620 134100 117880
rect 134400 117620 134600 117880
rect 134900 117620 135100 117880
rect 135400 117620 135600 117880
rect 135900 117620 136100 117880
rect 136400 117620 136600 117880
rect 136900 117620 137100 117880
rect 137400 117620 137600 117880
rect 137900 117620 138100 117880
rect 138400 117620 138600 117880
rect 138900 117620 139100 117880
rect 139400 117620 139600 117880
rect 139900 117620 140100 117880
rect 140400 117620 140600 117880
rect 140900 117620 141100 117880
rect 141400 117620 141600 117880
rect 141900 117620 142000 117880
rect 118000 117600 118120 117620
rect 118380 117600 118620 117620
rect 118880 117600 119120 117620
rect 119380 117600 119620 117620
rect 119880 117600 120120 117620
rect 120380 117600 120620 117620
rect 120880 117600 121120 117620
rect 121380 117600 121620 117620
rect 121880 117600 122120 117620
rect 122380 117600 122620 117620
rect 122880 117600 123120 117620
rect 123380 117600 123620 117620
rect 123880 117600 124120 117620
rect 124380 117600 124620 117620
rect 124880 117600 125120 117620
rect 125380 117600 125620 117620
rect 125880 117600 126120 117620
rect 126380 117600 126620 117620
rect 126880 117600 127120 117620
rect 127380 117600 127620 117620
rect 127880 117600 128120 117620
rect 128380 117600 128620 117620
rect 128880 117600 129120 117620
rect 129380 117600 129620 117620
rect 129880 117600 130120 117620
rect 130380 117600 130620 117620
rect 130880 117600 131120 117620
rect 131380 117600 131620 117620
rect 131880 117600 132120 117620
rect 132380 117600 132620 117620
rect 132880 117600 133120 117620
rect 133380 117600 133620 117620
rect 133880 117600 134120 117620
rect 134380 117600 134620 117620
rect 134880 117600 135120 117620
rect 135380 117600 135620 117620
rect 135880 117600 136120 117620
rect 136380 117600 136620 117620
rect 136880 117600 137120 117620
rect 137380 117600 137620 117620
rect 137880 117600 138120 117620
rect 138380 117600 138620 117620
rect 138880 117600 139120 117620
rect 139380 117600 139620 117620
rect 139880 117600 140120 117620
rect 140380 117600 140620 117620
rect 140880 117600 141120 117620
rect 141380 117600 141620 117620
rect 141880 117600 142000 117620
rect 118000 117400 142000 117600
rect 118000 117380 118120 117400
rect 118380 117380 118620 117400
rect 118880 117380 119120 117400
rect 119380 117380 119620 117400
rect 119880 117380 120120 117400
rect 120380 117380 120620 117400
rect 120880 117380 121120 117400
rect 121380 117380 121620 117400
rect 121880 117380 122120 117400
rect 122380 117380 122620 117400
rect 122880 117380 123120 117400
rect 123380 117380 123620 117400
rect 123880 117380 124120 117400
rect 124380 117380 124620 117400
rect 124880 117380 125120 117400
rect 125380 117380 125620 117400
rect 125880 117380 126120 117400
rect 126380 117380 126620 117400
rect 126880 117380 127120 117400
rect 127380 117380 127620 117400
rect 127880 117380 128120 117400
rect 128380 117380 128620 117400
rect 128880 117380 129120 117400
rect 129380 117380 129620 117400
rect 129880 117380 130120 117400
rect 130380 117380 130620 117400
rect 130880 117380 131120 117400
rect 131380 117380 131620 117400
rect 131880 117380 132120 117400
rect 132380 117380 132620 117400
rect 132880 117380 133120 117400
rect 133380 117380 133620 117400
rect 133880 117380 134120 117400
rect 134380 117380 134620 117400
rect 134880 117380 135120 117400
rect 135380 117380 135620 117400
rect 135880 117380 136120 117400
rect 136380 117380 136620 117400
rect 136880 117380 137120 117400
rect 137380 117380 137620 117400
rect 137880 117380 138120 117400
rect 138380 117380 138620 117400
rect 138880 117380 139120 117400
rect 139380 117380 139620 117400
rect 139880 117380 140120 117400
rect 140380 117380 140620 117400
rect 140880 117380 141120 117400
rect 141380 117380 141620 117400
rect 141880 117380 142000 117400
rect 118000 117120 118100 117380
rect 118400 117120 118600 117380
rect 118900 117120 119100 117380
rect 119400 117120 119600 117380
rect 119900 117120 120100 117380
rect 120400 117120 120600 117380
rect 120900 117120 121100 117380
rect 121400 117120 121600 117380
rect 121900 117120 122100 117380
rect 122400 117120 122600 117380
rect 122900 117120 123100 117380
rect 123400 117120 123600 117380
rect 123900 117120 124100 117380
rect 124400 117120 124600 117380
rect 124900 117120 125100 117380
rect 125400 117120 125600 117380
rect 125900 117120 126100 117380
rect 126400 117120 126600 117380
rect 126900 117120 127100 117380
rect 127400 117120 127600 117380
rect 127900 117120 128100 117380
rect 128400 117120 128600 117380
rect 128900 117120 129100 117380
rect 129400 117120 129600 117380
rect 129900 117120 130100 117380
rect 130400 117120 130600 117380
rect 130900 117120 131100 117380
rect 131400 117120 131600 117380
rect 131900 117120 132100 117380
rect 132400 117120 132600 117380
rect 132900 117120 133100 117380
rect 133400 117120 133600 117380
rect 133900 117120 134100 117380
rect 134400 117120 134600 117380
rect 134900 117120 135100 117380
rect 135400 117120 135600 117380
rect 135900 117120 136100 117380
rect 136400 117120 136600 117380
rect 136900 117120 137100 117380
rect 137400 117120 137600 117380
rect 137900 117120 138100 117380
rect 138400 117120 138600 117380
rect 138900 117120 139100 117380
rect 139400 117120 139600 117380
rect 139900 117120 140100 117380
rect 140400 117120 140600 117380
rect 140900 117120 141100 117380
rect 141400 117120 141600 117380
rect 141900 117120 142000 117380
rect 118000 117100 118120 117120
rect 118380 117100 118620 117120
rect 118880 117100 119120 117120
rect 119380 117100 119620 117120
rect 119880 117100 120120 117120
rect 120380 117100 120620 117120
rect 120880 117100 121120 117120
rect 121380 117100 121620 117120
rect 121880 117100 122120 117120
rect 122380 117100 122620 117120
rect 122880 117100 123120 117120
rect 123380 117100 123620 117120
rect 123880 117100 124120 117120
rect 124380 117100 124620 117120
rect 124880 117100 125120 117120
rect 125380 117100 125620 117120
rect 125880 117100 126120 117120
rect 126380 117100 126620 117120
rect 126880 117100 127120 117120
rect 127380 117100 127620 117120
rect 127880 117100 128120 117120
rect 128380 117100 128620 117120
rect 128880 117100 129120 117120
rect 129380 117100 129620 117120
rect 129880 117100 130120 117120
rect 130380 117100 130620 117120
rect 130880 117100 131120 117120
rect 131380 117100 131620 117120
rect 131880 117100 132120 117120
rect 132380 117100 132620 117120
rect 132880 117100 133120 117120
rect 133380 117100 133620 117120
rect 133880 117100 134120 117120
rect 134380 117100 134620 117120
rect 134880 117100 135120 117120
rect 135380 117100 135620 117120
rect 135880 117100 136120 117120
rect 136380 117100 136620 117120
rect 136880 117100 137120 117120
rect 137380 117100 137620 117120
rect 137880 117100 138120 117120
rect 138380 117100 138620 117120
rect 138880 117100 139120 117120
rect 139380 117100 139620 117120
rect 139880 117100 140120 117120
rect 140380 117100 140620 117120
rect 140880 117100 141120 117120
rect 141380 117100 141620 117120
rect 141880 117100 142000 117120
rect 118000 116900 142000 117100
rect 118000 116880 118120 116900
rect 118380 116880 118620 116900
rect 118880 116880 119120 116900
rect 119380 116880 119620 116900
rect 119880 116880 120120 116900
rect 120380 116880 120620 116900
rect 120880 116880 121120 116900
rect 121380 116880 121620 116900
rect 121880 116880 122120 116900
rect 122380 116880 122620 116900
rect 122880 116880 123120 116900
rect 123380 116880 123620 116900
rect 123880 116880 124120 116900
rect 124380 116880 124620 116900
rect 124880 116880 125120 116900
rect 125380 116880 125620 116900
rect 125880 116880 126120 116900
rect 126380 116880 126620 116900
rect 126880 116880 127120 116900
rect 127380 116880 127620 116900
rect 127880 116880 128120 116900
rect 128380 116880 128620 116900
rect 128880 116880 129120 116900
rect 129380 116880 129620 116900
rect 129880 116880 130120 116900
rect 130380 116880 130620 116900
rect 130880 116880 131120 116900
rect 131380 116880 131620 116900
rect 131880 116880 132120 116900
rect 132380 116880 132620 116900
rect 132880 116880 133120 116900
rect 133380 116880 133620 116900
rect 133880 116880 134120 116900
rect 134380 116880 134620 116900
rect 134880 116880 135120 116900
rect 135380 116880 135620 116900
rect 135880 116880 136120 116900
rect 136380 116880 136620 116900
rect 136880 116880 137120 116900
rect 137380 116880 137620 116900
rect 137880 116880 138120 116900
rect 138380 116880 138620 116900
rect 138880 116880 139120 116900
rect 139380 116880 139620 116900
rect 139880 116880 140120 116900
rect 140380 116880 140620 116900
rect 140880 116880 141120 116900
rect 141380 116880 141620 116900
rect 141880 116880 142000 116900
rect 118000 116620 118100 116880
rect 118400 116620 118600 116880
rect 118900 116620 119100 116880
rect 119400 116620 119600 116880
rect 119900 116620 120100 116880
rect 120400 116620 120600 116880
rect 120900 116620 121100 116880
rect 121400 116620 121600 116880
rect 121900 116620 122100 116880
rect 122400 116620 122600 116880
rect 122900 116620 123100 116880
rect 123400 116620 123600 116880
rect 123900 116620 124100 116880
rect 124400 116620 124600 116880
rect 124900 116620 125100 116880
rect 125400 116620 125600 116880
rect 125900 116620 126100 116880
rect 126400 116620 126600 116880
rect 126900 116620 127100 116880
rect 127400 116620 127600 116880
rect 127900 116620 128100 116880
rect 128400 116620 128600 116880
rect 128900 116620 129100 116880
rect 129400 116620 129600 116880
rect 129900 116620 130100 116880
rect 130400 116620 130600 116880
rect 130900 116620 131100 116880
rect 131400 116620 131600 116880
rect 131900 116620 132100 116880
rect 132400 116620 132600 116880
rect 132900 116620 133100 116880
rect 133400 116620 133600 116880
rect 133900 116620 134100 116880
rect 134400 116620 134600 116880
rect 134900 116620 135100 116880
rect 135400 116620 135600 116880
rect 135900 116620 136100 116880
rect 136400 116620 136600 116880
rect 136900 116620 137100 116880
rect 137400 116620 137600 116880
rect 137900 116620 138100 116880
rect 138400 116620 138600 116880
rect 138900 116620 139100 116880
rect 139400 116620 139600 116880
rect 139900 116620 140100 116880
rect 140400 116620 140600 116880
rect 140900 116620 141100 116880
rect 141400 116620 141600 116880
rect 141900 116620 142000 116880
rect 118000 116600 118120 116620
rect 118380 116600 118620 116620
rect 118880 116600 119120 116620
rect 119380 116600 119620 116620
rect 119880 116600 120120 116620
rect 120380 116600 120620 116620
rect 120880 116600 121120 116620
rect 121380 116600 121620 116620
rect 121880 116600 122120 116620
rect 122380 116600 122620 116620
rect 122880 116600 123120 116620
rect 123380 116600 123620 116620
rect 123880 116600 124120 116620
rect 124380 116600 124620 116620
rect 124880 116600 125120 116620
rect 125380 116600 125620 116620
rect 125880 116600 126120 116620
rect 126380 116600 126620 116620
rect 126880 116600 127120 116620
rect 127380 116600 127620 116620
rect 127880 116600 128120 116620
rect 128380 116600 128620 116620
rect 128880 116600 129120 116620
rect 129380 116600 129620 116620
rect 129880 116600 130120 116620
rect 130380 116600 130620 116620
rect 130880 116600 131120 116620
rect 131380 116600 131620 116620
rect 131880 116600 132120 116620
rect 132380 116600 132620 116620
rect 132880 116600 133120 116620
rect 133380 116600 133620 116620
rect 133880 116600 134120 116620
rect 134380 116600 134620 116620
rect 134880 116600 135120 116620
rect 135380 116600 135620 116620
rect 135880 116600 136120 116620
rect 136380 116600 136620 116620
rect 136880 116600 137120 116620
rect 137380 116600 137620 116620
rect 137880 116600 138120 116620
rect 138380 116600 138620 116620
rect 138880 116600 139120 116620
rect 139380 116600 139620 116620
rect 139880 116600 140120 116620
rect 140380 116600 140620 116620
rect 140880 116600 141120 116620
rect 141380 116600 141620 116620
rect 141880 116600 142000 116620
rect 118000 116400 142000 116600
rect 118000 116380 118120 116400
rect 118380 116380 118620 116400
rect 118880 116380 119120 116400
rect 119380 116380 119620 116400
rect 119880 116380 120120 116400
rect 120380 116380 120620 116400
rect 120880 116380 121120 116400
rect 121380 116380 121620 116400
rect 121880 116380 122120 116400
rect 122380 116380 122620 116400
rect 122880 116380 123120 116400
rect 123380 116380 123620 116400
rect 123880 116380 124120 116400
rect 124380 116380 124620 116400
rect 124880 116380 125120 116400
rect 125380 116380 125620 116400
rect 125880 116380 126120 116400
rect 126380 116380 126620 116400
rect 126880 116380 127120 116400
rect 127380 116380 127620 116400
rect 127880 116380 128120 116400
rect 128380 116380 128620 116400
rect 128880 116380 129120 116400
rect 129380 116380 129620 116400
rect 129880 116380 130120 116400
rect 130380 116380 130620 116400
rect 130880 116380 131120 116400
rect 131380 116380 131620 116400
rect 131880 116380 132120 116400
rect 132380 116380 132620 116400
rect 132880 116380 133120 116400
rect 133380 116380 133620 116400
rect 133880 116380 134120 116400
rect 134380 116380 134620 116400
rect 134880 116380 135120 116400
rect 135380 116380 135620 116400
rect 135880 116380 136120 116400
rect 136380 116380 136620 116400
rect 136880 116380 137120 116400
rect 137380 116380 137620 116400
rect 137880 116380 138120 116400
rect 138380 116380 138620 116400
rect 138880 116380 139120 116400
rect 139380 116380 139620 116400
rect 139880 116380 140120 116400
rect 140380 116380 140620 116400
rect 140880 116380 141120 116400
rect 141380 116380 141620 116400
rect 141880 116380 142000 116400
rect 118000 116120 118100 116380
rect 118400 116120 118600 116380
rect 118900 116120 119100 116380
rect 119400 116120 119600 116380
rect 119900 116120 120100 116380
rect 120400 116120 120600 116380
rect 120900 116120 121100 116380
rect 121400 116120 121600 116380
rect 121900 116120 122100 116380
rect 122400 116120 122600 116380
rect 122900 116120 123100 116380
rect 123400 116120 123600 116380
rect 123900 116120 124100 116380
rect 124400 116120 124600 116380
rect 124900 116120 125100 116380
rect 125400 116120 125600 116380
rect 125900 116120 126100 116380
rect 126400 116120 126600 116380
rect 126900 116120 127100 116380
rect 127400 116120 127600 116380
rect 127900 116120 128100 116380
rect 128400 116120 128600 116380
rect 128900 116120 129100 116380
rect 129400 116120 129600 116380
rect 129900 116120 130100 116380
rect 130400 116120 130600 116380
rect 130900 116120 131100 116380
rect 131400 116120 131600 116380
rect 131900 116120 132100 116380
rect 132400 116120 132600 116380
rect 132900 116120 133100 116380
rect 133400 116120 133600 116380
rect 133900 116120 134100 116380
rect 134400 116120 134600 116380
rect 134900 116120 135100 116380
rect 135400 116120 135600 116380
rect 135900 116120 136100 116380
rect 136400 116120 136600 116380
rect 136900 116120 137100 116380
rect 137400 116120 137600 116380
rect 137900 116120 138100 116380
rect 138400 116120 138600 116380
rect 138900 116120 139100 116380
rect 139400 116120 139600 116380
rect 139900 116120 140100 116380
rect 140400 116120 140600 116380
rect 140900 116120 141100 116380
rect 141400 116120 141600 116380
rect 141900 116120 142000 116380
rect 118000 116100 118120 116120
rect 118380 116100 118620 116120
rect 118880 116100 119120 116120
rect 119380 116100 119620 116120
rect 119880 116100 120120 116120
rect 120380 116100 120620 116120
rect 120880 116100 121120 116120
rect 121380 116100 121620 116120
rect 121880 116100 122120 116120
rect 122380 116100 122620 116120
rect 122880 116100 123120 116120
rect 123380 116100 123620 116120
rect 123880 116100 124120 116120
rect 124380 116100 124620 116120
rect 124880 116100 125120 116120
rect 125380 116100 125620 116120
rect 125880 116100 126120 116120
rect 126380 116100 126620 116120
rect 126880 116100 127120 116120
rect 127380 116100 127620 116120
rect 127880 116100 128120 116120
rect 128380 116100 128620 116120
rect 128880 116100 129120 116120
rect 129380 116100 129620 116120
rect 129880 116100 130120 116120
rect 130380 116100 130620 116120
rect 130880 116100 131120 116120
rect 131380 116100 131620 116120
rect 131880 116100 132120 116120
rect 132380 116100 132620 116120
rect 132880 116100 133120 116120
rect 133380 116100 133620 116120
rect 133880 116100 134120 116120
rect 134380 116100 134620 116120
rect 134880 116100 135120 116120
rect 135380 116100 135620 116120
rect 135880 116100 136120 116120
rect 136380 116100 136620 116120
rect 136880 116100 137120 116120
rect 137380 116100 137620 116120
rect 137880 116100 138120 116120
rect 138380 116100 138620 116120
rect 138880 116100 139120 116120
rect 139380 116100 139620 116120
rect 139880 116100 140120 116120
rect 140380 116100 140620 116120
rect 140880 116100 141120 116120
rect 141380 116100 141620 116120
rect 141880 116100 142000 116120
rect 118000 115900 142000 116100
rect 118000 115880 118120 115900
rect 118380 115880 118620 115900
rect 118880 115880 119120 115900
rect 119380 115880 119620 115900
rect 119880 115880 120120 115900
rect 120380 115880 120620 115900
rect 120880 115880 121120 115900
rect 121380 115880 121620 115900
rect 121880 115880 122120 115900
rect 122380 115880 122620 115900
rect 122880 115880 123120 115900
rect 123380 115880 123620 115900
rect 123880 115880 124120 115900
rect 124380 115880 124620 115900
rect 124880 115880 125120 115900
rect 125380 115880 125620 115900
rect 125880 115880 126120 115900
rect 126380 115880 126620 115900
rect 126880 115880 127120 115900
rect 127380 115880 127620 115900
rect 127880 115880 128120 115900
rect 128380 115880 128620 115900
rect 128880 115880 129120 115900
rect 129380 115880 129620 115900
rect 129880 115880 130120 115900
rect 130380 115880 130620 115900
rect 130880 115880 131120 115900
rect 131380 115880 131620 115900
rect 131880 115880 132120 115900
rect 132380 115880 132620 115900
rect 132880 115880 133120 115900
rect 133380 115880 133620 115900
rect 133880 115880 134120 115900
rect 134380 115880 134620 115900
rect 134880 115880 135120 115900
rect 135380 115880 135620 115900
rect 135880 115880 136120 115900
rect 136380 115880 136620 115900
rect 136880 115880 137120 115900
rect 137380 115880 137620 115900
rect 137880 115880 138120 115900
rect 138380 115880 138620 115900
rect 138880 115880 139120 115900
rect 139380 115880 139620 115900
rect 139880 115880 140120 115900
rect 140380 115880 140620 115900
rect 140880 115880 141120 115900
rect 141380 115880 141620 115900
rect 141880 115880 142000 115900
rect 118000 115620 118100 115880
rect 118400 115620 118600 115880
rect 118900 115620 119100 115880
rect 119400 115620 119600 115880
rect 119900 115620 120100 115880
rect 120400 115620 120600 115880
rect 120900 115620 121100 115880
rect 121400 115620 121600 115880
rect 121900 115620 122100 115880
rect 122400 115620 122600 115880
rect 122900 115620 123100 115880
rect 123400 115620 123600 115880
rect 123900 115620 124100 115880
rect 124400 115620 124600 115880
rect 124900 115620 125100 115880
rect 125400 115620 125600 115880
rect 125900 115620 126100 115880
rect 126400 115620 126600 115880
rect 126900 115620 127100 115880
rect 127400 115620 127600 115880
rect 127900 115620 128100 115880
rect 128400 115620 128600 115880
rect 128900 115620 129100 115880
rect 129400 115620 129600 115880
rect 129900 115620 130100 115880
rect 130400 115620 130600 115880
rect 130900 115620 131100 115880
rect 131400 115620 131600 115880
rect 131900 115620 132100 115880
rect 132400 115620 132600 115880
rect 132900 115620 133100 115880
rect 133400 115620 133600 115880
rect 133900 115620 134100 115880
rect 134400 115620 134600 115880
rect 134900 115620 135100 115880
rect 135400 115620 135600 115880
rect 135900 115620 136100 115880
rect 136400 115620 136600 115880
rect 136900 115620 137100 115880
rect 137400 115620 137600 115880
rect 137900 115620 138100 115880
rect 138400 115620 138600 115880
rect 138900 115620 139100 115880
rect 139400 115620 139600 115880
rect 139900 115620 140100 115880
rect 140400 115620 140600 115880
rect 140900 115620 141100 115880
rect 141400 115620 141600 115880
rect 141900 115620 142000 115880
rect 118000 115600 118120 115620
rect 118380 115600 118620 115620
rect 118880 115600 119120 115620
rect 119380 115600 119620 115620
rect 119880 115600 120120 115620
rect 120380 115600 120620 115620
rect 120880 115600 121120 115620
rect 121380 115600 121620 115620
rect 121880 115600 122120 115620
rect 122380 115600 122620 115620
rect 122880 115600 123120 115620
rect 123380 115600 123620 115620
rect 123880 115600 124120 115620
rect 124380 115600 124620 115620
rect 124880 115600 125120 115620
rect 125380 115600 125620 115620
rect 125880 115600 126120 115620
rect 126380 115600 126620 115620
rect 126880 115600 127120 115620
rect 127380 115600 127620 115620
rect 127880 115600 128120 115620
rect 128380 115600 128620 115620
rect 128880 115600 129120 115620
rect 129380 115600 129620 115620
rect 129880 115600 130120 115620
rect 130380 115600 130620 115620
rect 130880 115600 131120 115620
rect 131380 115600 131620 115620
rect 131880 115600 132120 115620
rect 132380 115600 132620 115620
rect 132880 115600 133120 115620
rect 133380 115600 133620 115620
rect 133880 115600 134120 115620
rect 134380 115600 134620 115620
rect 134880 115600 135120 115620
rect 135380 115600 135620 115620
rect 135880 115600 136120 115620
rect 136380 115600 136620 115620
rect 136880 115600 137120 115620
rect 137380 115600 137620 115620
rect 137880 115600 138120 115620
rect 138380 115600 138620 115620
rect 138880 115600 139120 115620
rect 139380 115600 139620 115620
rect 139880 115600 140120 115620
rect 140380 115600 140620 115620
rect 140880 115600 141120 115620
rect 141380 115600 141620 115620
rect 141880 115600 142000 115620
rect 118000 115400 142000 115600
rect 118000 115380 118120 115400
rect 118380 115380 118620 115400
rect 118880 115380 119120 115400
rect 119380 115380 119620 115400
rect 119880 115380 120120 115400
rect 120380 115380 120620 115400
rect 120880 115380 121120 115400
rect 121380 115380 121620 115400
rect 121880 115380 122120 115400
rect 122380 115380 122620 115400
rect 122880 115380 123120 115400
rect 123380 115380 123620 115400
rect 123880 115380 124120 115400
rect 124380 115380 124620 115400
rect 124880 115380 125120 115400
rect 125380 115380 125620 115400
rect 125880 115380 126120 115400
rect 126380 115380 126620 115400
rect 126880 115380 127120 115400
rect 127380 115380 127620 115400
rect 127880 115380 128120 115400
rect 128380 115380 128620 115400
rect 128880 115380 129120 115400
rect 129380 115380 129620 115400
rect 129880 115380 130120 115400
rect 130380 115380 130620 115400
rect 130880 115380 131120 115400
rect 131380 115380 131620 115400
rect 131880 115380 132120 115400
rect 132380 115380 132620 115400
rect 132880 115380 133120 115400
rect 133380 115380 133620 115400
rect 133880 115380 134120 115400
rect 134380 115380 134620 115400
rect 134880 115380 135120 115400
rect 135380 115380 135620 115400
rect 135880 115380 136120 115400
rect 136380 115380 136620 115400
rect 136880 115380 137120 115400
rect 137380 115380 137620 115400
rect 137880 115380 138120 115400
rect 138380 115380 138620 115400
rect 138880 115380 139120 115400
rect 139380 115380 139620 115400
rect 139880 115380 140120 115400
rect 140380 115380 140620 115400
rect 140880 115380 141120 115400
rect 141380 115380 141620 115400
rect 141880 115380 142000 115400
rect 118000 115120 118100 115380
rect 118400 115120 118600 115380
rect 118900 115120 119100 115380
rect 119400 115120 119600 115380
rect 119900 115120 120100 115380
rect 120400 115120 120600 115380
rect 120900 115120 121100 115380
rect 121400 115120 121600 115380
rect 121900 115120 122100 115380
rect 122400 115120 122600 115380
rect 122900 115120 123100 115380
rect 123400 115120 123600 115380
rect 123900 115120 124100 115380
rect 124400 115120 124600 115380
rect 124900 115120 125100 115380
rect 125400 115120 125600 115380
rect 125900 115120 126100 115380
rect 126400 115120 126600 115380
rect 126900 115120 127100 115380
rect 127400 115120 127600 115380
rect 127900 115120 128100 115380
rect 128400 115120 128600 115380
rect 128900 115120 129100 115380
rect 129400 115120 129600 115380
rect 129900 115120 130100 115380
rect 130400 115120 130600 115380
rect 130900 115120 131100 115380
rect 131400 115120 131600 115380
rect 131900 115120 132100 115380
rect 132400 115120 132600 115380
rect 132900 115120 133100 115380
rect 133400 115120 133600 115380
rect 133900 115120 134100 115380
rect 134400 115120 134600 115380
rect 134900 115120 135100 115380
rect 135400 115120 135600 115380
rect 135900 115120 136100 115380
rect 136400 115120 136600 115380
rect 136900 115120 137100 115380
rect 137400 115120 137600 115380
rect 137900 115120 138100 115380
rect 138400 115120 138600 115380
rect 138900 115120 139100 115380
rect 139400 115120 139600 115380
rect 139900 115120 140100 115380
rect 140400 115120 140600 115380
rect 140900 115120 141100 115380
rect 141400 115120 141600 115380
rect 141900 115120 142000 115380
rect 118000 115100 118120 115120
rect 118380 115100 118620 115120
rect 118880 115100 119120 115120
rect 119380 115100 119620 115120
rect 119880 115100 120120 115120
rect 120380 115100 120620 115120
rect 120880 115100 121120 115120
rect 121380 115100 121620 115120
rect 121880 115100 122120 115120
rect 122380 115100 122620 115120
rect 122880 115100 123120 115120
rect 123380 115100 123620 115120
rect 123880 115100 124120 115120
rect 124380 115100 124620 115120
rect 124880 115100 125120 115120
rect 125380 115100 125620 115120
rect 125880 115100 126120 115120
rect 126380 115100 126620 115120
rect 126880 115100 127120 115120
rect 127380 115100 127620 115120
rect 127880 115100 128120 115120
rect 128380 115100 128620 115120
rect 128880 115100 129120 115120
rect 129380 115100 129620 115120
rect 129880 115100 130120 115120
rect 130380 115100 130620 115120
rect 130880 115100 131120 115120
rect 131380 115100 131620 115120
rect 131880 115100 132120 115120
rect 132380 115100 132620 115120
rect 132880 115100 133120 115120
rect 133380 115100 133620 115120
rect 133880 115100 134120 115120
rect 134380 115100 134620 115120
rect 134880 115100 135120 115120
rect 135380 115100 135620 115120
rect 135880 115100 136120 115120
rect 136380 115100 136620 115120
rect 136880 115100 137120 115120
rect 137380 115100 137620 115120
rect 137880 115100 138120 115120
rect 138380 115100 138620 115120
rect 138880 115100 139120 115120
rect 139380 115100 139620 115120
rect 139880 115100 140120 115120
rect 140380 115100 140620 115120
rect 140880 115100 141120 115120
rect 141380 115100 141620 115120
rect 141880 115100 142000 115120
rect 118000 114900 142000 115100
rect 118000 114880 118120 114900
rect 118380 114880 118620 114900
rect 118880 114880 119120 114900
rect 119380 114880 119620 114900
rect 119880 114880 120120 114900
rect 120380 114880 120620 114900
rect 120880 114880 121120 114900
rect 121380 114880 121620 114900
rect 121880 114880 122120 114900
rect 122380 114880 122620 114900
rect 122880 114880 123120 114900
rect 123380 114880 123620 114900
rect 123880 114880 124120 114900
rect 124380 114880 124620 114900
rect 124880 114880 125120 114900
rect 125380 114880 125620 114900
rect 125880 114880 126120 114900
rect 126380 114880 126620 114900
rect 126880 114880 127120 114900
rect 127380 114880 127620 114900
rect 127880 114880 128120 114900
rect 128380 114880 128620 114900
rect 128880 114880 129120 114900
rect 129380 114880 129620 114900
rect 129880 114880 130120 114900
rect 130380 114880 130620 114900
rect 130880 114880 131120 114900
rect 131380 114880 131620 114900
rect 131880 114880 132120 114900
rect 132380 114880 132620 114900
rect 132880 114880 133120 114900
rect 133380 114880 133620 114900
rect 133880 114880 134120 114900
rect 134380 114880 134620 114900
rect 134880 114880 135120 114900
rect 135380 114880 135620 114900
rect 135880 114880 136120 114900
rect 136380 114880 136620 114900
rect 136880 114880 137120 114900
rect 137380 114880 137620 114900
rect 137880 114880 138120 114900
rect 138380 114880 138620 114900
rect 138880 114880 139120 114900
rect 139380 114880 139620 114900
rect 139880 114880 140120 114900
rect 140380 114880 140620 114900
rect 140880 114880 141120 114900
rect 141380 114880 141620 114900
rect 141880 114880 142000 114900
rect 118000 114620 118100 114880
rect 118400 114620 118600 114880
rect 118900 114620 119100 114880
rect 119400 114620 119600 114880
rect 119900 114620 120100 114880
rect 120400 114620 120600 114880
rect 120900 114620 121100 114880
rect 121400 114620 121600 114880
rect 121900 114620 122100 114880
rect 122400 114620 122600 114880
rect 122900 114620 123100 114880
rect 123400 114620 123600 114880
rect 123900 114620 124100 114880
rect 124400 114620 124600 114880
rect 124900 114620 125100 114880
rect 125400 114620 125600 114880
rect 125900 114620 126100 114880
rect 126400 114620 126600 114880
rect 126900 114620 127100 114880
rect 127400 114620 127600 114880
rect 127900 114620 128100 114880
rect 128400 114620 128600 114880
rect 128900 114620 129100 114880
rect 129400 114620 129600 114880
rect 129900 114620 130100 114880
rect 130400 114620 130600 114880
rect 130900 114620 131100 114880
rect 131400 114620 131600 114880
rect 131900 114620 132100 114880
rect 132400 114620 132600 114880
rect 132900 114620 133100 114880
rect 133400 114620 133600 114880
rect 133900 114620 134100 114880
rect 134400 114620 134600 114880
rect 134900 114620 135100 114880
rect 135400 114620 135600 114880
rect 135900 114620 136100 114880
rect 136400 114620 136600 114880
rect 136900 114620 137100 114880
rect 137400 114620 137600 114880
rect 137900 114620 138100 114880
rect 138400 114620 138600 114880
rect 138900 114620 139100 114880
rect 139400 114620 139600 114880
rect 139900 114620 140100 114880
rect 140400 114620 140600 114880
rect 140900 114620 141100 114880
rect 141400 114620 141600 114880
rect 141900 114620 142000 114880
rect 118000 114600 118120 114620
rect 118380 114600 118620 114620
rect 118880 114600 119120 114620
rect 119380 114600 119620 114620
rect 119880 114600 120120 114620
rect 120380 114600 120620 114620
rect 120880 114600 121120 114620
rect 121380 114600 121620 114620
rect 121880 114600 122120 114620
rect 122380 114600 122620 114620
rect 122880 114600 123120 114620
rect 123380 114600 123620 114620
rect 123880 114600 124120 114620
rect 124380 114600 124620 114620
rect 124880 114600 125120 114620
rect 125380 114600 125620 114620
rect 125880 114600 126120 114620
rect 126380 114600 126620 114620
rect 126880 114600 127120 114620
rect 127380 114600 127620 114620
rect 127880 114600 128120 114620
rect 128380 114600 128620 114620
rect 128880 114600 129120 114620
rect 129380 114600 129620 114620
rect 129880 114600 130120 114620
rect 130380 114600 130620 114620
rect 130880 114600 131120 114620
rect 131380 114600 131620 114620
rect 131880 114600 132120 114620
rect 132380 114600 132620 114620
rect 132880 114600 133120 114620
rect 133380 114600 133620 114620
rect 133880 114600 134120 114620
rect 134380 114600 134620 114620
rect 134880 114600 135120 114620
rect 135380 114600 135620 114620
rect 135880 114600 136120 114620
rect 136380 114600 136620 114620
rect 136880 114600 137120 114620
rect 137380 114600 137620 114620
rect 137880 114600 138120 114620
rect 138380 114600 138620 114620
rect 138880 114600 139120 114620
rect 139380 114600 139620 114620
rect 139880 114600 140120 114620
rect 140380 114600 140620 114620
rect 140880 114600 141120 114620
rect 141380 114600 141620 114620
rect 141880 114600 142000 114620
rect 118000 114400 142000 114600
rect 118000 114380 118120 114400
rect 118380 114380 118620 114400
rect 118880 114380 119120 114400
rect 119380 114380 119620 114400
rect 119880 114380 120120 114400
rect 120380 114380 120620 114400
rect 120880 114380 121120 114400
rect 121380 114380 121620 114400
rect 121880 114380 122120 114400
rect 122380 114380 122620 114400
rect 122880 114380 123120 114400
rect 123380 114380 123620 114400
rect 123880 114380 124120 114400
rect 124380 114380 124620 114400
rect 124880 114380 125120 114400
rect 125380 114380 125620 114400
rect 125880 114380 126120 114400
rect 126380 114380 126620 114400
rect 126880 114380 127120 114400
rect 127380 114380 127620 114400
rect 127880 114380 128120 114400
rect 128380 114380 128620 114400
rect 128880 114380 129120 114400
rect 129380 114380 129620 114400
rect 129880 114380 130120 114400
rect 130380 114380 130620 114400
rect 130880 114380 131120 114400
rect 131380 114380 131620 114400
rect 131880 114380 132120 114400
rect 132380 114380 132620 114400
rect 132880 114380 133120 114400
rect 133380 114380 133620 114400
rect 133880 114380 134120 114400
rect 134380 114380 134620 114400
rect 134880 114380 135120 114400
rect 135380 114380 135620 114400
rect 135880 114380 136120 114400
rect 136380 114380 136620 114400
rect 136880 114380 137120 114400
rect 137380 114380 137620 114400
rect 137880 114380 138120 114400
rect 138380 114380 138620 114400
rect 138880 114380 139120 114400
rect 139380 114380 139620 114400
rect 139880 114380 140120 114400
rect 140380 114380 140620 114400
rect 140880 114380 141120 114400
rect 141380 114380 141620 114400
rect 141880 114380 142000 114400
rect 118000 114120 118100 114380
rect 118400 114120 118600 114380
rect 118900 114120 119100 114380
rect 119400 114120 119600 114380
rect 119900 114120 120100 114380
rect 120400 114120 120600 114380
rect 120900 114120 121100 114380
rect 121400 114120 121600 114380
rect 121900 114120 122100 114380
rect 122400 114120 122600 114380
rect 122900 114120 123100 114380
rect 123400 114120 123600 114380
rect 123900 114120 124100 114380
rect 124400 114120 124600 114380
rect 124900 114120 125100 114380
rect 125400 114120 125600 114380
rect 125900 114120 126100 114380
rect 126400 114120 126600 114380
rect 126900 114120 127100 114380
rect 127400 114120 127600 114380
rect 127900 114120 128100 114380
rect 128400 114120 128600 114380
rect 128900 114120 129100 114380
rect 129400 114120 129600 114380
rect 129900 114120 130100 114380
rect 130400 114120 130600 114380
rect 130900 114120 131100 114380
rect 131400 114120 131600 114380
rect 131900 114120 132100 114380
rect 132400 114120 132600 114380
rect 132900 114120 133100 114380
rect 133400 114120 133600 114380
rect 133900 114120 134100 114380
rect 134400 114120 134600 114380
rect 134900 114120 135100 114380
rect 135400 114120 135600 114380
rect 135900 114120 136100 114380
rect 136400 114120 136600 114380
rect 136900 114120 137100 114380
rect 137400 114120 137600 114380
rect 137900 114120 138100 114380
rect 138400 114120 138600 114380
rect 138900 114120 139100 114380
rect 139400 114120 139600 114380
rect 139900 114120 140100 114380
rect 140400 114120 140600 114380
rect 140900 114120 141100 114380
rect 141400 114120 141600 114380
rect 141900 114120 142000 114380
rect 118000 114100 118120 114120
rect 118380 114100 118620 114120
rect 118880 114100 119120 114120
rect 119380 114100 119620 114120
rect 119880 114100 120120 114120
rect 120380 114100 120620 114120
rect 120880 114100 121120 114120
rect 121380 114100 121620 114120
rect 121880 114100 122120 114120
rect 122380 114100 122620 114120
rect 122880 114100 123120 114120
rect 123380 114100 123620 114120
rect 123880 114100 124120 114120
rect 124380 114100 124620 114120
rect 124880 114100 125120 114120
rect 125380 114100 125620 114120
rect 125880 114100 126120 114120
rect 126380 114100 126620 114120
rect 126880 114100 127120 114120
rect 127380 114100 127620 114120
rect 127880 114100 128120 114120
rect 128380 114100 128620 114120
rect 128880 114100 129120 114120
rect 129380 114100 129620 114120
rect 129880 114100 130120 114120
rect 130380 114100 130620 114120
rect 130880 114100 131120 114120
rect 131380 114100 131620 114120
rect 131880 114100 132120 114120
rect 132380 114100 132620 114120
rect 132880 114100 133120 114120
rect 133380 114100 133620 114120
rect 133880 114100 134120 114120
rect 134380 114100 134620 114120
rect 134880 114100 135120 114120
rect 135380 114100 135620 114120
rect 135880 114100 136120 114120
rect 136380 114100 136620 114120
rect 136880 114100 137120 114120
rect 137380 114100 137620 114120
rect 137880 114100 138120 114120
rect 138380 114100 138620 114120
rect 138880 114100 139120 114120
rect 139380 114100 139620 114120
rect 139880 114100 140120 114120
rect 140380 114100 140620 114120
rect 140880 114100 141120 114120
rect 141380 114100 141620 114120
rect 141880 114100 142000 114120
rect 118000 114000 142000 114100
rect 162000 121900 184000 122000
rect 162000 121880 162120 121900
rect 162380 121880 162620 121900
rect 162880 121880 163120 121900
rect 163380 121880 163620 121900
rect 163880 121880 164120 121900
rect 164380 121880 164620 121900
rect 164880 121880 165120 121900
rect 165380 121880 165620 121900
rect 165880 121880 166120 121900
rect 166380 121880 166620 121900
rect 166880 121880 167120 121900
rect 167380 121880 167620 121900
rect 167880 121880 168120 121900
rect 168380 121880 168620 121900
rect 168880 121880 169120 121900
rect 169380 121880 169620 121900
rect 169880 121880 170120 121900
rect 170380 121880 170620 121900
rect 170880 121880 171120 121900
rect 171380 121880 171620 121900
rect 171880 121880 172120 121900
rect 172380 121880 172620 121900
rect 172880 121880 173120 121900
rect 173380 121880 173620 121900
rect 173880 121880 174120 121900
rect 174380 121880 174620 121900
rect 174880 121880 175120 121900
rect 175380 121880 175620 121900
rect 175880 121880 176120 121900
rect 176380 121880 176620 121900
rect 176880 121880 177120 121900
rect 177380 121880 177620 121900
rect 177880 121880 178120 121900
rect 178380 121880 178620 121900
rect 178880 121880 179120 121900
rect 179380 121880 179620 121900
rect 179880 121880 180120 121900
rect 180380 121880 180620 121900
rect 180880 121880 181120 121900
rect 181380 121880 181620 121900
rect 181880 121880 182120 121900
rect 182380 121880 182620 121900
rect 182880 121880 183120 121900
rect 183380 121880 183620 121900
rect 183880 121880 184000 121900
rect 162000 121620 162100 121880
rect 162400 121620 162600 121880
rect 162900 121620 163100 121880
rect 163400 121620 163600 121880
rect 163900 121620 164100 121880
rect 164400 121620 164600 121880
rect 164900 121620 165100 121880
rect 165400 121620 165600 121880
rect 165900 121620 166100 121880
rect 166400 121620 166600 121880
rect 166900 121620 167100 121880
rect 167400 121620 167600 121880
rect 167900 121620 168100 121880
rect 168400 121620 168600 121880
rect 168900 121620 169100 121880
rect 169400 121620 169600 121880
rect 169900 121620 170100 121880
rect 170400 121620 170600 121880
rect 170900 121620 171100 121880
rect 171400 121620 171600 121880
rect 171900 121620 172100 121880
rect 172400 121620 172600 121880
rect 172900 121620 173100 121880
rect 173400 121620 173600 121880
rect 173900 121620 174100 121880
rect 174400 121620 174600 121880
rect 174900 121620 175100 121880
rect 175400 121620 175600 121880
rect 175900 121620 176100 121880
rect 176400 121620 176600 121880
rect 176900 121620 177100 121880
rect 177400 121620 177600 121880
rect 177900 121620 178100 121880
rect 178400 121620 178600 121880
rect 178900 121620 179100 121880
rect 179400 121620 179600 121880
rect 179900 121620 180100 121880
rect 180400 121620 180600 121880
rect 180900 121620 181100 121880
rect 181400 121620 181600 121880
rect 181900 121620 182100 121880
rect 182400 121620 182600 121880
rect 182900 121620 183100 121880
rect 183400 121620 183600 121880
rect 183900 121620 184000 121880
rect 162000 121600 162120 121620
rect 162380 121600 162620 121620
rect 162880 121600 163120 121620
rect 163380 121600 163620 121620
rect 163880 121600 164120 121620
rect 164380 121600 164620 121620
rect 164880 121600 165120 121620
rect 165380 121600 165620 121620
rect 165880 121600 166120 121620
rect 166380 121600 166620 121620
rect 166880 121600 167120 121620
rect 167380 121600 167620 121620
rect 167880 121600 168120 121620
rect 168380 121600 168620 121620
rect 168880 121600 169120 121620
rect 169380 121600 169620 121620
rect 169880 121600 170120 121620
rect 170380 121600 170620 121620
rect 170880 121600 171120 121620
rect 171380 121600 171620 121620
rect 171880 121600 172120 121620
rect 172380 121600 172620 121620
rect 172880 121600 173120 121620
rect 173380 121600 173620 121620
rect 173880 121600 174120 121620
rect 174380 121600 174620 121620
rect 174880 121600 175120 121620
rect 175380 121600 175620 121620
rect 175880 121600 176120 121620
rect 176380 121600 176620 121620
rect 176880 121600 177120 121620
rect 177380 121600 177620 121620
rect 177880 121600 178120 121620
rect 178380 121600 178620 121620
rect 178880 121600 179120 121620
rect 179380 121600 179620 121620
rect 179880 121600 180120 121620
rect 180380 121600 180620 121620
rect 180880 121600 181120 121620
rect 181380 121600 181620 121620
rect 181880 121600 182120 121620
rect 182380 121600 182620 121620
rect 182880 121600 183120 121620
rect 183380 121600 183620 121620
rect 183880 121600 184000 121620
rect 162000 121400 184000 121600
rect 162000 121380 162120 121400
rect 162380 121380 162620 121400
rect 162880 121380 163120 121400
rect 163380 121380 163620 121400
rect 163880 121380 164120 121400
rect 164380 121380 164620 121400
rect 164880 121380 165120 121400
rect 165380 121380 165620 121400
rect 165880 121380 166120 121400
rect 166380 121380 166620 121400
rect 166880 121380 167120 121400
rect 167380 121380 167620 121400
rect 167880 121380 168120 121400
rect 168380 121380 168620 121400
rect 168880 121380 169120 121400
rect 169380 121380 169620 121400
rect 169880 121380 170120 121400
rect 170380 121380 170620 121400
rect 170880 121380 171120 121400
rect 171380 121380 171620 121400
rect 171880 121380 172120 121400
rect 172380 121380 172620 121400
rect 172880 121380 173120 121400
rect 173380 121380 173620 121400
rect 173880 121380 174120 121400
rect 174380 121380 174620 121400
rect 174880 121380 175120 121400
rect 175380 121380 175620 121400
rect 175880 121380 176120 121400
rect 176380 121380 176620 121400
rect 176880 121380 177120 121400
rect 177380 121380 177620 121400
rect 177880 121380 178120 121400
rect 178380 121380 178620 121400
rect 178880 121380 179120 121400
rect 179380 121380 179620 121400
rect 179880 121380 180120 121400
rect 180380 121380 180620 121400
rect 180880 121380 181120 121400
rect 181380 121380 181620 121400
rect 181880 121380 182120 121400
rect 182380 121380 182620 121400
rect 182880 121380 183120 121400
rect 183380 121380 183620 121400
rect 183880 121380 184000 121400
rect 162000 121120 162100 121380
rect 162400 121120 162600 121380
rect 162900 121120 163100 121380
rect 163400 121120 163600 121380
rect 163900 121120 164100 121380
rect 164400 121120 164600 121380
rect 164900 121120 165100 121380
rect 165400 121120 165600 121380
rect 165900 121120 166100 121380
rect 166400 121120 166600 121380
rect 166900 121120 167100 121380
rect 167400 121120 167600 121380
rect 167900 121120 168100 121380
rect 168400 121120 168600 121380
rect 168900 121120 169100 121380
rect 169400 121120 169600 121380
rect 169900 121120 170100 121380
rect 170400 121120 170600 121380
rect 170900 121120 171100 121380
rect 171400 121120 171600 121380
rect 171900 121120 172100 121380
rect 172400 121120 172600 121380
rect 172900 121120 173100 121380
rect 173400 121120 173600 121380
rect 173900 121120 174100 121380
rect 174400 121120 174600 121380
rect 174900 121120 175100 121380
rect 175400 121120 175600 121380
rect 175900 121120 176100 121380
rect 176400 121120 176600 121380
rect 176900 121120 177100 121380
rect 177400 121120 177600 121380
rect 177900 121120 178100 121380
rect 178400 121120 178600 121380
rect 178900 121120 179100 121380
rect 179400 121120 179600 121380
rect 179900 121120 180100 121380
rect 180400 121120 180600 121380
rect 180900 121120 181100 121380
rect 181400 121120 181600 121380
rect 181900 121120 182100 121380
rect 182400 121120 182600 121380
rect 182900 121120 183100 121380
rect 183400 121120 183600 121380
rect 183900 121120 184000 121380
rect 162000 121100 162120 121120
rect 162380 121100 162620 121120
rect 162880 121100 163120 121120
rect 163380 121100 163620 121120
rect 163880 121100 164120 121120
rect 164380 121100 164620 121120
rect 164880 121100 165120 121120
rect 165380 121100 165620 121120
rect 165880 121100 166120 121120
rect 166380 121100 166620 121120
rect 166880 121100 167120 121120
rect 167380 121100 167620 121120
rect 167880 121100 168120 121120
rect 168380 121100 168620 121120
rect 168880 121100 169120 121120
rect 169380 121100 169620 121120
rect 169880 121100 170120 121120
rect 170380 121100 170620 121120
rect 170880 121100 171120 121120
rect 171380 121100 171620 121120
rect 171880 121100 172120 121120
rect 172380 121100 172620 121120
rect 172880 121100 173120 121120
rect 173380 121100 173620 121120
rect 173880 121100 174120 121120
rect 174380 121100 174620 121120
rect 174880 121100 175120 121120
rect 175380 121100 175620 121120
rect 175880 121100 176120 121120
rect 176380 121100 176620 121120
rect 176880 121100 177120 121120
rect 177380 121100 177620 121120
rect 177880 121100 178120 121120
rect 178380 121100 178620 121120
rect 178880 121100 179120 121120
rect 179380 121100 179620 121120
rect 179880 121100 180120 121120
rect 180380 121100 180620 121120
rect 180880 121100 181120 121120
rect 181380 121100 181620 121120
rect 181880 121100 182120 121120
rect 182380 121100 182620 121120
rect 182880 121100 183120 121120
rect 183380 121100 183620 121120
rect 183880 121100 184000 121120
rect 162000 120900 184000 121100
rect 162000 120880 162120 120900
rect 162380 120880 162620 120900
rect 162880 120880 163120 120900
rect 163380 120880 163620 120900
rect 163880 120880 164120 120900
rect 164380 120880 164620 120900
rect 164880 120880 165120 120900
rect 165380 120880 165620 120900
rect 165880 120880 166120 120900
rect 166380 120880 166620 120900
rect 166880 120880 167120 120900
rect 167380 120880 167620 120900
rect 167880 120880 168120 120900
rect 168380 120880 168620 120900
rect 168880 120880 169120 120900
rect 169380 120880 169620 120900
rect 169880 120880 170120 120900
rect 170380 120880 170620 120900
rect 170880 120880 171120 120900
rect 171380 120880 171620 120900
rect 171880 120880 172120 120900
rect 172380 120880 172620 120900
rect 172880 120880 173120 120900
rect 173380 120880 173620 120900
rect 173880 120880 174120 120900
rect 174380 120880 174620 120900
rect 174880 120880 175120 120900
rect 175380 120880 175620 120900
rect 175880 120880 176120 120900
rect 176380 120880 176620 120900
rect 176880 120880 177120 120900
rect 177380 120880 177620 120900
rect 177880 120880 178120 120900
rect 178380 120880 178620 120900
rect 178880 120880 179120 120900
rect 179380 120880 179620 120900
rect 179880 120880 180120 120900
rect 180380 120880 180620 120900
rect 180880 120880 181120 120900
rect 181380 120880 181620 120900
rect 181880 120880 182120 120900
rect 182380 120880 182620 120900
rect 182880 120880 183120 120900
rect 183380 120880 183620 120900
rect 183880 120880 184000 120900
rect 162000 120620 162100 120880
rect 162400 120620 162600 120880
rect 162900 120620 163100 120880
rect 163400 120620 163600 120880
rect 163900 120620 164100 120880
rect 164400 120620 164600 120880
rect 164900 120620 165100 120880
rect 165400 120620 165600 120880
rect 165900 120620 166100 120880
rect 166400 120620 166600 120880
rect 166900 120620 167100 120880
rect 167400 120620 167600 120880
rect 167900 120620 168100 120880
rect 168400 120620 168600 120880
rect 168900 120620 169100 120880
rect 169400 120620 169600 120880
rect 169900 120620 170100 120880
rect 170400 120620 170600 120880
rect 170900 120620 171100 120880
rect 171400 120620 171600 120880
rect 171900 120620 172100 120880
rect 172400 120620 172600 120880
rect 172900 120620 173100 120880
rect 173400 120620 173600 120880
rect 173900 120620 174100 120880
rect 174400 120620 174600 120880
rect 174900 120620 175100 120880
rect 175400 120620 175600 120880
rect 175900 120620 176100 120880
rect 176400 120620 176600 120880
rect 176900 120620 177100 120880
rect 177400 120620 177600 120880
rect 177900 120620 178100 120880
rect 178400 120620 178600 120880
rect 178900 120620 179100 120880
rect 179400 120620 179600 120880
rect 179900 120620 180100 120880
rect 180400 120620 180600 120880
rect 180900 120620 181100 120880
rect 181400 120620 181600 120880
rect 181900 120620 182100 120880
rect 182400 120620 182600 120880
rect 182900 120620 183100 120880
rect 183400 120620 183600 120880
rect 183900 120620 184000 120880
rect 162000 120600 162120 120620
rect 162380 120600 162620 120620
rect 162880 120600 163120 120620
rect 163380 120600 163620 120620
rect 163880 120600 164120 120620
rect 164380 120600 164620 120620
rect 164880 120600 165120 120620
rect 165380 120600 165620 120620
rect 165880 120600 166120 120620
rect 166380 120600 166620 120620
rect 166880 120600 167120 120620
rect 167380 120600 167620 120620
rect 167880 120600 168120 120620
rect 168380 120600 168620 120620
rect 168880 120600 169120 120620
rect 169380 120600 169620 120620
rect 169880 120600 170120 120620
rect 170380 120600 170620 120620
rect 170880 120600 171120 120620
rect 171380 120600 171620 120620
rect 171880 120600 172120 120620
rect 172380 120600 172620 120620
rect 172880 120600 173120 120620
rect 173380 120600 173620 120620
rect 173880 120600 174120 120620
rect 174380 120600 174620 120620
rect 174880 120600 175120 120620
rect 175380 120600 175620 120620
rect 175880 120600 176120 120620
rect 176380 120600 176620 120620
rect 176880 120600 177120 120620
rect 177380 120600 177620 120620
rect 177880 120600 178120 120620
rect 178380 120600 178620 120620
rect 178880 120600 179120 120620
rect 179380 120600 179620 120620
rect 179880 120600 180120 120620
rect 180380 120600 180620 120620
rect 180880 120600 181120 120620
rect 181380 120600 181620 120620
rect 181880 120600 182120 120620
rect 182380 120600 182620 120620
rect 182880 120600 183120 120620
rect 183380 120600 183620 120620
rect 183880 120600 184000 120620
rect 162000 120400 184000 120600
rect 162000 120380 162120 120400
rect 162380 120380 162620 120400
rect 162880 120380 163120 120400
rect 163380 120380 163620 120400
rect 163880 120380 164120 120400
rect 164380 120380 164620 120400
rect 164880 120380 165120 120400
rect 165380 120380 165620 120400
rect 165880 120380 166120 120400
rect 166380 120380 166620 120400
rect 166880 120380 167120 120400
rect 167380 120380 167620 120400
rect 167880 120380 168120 120400
rect 168380 120380 168620 120400
rect 168880 120380 169120 120400
rect 169380 120380 169620 120400
rect 169880 120380 170120 120400
rect 170380 120380 170620 120400
rect 170880 120380 171120 120400
rect 171380 120380 171620 120400
rect 171880 120380 172120 120400
rect 172380 120380 172620 120400
rect 172880 120380 173120 120400
rect 173380 120380 173620 120400
rect 173880 120380 174120 120400
rect 174380 120380 174620 120400
rect 174880 120380 175120 120400
rect 175380 120380 175620 120400
rect 175880 120380 176120 120400
rect 176380 120380 176620 120400
rect 176880 120380 177120 120400
rect 177380 120380 177620 120400
rect 177880 120380 178120 120400
rect 178380 120380 178620 120400
rect 178880 120380 179120 120400
rect 179380 120380 179620 120400
rect 179880 120380 180120 120400
rect 180380 120380 180620 120400
rect 180880 120380 181120 120400
rect 181380 120380 181620 120400
rect 181880 120380 182120 120400
rect 182380 120380 182620 120400
rect 182880 120380 183120 120400
rect 183380 120380 183620 120400
rect 183880 120380 184000 120400
rect 162000 120120 162100 120380
rect 162400 120120 162600 120380
rect 162900 120120 163100 120380
rect 163400 120120 163600 120380
rect 163900 120120 164100 120380
rect 164400 120120 164600 120380
rect 164900 120120 165100 120380
rect 165400 120120 165600 120380
rect 165900 120120 166100 120380
rect 166400 120120 166600 120380
rect 166900 120120 167100 120380
rect 167400 120120 167600 120380
rect 167900 120120 168100 120380
rect 168400 120120 168600 120380
rect 168900 120120 169100 120380
rect 169400 120120 169600 120380
rect 169900 120120 170100 120380
rect 170400 120120 170600 120380
rect 170900 120120 171100 120380
rect 171400 120120 171600 120380
rect 171900 120120 172100 120380
rect 172400 120120 172600 120380
rect 172900 120120 173100 120380
rect 173400 120120 173600 120380
rect 173900 120120 174100 120380
rect 174400 120120 174600 120380
rect 174900 120120 175100 120380
rect 175400 120120 175600 120380
rect 175900 120120 176100 120380
rect 176400 120120 176600 120380
rect 176900 120120 177100 120380
rect 177400 120120 177600 120380
rect 177900 120120 178100 120380
rect 178400 120120 178600 120380
rect 178900 120120 179100 120380
rect 179400 120120 179600 120380
rect 179900 120120 180100 120380
rect 180400 120120 180600 120380
rect 180900 120120 181100 120380
rect 181400 120120 181600 120380
rect 181900 120120 182100 120380
rect 182400 120120 182600 120380
rect 182900 120120 183100 120380
rect 183400 120120 183600 120380
rect 183900 120120 184000 120380
rect 162000 120100 162120 120120
rect 162380 120100 162620 120120
rect 162880 120100 163120 120120
rect 163380 120100 163620 120120
rect 163880 120100 164120 120120
rect 164380 120100 164620 120120
rect 164880 120100 165120 120120
rect 165380 120100 165620 120120
rect 165880 120100 166120 120120
rect 166380 120100 166620 120120
rect 166880 120100 167120 120120
rect 167380 120100 167620 120120
rect 167880 120100 168120 120120
rect 168380 120100 168620 120120
rect 168880 120100 169120 120120
rect 169380 120100 169620 120120
rect 169880 120100 170120 120120
rect 170380 120100 170620 120120
rect 170880 120100 171120 120120
rect 171380 120100 171620 120120
rect 171880 120100 172120 120120
rect 172380 120100 172620 120120
rect 172880 120100 173120 120120
rect 173380 120100 173620 120120
rect 173880 120100 174120 120120
rect 174380 120100 174620 120120
rect 174880 120100 175120 120120
rect 175380 120100 175620 120120
rect 175880 120100 176120 120120
rect 176380 120100 176620 120120
rect 176880 120100 177120 120120
rect 177380 120100 177620 120120
rect 177880 120100 178120 120120
rect 178380 120100 178620 120120
rect 178880 120100 179120 120120
rect 179380 120100 179620 120120
rect 179880 120100 180120 120120
rect 180380 120100 180620 120120
rect 180880 120100 181120 120120
rect 181380 120100 181620 120120
rect 181880 120100 182120 120120
rect 182380 120100 182620 120120
rect 182880 120100 183120 120120
rect 183380 120100 183620 120120
rect 183880 120100 184000 120120
rect 162000 119900 184000 120100
rect 162000 119880 162120 119900
rect 162380 119880 162620 119900
rect 162880 119880 163120 119900
rect 163380 119880 163620 119900
rect 163880 119880 164120 119900
rect 164380 119880 164620 119900
rect 164880 119880 165120 119900
rect 165380 119880 165620 119900
rect 165880 119880 166120 119900
rect 166380 119880 166620 119900
rect 166880 119880 167120 119900
rect 167380 119880 167620 119900
rect 167880 119880 168120 119900
rect 168380 119880 168620 119900
rect 168880 119880 169120 119900
rect 169380 119880 169620 119900
rect 169880 119880 170120 119900
rect 170380 119880 170620 119900
rect 170880 119880 171120 119900
rect 171380 119880 171620 119900
rect 171880 119880 172120 119900
rect 172380 119880 172620 119900
rect 172880 119880 173120 119900
rect 173380 119880 173620 119900
rect 173880 119880 174120 119900
rect 174380 119880 174620 119900
rect 174880 119880 175120 119900
rect 175380 119880 175620 119900
rect 175880 119880 176120 119900
rect 176380 119880 176620 119900
rect 176880 119880 177120 119900
rect 177380 119880 177620 119900
rect 177880 119880 178120 119900
rect 178380 119880 178620 119900
rect 178880 119880 179120 119900
rect 179380 119880 179620 119900
rect 179880 119880 180120 119900
rect 180380 119880 180620 119900
rect 180880 119880 181120 119900
rect 181380 119880 181620 119900
rect 181880 119880 182120 119900
rect 182380 119880 182620 119900
rect 182880 119880 183120 119900
rect 183380 119880 183620 119900
rect 183880 119880 184000 119900
rect 162000 119620 162100 119880
rect 162400 119620 162600 119880
rect 162900 119620 163100 119880
rect 163400 119620 163600 119880
rect 163900 119620 164100 119880
rect 164400 119620 164600 119880
rect 164900 119620 165100 119880
rect 165400 119620 165600 119880
rect 165900 119620 166100 119880
rect 166400 119620 166600 119880
rect 166900 119620 167100 119880
rect 167400 119620 167600 119880
rect 167900 119620 168100 119880
rect 168400 119620 168600 119880
rect 168900 119620 169100 119880
rect 169400 119620 169600 119880
rect 169900 119620 170100 119880
rect 170400 119620 170600 119880
rect 170900 119620 171100 119880
rect 171400 119620 171600 119880
rect 171900 119620 172100 119880
rect 172400 119620 172600 119880
rect 172900 119620 173100 119880
rect 173400 119620 173600 119880
rect 173900 119620 174100 119880
rect 174400 119620 174600 119880
rect 174900 119620 175100 119880
rect 175400 119620 175600 119880
rect 175900 119620 176100 119880
rect 176400 119620 176600 119880
rect 176900 119620 177100 119880
rect 177400 119620 177600 119880
rect 177900 119620 178100 119880
rect 178400 119620 178600 119880
rect 178900 119620 179100 119880
rect 179400 119620 179600 119880
rect 179900 119620 180100 119880
rect 180400 119620 180600 119880
rect 180900 119620 181100 119880
rect 181400 119620 181600 119880
rect 181900 119620 182100 119880
rect 182400 119620 182600 119880
rect 182900 119620 183100 119880
rect 183400 119620 183600 119880
rect 183900 119620 184000 119880
rect 162000 119600 162120 119620
rect 162380 119600 162620 119620
rect 162880 119600 163120 119620
rect 163380 119600 163620 119620
rect 163880 119600 164120 119620
rect 164380 119600 164620 119620
rect 164880 119600 165120 119620
rect 165380 119600 165620 119620
rect 165880 119600 166120 119620
rect 166380 119600 166620 119620
rect 166880 119600 167120 119620
rect 167380 119600 167620 119620
rect 167880 119600 168120 119620
rect 168380 119600 168620 119620
rect 168880 119600 169120 119620
rect 169380 119600 169620 119620
rect 169880 119600 170120 119620
rect 170380 119600 170620 119620
rect 170880 119600 171120 119620
rect 171380 119600 171620 119620
rect 171880 119600 172120 119620
rect 172380 119600 172620 119620
rect 172880 119600 173120 119620
rect 173380 119600 173620 119620
rect 173880 119600 174120 119620
rect 174380 119600 174620 119620
rect 174880 119600 175120 119620
rect 175380 119600 175620 119620
rect 175880 119600 176120 119620
rect 176380 119600 176620 119620
rect 176880 119600 177120 119620
rect 177380 119600 177620 119620
rect 177880 119600 178120 119620
rect 178380 119600 178620 119620
rect 178880 119600 179120 119620
rect 179380 119600 179620 119620
rect 179880 119600 180120 119620
rect 180380 119600 180620 119620
rect 180880 119600 181120 119620
rect 181380 119600 181620 119620
rect 181880 119600 182120 119620
rect 182380 119600 182620 119620
rect 182880 119600 183120 119620
rect 183380 119600 183620 119620
rect 183880 119600 184000 119620
rect 162000 119400 184000 119600
rect 162000 119380 162120 119400
rect 162380 119380 162620 119400
rect 162880 119380 163120 119400
rect 163380 119380 163620 119400
rect 163880 119380 164120 119400
rect 164380 119380 164620 119400
rect 164880 119380 165120 119400
rect 165380 119380 165620 119400
rect 165880 119380 166120 119400
rect 166380 119380 166620 119400
rect 166880 119380 167120 119400
rect 167380 119380 167620 119400
rect 167880 119380 168120 119400
rect 168380 119380 168620 119400
rect 168880 119380 169120 119400
rect 169380 119380 169620 119400
rect 169880 119380 170120 119400
rect 170380 119380 170620 119400
rect 170880 119380 171120 119400
rect 171380 119380 171620 119400
rect 171880 119380 172120 119400
rect 172380 119380 172620 119400
rect 172880 119380 173120 119400
rect 173380 119380 173620 119400
rect 173880 119380 174120 119400
rect 174380 119380 174620 119400
rect 174880 119380 175120 119400
rect 175380 119380 175620 119400
rect 175880 119380 176120 119400
rect 176380 119380 176620 119400
rect 176880 119380 177120 119400
rect 177380 119380 177620 119400
rect 177880 119380 178120 119400
rect 178380 119380 178620 119400
rect 178880 119380 179120 119400
rect 179380 119380 179620 119400
rect 179880 119380 180120 119400
rect 180380 119380 180620 119400
rect 180880 119380 181120 119400
rect 181380 119380 181620 119400
rect 181880 119380 182120 119400
rect 182380 119380 182620 119400
rect 182880 119380 183120 119400
rect 183380 119380 183620 119400
rect 183880 119380 184000 119400
rect 162000 119120 162100 119380
rect 162400 119120 162600 119380
rect 162900 119120 163100 119380
rect 163400 119120 163600 119380
rect 163900 119120 164100 119380
rect 164400 119120 164600 119380
rect 164900 119120 165100 119380
rect 165400 119120 165600 119380
rect 165900 119120 166100 119380
rect 166400 119120 166600 119380
rect 166900 119120 167100 119380
rect 167400 119120 167600 119380
rect 167900 119120 168100 119380
rect 168400 119120 168600 119380
rect 168900 119120 169100 119380
rect 169400 119120 169600 119380
rect 169900 119120 170100 119380
rect 170400 119120 170600 119380
rect 170900 119120 171100 119380
rect 171400 119120 171600 119380
rect 171900 119120 172100 119380
rect 172400 119120 172600 119380
rect 172900 119120 173100 119380
rect 173400 119120 173600 119380
rect 173900 119120 174100 119380
rect 174400 119120 174600 119380
rect 174900 119120 175100 119380
rect 175400 119120 175600 119380
rect 175900 119120 176100 119380
rect 176400 119120 176600 119380
rect 176900 119120 177100 119380
rect 177400 119120 177600 119380
rect 177900 119120 178100 119380
rect 178400 119120 178600 119380
rect 178900 119120 179100 119380
rect 179400 119120 179600 119380
rect 179900 119120 180100 119380
rect 180400 119120 180600 119380
rect 180900 119120 181100 119380
rect 181400 119120 181600 119380
rect 181900 119120 182100 119380
rect 182400 119120 182600 119380
rect 182900 119120 183100 119380
rect 183400 119120 183600 119380
rect 183900 119120 184000 119380
rect 162000 119100 162120 119120
rect 162380 119100 162620 119120
rect 162880 119100 163120 119120
rect 163380 119100 163620 119120
rect 163880 119100 164120 119120
rect 164380 119100 164620 119120
rect 164880 119100 165120 119120
rect 165380 119100 165620 119120
rect 165880 119100 166120 119120
rect 166380 119100 166620 119120
rect 166880 119100 167120 119120
rect 167380 119100 167620 119120
rect 167880 119100 168120 119120
rect 168380 119100 168620 119120
rect 168880 119100 169120 119120
rect 169380 119100 169620 119120
rect 169880 119100 170120 119120
rect 170380 119100 170620 119120
rect 170880 119100 171120 119120
rect 171380 119100 171620 119120
rect 171880 119100 172120 119120
rect 172380 119100 172620 119120
rect 172880 119100 173120 119120
rect 173380 119100 173620 119120
rect 173880 119100 174120 119120
rect 174380 119100 174620 119120
rect 174880 119100 175120 119120
rect 175380 119100 175620 119120
rect 175880 119100 176120 119120
rect 176380 119100 176620 119120
rect 176880 119100 177120 119120
rect 177380 119100 177620 119120
rect 177880 119100 178120 119120
rect 178380 119100 178620 119120
rect 178880 119100 179120 119120
rect 179380 119100 179620 119120
rect 179880 119100 180120 119120
rect 180380 119100 180620 119120
rect 180880 119100 181120 119120
rect 181380 119100 181620 119120
rect 181880 119100 182120 119120
rect 182380 119100 182620 119120
rect 182880 119100 183120 119120
rect 183380 119100 183620 119120
rect 183880 119100 184000 119120
rect 162000 118900 184000 119100
rect 162000 118880 162120 118900
rect 162380 118880 162620 118900
rect 162880 118880 163120 118900
rect 163380 118880 163620 118900
rect 163880 118880 164120 118900
rect 164380 118880 164620 118900
rect 164880 118880 165120 118900
rect 165380 118880 165620 118900
rect 165880 118880 166120 118900
rect 166380 118880 166620 118900
rect 166880 118880 167120 118900
rect 167380 118880 167620 118900
rect 167880 118880 168120 118900
rect 168380 118880 168620 118900
rect 168880 118880 169120 118900
rect 169380 118880 169620 118900
rect 169880 118880 170120 118900
rect 170380 118880 170620 118900
rect 170880 118880 171120 118900
rect 171380 118880 171620 118900
rect 171880 118880 172120 118900
rect 172380 118880 172620 118900
rect 172880 118880 173120 118900
rect 173380 118880 173620 118900
rect 173880 118880 174120 118900
rect 174380 118880 174620 118900
rect 174880 118880 175120 118900
rect 175380 118880 175620 118900
rect 175880 118880 176120 118900
rect 176380 118880 176620 118900
rect 176880 118880 177120 118900
rect 177380 118880 177620 118900
rect 177880 118880 178120 118900
rect 178380 118880 178620 118900
rect 178880 118880 179120 118900
rect 179380 118880 179620 118900
rect 179880 118880 180120 118900
rect 180380 118880 180620 118900
rect 180880 118880 181120 118900
rect 181380 118880 181620 118900
rect 181880 118880 182120 118900
rect 182380 118880 182620 118900
rect 182880 118880 183120 118900
rect 183380 118880 183620 118900
rect 183880 118880 184000 118900
rect 162000 118620 162100 118880
rect 162400 118620 162600 118880
rect 162900 118620 163100 118880
rect 163400 118620 163600 118880
rect 163900 118620 164100 118880
rect 164400 118620 164600 118880
rect 164900 118620 165100 118880
rect 165400 118620 165600 118880
rect 165900 118620 166100 118880
rect 166400 118620 166600 118880
rect 166900 118620 167100 118880
rect 167400 118620 167600 118880
rect 167900 118620 168100 118880
rect 168400 118620 168600 118880
rect 168900 118620 169100 118880
rect 169400 118620 169600 118880
rect 169900 118620 170100 118880
rect 170400 118620 170600 118880
rect 170900 118620 171100 118880
rect 171400 118620 171600 118880
rect 171900 118620 172100 118880
rect 172400 118620 172600 118880
rect 172900 118620 173100 118880
rect 173400 118620 173600 118880
rect 173900 118620 174100 118880
rect 174400 118620 174600 118880
rect 174900 118620 175100 118880
rect 175400 118620 175600 118880
rect 175900 118620 176100 118880
rect 176400 118620 176600 118880
rect 176900 118620 177100 118880
rect 177400 118620 177600 118880
rect 177900 118620 178100 118880
rect 178400 118620 178600 118880
rect 178900 118620 179100 118880
rect 179400 118620 179600 118880
rect 179900 118620 180100 118880
rect 180400 118620 180600 118880
rect 180900 118620 181100 118880
rect 181400 118620 181600 118880
rect 181900 118620 182100 118880
rect 182400 118620 182600 118880
rect 182900 118620 183100 118880
rect 183400 118620 183600 118880
rect 183900 118620 184000 118880
rect 162000 118600 162120 118620
rect 162380 118600 162620 118620
rect 162880 118600 163120 118620
rect 163380 118600 163620 118620
rect 163880 118600 164120 118620
rect 164380 118600 164620 118620
rect 164880 118600 165120 118620
rect 165380 118600 165620 118620
rect 165880 118600 166120 118620
rect 166380 118600 166620 118620
rect 166880 118600 167120 118620
rect 167380 118600 167620 118620
rect 167880 118600 168120 118620
rect 168380 118600 168620 118620
rect 168880 118600 169120 118620
rect 169380 118600 169620 118620
rect 169880 118600 170120 118620
rect 170380 118600 170620 118620
rect 170880 118600 171120 118620
rect 171380 118600 171620 118620
rect 171880 118600 172120 118620
rect 172380 118600 172620 118620
rect 172880 118600 173120 118620
rect 173380 118600 173620 118620
rect 173880 118600 174120 118620
rect 174380 118600 174620 118620
rect 174880 118600 175120 118620
rect 175380 118600 175620 118620
rect 175880 118600 176120 118620
rect 176380 118600 176620 118620
rect 176880 118600 177120 118620
rect 177380 118600 177620 118620
rect 177880 118600 178120 118620
rect 178380 118600 178620 118620
rect 178880 118600 179120 118620
rect 179380 118600 179620 118620
rect 179880 118600 180120 118620
rect 180380 118600 180620 118620
rect 180880 118600 181120 118620
rect 181380 118600 181620 118620
rect 181880 118600 182120 118620
rect 182380 118600 182620 118620
rect 182880 118600 183120 118620
rect 183380 118600 183620 118620
rect 183880 118600 184000 118620
rect 162000 118400 184000 118600
rect 162000 118380 162120 118400
rect 162380 118380 162620 118400
rect 162880 118380 163120 118400
rect 163380 118380 163620 118400
rect 163880 118380 164120 118400
rect 164380 118380 164620 118400
rect 164880 118380 165120 118400
rect 165380 118380 165620 118400
rect 165880 118380 166120 118400
rect 166380 118380 166620 118400
rect 166880 118380 167120 118400
rect 167380 118380 167620 118400
rect 167880 118380 168120 118400
rect 168380 118380 168620 118400
rect 168880 118380 169120 118400
rect 169380 118380 169620 118400
rect 169880 118380 170120 118400
rect 170380 118380 170620 118400
rect 170880 118380 171120 118400
rect 171380 118380 171620 118400
rect 171880 118380 172120 118400
rect 172380 118380 172620 118400
rect 172880 118380 173120 118400
rect 173380 118380 173620 118400
rect 173880 118380 174120 118400
rect 174380 118380 174620 118400
rect 174880 118380 175120 118400
rect 175380 118380 175620 118400
rect 175880 118380 176120 118400
rect 176380 118380 176620 118400
rect 176880 118380 177120 118400
rect 177380 118380 177620 118400
rect 177880 118380 178120 118400
rect 178380 118380 178620 118400
rect 178880 118380 179120 118400
rect 179380 118380 179620 118400
rect 179880 118380 180120 118400
rect 180380 118380 180620 118400
rect 180880 118380 181120 118400
rect 181380 118380 181620 118400
rect 181880 118380 182120 118400
rect 182380 118380 182620 118400
rect 182880 118380 183120 118400
rect 183380 118380 183620 118400
rect 183880 118380 184000 118400
rect 162000 118120 162100 118380
rect 162400 118120 162600 118380
rect 162900 118120 163100 118380
rect 163400 118120 163600 118380
rect 163900 118120 164100 118380
rect 164400 118120 164600 118380
rect 164900 118120 165100 118380
rect 165400 118120 165600 118380
rect 165900 118120 166100 118380
rect 166400 118120 166600 118380
rect 166900 118120 167100 118380
rect 167400 118120 167600 118380
rect 167900 118120 168100 118380
rect 168400 118120 168600 118380
rect 168900 118120 169100 118380
rect 169400 118120 169600 118380
rect 169900 118120 170100 118380
rect 170400 118120 170600 118380
rect 170900 118120 171100 118380
rect 171400 118120 171600 118380
rect 171900 118120 172100 118380
rect 172400 118120 172600 118380
rect 172900 118120 173100 118380
rect 173400 118120 173600 118380
rect 173900 118120 174100 118380
rect 174400 118120 174600 118380
rect 174900 118120 175100 118380
rect 175400 118120 175600 118380
rect 175900 118120 176100 118380
rect 176400 118120 176600 118380
rect 176900 118120 177100 118380
rect 177400 118120 177600 118380
rect 177900 118120 178100 118380
rect 178400 118120 178600 118380
rect 178900 118120 179100 118380
rect 179400 118120 179600 118380
rect 179900 118120 180100 118380
rect 180400 118120 180600 118380
rect 180900 118120 181100 118380
rect 181400 118120 181600 118380
rect 181900 118120 182100 118380
rect 182400 118120 182600 118380
rect 182900 118120 183100 118380
rect 183400 118120 183600 118380
rect 183900 118120 184000 118380
rect 162000 118100 162120 118120
rect 162380 118100 162620 118120
rect 162880 118100 163120 118120
rect 163380 118100 163620 118120
rect 163880 118100 164120 118120
rect 164380 118100 164620 118120
rect 164880 118100 165120 118120
rect 165380 118100 165620 118120
rect 165880 118100 166120 118120
rect 166380 118100 166620 118120
rect 166880 118100 167120 118120
rect 167380 118100 167620 118120
rect 167880 118100 168120 118120
rect 168380 118100 168620 118120
rect 168880 118100 169120 118120
rect 169380 118100 169620 118120
rect 169880 118100 170120 118120
rect 170380 118100 170620 118120
rect 170880 118100 171120 118120
rect 171380 118100 171620 118120
rect 171880 118100 172120 118120
rect 172380 118100 172620 118120
rect 172880 118100 173120 118120
rect 173380 118100 173620 118120
rect 173880 118100 174120 118120
rect 174380 118100 174620 118120
rect 174880 118100 175120 118120
rect 175380 118100 175620 118120
rect 175880 118100 176120 118120
rect 176380 118100 176620 118120
rect 176880 118100 177120 118120
rect 177380 118100 177620 118120
rect 177880 118100 178120 118120
rect 178380 118100 178620 118120
rect 178880 118100 179120 118120
rect 179380 118100 179620 118120
rect 179880 118100 180120 118120
rect 180380 118100 180620 118120
rect 180880 118100 181120 118120
rect 181380 118100 181620 118120
rect 181880 118100 182120 118120
rect 182380 118100 182620 118120
rect 182880 118100 183120 118120
rect 183380 118100 183620 118120
rect 183880 118100 184000 118120
rect 162000 117900 184000 118100
rect 162000 117880 162120 117900
rect 162380 117880 162620 117900
rect 162880 117880 163120 117900
rect 163380 117880 163620 117900
rect 163880 117880 164120 117900
rect 164380 117880 164620 117900
rect 164880 117880 165120 117900
rect 165380 117880 165620 117900
rect 165880 117880 166120 117900
rect 166380 117880 166620 117900
rect 166880 117880 167120 117900
rect 167380 117880 167620 117900
rect 167880 117880 168120 117900
rect 168380 117880 168620 117900
rect 168880 117880 169120 117900
rect 169380 117880 169620 117900
rect 169880 117880 170120 117900
rect 170380 117880 170620 117900
rect 170880 117880 171120 117900
rect 171380 117880 171620 117900
rect 171880 117880 172120 117900
rect 172380 117880 172620 117900
rect 172880 117880 173120 117900
rect 173380 117880 173620 117900
rect 173880 117880 174120 117900
rect 174380 117880 174620 117900
rect 174880 117880 175120 117900
rect 175380 117880 175620 117900
rect 175880 117880 176120 117900
rect 176380 117880 176620 117900
rect 176880 117880 177120 117900
rect 177380 117880 177620 117900
rect 177880 117880 178120 117900
rect 178380 117880 178620 117900
rect 178880 117880 179120 117900
rect 179380 117880 179620 117900
rect 179880 117880 180120 117900
rect 180380 117880 180620 117900
rect 180880 117880 181120 117900
rect 181380 117880 181620 117900
rect 181880 117880 182120 117900
rect 182380 117880 182620 117900
rect 182880 117880 183120 117900
rect 183380 117880 183620 117900
rect 183880 117880 184000 117900
rect 162000 117620 162100 117880
rect 162400 117620 162600 117880
rect 162900 117620 163100 117880
rect 163400 117620 163600 117880
rect 163900 117620 164100 117880
rect 164400 117620 164600 117880
rect 164900 117620 165100 117880
rect 165400 117620 165600 117880
rect 165900 117620 166100 117880
rect 166400 117620 166600 117880
rect 166900 117620 167100 117880
rect 167400 117620 167600 117880
rect 167900 117620 168100 117880
rect 168400 117620 168600 117880
rect 168900 117620 169100 117880
rect 169400 117620 169600 117880
rect 169900 117620 170100 117880
rect 170400 117620 170600 117880
rect 170900 117620 171100 117880
rect 171400 117620 171600 117880
rect 171900 117620 172100 117880
rect 172400 117620 172600 117880
rect 172900 117620 173100 117880
rect 173400 117620 173600 117880
rect 173900 117620 174100 117880
rect 174400 117620 174600 117880
rect 174900 117620 175100 117880
rect 175400 117620 175600 117880
rect 175900 117620 176100 117880
rect 176400 117620 176600 117880
rect 176900 117620 177100 117880
rect 177400 117620 177600 117880
rect 177900 117620 178100 117880
rect 178400 117620 178600 117880
rect 178900 117620 179100 117880
rect 179400 117620 179600 117880
rect 179900 117620 180100 117880
rect 180400 117620 180600 117880
rect 180900 117620 181100 117880
rect 181400 117620 181600 117880
rect 181900 117620 182100 117880
rect 182400 117620 182600 117880
rect 182900 117620 183100 117880
rect 183400 117620 183600 117880
rect 183900 117620 184000 117880
rect 162000 117600 162120 117620
rect 162380 117600 162620 117620
rect 162880 117600 163120 117620
rect 163380 117600 163620 117620
rect 163880 117600 164120 117620
rect 164380 117600 164620 117620
rect 164880 117600 165120 117620
rect 165380 117600 165620 117620
rect 165880 117600 166120 117620
rect 166380 117600 166620 117620
rect 166880 117600 167120 117620
rect 167380 117600 167620 117620
rect 167880 117600 168120 117620
rect 168380 117600 168620 117620
rect 168880 117600 169120 117620
rect 169380 117600 169620 117620
rect 169880 117600 170120 117620
rect 170380 117600 170620 117620
rect 170880 117600 171120 117620
rect 171380 117600 171620 117620
rect 171880 117600 172120 117620
rect 172380 117600 172620 117620
rect 172880 117600 173120 117620
rect 173380 117600 173620 117620
rect 173880 117600 174120 117620
rect 174380 117600 174620 117620
rect 174880 117600 175120 117620
rect 175380 117600 175620 117620
rect 175880 117600 176120 117620
rect 176380 117600 176620 117620
rect 176880 117600 177120 117620
rect 177380 117600 177620 117620
rect 177880 117600 178120 117620
rect 178380 117600 178620 117620
rect 178880 117600 179120 117620
rect 179380 117600 179620 117620
rect 179880 117600 180120 117620
rect 180380 117600 180620 117620
rect 180880 117600 181120 117620
rect 181380 117600 181620 117620
rect 181880 117600 182120 117620
rect 182380 117600 182620 117620
rect 182880 117600 183120 117620
rect 183380 117600 183620 117620
rect 183880 117600 184000 117620
rect 162000 117400 184000 117600
rect 162000 117380 162120 117400
rect 162380 117380 162620 117400
rect 162880 117380 163120 117400
rect 163380 117380 163620 117400
rect 163880 117380 164120 117400
rect 164380 117380 164620 117400
rect 164880 117380 165120 117400
rect 165380 117380 165620 117400
rect 165880 117380 166120 117400
rect 166380 117380 166620 117400
rect 166880 117380 167120 117400
rect 167380 117380 167620 117400
rect 167880 117380 168120 117400
rect 168380 117380 168620 117400
rect 168880 117380 169120 117400
rect 169380 117380 169620 117400
rect 169880 117380 170120 117400
rect 170380 117380 170620 117400
rect 170880 117380 171120 117400
rect 171380 117380 171620 117400
rect 171880 117380 172120 117400
rect 172380 117380 172620 117400
rect 172880 117380 173120 117400
rect 173380 117380 173620 117400
rect 173880 117380 174120 117400
rect 174380 117380 174620 117400
rect 174880 117380 175120 117400
rect 175380 117380 175620 117400
rect 175880 117380 176120 117400
rect 176380 117380 176620 117400
rect 176880 117380 177120 117400
rect 177380 117380 177620 117400
rect 177880 117380 178120 117400
rect 178380 117380 178620 117400
rect 178880 117380 179120 117400
rect 179380 117380 179620 117400
rect 179880 117380 180120 117400
rect 180380 117380 180620 117400
rect 180880 117380 181120 117400
rect 181380 117380 181620 117400
rect 181880 117380 182120 117400
rect 182380 117380 182620 117400
rect 182880 117380 183120 117400
rect 183380 117380 183620 117400
rect 183880 117380 184000 117400
rect 162000 117120 162100 117380
rect 162400 117120 162600 117380
rect 162900 117120 163100 117380
rect 163400 117120 163600 117380
rect 163900 117120 164100 117380
rect 164400 117120 164600 117380
rect 164900 117120 165100 117380
rect 165400 117120 165600 117380
rect 165900 117120 166100 117380
rect 166400 117120 166600 117380
rect 166900 117120 167100 117380
rect 167400 117120 167600 117380
rect 167900 117120 168100 117380
rect 168400 117120 168600 117380
rect 168900 117120 169100 117380
rect 169400 117120 169600 117380
rect 169900 117120 170100 117380
rect 170400 117120 170600 117380
rect 170900 117120 171100 117380
rect 171400 117120 171600 117380
rect 171900 117120 172100 117380
rect 172400 117120 172600 117380
rect 172900 117120 173100 117380
rect 173400 117120 173600 117380
rect 173900 117120 174100 117380
rect 174400 117120 174600 117380
rect 174900 117120 175100 117380
rect 175400 117120 175600 117380
rect 175900 117120 176100 117380
rect 176400 117120 176600 117380
rect 176900 117120 177100 117380
rect 177400 117120 177600 117380
rect 177900 117120 178100 117380
rect 178400 117120 178600 117380
rect 178900 117120 179100 117380
rect 179400 117120 179600 117380
rect 179900 117120 180100 117380
rect 180400 117120 180600 117380
rect 180900 117120 181100 117380
rect 181400 117120 181600 117380
rect 181900 117120 182100 117380
rect 182400 117120 182600 117380
rect 182900 117120 183100 117380
rect 183400 117120 183600 117380
rect 183900 117120 184000 117380
rect 162000 117100 162120 117120
rect 162380 117100 162620 117120
rect 162880 117100 163120 117120
rect 163380 117100 163620 117120
rect 163880 117100 164120 117120
rect 164380 117100 164620 117120
rect 164880 117100 165120 117120
rect 165380 117100 165620 117120
rect 165880 117100 166120 117120
rect 166380 117100 166620 117120
rect 166880 117100 167120 117120
rect 167380 117100 167620 117120
rect 167880 117100 168120 117120
rect 168380 117100 168620 117120
rect 168880 117100 169120 117120
rect 169380 117100 169620 117120
rect 169880 117100 170120 117120
rect 170380 117100 170620 117120
rect 170880 117100 171120 117120
rect 171380 117100 171620 117120
rect 171880 117100 172120 117120
rect 172380 117100 172620 117120
rect 172880 117100 173120 117120
rect 173380 117100 173620 117120
rect 173880 117100 174120 117120
rect 174380 117100 174620 117120
rect 174880 117100 175120 117120
rect 175380 117100 175620 117120
rect 175880 117100 176120 117120
rect 176380 117100 176620 117120
rect 176880 117100 177120 117120
rect 177380 117100 177620 117120
rect 177880 117100 178120 117120
rect 178380 117100 178620 117120
rect 178880 117100 179120 117120
rect 179380 117100 179620 117120
rect 179880 117100 180120 117120
rect 180380 117100 180620 117120
rect 180880 117100 181120 117120
rect 181380 117100 181620 117120
rect 181880 117100 182120 117120
rect 182380 117100 182620 117120
rect 182880 117100 183120 117120
rect 183380 117100 183620 117120
rect 183880 117100 184000 117120
rect 162000 116900 184000 117100
rect 162000 116880 162120 116900
rect 162380 116880 162620 116900
rect 162880 116880 163120 116900
rect 163380 116880 163620 116900
rect 163880 116880 164120 116900
rect 164380 116880 164620 116900
rect 164880 116880 165120 116900
rect 165380 116880 165620 116900
rect 165880 116880 166120 116900
rect 166380 116880 166620 116900
rect 166880 116880 167120 116900
rect 167380 116880 167620 116900
rect 167880 116880 168120 116900
rect 168380 116880 168620 116900
rect 168880 116880 169120 116900
rect 169380 116880 169620 116900
rect 169880 116880 170120 116900
rect 170380 116880 170620 116900
rect 170880 116880 171120 116900
rect 171380 116880 171620 116900
rect 171880 116880 172120 116900
rect 172380 116880 172620 116900
rect 172880 116880 173120 116900
rect 173380 116880 173620 116900
rect 173880 116880 174120 116900
rect 174380 116880 174620 116900
rect 174880 116880 175120 116900
rect 175380 116880 175620 116900
rect 175880 116880 176120 116900
rect 176380 116880 176620 116900
rect 176880 116880 177120 116900
rect 177380 116880 177620 116900
rect 177880 116880 178120 116900
rect 178380 116880 178620 116900
rect 178880 116880 179120 116900
rect 179380 116880 179620 116900
rect 179880 116880 180120 116900
rect 180380 116880 180620 116900
rect 180880 116880 181120 116900
rect 181380 116880 181620 116900
rect 181880 116880 182120 116900
rect 182380 116880 182620 116900
rect 182880 116880 183120 116900
rect 183380 116880 183620 116900
rect 183880 116880 184000 116900
rect 162000 116620 162100 116880
rect 162400 116620 162600 116880
rect 162900 116620 163100 116880
rect 163400 116620 163600 116880
rect 163900 116620 164100 116880
rect 164400 116620 164600 116880
rect 164900 116620 165100 116880
rect 165400 116620 165600 116880
rect 165900 116620 166100 116880
rect 166400 116620 166600 116880
rect 166900 116620 167100 116880
rect 167400 116620 167600 116880
rect 167900 116620 168100 116880
rect 168400 116620 168600 116880
rect 168900 116620 169100 116880
rect 169400 116620 169600 116880
rect 169900 116620 170100 116880
rect 170400 116620 170600 116880
rect 170900 116620 171100 116880
rect 171400 116620 171600 116880
rect 171900 116620 172100 116880
rect 172400 116620 172600 116880
rect 172900 116620 173100 116880
rect 173400 116620 173600 116880
rect 173900 116620 174100 116880
rect 174400 116620 174600 116880
rect 174900 116620 175100 116880
rect 175400 116620 175600 116880
rect 175900 116620 176100 116880
rect 176400 116620 176600 116880
rect 176900 116620 177100 116880
rect 177400 116620 177600 116880
rect 177900 116620 178100 116880
rect 178400 116620 178600 116880
rect 178900 116620 179100 116880
rect 179400 116620 179600 116880
rect 179900 116620 180100 116880
rect 180400 116620 180600 116880
rect 180900 116620 181100 116880
rect 181400 116620 181600 116880
rect 181900 116620 182100 116880
rect 182400 116620 182600 116880
rect 182900 116620 183100 116880
rect 183400 116620 183600 116880
rect 183900 116620 184000 116880
rect 162000 116600 162120 116620
rect 162380 116600 162620 116620
rect 162880 116600 163120 116620
rect 163380 116600 163620 116620
rect 163880 116600 164120 116620
rect 164380 116600 164620 116620
rect 164880 116600 165120 116620
rect 165380 116600 165620 116620
rect 165880 116600 166120 116620
rect 166380 116600 166620 116620
rect 166880 116600 167120 116620
rect 167380 116600 167620 116620
rect 167880 116600 168120 116620
rect 168380 116600 168620 116620
rect 168880 116600 169120 116620
rect 169380 116600 169620 116620
rect 169880 116600 170120 116620
rect 170380 116600 170620 116620
rect 170880 116600 171120 116620
rect 171380 116600 171620 116620
rect 171880 116600 172120 116620
rect 172380 116600 172620 116620
rect 172880 116600 173120 116620
rect 173380 116600 173620 116620
rect 173880 116600 174120 116620
rect 174380 116600 174620 116620
rect 174880 116600 175120 116620
rect 175380 116600 175620 116620
rect 175880 116600 176120 116620
rect 176380 116600 176620 116620
rect 176880 116600 177120 116620
rect 177380 116600 177620 116620
rect 177880 116600 178120 116620
rect 178380 116600 178620 116620
rect 178880 116600 179120 116620
rect 179380 116600 179620 116620
rect 179880 116600 180120 116620
rect 180380 116600 180620 116620
rect 180880 116600 181120 116620
rect 181380 116600 181620 116620
rect 181880 116600 182120 116620
rect 182380 116600 182620 116620
rect 182880 116600 183120 116620
rect 183380 116600 183620 116620
rect 183880 116600 184000 116620
rect 162000 116400 184000 116600
rect 162000 116380 162120 116400
rect 162380 116380 162620 116400
rect 162880 116380 163120 116400
rect 163380 116380 163620 116400
rect 163880 116380 164120 116400
rect 164380 116380 164620 116400
rect 164880 116380 165120 116400
rect 165380 116380 165620 116400
rect 165880 116380 166120 116400
rect 166380 116380 166620 116400
rect 166880 116380 167120 116400
rect 167380 116380 167620 116400
rect 167880 116380 168120 116400
rect 168380 116380 168620 116400
rect 168880 116380 169120 116400
rect 169380 116380 169620 116400
rect 169880 116380 170120 116400
rect 170380 116380 170620 116400
rect 170880 116380 171120 116400
rect 171380 116380 171620 116400
rect 171880 116380 172120 116400
rect 172380 116380 172620 116400
rect 172880 116380 173120 116400
rect 173380 116380 173620 116400
rect 173880 116380 174120 116400
rect 174380 116380 174620 116400
rect 174880 116380 175120 116400
rect 175380 116380 175620 116400
rect 175880 116380 176120 116400
rect 176380 116380 176620 116400
rect 176880 116380 177120 116400
rect 177380 116380 177620 116400
rect 177880 116380 178120 116400
rect 178380 116380 178620 116400
rect 178880 116380 179120 116400
rect 179380 116380 179620 116400
rect 179880 116380 180120 116400
rect 180380 116380 180620 116400
rect 180880 116380 181120 116400
rect 181380 116380 181620 116400
rect 181880 116380 182120 116400
rect 182380 116380 182620 116400
rect 182880 116380 183120 116400
rect 183380 116380 183620 116400
rect 183880 116380 184000 116400
rect 162000 116120 162100 116380
rect 162400 116120 162600 116380
rect 162900 116120 163100 116380
rect 163400 116120 163600 116380
rect 163900 116120 164100 116380
rect 164400 116120 164600 116380
rect 164900 116120 165100 116380
rect 165400 116120 165600 116380
rect 165900 116120 166100 116380
rect 166400 116120 166600 116380
rect 166900 116120 167100 116380
rect 167400 116120 167600 116380
rect 167900 116120 168100 116380
rect 168400 116120 168600 116380
rect 168900 116120 169100 116380
rect 169400 116120 169600 116380
rect 169900 116120 170100 116380
rect 170400 116120 170600 116380
rect 170900 116120 171100 116380
rect 171400 116120 171600 116380
rect 171900 116120 172100 116380
rect 172400 116120 172600 116380
rect 172900 116120 173100 116380
rect 173400 116120 173600 116380
rect 173900 116120 174100 116380
rect 174400 116120 174600 116380
rect 174900 116120 175100 116380
rect 175400 116120 175600 116380
rect 175900 116120 176100 116380
rect 176400 116120 176600 116380
rect 176900 116120 177100 116380
rect 177400 116120 177600 116380
rect 177900 116120 178100 116380
rect 178400 116120 178600 116380
rect 178900 116120 179100 116380
rect 179400 116120 179600 116380
rect 179900 116120 180100 116380
rect 180400 116120 180600 116380
rect 180900 116120 181100 116380
rect 181400 116120 181600 116380
rect 181900 116120 182100 116380
rect 182400 116120 182600 116380
rect 182900 116120 183100 116380
rect 183400 116120 183600 116380
rect 183900 116120 184000 116380
rect 162000 116100 162120 116120
rect 162380 116100 162620 116120
rect 162880 116100 163120 116120
rect 163380 116100 163620 116120
rect 163880 116100 164120 116120
rect 164380 116100 164620 116120
rect 164880 116100 165120 116120
rect 165380 116100 165620 116120
rect 165880 116100 166120 116120
rect 166380 116100 166620 116120
rect 166880 116100 167120 116120
rect 167380 116100 167620 116120
rect 167880 116100 168120 116120
rect 168380 116100 168620 116120
rect 168880 116100 169120 116120
rect 169380 116100 169620 116120
rect 169880 116100 170120 116120
rect 170380 116100 170620 116120
rect 170880 116100 171120 116120
rect 171380 116100 171620 116120
rect 171880 116100 172120 116120
rect 172380 116100 172620 116120
rect 172880 116100 173120 116120
rect 173380 116100 173620 116120
rect 173880 116100 174120 116120
rect 174380 116100 174620 116120
rect 174880 116100 175120 116120
rect 175380 116100 175620 116120
rect 175880 116100 176120 116120
rect 176380 116100 176620 116120
rect 176880 116100 177120 116120
rect 177380 116100 177620 116120
rect 177880 116100 178120 116120
rect 178380 116100 178620 116120
rect 178880 116100 179120 116120
rect 179380 116100 179620 116120
rect 179880 116100 180120 116120
rect 180380 116100 180620 116120
rect 180880 116100 181120 116120
rect 181380 116100 181620 116120
rect 181880 116100 182120 116120
rect 182380 116100 182620 116120
rect 182880 116100 183120 116120
rect 183380 116100 183620 116120
rect 183880 116100 184000 116120
rect 162000 115900 184000 116100
rect 162000 115880 162120 115900
rect 162380 115880 162620 115900
rect 162880 115880 163120 115900
rect 163380 115880 163620 115900
rect 163880 115880 164120 115900
rect 164380 115880 164620 115900
rect 164880 115880 165120 115900
rect 165380 115880 165620 115900
rect 165880 115880 166120 115900
rect 166380 115880 166620 115900
rect 166880 115880 167120 115900
rect 167380 115880 167620 115900
rect 167880 115880 168120 115900
rect 168380 115880 168620 115900
rect 168880 115880 169120 115900
rect 169380 115880 169620 115900
rect 169880 115880 170120 115900
rect 170380 115880 170620 115900
rect 170880 115880 171120 115900
rect 171380 115880 171620 115900
rect 171880 115880 172120 115900
rect 172380 115880 172620 115900
rect 172880 115880 173120 115900
rect 173380 115880 173620 115900
rect 173880 115880 174120 115900
rect 174380 115880 174620 115900
rect 174880 115880 175120 115900
rect 175380 115880 175620 115900
rect 175880 115880 176120 115900
rect 176380 115880 176620 115900
rect 176880 115880 177120 115900
rect 177380 115880 177620 115900
rect 177880 115880 178120 115900
rect 178380 115880 178620 115900
rect 178880 115880 179120 115900
rect 179380 115880 179620 115900
rect 179880 115880 180120 115900
rect 180380 115880 180620 115900
rect 180880 115880 181120 115900
rect 181380 115880 181620 115900
rect 181880 115880 182120 115900
rect 182380 115880 182620 115900
rect 182880 115880 183120 115900
rect 183380 115880 183620 115900
rect 183880 115880 184000 115900
rect 162000 115620 162100 115880
rect 162400 115620 162600 115880
rect 162900 115620 163100 115880
rect 163400 115620 163600 115880
rect 163900 115620 164100 115880
rect 164400 115620 164600 115880
rect 164900 115620 165100 115880
rect 165400 115620 165600 115880
rect 165900 115620 166100 115880
rect 166400 115620 166600 115880
rect 166900 115620 167100 115880
rect 167400 115620 167600 115880
rect 167900 115620 168100 115880
rect 168400 115620 168600 115880
rect 168900 115620 169100 115880
rect 169400 115620 169600 115880
rect 169900 115620 170100 115880
rect 170400 115620 170600 115880
rect 170900 115620 171100 115880
rect 171400 115620 171600 115880
rect 171900 115620 172100 115880
rect 172400 115620 172600 115880
rect 172900 115620 173100 115880
rect 173400 115620 173600 115880
rect 173900 115620 174100 115880
rect 174400 115620 174600 115880
rect 174900 115620 175100 115880
rect 175400 115620 175600 115880
rect 175900 115620 176100 115880
rect 176400 115620 176600 115880
rect 176900 115620 177100 115880
rect 177400 115620 177600 115880
rect 177900 115620 178100 115880
rect 178400 115620 178600 115880
rect 178900 115620 179100 115880
rect 179400 115620 179600 115880
rect 179900 115620 180100 115880
rect 180400 115620 180600 115880
rect 180900 115620 181100 115880
rect 181400 115620 181600 115880
rect 181900 115620 182100 115880
rect 182400 115620 182600 115880
rect 182900 115620 183100 115880
rect 183400 115620 183600 115880
rect 183900 115620 184000 115880
rect 162000 115600 162120 115620
rect 162380 115600 162620 115620
rect 162880 115600 163120 115620
rect 163380 115600 163620 115620
rect 163880 115600 164120 115620
rect 164380 115600 164620 115620
rect 164880 115600 165120 115620
rect 165380 115600 165620 115620
rect 165880 115600 166120 115620
rect 166380 115600 166620 115620
rect 166880 115600 167120 115620
rect 167380 115600 167620 115620
rect 167880 115600 168120 115620
rect 168380 115600 168620 115620
rect 168880 115600 169120 115620
rect 169380 115600 169620 115620
rect 169880 115600 170120 115620
rect 170380 115600 170620 115620
rect 170880 115600 171120 115620
rect 171380 115600 171620 115620
rect 171880 115600 172120 115620
rect 172380 115600 172620 115620
rect 172880 115600 173120 115620
rect 173380 115600 173620 115620
rect 173880 115600 174120 115620
rect 174380 115600 174620 115620
rect 174880 115600 175120 115620
rect 175380 115600 175620 115620
rect 175880 115600 176120 115620
rect 176380 115600 176620 115620
rect 176880 115600 177120 115620
rect 177380 115600 177620 115620
rect 177880 115600 178120 115620
rect 178380 115600 178620 115620
rect 178880 115600 179120 115620
rect 179380 115600 179620 115620
rect 179880 115600 180120 115620
rect 180380 115600 180620 115620
rect 180880 115600 181120 115620
rect 181380 115600 181620 115620
rect 181880 115600 182120 115620
rect 182380 115600 182620 115620
rect 182880 115600 183120 115620
rect 183380 115600 183620 115620
rect 183880 115600 184000 115620
rect 162000 115400 184000 115600
rect 162000 115380 162120 115400
rect 162380 115380 162620 115400
rect 162880 115380 163120 115400
rect 163380 115380 163620 115400
rect 163880 115380 164120 115400
rect 164380 115380 164620 115400
rect 164880 115380 165120 115400
rect 165380 115380 165620 115400
rect 165880 115380 166120 115400
rect 166380 115380 166620 115400
rect 166880 115380 167120 115400
rect 167380 115380 167620 115400
rect 167880 115380 168120 115400
rect 168380 115380 168620 115400
rect 168880 115380 169120 115400
rect 169380 115380 169620 115400
rect 169880 115380 170120 115400
rect 170380 115380 170620 115400
rect 170880 115380 171120 115400
rect 171380 115380 171620 115400
rect 171880 115380 172120 115400
rect 172380 115380 172620 115400
rect 172880 115380 173120 115400
rect 173380 115380 173620 115400
rect 173880 115380 174120 115400
rect 174380 115380 174620 115400
rect 174880 115380 175120 115400
rect 175380 115380 175620 115400
rect 175880 115380 176120 115400
rect 176380 115380 176620 115400
rect 176880 115380 177120 115400
rect 177380 115380 177620 115400
rect 177880 115380 178120 115400
rect 178380 115380 178620 115400
rect 178880 115380 179120 115400
rect 179380 115380 179620 115400
rect 179880 115380 180120 115400
rect 180380 115380 180620 115400
rect 180880 115380 181120 115400
rect 181380 115380 181620 115400
rect 181880 115380 182120 115400
rect 182380 115380 182620 115400
rect 182880 115380 183120 115400
rect 183380 115380 183620 115400
rect 183880 115380 184000 115400
rect 162000 115120 162100 115380
rect 162400 115120 162600 115380
rect 162900 115120 163100 115380
rect 163400 115120 163600 115380
rect 163900 115120 164100 115380
rect 164400 115120 164600 115380
rect 164900 115120 165100 115380
rect 165400 115120 165600 115380
rect 165900 115120 166100 115380
rect 166400 115120 166600 115380
rect 166900 115120 167100 115380
rect 167400 115120 167600 115380
rect 167900 115120 168100 115380
rect 168400 115120 168600 115380
rect 168900 115120 169100 115380
rect 169400 115120 169600 115380
rect 169900 115120 170100 115380
rect 170400 115120 170600 115380
rect 170900 115120 171100 115380
rect 171400 115120 171600 115380
rect 171900 115120 172100 115380
rect 172400 115120 172600 115380
rect 172900 115120 173100 115380
rect 173400 115120 173600 115380
rect 173900 115120 174100 115380
rect 174400 115120 174600 115380
rect 174900 115120 175100 115380
rect 175400 115120 175600 115380
rect 175900 115120 176100 115380
rect 176400 115120 176600 115380
rect 176900 115120 177100 115380
rect 177400 115120 177600 115380
rect 177900 115120 178100 115380
rect 178400 115120 178600 115380
rect 178900 115120 179100 115380
rect 179400 115120 179600 115380
rect 179900 115120 180100 115380
rect 180400 115120 180600 115380
rect 180900 115120 181100 115380
rect 181400 115120 181600 115380
rect 181900 115120 182100 115380
rect 182400 115120 182600 115380
rect 182900 115120 183100 115380
rect 183400 115120 183600 115380
rect 183900 115120 184000 115380
rect 162000 115100 162120 115120
rect 162380 115100 162620 115120
rect 162880 115100 163120 115120
rect 163380 115100 163620 115120
rect 163880 115100 164120 115120
rect 164380 115100 164620 115120
rect 164880 115100 165120 115120
rect 165380 115100 165620 115120
rect 165880 115100 166120 115120
rect 166380 115100 166620 115120
rect 166880 115100 167120 115120
rect 167380 115100 167620 115120
rect 167880 115100 168120 115120
rect 168380 115100 168620 115120
rect 168880 115100 169120 115120
rect 169380 115100 169620 115120
rect 169880 115100 170120 115120
rect 170380 115100 170620 115120
rect 170880 115100 171120 115120
rect 171380 115100 171620 115120
rect 171880 115100 172120 115120
rect 172380 115100 172620 115120
rect 172880 115100 173120 115120
rect 173380 115100 173620 115120
rect 173880 115100 174120 115120
rect 174380 115100 174620 115120
rect 174880 115100 175120 115120
rect 175380 115100 175620 115120
rect 175880 115100 176120 115120
rect 176380 115100 176620 115120
rect 176880 115100 177120 115120
rect 177380 115100 177620 115120
rect 177880 115100 178120 115120
rect 178380 115100 178620 115120
rect 178880 115100 179120 115120
rect 179380 115100 179620 115120
rect 179880 115100 180120 115120
rect 180380 115100 180620 115120
rect 180880 115100 181120 115120
rect 181380 115100 181620 115120
rect 181880 115100 182120 115120
rect 182380 115100 182620 115120
rect 182880 115100 183120 115120
rect 183380 115100 183620 115120
rect 183880 115100 184000 115120
rect 162000 114900 184000 115100
rect 162000 114880 162120 114900
rect 162380 114880 162620 114900
rect 162880 114880 163120 114900
rect 163380 114880 163620 114900
rect 163880 114880 164120 114900
rect 164380 114880 164620 114900
rect 164880 114880 165120 114900
rect 165380 114880 165620 114900
rect 165880 114880 166120 114900
rect 166380 114880 166620 114900
rect 166880 114880 167120 114900
rect 167380 114880 167620 114900
rect 167880 114880 168120 114900
rect 168380 114880 168620 114900
rect 168880 114880 169120 114900
rect 169380 114880 169620 114900
rect 169880 114880 170120 114900
rect 170380 114880 170620 114900
rect 170880 114880 171120 114900
rect 171380 114880 171620 114900
rect 171880 114880 172120 114900
rect 172380 114880 172620 114900
rect 172880 114880 173120 114900
rect 173380 114880 173620 114900
rect 173880 114880 174120 114900
rect 174380 114880 174620 114900
rect 174880 114880 175120 114900
rect 175380 114880 175620 114900
rect 175880 114880 176120 114900
rect 176380 114880 176620 114900
rect 176880 114880 177120 114900
rect 177380 114880 177620 114900
rect 177880 114880 178120 114900
rect 178380 114880 178620 114900
rect 178880 114880 179120 114900
rect 179380 114880 179620 114900
rect 179880 114880 180120 114900
rect 180380 114880 180620 114900
rect 180880 114880 181120 114900
rect 181380 114880 181620 114900
rect 181880 114880 182120 114900
rect 182380 114880 182620 114900
rect 182880 114880 183120 114900
rect 183380 114880 183620 114900
rect 183880 114880 184000 114900
rect 162000 114620 162100 114880
rect 162400 114620 162600 114880
rect 162900 114620 163100 114880
rect 163400 114620 163600 114880
rect 163900 114620 164100 114880
rect 164400 114620 164600 114880
rect 164900 114620 165100 114880
rect 165400 114620 165600 114880
rect 165900 114620 166100 114880
rect 166400 114620 166600 114880
rect 166900 114620 167100 114880
rect 167400 114620 167600 114880
rect 167900 114620 168100 114880
rect 168400 114620 168600 114880
rect 168900 114620 169100 114880
rect 169400 114620 169600 114880
rect 169900 114620 170100 114880
rect 170400 114620 170600 114880
rect 170900 114620 171100 114880
rect 171400 114620 171600 114880
rect 171900 114620 172100 114880
rect 172400 114620 172600 114880
rect 172900 114620 173100 114880
rect 173400 114620 173600 114880
rect 173900 114620 174100 114880
rect 174400 114620 174600 114880
rect 174900 114620 175100 114880
rect 175400 114620 175600 114880
rect 175900 114620 176100 114880
rect 176400 114620 176600 114880
rect 176900 114620 177100 114880
rect 177400 114620 177600 114880
rect 177900 114620 178100 114880
rect 178400 114620 178600 114880
rect 178900 114620 179100 114880
rect 179400 114620 179600 114880
rect 179900 114620 180100 114880
rect 180400 114620 180600 114880
rect 180900 114620 181100 114880
rect 181400 114620 181600 114880
rect 181900 114620 182100 114880
rect 182400 114620 182600 114880
rect 182900 114620 183100 114880
rect 183400 114620 183600 114880
rect 183900 114620 184000 114880
rect 162000 114600 162120 114620
rect 162380 114600 162620 114620
rect 162880 114600 163120 114620
rect 163380 114600 163620 114620
rect 163880 114600 164120 114620
rect 164380 114600 164620 114620
rect 164880 114600 165120 114620
rect 165380 114600 165620 114620
rect 165880 114600 166120 114620
rect 166380 114600 166620 114620
rect 166880 114600 167120 114620
rect 167380 114600 167620 114620
rect 167880 114600 168120 114620
rect 168380 114600 168620 114620
rect 168880 114600 169120 114620
rect 169380 114600 169620 114620
rect 169880 114600 170120 114620
rect 170380 114600 170620 114620
rect 170880 114600 171120 114620
rect 171380 114600 171620 114620
rect 171880 114600 172120 114620
rect 172380 114600 172620 114620
rect 172880 114600 173120 114620
rect 173380 114600 173620 114620
rect 173880 114600 174120 114620
rect 174380 114600 174620 114620
rect 174880 114600 175120 114620
rect 175380 114600 175620 114620
rect 175880 114600 176120 114620
rect 176380 114600 176620 114620
rect 176880 114600 177120 114620
rect 177380 114600 177620 114620
rect 177880 114600 178120 114620
rect 178380 114600 178620 114620
rect 178880 114600 179120 114620
rect 179380 114600 179620 114620
rect 179880 114600 180120 114620
rect 180380 114600 180620 114620
rect 180880 114600 181120 114620
rect 181380 114600 181620 114620
rect 181880 114600 182120 114620
rect 182380 114600 182620 114620
rect 182880 114600 183120 114620
rect 183380 114600 183620 114620
rect 183880 114600 184000 114620
rect 162000 114400 184000 114600
rect 162000 114380 162120 114400
rect 162380 114380 162620 114400
rect 162880 114380 163120 114400
rect 163380 114380 163620 114400
rect 163880 114380 164120 114400
rect 164380 114380 164620 114400
rect 164880 114380 165120 114400
rect 165380 114380 165620 114400
rect 165880 114380 166120 114400
rect 166380 114380 166620 114400
rect 166880 114380 167120 114400
rect 167380 114380 167620 114400
rect 167880 114380 168120 114400
rect 168380 114380 168620 114400
rect 168880 114380 169120 114400
rect 169380 114380 169620 114400
rect 169880 114380 170120 114400
rect 170380 114380 170620 114400
rect 170880 114380 171120 114400
rect 171380 114380 171620 114400
rect 171880 114380 172120 114400
rect 172380 114380 172620 114400
rect 172880 114380 173120 114400
rect 173380 114380 173620 114400
rect 173880 114380 174120 114400
rect 174380 114380 174620 114400
rect 174880 114380 175120 114400
rect 175380 114380 175620 114400
rect 175880 114380 176120 114400
rect 176380 114380 176620 114400
rect 176880 114380 177120 114400
rect 177380 114380 177620 114400
rect 177880 114380 178120 114400
rect 178380 114380 178620 114400
rect 178880 114380 179120 114400
rect 179380 114380 179620 114400
rect 179880 114380 180120 114400
rect 180380 114380 180620 114400
rect 180880 114380 181120 114400
rect 181380 114380 181620 114400
rect 181880 114380 182120 114400
rect 182380 114380 182620 114400
rect 182880 114380 183120 114400
rect 183380 114380 183620 114400
rect 183880 114380 184000 114400
rect 162000 114120 162100 114380
rect 162400 114120 162600 114380
rect 162900 114120 163100 114380
rect 163400 114120 163600 114380
rect 163900 114120 164100 114380
rect 164400 114120 164600 114380
rect 164900 114120 165100 114380
rect 165400 114120 165600 114380
rect 165900 114120 166100 114380
rect 166400 114120 166600 114380
rect 166900 114120 167100 114380
rect 167400 114120 167600 114380
rect 167900 114120 168100 114380
rect 168400 114120 168600 114380
rect 168900 114120 169100 114380
rect 169400 114120 169600 114380
rect 169900 114120 170100 114380
rect 170400 114120 170600 114380
rect 170900 114120 171100 114380
rect 171400 114120 171600 114380
rect 171900 114120 172100 114380
rect 172400 114120 172600 114380
rect 172900 114120 173100 114380
rect 173400 114120 173600 114380
rect 173900 114120 174100 114380
rect 174400 114120 174600 114380
rect 174900 114120 175100 114380
rect 175400 114120 175600 114380
rect 175900 114120 176100 114380
rect 176400 114120 176600 114380
rect 176900 114120 177100 114380
rect 177400 114120 177600 114380
rect 177900 114120 178100 114380
rect 178400 114120 178600 114380
rect 178900 114120 179100 114380
rect 179400 114120 179600 114380
rect 179900 114120 180100 114380
rect 180400 114120 180600 114380
rect 180900 114120 181100 114380
rect 181400 114120 181600 114380
rect 181900 114120 182100 114380
rect 182400 114120 182600 114380
rect 182900 114120 183100 114380
rect 183400 114120 183600 114380
rect 183900 114120 184000 114380
rect 162000 114100 162120 114120
rect 162380 114100 162620 114120
rect 162880 114100 163120 114120
rect 163380 114100 163620 114120
rect 163880 114100 164120 114120
rect 164380 114100 164620 114120
rect 164880 114100 165120 114120
rect 165380 114100 165620 114120
rect 165880 114100 166120 114120
rect 166380 114100 166620 114120
rect 166880 114100 167120 114120
rect 167380 114100 167620 114120
rect 167880 114100 168120 114120
rect 168380 114100 168620 114120
rect 168880 114100 169120 114120
rect 169380 114100 169620 114120
rect 169880 114100 170120 114120
rect 170380 114100 170620 114120
rect 170880 114100 171120 114120
rect 171380 114100 171620 114120
rect 171880 114100 172120 114120
rect 172380 114100 172620 114120
rect 172880 114100 173120 114120
rect 173380 114100 173620 114120
rect 173880 114100 174120 114120
rect 174380 114100 174620 114120
rect 174880 114100 175120 114120
rect 175380 114100 175620 114120
rect 175880 114100 176120 114120
rect 176380 114100 176620 114120
rect 176880 114100 177120 114120
rect 177380 114100 177620 114120
rect 177880 114100 178120 114120
rect 178380 114100 178620 114120
rect 178880 114100 179120 114120
rect 179380 114100 179620 114120
rect 179880 114100 180120 114120
rect 180380 114100 180620 114120
rect 180880 114100 181120 114120
rect 181380 114100 181620 114120
rect 181880 114100 182120 114120
rect 182380 114100 182620 114120
rect 182880 114100 183120 114120
rect 183380 114100 183620 114120
rect 183880 114100 184000 114120
rect 162000 114000 184000 114100
rect 214000 121900 232000 122000
rect 214000 121880 214120 121900
rect 214380 121880 214620 121900
rect 214880 121880 215120 121900
rect 215380 121880 215620 121900
rect 215880 121880 216120 121900
rect 216380 121880 216620 121900
rect 216880 121880 217120 121900
rect 217380 121880 217620 121900
rect 217880 121880 218120 121900
rect 218380 121880 218620 121900
rect 218880 121880 219120 121900
rect 219380 121880 219620 121900
rect 219880 121880 220120 121900
rect 220380 121880 220620 121900
rect 220880 121880 221120 121900
rect 221380 121880 221620 121900
rect 221880 121880 222120 121900
rect 222380 121880 222620 121900
rect 222880 121880 223120 121900
rect 223380 121880 223620 121900
rect 223880 121880 224120 121900
rect 224380 121880 224620 121900
rect 224880 121880 225120 121900
rect 225380 121880 225620 121900
rect 225880 121880 226120 121900
rect 226380 121880 226620 121900
rect 226880 121880 227120 121900
rect 227380 121880 227620 121900
rect 227880 121880 228120 121900
rect 228380 121880 228620 121900
rect 228880 121880 229120 121900
rect 229380 121880 229620 121900
rect 229880 121880 230120 121900
rect 230380 121880 230620 121900
rect 230880 121880 231120 121900
rect 231380 121880 231620 121900
rect 231880 121880 232000 121900
rect 214000 121620 214100 121880
rect 214400 121620 214600 121880
rect 214900 121620 215100 121880
rect 215400 121620 215600 121880
rect 215900 121620 216100 121880
rect 216400 121620 216600 121880
rect 216900 121620 217100 121880
rect 217400 121620 217600 121880
rect 217900 121620 218100 121880
rect 218400 121620 218600 121880
rect 218900 121620 219100 121880
rect 219400 121620 219600 121880
rect 219900 121620 220100 121880
rect 220400 121620 220600 121880
rect 220900 121620 221100 121880
rect 221400 121620 221600 121880
rect 221900 121620 222100 121880
rect 222400 121620 222600 121880
rect 222900 121620 223100 121880
rect 223400 121620 223600 121880
rect 223900 121620 224100 121880
rect 224400 121620 224600 121880
rect 224900 121620 225100 121880
rect 225400 121620 225600 121880
rect 225900 121620 226100 121880
rect 226400 121620 226600 121880
rect 226900 121620 227100 121880
rect 227400 121620 227600 121880
rect 227900 121620 228100 121880
rect 228400 121620 228600 121880
rect 228900 121620 229100 121880
rect 229400 121620 229600 121880
rect 229900 121620 230100 121880
rect 230400 121620 230600 121880
rect 230900 121620 231100 121880
rect 231400 121620 231600 121880
rect 231900 121620 232000 121880
rect 214000 121600 214120 121620
rect 214380 121600 214620 121620
rect 214880 121600 215120 121620
rect 215380 121600 215620 121620
rect 215880 121600 216120 121620
rect 216380 121600 216620 121620
rect 216880 121600 217120 121620
rect 217380 121600 217620 121620
rect 217880 121600 218120 121620
rect 218380 121600 218620 121620
rect 218880 121600 219120 121620
rect 219380 121600 219620 121620
rect 219880 121600 220120 121620
rect 220380 121600 220620 121620
rect 220880 121600 221120 121620
rect 221380 121600 221620 121620
rect 221880 121600 222120 121620
rect 222380 121600 222620 121620
rect 222880 121600 223120 121620
rect 223380 121600 223620 121620
rect 223880 121600 224120 121620
rect 224380 121600 224620 121620
rect 224880 121600 225120 121620
rect 225380 121600 225620 121620
rect 225880 121600 226120 121620
rect 226380 121600 226620 121620
rect 226880 121600 227120 121620
rect 227380 121600 227620 121620
rect 227880 121600 228120 121620
rect 228380 121600 228620 121620
rect 228880 121600 229120 121620
rect 229380 121600 229620 121620
rect 229880 121600 230120 121620
rect 230380 121600 230620 121620
rect 230880 121600 231120 121620
rect 231380 121600 231620 121620
rect 231880 121600 232000 121620
rect 214000 121400 232000 121600
rect 214000 121380 214120 121400
rect 214380 121380 214620 121400
rect 214880 121380 215120 121400
rect 215380 121380 215620 121400
rect 215880 121380 216120 121400
rect 216380 121380 216620 121400
rect 216880 121380 217120 121400
rect 217380 121380 217620 121400
rect 217880 121380 218120 121400
rect 218380 121380 218620 121400
rect 218880 121380 219120 121400
rect 219380 121380 219620 121400
rect 219880 121380 220120 121400
rect 220380 121380 220620 121400
rect 220880 121380 221120 121400
rect 221380 121380 221620 121400
rect 221880 121380 222120 121400
rect 222380 121380 222620 121400
rect 222880 121380 223120 121400
rect 223380 121380 223620 121400
rect 223880 121380 224120 121400
rect 224380 121380 224620 121400
rect 224880 121380 225120 121400
rect 225380 121380 225620 121400
rect 225880 121380 226120 121400
rect 226380 121380 226620 121400
rect 226880 121380 227120 121400
rect 227380 121380 227620 121400
rect 227880 121380 228120 121400
rect 228380 121380 228620 121400
rect 228880 121380 229120 121400
rect 229380 121380 229620 121400
rect 229880 121380 230120 121400
rect 230380 121380 230620 121400
rect 230880 121380 231120 121400
rect 231380 121380 231620 121400
rect 231880 121380 232000 121400
rect 214000 121120 214100 121380
rect 214400 121120 214600 121380
rect 214900 121120 215100 121380
rect 215400 121120 215600 121380
rect 215900 121120 216100 121380
rect 216400 121120 216600 121380
rect 216900 121120 217100 121380
rect 217400 121120 217600 121380
rect 217900 121120 218100 121380
rect 218400 121120 218600 121380
rect 218900 121120 219100 121380
rect 219400 121120 219600 121380
rect 219900 121120 220100 121380
rect 220400 121120 220600 121380
rect 220900 121120 221100 121380
rect 221400 121120 221600 121380
rect 221900 121120 222100 121380
rect 222400 121120 222600 121380
rect 222900 121120 223100 121380
rect 223400 121120 223600 121380
rect 223900 121120 224100 121380
rect 224400 121120 224600 121380
rect 224900 121120 225100 121380
rect 225400 121120 225600 121380
rect 225900 121120 226100 121380
rect 226400 121120 226600 121380
rect 226900 121120 227100 121380
rect 227400 121120 227600 121380
rect 227900 121120 228100 121380
rect 228400 121120 228600 121380
rect 228900 121120 229100 121380
rect 229400 121120 229600 121380
rect 229900 121120 230100 121380
rect 230400 121120 230600 121380
rect 230900 121120 231100 121380
rect 231400 121120 231600 121380
rect 231900 121120 232000 121380
rect 214000 121100 214120 121120
rect 214380 121100 214620 121120
rect 214880 121100 215120 121120
rect 215380 121100 215620 121120
rect 215880 121100 216120 121120
rect 216380 121100 216620 121120
rect 216880 121100 217120 121120
rect 217380 121100 217620 121120
rect 217880 121100 218120 121120
rect 218380 121100 218620 121120
rect 218880 121100 219120 121120
rect 219380 121100 219620 121120
rect 219880 121100 220120 121120
rect 220380 121100 220620 121120
rect 220880 121100 221120 121120
rect 221380 121100 221620 121120
rect 221880 121100 222120 121120
rect 222380 121100 222620 121120
rect 222880 121100 223120 121120
rect 223380 121100 223620 121120
rect 223880 121100 224120 121120
rect 224380 121100 224620 121120
rect 224880 121100 225120 121120
rect 225380 121100 225620 121120
rect 225880 121100 226120 121120
rect 226380 121100 226620 121120
rect 226880 121100 227120 121120
rect 227380 121100 227620 121120
rect 227880 121100 228120 121120
rect 228380 121100 228620 121120
rect 228880 121100 229120 121120
rect 229380 121100 229620 121120
rect 229880 121100 230120 121120
rect 230380 121100 230620 121120
rect 230880 121100 231120 121120
rect 231380 121100 231620 121120
rect 231880 121100 232000 121120
rect 214000 120900 232000 121100
rect 214000 120880 214120 120900
rect 214380 120880 214620 120900
rect 214880 120880 215120 120900
rect 215380 120880 215620 120900
rect 215880 120880 216120 120900
rect 216380 120880 216620 120900
rect 216880 120880 217120 120900
rect 217380 120880 217620 120900
rect 217880 120880 218120 120900
rect 218380 120880 218620 120900
rect 218880 120880 219120 120900
rect 219380 120880 219620 120900
rect 219880 120880 220120 120900
rect 220380 120880 220620 120900
rect 220880 120880 221120 120900
rect 221380 120880 221620 120900
rect 221880 120880 222120 120900
rect 222380 120880 222620 120900
rect 222880 120880 223120 120900
rect 223380 120880 223620 120900
rect 223880 120880 224120 120900
rect 224380 120880 224620 120900
rect 224880 120880 225120 120900
rect 225380 120880 225620 120900
rect 225880 120880 226120 120900
rect 226380 120880 226620 120900
rect 226880 120880 227120 120900
rect 227380 120880 227620 120900
rect 227880 120880 228120 120900
rect 228380 120880 228620 120900
rect 228880 120880 229120 120900
rect 229380 120880 229620 120900
rect 229880 120880 230120 120900
rect 230380 120880 230620 120900
rect 230880 120880 231120 120900
rect 231380 120880 231620 120900
rect 231880 120880 232000 120900
rect 214000 120620 214100 120880
rect 214400 120620 214600 120880
rect 214900 120620 215100 120880
rect 215400 120620 215600 120880
rect 215900 120620 216100 120880
rect 216400 120620 216600 120880
rect 216900 120620 217100 120880
rect 217400 120620 217600 120880
rect 217900 120620 218100 120880
rect 218400 120620 218600 120880
rect 218900 120620 219100 120880
rect 219400 120620 219600 120880
rect 219900 120620 220100 120880
rect 220400 120620 220600 120880
rect 220900 120620 221100 120880
rect 221400 120620 221600 120880
rect 221900 120620 222100 120880
rect 222400 120620 222600 120880
rect 222900 120620 223100 120880
rect 223400 120620 223600 120880
rect 223900 120620 224100 120880
rect 224400 120620 224600 120880
rect 224900 120620 225100 120880
rect 225400 120620 225600 120880
rect 225900 120620 226100 120880
rect 226400 120620 226600 120880
rect 226900 120620 227100 120880
rect 227400 120620 227600 120880
rect 227900 120620 228100 120880
rect 228400 120620 228600 120880
rect 228900 120620 229100 120880
rect 229400 120620 229600 120880
rect 229900 120620 230100 120880
rect 230400 120620 230600 120880
rect 230900 120620 231100 120880
rect 231400 120620 231600 120880
rect 231900 120620 232000 120880
rect 214000 120600 214120 120620
rect 214380 120600 214620 120620
rect 214880 120600 215120 120620
rect 215380 120600 215620 120620
rect 215880 120600 216120 120620
rect 216380 120600 216620 120620
rect 216880 120600 217120 120620
rect 217380 120600 217620 120620
rect 217880 120600 218120 120620
rect 218380 120600 218620 120620
rect 218880 120600 219120 120620
rect 219380 120600 219620 120620
rect 219880 120600 220120 120620
rect 220380 120600 220620 120620
rect 220880 120600 221120 120620
rect 221380 120600 221620 120620
rect 221880 120600 222120 120620
rect 222380 120600 222620 120620
rect 222880 120600 223120 120620
rect 223380 120600 223620 120620
rect 223880 120600 224120 120620
rect 224380 120600 224620 120620
rect 224880 120600 225120 120620
rect 225380 120600 225620 120620
rect 225880 120600 226120 120620
rect 226380 120600 226620 120620
rect 226880 120600 227120 120620
rect 227380 120600 227620 120620
rect 227880 120600 228120 120620
rect 228380 120600 228620 120620
rect 228880 120600 229120 120620
rect 229380 120600 229620 120620
rect 229880 120600 230120 120620
rect 230380 120600 230620 120620
rect 230880 120600 231120 120620
rect 231380 120600 231620 120620
rect 231880 120600 232000 120620
rect 214000 120400 232000 120600
rect 214000 120380 214120 120400
rect 214380 120380 214620 120400
rect 214880 120380 215120 120400
rect 215380 120380 215620 120400
rect 215880 120380 216120 120400
rect 216380 120380 216620 120400
rect 216880 120380 217120 120400
rect 217380 120380 217620 120400
rect 217880 120380 218120 120400
rect 218380 120380 218620 120400
rect 218880 120380 219120 120400
rect 219380 120380 219620 120400
rect 219880 120380 220120 120400
rect 220380 120380 220620 120400
rect 220880 120380 221120 120400
rect 221380 120380 221620 120400
rect 221880 120380 222120 120400
rect 222380 120380 222620 120400
rect 222880 120380 223120 120400
rect 223380 120380 223620 120400
rect 223880 120380 224120 120400
rect 224380 120380 224620 120400
rect 224880 120380 225120 120400
rect 225380 120380 225620 120400
rect 225880 120380 226120 120400
rect 226380 120380 226620 120400
rect 226880 120380 227120 120400
rect 227380 120380 227620 120400
rect 227880 120380 228120 120400
rect 228380 120380 228620 120400
rect 228880 120380 229120 120400
rect 229380 120380 229620 120400
rect 229880 120380 230120 120400
rect 230380 120380 230620 120400
rect 230880 120380 231120 120400
rect 231380 120380 231620 120400
rect 231880 120380 232000 120400
rect 214000 120120 214100 120380
rect 214400 120120 214600 120380
rect 214900 120120 215100 120380
rect 215400 120120 215600 120380
rect 215900 120120 216100 120380
rect 216400 120120 216600 120380
rect 216900 120120 217100 120380
rect 217400 120120 217600 120380
rect 217900 120120 218100 120380
rect 218400 120120 218600 120380
rect 218900 120120 219100 120380
rect 219400 120120 219600 120380
rect 219900 120120 220100 120380
rect 220400 120120 220600 120380
rect 220900 120120 221100 120380
rect 221400 120120 221600 120380
rect 221900 120120 222100 120380
rect 222400 120120 222600 120380
rect 222900 120120 223100 120380
rect 223400 120120 223600 120380
rect 223900 120120 224100 120380
rect 224400 120120 224600 120380
rect 224900 120120 225100 120380
rect 225400 120120 225600 120380
rect 225900 120120 226100 120380
rect 226400 120120 226600 120380
rect 226900 120120 227100 120380
rect 227400 120120 227600 120380
rect 227900 120120 228100 120380
rect 228400 120120 228600 120380
rect 228900 120120 229100 120380
rect 229400 120120 229600 120380
rect 229900 120120 230100 120380
rect 230400 120120 230600 120380
rect 230900 120120 231100 120380
rect 231400 120120 231600 120380
rect 231900 120120 232000 120380
rect 214000 120100 214120 120120
rect 214380 120100 214620 120120
rect 214880 120100 215120 120120
rect 215380 120100 215620 120120
rect 215880 120100 216120 120120
rect 216380 120100 216620 120120
rect 216880 120100 217120 120120
rect 217380 120100 217620 120120
rect 217880 120100 218120 120120
rect 218380 120100 218620 120120
rect 218880 120100 219120 120120
rect 219380 120100 219620 120120
rect 219880 120100 220120 120120
rect 220380 120100 220620 120120
rect 220880 120100 221120 120120
rect 221380 120100 221620 120120
rect 221880 120100 222120 120120
rect 222380 120100 222620 120120
rect 222880 120100 223120 120120
rect 223380 120100 223620 120120
rect 223880 120100 224120 120120
rect 224380 120100 224620 120120
rect 224880 120100 225120 120120
rect 225380 120100 225620 120120
rect 225880 120100 226120 120120
rect 226380 120100 226620 120120
rect 226880 120100 227120 120120
rect 227380 120100 227620 120120
rect 227880 120100 228120 120120
rect 228380 120100 228620 120120
rect 228880 120100 229120 120120
rect 229380 120100 229620 120120
rect 229880 120100 230120 120120
rect 230380 120100 230620 120120
rect 230880 120100 231120 120120
rect 231380 120100 231620 120120
rect 231880 120100 232000 120120
rect 214000 119900 232000 120100
rect 214000 119880 214120 119900
rect 214380 119880 214620 119900
rect 214880 119880 215120 119900
rect 215380 119880 215620 119900
rect 215880 119880 216120 119900
rect 216380 119880 216620 119900
rect 216880 119880 217120 119900
rect 217380 119880 217620 119900
rect 217880 119880 218120 119900
rect 218380 119880 218620 119900
rect 218880 119880 219120 119900
rect 219380 119880 219620 119900
rect 219880 119880 220120 119900
rect 220380 119880 220620 119900
rect 220880 119880 221120 119900
rect 221380 119880 221620 119900
rect 221880 119880 222120 119900
rect 222380 119880 222620 119900
rect 222880 119880 223120 119900
rect 223380 119880 223620 119900
rect 223880 119880 224120 119900
rect 224380 119880 224620 119900
rect 224880 119880 225120 119900
rect 225380 119880 225620 119900
rect 225880 119880 226120 119900
rect 226380 119880 226620 119900
rect 226880 119880 227120 119900
rect 227380 119880 227620 119900
rect 227880 119880 228120 119900
rect 228380 119880 228620 119900
rect 228880 119880 229120 119900
rect 229380 119880 229620 119900
rect 229880 119880 230120 119900
rect 230380 119880 230620 119900
rect 230880 119880 231120 119900
rect 231380 119880 231620 119900
rect 231880 119880 232000 119900
rect 214000 119620 214100 119880
rect 214400 119620 214600 119880
rect 214900 119620 215100 119880
rect 215400 119620 215600 119880
rect 215900 119620 216100 119880
rect 216400 119620 216600 119880
rect 216900 119620 217100 119880
rect 217400 119620 217600 119880
rect 217900 119620 218100 119880
rect 218400 119620 218600 119880
rect 218900 119620 219100 119880
rect 219400 119620 219600 119880
rect 219900 119620 220100 119880
rect 220400 119620 220600 119880
rect 220900 119620 221100 119880
rect 221400 119620 221600 119880
rect 221900 119620 222100 119880
rect 222400 119620 222600 119880
rect 222900 119620 223100 119880
rect 223400 119620 223600 119880
rect 223900 119620 224100 119880
rect 224400 119620 224600 119880
rect 224900 119620 225100 119880
rect 225400 119620 225600 119880
rect 225900 119620 226100 119880
rect 226400 119620 226600 119880
rect 226900 119620 227100 119880
rect 227400 119620 227600 119880
rect 227900 119620 228100 119880
rect 228400 119620 228600 119880
rect 228900 119620 229100 119880
rect 229400 119620 229600 119880
rect 229900 119620 230100 119880
rect 230400 119620 230600 119880
rect 230900 119620 231100 119880
rect 231400 119620 231600 119880
rect 231900 119620 232000 119880
rect 214000 119600 214120 119620
rect 214380 119600 214620 119620
rect 214880 119600 215120 119620
rect 215380 119600 215620 119620
rect 215880 119600 216120 119620
rect 216380 119600 216620 119620
rect 216880 119600 217120 119620
rect 217380 119600 217620 119620
rect 217880 119600 218120 119620
rect 218380 119600 218620 119620
rect 218880 119600 219120 119620
rect 219380 119600 219620 119620
rect 219880 119600 220120 119620
rect 220380 119600 220620 119620
rect 220880 119600 221120 119620
rect 221380 119600 221620 119620
rect 221880 119600 222120 119620
rect 222380 119600 222620 119620
rect 222880 119600 223120 119620
rect 223380 119600 223620 119620
rect 223880 119600 224120 119620
rect 224380 119600 224620 119620
rect 224880 119600 225120 119620
rect 225380 119600 225620 119620
rect 225880 119600 226120 119620
rect 226380 119600 226620 119620
rect 226880 119600 227120 119620
rect 227380 119600 227620 119620
rect 227880 119600 228120 119620
rect 228380 119600 228620 119620
rect 228880 119600 229120 119620
rect 229380 119600 229620 119620
rect 229880 119600 230120 119620
rect 230380 119600 230620 119620
rect 230880 119600 231120 119620
rect 231380 119600 231620 119620
rect 231880 119600 232000 119620
rect 214000 119400 232000 119600
rect 214000 119380 214120 119400
rect 214380 119380 214620 119400
rect 214880 119380 215120 119400
rect 215380 119380 215620 119400
rect 215880 119380 216120 119400
rect 216380 119380 216620 119400
rect 216880 119380 217120 119400
rect 217380 119380 217620 119400
rect 217880 119380 218120 119400
rect 218380 119380 218620 119400
rect 218880 119380 219120 119400
rect 219380 119380 219620 119400
rect 219880 119380 220120 119400
rect 220380 119380 220620 119400
rect 220880 119380 221120 119400
rect 221380 119380 221620 119400
rect 221880 119380 222120 119400
rect 222380 119380 222620 119400
rect 222880 119380 223120 119400
rect 223380 119380 223620 119400
rect 223880 119380 224120 119400
rect 224380 119380 224620 119400
rect 224880 119380 225120 119400
rect 225380 119380 225620 119400
rect 225880 119380 226120 119400
rect 226380 119380 226620 119400
rect 226880 119380 227120 119400
rect 227380 119380 227620 119400
rect 227880 119380 228120 119400
rect 228380 119380 228620 119400
rect 228880 119380 229120 119400
rect 229380 119380 229620 119400
rect 229880 119380 230120 119400
rect 230380 119380 230620 119400
rect 230880 119380 231120 119400
rect 231380 119380 231620 119400
rect 231880 119380 232000 119400
rect 214000 119120 214100 119380
rect 214400 119120 214600 119380
rect 214900 119120 215100 119380
rect 215400 119120 215600 119380
rect 215900 119120 216100 119380
rect 216400 119120 216600 119380
rect 216900 119120 217100 119380
rect 217400 119120 217600 119380
rect 217900 119120 218100 119380
rect 218400 119120 218600 119380
rect 218900 119120 219100 119380
rect 219400 119120 219600 119380
rect 219900 119120 220100 119380
rect 220400 119120 220600 119380
rect 220900 119120 221100 119380
rect 221400 119120 221600 119380
rect 221900 119120 222100 119380
rect 222400 119120 222600 119380
rect 222900 119120 223100 119380
rect 223400 119120 223600 119380
rect 223900 119120 224100 119380
rect 224400 119120 224600 119380
rect 224900 119120 225100 119380
rect 225400 119120 225600 119380
rect 225900 119120 226100 119380
rect 226400 119120 226600 119380
rect 226900 119120 227100 119380
rect 227400 119120 227600 119380
rect 227900 119120 228100 119380
rect 228400 119120 228600 119380
rect 228900 119120 229100 119380
rect 229400 119120 229600 119380
rect 229900 119120 230100 119380
rect 230400 119120 230600 119380
rect 230900 119120 231100 119380
rect 231400 119120 231600 119380
rect 231900 119120 232000 119380
rect 214000 119100 214120 119120
rect 214380 119100 214620 119120
rect 214880 119100 215120 119120
rect 215380 119100 215620 119120
rect 215880 119100 216120 119120
rect 216380 119100 216620 119120
rect 216880 119100 217120 119120
rect 217380 119100 217620 119120
rect 217880 119100 218120 119120
rect 218380 119100 218620 119120
rect 218880 119100 219120 119120
rect 219380 119100 219620 119120
rect 219880 119100 220120 119120
rect 220380 119100 220620 119120
rect 220880 119100 221120 119120
rect 221380 119100 221620 119120
rect 221880 119100 222120 119120
rect 222380 119100 222620 119120
rect 222880 119100 223120 119120
rect 223380 119100 223620 119120
rect 223880 119100 224120 119120
rect 224380 119100 224620 119120
rect 224880 119100 225120 119120
rect 225380 119100 225620 119120
rect 225880 119100 226120 119120
rect 226380 119100 226620 119120
rect 226880 119100 227120 119120
rect 227380 119100 227620 119120
rect 227880 119100 228120 119120
rect 228380 119100 228620 119120
rect 228880 119100 229120 119120
rect 229380 119100 229620 119120
rect 229880 119100 230120 119120
rect 230380 119100 230620 119120
rect 230880 119100 231120 119120
rect 231380 119100 231620 119120
rect 231880 119100 232000 119120
rect 214000 118900 232000 119100
rect 214000 118880 214120 118900
rect 214380 118880 214620 118900
rect 214880 118880 215120 118900
rect 215380 118880 215620 118900
rect 215880 118880 216120 118900
rect 216380 118880 216620 118900
rect 216880 118880 217120 118900
rect 217380 118880 217620 118900
rect 217880 118880 218120 118900
rect 218380 118880 218620 118900
rect 218880 118880 219120 118900
rect 219380 118880 219620 118900
rect 219880 118880 220120 118900
rect 220380 118880 220620 118900
rect 220880 118880 221120 118900
rect 221380 118880 221620 118900
rect 221880 118880 222120 118900
rect 222380 118880 222620 118900
rect 222880 118880 223120 118900
rect 223380 118880 223620 118900
rect 223880 118880 224120 118900
rect 224380 118880 224620 118900
rect 224880 118880 225120 118900
rect 225380 118880 225620 118900
rect 225880 118880 226120 118900
rect 226380 118880 226620 118900
rect 226880 118880 227120 118900
rect 227380 118880 227620 118900
rect 227880 118880 228120 118900
rect 228380 118880 228620 118900
rect 228880 118880 229120 118900
rect 229380 118880 229620 118900
rect 229880 118880 230120 118900
rect 230380 118880 230620 118900
rect 230880 118880 231120 118900
rect 231380 118880 231620 118900
rect 231880 118880 232000 118900
rect 214000 118620 214100 118880
rect 214400 118620 214600 118880
rect 214900 118620 215100 118880
rect 215400 118620 215600 118880
rect 215900 118620 216100 118880
rect 216400 118620 216600 118880
rect 216900 118620 217100 118880
rect 217400 118620 217600 118880
rect 217900 118620 218100 118880
rect 218400 118620 218600 118880
rect 218900 118620 219100 118880
rect 219400 118620 219600 118880
rect 219900 118620 220100 118880
rect 220400 118620 220600 118880
rect 220900 118620 221100 118880
rect 221400 118620 221600 118880
rect 221900 118620 222100 118880
rect 222400 118620 222600 118880
rect 222900 118620 223100 118880
rect 223400 118620 223600 118880
rect 223900 118620 224100 118880
rect 224400 118620 224600 118880
rect 224900 118620 225100 118880
rect 225400 118620 225600 118880
rect 225900 118620 226100 118880
rect 226400 118620 226600 118880
rect 226900 118620 227100 118880
rect 227400 118620 227600 118880
rect 227900 118620 228100 118880
rect 228400 118620 228600 118880
rect 228900 118620 229100 118880
rect 229400 118620 229600 118880
rect 229900 118620 230100 118880
rect 230400 118620 230600 118880
rect 230900 118620 231100 118880
rect 231400 118620 231600 118880
rect 231900 118620 232000 118880
rect 214000 118600 214120 118620
rect 214380 118600 214620 118620
rect 214880 118600 215120 118620
rect 215380 118600 215620 118620
rect 215880 118600 216120 118620
rect 216380 118600 216620 118620
rect 216880 118600 217120 118620
rect 217380 118600 217620 118620
rect 217880 118600 218120 118620
rect 218380 118600 218620 118620
rect 218880 118600 219120 118620
rect 219380 118600 219620 118620
rect 219880 118600 220120 118620
rect 220380 118600 220620 118620
rect 220880 118600 221120 118620
rect 221380 118600 221620 118620
rect 221880 118600 222120 118620
rect 222380 118600 222620 118620
rect 222880 118600 223120 118620
rect 223380 118600 223620 118620
rect 223880 118600 224120 118620
rect 224380 118600 224620 118620
rect 224880 118600 225120 118620
rect 225380 118600 225620 118620
rect 225880 118600 226120 118620
rect 226380 118600 226620 118620
rect 226880 118600 227120 118620
rect 227380 118600 227620 118620
rect 227880 118600 228120 118620
rect 228380 118600 228620 118620
rect 228880 118600 229120 118620
rect 229380 118600 229620 118620
rect 229880 118600 230120 118620
rect 230380 118600 230620 118620
rect 230880 118600 231120 118620
rect 231380 118600 231620 118620
rect 231880 118600 232000 118620
rect 214000 118400 232000 118600
rect 214000 118380 214120 118400
rect 214380 118380 214620 118400
rect 214880 118380 215120 118400
rect 215380 118380 215620 118400
rect 215880 118380 216120 118400
rect 216380 118380 216620 118400
rect 216880 118380 217120 118400
rect 217380 118380 217620 118400
rect 217880 118380 218120 118400
rect 218380 118380 218620 118400
rect 218880 118380 219120 118400
rect 219380 118380 219620 118400
rect 219880 118380 220120 118400
rect 220380 118380 220620 118400
rect 220880 118380 221120 118400
rect 221380 118380 221620 118400
rect 221880 118380 222120 118400
rect 222380 118380 222620 118400
rect 222880 118380 223120 118400
rect 223380 118380 223620 118400
rect 223880 118380 224120 118400
rect 224380 118380 224620 118400
rect 224880 118380 225120 118400
rect 225380 118380 225620 118400
rect 225880 118380 226120 118400
rect 226380 118380 226620 118400
rect 226880 118380 227120 118400
rect 227380 118380 227620 118400
rect 227880 118380 228120 118400
rect 228380 118380 228620 118400
rect 228880 118380 229120 118400
rect 229380 118380 229620 118400
rect 229880 118380 230120 118400
rect 230380 118380 230620 118400
rect 230880 118380 231120 118400
rect 231380 118380 231620 118400
rect 231880 118380 232000 118400
rect 214000 118120 214100 118380
rect 214400 118120 214600 118380
rect 214900 118120 215100 118380
rect 215400 118120 215600 118380
rect 215900 118120 216100 118380
rect 216400 118120 216600 118380
rect 216900 118120 217100 118380
rect 217400 118120 217600 118380
rect 217900 118120 218100 118380
rect 218400 118120 218600 118380
rect 218900 118120 219100 118380
rect 219400 118120 219600 118380
rect 219900 118120 220100 118380
rect 220400 118120 220600 118380
rect 220900 118120 221100 118380
rect 221400 118120 221600 118380
rect 221900 118120 222100 118380
rect 222400 118120 222600 118380
rect 222900 118120 223100 118380
rect 223400 118120 223600 118380
rect 223900 118120 224100 118380
rect 224400 118120 224600 118380
rect 224900 118120 225100 118380
rect 225400 118120 225600 118380
rect 225900 118120 226100 118380
rect 226400 118120 226600 118380
rect 226900 118120 227100 118380
rect 227400 118120 227600 118380
rect 227900 118120 228100 118380
rect 228400 118120 228600 118380
rect 228900 118120 229100 118380
rect 229400 118120 229600 118380
rect 229900 118120 230100 118380
rect 230400 118120 230600 118380
rect 230900 118120 231100 118380
rect 231400 118120 231600 118380
rect 231900 118120 232000 118380
rect 214000 118100 214120 118120
rect 214380 118100 214620 118120
rect 214880 118100 215120 118120
rect 215380 118100 215620 118120
rect 215880 118100 216120 118120
rect 216380 118100 216620 118120
rect 216880 118100 217120 118120
rect 217380 118100 217620 118120
rect 217880 118100 218120 118120
rect 218380 118100 218620 118120
rect 218880 118100 219120 118120
rect 219380 118100 219620 118120
rect 219880 118100 220120 118120
rect 220380 118100 220620 118120
rect 220880 118100 221120 118120
rect 221380 118100 221620 118120
rect 221880 118100 222120 118120
rect 222380 118100 222620 118120
rect 222880 118100 223120 118120
rect 223380 118100 223620 118120
rect 223880 118100 224120 118120
rect 224380 118100 224620 118120
rect 224880 118100 225120 118120
rect 225380 118100 225620 118120
rect 225880 118100 226120 118120
rect 226380 118100 226620 118120
rect 226880 118100 227120 118120
rect 227380 118100 227620 118120
rect 227880 118100 228120 118120
rect 228380 118100 228620 118120
rect 228880 118100 229120 118120
rect 229380 118100 229620 118120
rect 229880 118100 230120 118120
rect 230380 118100 230620 118120
rect 230880 118100 231120 118120
rect 231380 118100 231620 118120
rect 231880 118100 232000 118120
rect 214000 117900 232000 118100
rect 214000 117880 214120 117900
rect 214380 117880 214620 117900
rect 214880 117880 215120 117900
rect 215380 117880 215620 117900
rect 215880 117880 216120 117900
rect 216380 117880 216620 117900
rect 216880 117880 217120 117900
rect 217380 117880 217620 117900
rect 217880 117880 218120 117900
rect 218380 117880 218620 117900
rect 218880 117880 219120 117900
rect 219380 117880 219620 117900
rect 219880 117880 220120 117900
rect 220380 117880 220620 117900
rect 220880 117880 221120 117900
rect 221380 117880 221620 117900
rect 221880 117880 222120 117900
rect 222380 117880 222620 117900
rect 222880 117880 223120 117900
rect 223380 117880 223620 117900
rect 223880 117880 224120 117900
rect 224380 117880 224620 117900
rect 224880 117880 225120 117900
rect 225380 117880 225620 117900
rect 225880 117880 226120 117900
rect 226380 117880 226620 117900
rect 226880 117880 227120 117900
rect 227380 117880 227620 117900
rect 227880 117880 228120 117900
rect 228380 117880 228620 117900
rect 228880 117880 229120 117900
rect 229380 117880 229620 117900
rect 229880 117880 230120 117900
rect 230380 117880 230620 117900
rect 230880 117880 231120 117900
rect 231380 117880 231620 117900
rect 231880 117880 232000 117900
rect 214000 117620 214100 117880
rect 214400 117620 214600 117880
rect 214900 117620 215100 117880
rect 215400 117620 215600 117880
rect 215900 117620 216100 117880
rect 216400 117620 216600 117880
rect 216900 117620 217100 117880
rect 217400 117620 217600 117880
rect 217900 117620 218100 117880
rect 218400 117620 218600 117880
rect 218900 117620 219100 117880
rect 219400 117620 219600 117880
rect 219900 117620 220100 117880
rect 220400 117620 220600 117880
rect 220900 117620 221100 117880
rect 221400 117620 221600 117880
rect 221900 117620 222100 117880
rect 222400 117620 222600 117880
rect 222900 117620 223100 117880
rect 223400 117620 223600 117880
rect 223900 117620 224100 117880
rect 224400 117620 224600 117880
rect 224900 117620 225100 117880
rect 225400 117620 225600 117880
rect 225900 117620 226100 117880
rect 226400 117620 226600 117880
rect 226900 117620 227100 117880
rect 227400 117620 227600 117880
rect 227900 117620 228100 117880
rect 228400 117620 228600 117880
rect 228900 117620 229100 117880
rect 229400 117620 229600 117880
rect 229900 117620 230100 117880
rect 230400 117620 230600 117880
rect 230900 117620 231100 117880
rect 231400 117620 231600 117880
rect 231900 117620 232000 117880
rect 214000 117600 214120 117620
rect 214380 117600 214620 117620
rect 214880 117600 215120 117620
rect 215380 117600 215620 117620
rect 215880 117600 216120 117620
rect 216380 117600 216620 117620
rect 216880 117600 217120 117620
rect 217380 117600 217620 117620
rect 217880 117600 218120 117620
rect 218380 117600 218620 117620
rect 218880 117600 219120 117620
rect 219380 117600 219620 117620
rect 219880 117600 220120 117620
rect 220380 117600 220620 117620
rect 220880 117600 221120 117620
rect 221380 117600 221620 117620
rect 221880 117600 222120 117620
rect 222380 117600 222620 117620
rect 222880 117600 223120 117620
rect 223380 117600 223620 117620
rect 223880 117600 224120 117620
rect 224380 117600 224620 117620
rect 224880 117600 225120 117620
rect 225380 117600 225620 117620
rect 225880 117600 226120 117620
rect 226380 117600 226620 117620
rect 226880 117600 227120 117620
rect 227380 117600 227620 117620
rect 227880 117600 228120 117620
rect 228380 117600 228620 117620
rect 228880 117600 229120 117620
rect 229380 117600 229620 117620
rect 229880 117600 230120 117620
rect 230380 117600 230620 117620
rect 230880 117600 231120 117620
rect 231380 117600 231620 117620
rect 231880 117600 232000 117620
rect 214000 117400 232000 117600
rect 214000 117380 214120 117400
rect 214380 117380 214620 117400
rect 214880 117380 215120 117400
rect 215380 117380 215620 117400
rect 215880 117380 216120 117400
rect 216380 117380 216620 117400
rect 216880 117380 217120 117400
rect 217380 117380 217620 117400
rect 217880 117380 218120 117400
rect 218380 117380 218620 117400
rect 218880 117380 219120 117400
rect 219380 117380 219620 117400
rect 219880 117380 220120 117400
rect 220380 117380 220620 117400
rect 220880 117380 221120 117400
rect 221380 117380 221620 117400
rect 221880 117380 222120 117400
rect 222380 117380 222620 117400
rect 222880 117380 223120 117400
rect 223380 117380 223620 117400
rect 223880 117380 224120 117400
rect 224380 117380 224620 117400
rect 224880 117380 225120 117400
rect 225380 117380 225620 117400
rect 225880 117380 226120 117400
rect 226380 117380 226620 117400
rect 226880 117380 227120 117400
rect 227380 117380 227620 117400
rect 227880 117380 228120 117400
rect 228380 117380 228620 117400
rect 228880 117380 229120 117400
rect 229380 117380 229620 117400
rect 229880 117380 230120 117400
rect 230380 117380 230620 117400
rect 230880 117380 231120 117400
rect 231380 117380 231620 117400
rect 231880 117380 232000 117400
rect 214000 117120 214100 117380
rect 214400 117120 214600 117380
rect 214900 117120 215100 117380
rect 215400 117120 215600 117380
rect 215900 117120 216100 117380
rect 216400 117120 216600 117380
rect 216900 117120 217100 117380
rect 217400 117120 217600 117380
rect 217900 117120 218100 117380
rect 218400 117120 218600 117380
rect 218900 117120 219100 117380
rect 219400 117120 219600 117380
rect 219900 117120 220100 117380
rect 220400 117120 220600 117380
rect 220900 117120 221100 117380
rect 221400 117120 221600 117380
rect 221900 117120 222100 117380
rect 222400 117120 222600 117380
rect 222900 117120 223100 117380
rect 223400 117120 223600 117380
rect 223900 117120 224100 117380
rect 224400 117120 224600 117380
rect 224900 117120 225100 117380
rect 225400 117120 225600 117380
rect 225900 117120 226100 117380
rect 226400 117120 226600 117380
rect 226900 117120 227100 117380
rect 227400 117120 227600 117380
rect 227900 117120 228100 117380
rect 228400 117120 228600 117380
rect 228900 117120 229100 117380
rect 229400 117120 229600 117380
rect 229900 117120 230100 117380
rect 230400 117120 230600 117380
rect 230900 117120 231100 117380
rect 231400 117120 231600 117380
rect 231900 117120 232000 117380
rect 214000 117100 214120 117120
rect 214380 117100 214620 117120
rect 214880 117100 215120 117120
rect 215380 117100 215620 117120
rect 215880 117100 216120 117120
rect 216380 117100 216620 117120
rect 216880 117100 217120 117120
rect 217380 117100 217620 117120
rect 217880 117100 218120 117120
rect 218380 117100 218620 117120
rect 218880 117100 219120 117120
rect 219380 117100 219620 117120
rect 219880 117100 220120 117120
rect 220380 117100 220620 117120
rect 220880 117100 221120 117120
rect 221380 117100 221620 117120
rect 221880 117100 222120 117120
rect 222380 117100 222620 117120
rect 222880 117100 223120 117120
rect 223380 117100 223620 117120
rect 223880 117100 224120 117120
rect 224380 117100 224620 117120
rect 224880 117100 225120 117120
rect 225380 117100 225620 117120
rect 225880 117100 226120 117120
rect 226380 117100 226620 117120
rect 226880 117100 227120 117120
rect 227380 117100 227620 117120
rect 227880 117100 228120 117120
rect 228380 117100 228620 117120
rect 228880 117100 229120 117120
rect 229380 117100 229620 117120
rect 229880 117100 230120 117120
rect 230380 117100 230620 117120
rect 230880 117100 231120 117120
rect 231380 117100 231620 117120
rect 231880 117100 232000 117120
rect 214000 116900 232000 117100
rect 214000 116880 214120 116900
rect 214380 116880 214620 116900
rect 214880 116880 215120 116900
rect 215380 116880 215620 116900
rect 215880 116880 216120 116900
rect 216380 116880 216620 116900
rect 216880 116880 217120 116900
rect 217380 116880 217620 116900
rect 217880 116880 218120 116900
rect 218380 116880 218620 116900
rect 218880 116880 219120 116900
rect 219380 116880 219620 116900
rect 219880 116880 220120 116900
rect 220380 116880 220620 116900
rect 220880 116880 221120 116900
rect 221380 116880 221620 116900
rect 221880 116880 222120 116900
rect 222380 116880 222620 116900
rect 222880 116880 223120 116900
rect 223380 116880 223620 116900
rect 223880 116880 224120 116900
rect 224380 116880 224620 116900
rect 224880 116880 225120 116900
rect 225380 116880 225620 116900
rect 225880 116880 226120 116900
rect 226380 116880 226620 116900
rect 226880 116880 227120 116900
rect 227380 116880 227620 116900
rect 227880 116880 228120 116900
rect 228380 116880 228620 116900
rect 228880 116880 229120 116900
rect 229380 116880 229620 116900
rect 229880 116880 230120 116900
rect 230380 116880 230620 116900
rect 230880 116880 231120 116900
rect 231380 116880 231620 116900
rect 231880 116880 232000 116900
rect 214000 116620 214100 116880
rect 214400 116620 214600 116880
rect 214900 116620 215100 116880
rect 215400 116620 215600 116880
rect 215900 116620 216100 116880
rect 216400 116620 216600 116880
rect 216900 116620 217100 116880
rect 217400 116620 217600 116880
rect 217900 116620 218100 116880
rect 218400 116620 218600 116880
rect 218900 116620 219100 116880
rect 219400 116620 219600 116880
rect 219900 116620 220100 116880
rect 220400 116620 220600 116880
rect 220900 116620 221100 116880
rect 221400 116620 221600 116880
rect 221900 116620 222100 116880
rect 222400 116620 222600 116880
rect 222900 116620 223100 116880
rect 223400 116620 223600 116880
rect 223900 116620 224100 116880
rect 224400 116620 224600 116880
rect 224900 116620 225100 116880
rect 225400 116620 225600 116880
rect 225900 116620 226100 116880
rect 226400 116620 226600 116880
rect 226900 116620 227100 116880
rect 227400 116620 227600 116880
rect 227900 116620 228100 116880
rect 228400 116620 228600 116880
rect 228900 116620 229100 116880
rect 229400 116620 229600 116880
rect 229900 116620 230100 116880
rect 230400 116620 230600 116880
rect 230900 116620 231100 116880
rect 231400 116620 231600 116880
rect 231900 116620 232000 116880
rect 214000 116600 214120 116620
rect 214380 116600 214620 116620
rect 214880 116600 215120 116620
rect 215380 116600 215620 116620
rect 215880 116600 216120 116620
rect 216380 116600 216620 116620
rect 216880 116600 217120 116620
rect 217380 116600 217620 116620
rect 217880 116600 218120 116620
rect 218380 116600 218620 116620
rect 218880 116600 219120 116620
rect 219380 116600 219620 116620
rect 219880 116600 220120 116620
rect 220380 116600 220620 116620
rect 220880 116600 221120 116620
rect 221380 116600 221620 116620
rect 221880 116600 222120 116620
rect 222380 116600 222620 116620
rect 222880 116600 223120 116620
rect 223380 116600 223620 116620
rect 223880 116600 224120 116620
rect 224380 116600 224620 116620
rect 224880 116600 225120 116620
rect 225380 116600 225620 116620
rect 225880 116600 226120 116620
rect 226380 116600 226620 116620
rect 226880 116600 227120 116620
rect 227380 116600 227620 116620
rect 227880 116600 228120 116620
rect 228380 116600 228620 116620
rect 228880 116600 229120 116620
rect 229380 116600 229620 116620
rect 229880 116600 230120 116620
rect 230380 116600 230620 116620
rect 230880 116600 231120 116620
rect 231380 116600 231620 116620
rect 231880 116600 232000 116620
rect 214000 116400 232000 116600
rect 214000 116380 214120 116400
rect 214380 116380 214620 116400
rect 214880 116380 215120 116400
rect 215380 116380 215620 116400
rect 215880 116380 216120 116400
rect 216380 116380 216620 116400
rect 216880 116380 217120 116400
rect 217380 116380 217620 116400
rect 217880 116380 218120 116400
rect 218380 116380 218620 116400
rect 218880 116380 219120 116400
rect 219380 116380 219620 116400
rect 219880 116380 220120 116400
rect 220380 116380 220620 116400
rect 220880 116380 221120 116400
rect 221380 116380 221620 116400
rect 221880 116380 222120 116400
rect 222380 116380 222620 116400
rect 222880 116380 223120 116400
rect 223380 116380 223620 116400
rect 223880 116380 224120 116400
rect 224380 116380 224620 116400
rect 224880 116380 225120 116400
rect 225380 116380 225620 116400
rect 225880 116380 226120 116400
rect 226380 116380 226620 116400
rect 226880 116380 227120 116400
rect 227380 116380 227620 116400
rect 227880 116380 228120 116400
rect 228380 116380 228620 116400
rect 228880 116380 229120 116400
rect 229380 116380 229620 116400
rect 229880 116380 230120 116400
rect 230380 116380 230620 116400
rect 230880 116380 231120 116400
rect 231380 116380 231620 116400
rect 231880 116380 232000 116400
rect 214000 116120 214100 116380
rect 214400 116120 214600 116380
rect 214900 116120 215100 116380
rect 215400 116120 215600 116380
rect 215900 116120 216100 116380
rect 216400 116120 216600 116380
rect 216900 116120 217100 116380
rect 217400 116120 217600 116380
rect 217900 116120 218100 116380
rect 218400 116120 218600 116380
rect 218900 116120 219100 116380
rect 219400 116120 219600 116380
rect 219900 116120 220100 116380
rect 220400 116120 220600 116380
rect 220900 116120 221100 116380
rect 221400 116120 221600 116380
rect 221900 116120 222100 116380
rect 222400 116120 222600 116380
rect 222900 116120 223100 116380
rect 223400 116120 223600 116380
rect 223900 116120 224100 116380
rect 224400 116120 224600 116380
rect 224900 116120 225100 116380
rect 225400 116120 225600 116380
rect 225900 116120 226100 116380
rect 226400 116120 226600 116380
rect 226900 116120 227100 116380
rect 227400 116120 227600 116380
rect 227900 116120 228100 116380
rect 228400 116120 228600 116380
rect 228900 116120 229100 116380
rect 229400 116120 229600 116380
rect 229900 116120 230100 116380
rect 230400 116120 230600 116380
rect 230900 116120 231100 116380
rect 231400 116120 231600 116380
rect 231900 116120 232000 116380
rect 214000 116100 214120 116120
rect 214380 116100 214620 116120
rect 214880 116100 215120 116120
rect 215380 116100 215620 116120
rect 215880 116100 216120 116120
rect 216380 116100 216620 116120
rect 216880 116100 217120 116120
rect 217380 116100 217620 116120
rect 217880 116100 218120 116120
rect 218380 116100 218620 116120
rect 218880 116100 219120 116120
rect 219380 116100 219620 116120
rect 219880 116100 220120 116120
rect 220380 116100 220620 116120
rect 220880 116100 221120 116120
rect 221380 116100 221620 116120
rect 221880 116100 222120 116120
rect 222380 116100 222620 116120
rect 222880 116100 223120 116120
rect 223380 116100 223620 116120
rect 223880 116100 224120 116120
rect 224380 116100 224620 116120
rect 224880 116100 225120 116120
rect 225380 116100 225620 116120
rect 225880 116100 226120 116120
rect 226380 116100 226620 116120
rect 226880 116100 227120 116120
rect 227380 116100 227620 116120
rect 227880 116100 228120 116120
rect 228380 116100 228620 116120
rect 228880 116100 229120 116120
rect 229380 116100 229620 116120
rect 229880 116100 230120 116120
rect 230380 116100 230620 116120
rect 230880 116100 231120 116120
rect 231380 116100 231620 116120
rect 231880 116100 232000 116120
rect 214000 115900 232000 116100
rect 214000 115880 214120 115900
rect 214380 115880 214620 115900
rect 214880 115880 215120 115900
rect 215380 115880 215620 115900
rect 215880 115880 216120 115900
rect 216380 115880 216620 115900
rect 216880 115880 217120 115900
rect 217380 115880 217620 115900
rect 217880 115880 218120 115900
rect 218380 115880 218620 115900
rect 218880 115880 219120 115900
rect 219380 115880 219620 115900
rect 219880 115880 220120 115900
rect 220380 115880 220620 115900
rect 220880 115880 221120 115900
rect 221380 115880 221620 115900
rect 221880 115880 222120 115900
rect 222380 115880 222620 115900
rect 222880 115880 223120 115900
rect 223380 115880 223620 115900
rect 223880 115880 224120 115900
rect 224380 115880 224620 115900
rect 224880 115880 225120 115900
rect 225380 115880 225620 115900
rect 225880 115880 226120 115900
rect 226380 115880 226620 115900
rect 226880 115880 227120 115900
rect 227380 115880 227620 115900
rect 227880 115880 228120 115900
rect 228380 115880 228620 115900
rect 228880 115880 229120 115900
rect 229380 115880 229620 115900
rect 229880 115880 230120 115900
rect 230380 115880 230620 115900
rect 230880 115880 231120 115900
rect 231380 115880 231620 115900
rect 231880 115880 232000 115900
rect 214000 115620 214100 115880
rect 214400 115620 214600 115880
rect 214900 115620 215100 115880
rect 215400 115620 215600 115880
rect 215900 115620 216100 115880
rect 216400 115620 216600 115880
rect 216900 115620 217100 115880
rect 217400 115620 217600 115880
rect 217900 115620 218100 115880
rect 218400 115620 218600 115880
rect 218900 115620 219100 115880
rect 219400 115620 219600 115880
rect 219900 115620 220100 115880
rect 220400 115620 220600 115880
rect 220900 115620 221100 115880
rect 221400 115620 221600 115880
rect 221900 115620 222100 115880
rect 222400 115620 222600 115880
rect 222900 115620 223100 115880
rect 223400 115620 223600 115880
rect 223900 115620 224100 115880
rect 224400 115620 224600 115880
rect 224900 115620 225100 115880
rect 225400 115620 225600 115880
rect 225900 115620 226100 115880
rect 226400 115620 226600 115880
rect 226900 115620 227100 115880
rect 227400 115620 227600 115880
rect 227900 115620 228100 115880
rect 228400 115620 228600 115880
rect 228900 115620 229100 115880
rect 229400 115620 229600 115880
rect 229900 115620 230100 115880
rect 230400 115620 230600 115880
rect 230900 115620 231100 115880
rect 231400 115620 231600 115880
rect 231900 115620 232000 115880
rect 214000 115600 214120 115620
rect 214380 115600 214620 115620
rect 214880 115600 215120 115620
rect 215380 115600 215620 115620
rect 215880 115600 216120 115620
rect 216380 115600 216620 115620
rect 216880 115600 217120 115620
rect 217380 115600 217620 115620
rect 217880 115600 218120 115620
rect 218380 115600 218620 115620
rect 218880 115600 219120 115620
rect 219380 115600 219620 115620
rect 219880 115600 220120 115620
rect 220380 115600 220620 115620
rect 220880 115600 221120 115620
rect 221380 115600 221620 115620
rect 221880 115600 222120 115620
rect 222380 115600 222620 115620
rect 222880 115600 223120 115620
rect 223380 115600 223620 115620
rect 223880 115600 224120 115620
rect 224380 115600 224620 115620
rect 224880 115600 225120 115620
rect 225380 115600 225620 115620
rect 225880 115600 226120 115620
rect 226380 115600 226620 115620
rect 226880 115600 227120 115620
rect 227380 115600 227620 115620
rect 227880 115600 228120 115620
rect 228380 115600 228620 115620
rect 228880 115600 229120 115620
rect 229380 115600 229620 115620
rect 229880 115600 230120 115620
rect 230380 115600 230620 115620
rect 230880 115600 231120 115620
rect 231380 115600 231620 115620
rect 231880 115600 232000 115620
rect 214000 115400 232000 115600
rect 214000 115380 214120 115400
rect 214380 115380 214620 115400
rect 214880 115380 215120 115400
rect 215380 115380 215620 115400
rect 215880 115380 216120 115400
rect 216380 115380 216620 115400
rect 216880 115380 217120 115400
rect 217380 115380 217620 115400
rect 217880 115380 218120 115400
rect 218380 115380 218620 115400
rect 218880 115380 219120 115400
rect 219380 115380 219620 115400
rect 219880 115380 220120 115400
rect 220380 115380 220620 115400
rect 220880 115380 221120 115400
rect 221380 115380 221620 115400
rect 221880 115380 222120 115400
rect 222380 115380 222620 115400
rect 222880 115380 223120 115400
rect 223380 115380 223620 115400
rect 223880 115380 224120 115400
rect 224380 115380 224620 115400
rect 224880 115380 225120 115400
rect 225380 115380 225620 115400
rect 225880 115380 226120 115400
rect 226380 115380 226620 115400
rect 226880 115380 227120 115400
rect 227380 115380 227620 115400
rect 227880 115380 228120 115400
rect 228380 115380 228620 115400
rect 228880 115380 229120 115400
rect 229380 115380 229620 115400
rect 229880 115380 230120 115400
rect 230380 115380 230620 115400
rect 230880 115380 231120 115400
rect 231380 115380 231620 115400
rect 231880 115380 232000 115400
rect 214000 115120 214100 115380
rect 214400 115120 214600 115380
rect 214900 115120 215100 115380
rect 215400 115120 215600 115380
rect 215900 115120 216100 115380
rect 216400 115120 216600 115380
rect 216900 115120 217100 115380
rect 217400 115120 217600 115380
rect 217900 115120 218100 115380
rect 218400 115120 218600 115380
rect 218900 115120 219100 115380
rect 219400 115120 219600 115380
rect 219900 115120 220100 115380
rect 220400 115120 220600 115380
rect 220900 115120 221100 115380
rect 221400 115120 221600 115380
rect 221900 115120 222100 115380
rect 222400 115120 222600 115380
rect 222900 115120 223100 115380
rect 223400 115120 223600 115380
rect 223900 115120 224100 115380
rect 224400 115120 224600 115380
rect 224900 115120 225100 115380
rect 225400 115120 225600 115380
rect 225900 115120 226100 115380
rect 226400 115120 226600 115380
rect 226900 115120 227100 115380
rect 227400 115120 227600 115380
rect 227900 115120 228100 115380
rect 228400 115120 228600 115380
rect 228900 115120 229100 115380
rect 229400 115120 229600 115380
rect 229900 115120 230100 115380
rect 230400 115120 230600 115380
rect 230900 115120 231100 115380
rect 231400 115120 231600 115380
rect 231900 115120 232000 115380
rect 214000 115100 214120 115120
rect 214380 115100 214620 115120
rect 214880 115100 215120 115120
rect 215380 115100 215620 115120
rect 215880 115100 216120 115120
rect 216380 115100 216620 115120
rect 216880 115100 217120 115120
rect 217380 115100 217620 115120
rect 217880 115100 218120 115120
rect 218380 115100 218620 115120
rect 218880 115100 219120 115120
rect 219380 115100 219620 115120
rect 219880 115100 220120 115120
rect 220380 115100 220620 115120
rect 220880 115100 221120 115120
rect 221380 115100 221620 115120
rect 221880 115100 222120 115120
rect 222380 115100 222620 115120
rect 222880 115100 223120 115120
rect 223380 115100 223620 115120
rect 223880 115100 224120 115120
rect 224380 115100 224620 115120
rect 224880 115100 225120 115120
rect 225380 115100 225620 115120
rect 225880 115100 226120 115120
rect 226380 115100 226620 115120
rect 226880 115100 227120 115120
rect 227380 115100 227620 115120
rect 227880 115100 228120 115120
rect 228380 115100 228620 115120
rect 228880 115100 229120 115120
rect 229380 115100 229620 115120
rect 229880 115100 230120 115120
rect 230380 115100 230620 115120
rect 230880 115100 231120 115120
rect 231380 115100 231620 115120
rect 231880 115100 232000 115120
rect 214000 114900 232000 115100
rect 214000 114880 214120 114900
rect 214380 114880 214620 114900
rect 214880 114880 215120 114900
rect 215380 114880 215620 114900
rect 215880 114880 216120 114900
rect 216380 114880 216620 114900
rect 216880 114880 217120 114900
rect 217380 114880 217620 114900
rect 217880 114880 218120 114900
rect 218380 114880 218620 114900
rect 218880 114880 219120 114900
rect 219380 114880 219620 114900
rect 219880 114880 220120 114900
rect 220380 114880 220620 114900
rect 220880 114880 221120 114900
rect 221380 114880 221620 114900
rect 221880 114880 222120 114900
rect 222380 114880 222620 114900
rect 222880 114880 223120 114900
rect 223380 114880 223620 114900
rect 223880 114880 224120 114900
rect 224380 114880 224620 114900
rect 224880 114880 225120 114900
rect 225380 114880 225620 114900
rect 225880 114880 226120 114900
rect 226380 114880 226620 114900
rect 226880 114880 227120 114900
rect 227380 114880 227620 114900
rect 227880 114880 228120 114900
rect 228380 114880 228620 114900
rect 228880 114880 229120 114900
rect 229380 114880 229620 114900
rect 229880 114880 230120 114900
rect 230380 114880 230620 114900
rect 230880 114880 231120 114900
rect 231380 114880 231620 114900
rect 231880 114880 232000 114900
rect 214000 114620 214100 114880
rect 214400 114620 214600 114880
rect 214900 114620 215100 114880
rect 215400 114620 215600 114880
rect 215900 114620 216100 114880
rect 216400 114620 216600 114880
rect 216900 114620 217100 114880
rect 217400 114620 217600 114880
rect 217900 114620 218100 114880
rect 218400 114620 218600 114880
rect 218900 114620 219100 114880
rect 219400 114620 219600 114880
rect 219900 114620 220100 114880
rect 220400 114620 220600 114880
rect 220900 114620 221100 114880
rect 221400 114620 221600 114880
rect 221900 114620 222100 114880
rect 222400 114620 222600 114880
rect 222900 114620 223100 114880
rect 223400 114620 223600 114880
rect 223900 114620 224100 114880
rect 224400 114620 224600 114880
rect 224900 114620 225100 114880
rect 225400 114620 225600 114880
rect 225900 114620 226100 114880
rect 226400 114620 226600 114880
rect 226900 114620 227100 114880
rect 227400 114620 227600 114880
rect 227900 114620 228100 114880
rect 228400 114620 228600 114880
rect 228900 114620 229100 114880
rect 229400 114620 229600 114880
rect 229900 114620 230100 114880
rect 230400 114620 230600 114880
rect 230900 114620 231100 114880
rect 231400 114620 231600 114880
rect 231900 114620 232000 114880
rect 214000 114600 214120 114620
rect 214380 114600 214620 114620
rect 214880 114600 215120 114620
rect 215380 114600 215620 114620
rect 215880 114600 216120 114620
rect 216380 114600 216620 114620
rect 216880 114600 217120 114620
rect 217380 114600 217620 114620
rect 217880 114600 218120 114620
rect 218380 114600 218620 114620
rect 218880 114600 219120 114620
rect 219380 114600 219620 114620
rect 219880 114600 220120 114620
rect 220380 114600 220620 114620
rect 220880 114600 221120 114620
rect 221380 114600 221620 114620
rect 221880 114600 222120 114620
rect 222380 114600 222620 114620
rect 222880 114600 223120 114620
rect 223380 114600 223620 114620
rect 223880 114600 224120 114620
rect 224380 114600 224620 114620
rect 224880 114600 225120 114620
rect 225380 114600 225620 114620
rect 225880 114600 226120 114620
rect 226380 114600 226620 114620
rect 226880 114600 227120 114620
rect 227380 114600 227620 114620
rect 227880 114600 228120 114620
rect 228380 114600 228620 114620
rect 228880 114600 229120 114620
rect 229380 114600 229620 114620
rect 229880 114600 230120 114620
rect 230380 114600 230620 114620
rect 230880 114600 231120 114620
rect 231380 114600 231620 114620
rect 231880 114600 232000 114620
rect 214000 114400 232000 114600
rect 214000 114380 214120 114400
rect 214380 114380 214620 114400
rect 214880 114380 215120 114400
rect 215380 114380 215620 114400
rect 215880 114380 216120 114400
rect 216380 114380 216620 114400
rect 216880 114380 217120 114400
rect 217380 114380 217620 114400
rect 217880 114380 218120 114400
rect 218380 114380 218620 114400
rect 218880 114380 219120 114400
rect 219380 114380 219620 114400
rect 219880 114380 220120 114400
rect 220380 114380 220620 114400
rect 220880 114380 221120 114400
rect 221380 114380 221620 114400
rect 221880 114380 222120 114400
rect 222380 114380 222620 114400
rect 222880 114380 223120 114400
rect 223380 114380 223620 114400
rect 223880 114380 224120 114400
rect 224380 114380 224620 114400
rect 224880 114380 225120 114400
rect 225380 114380 225620 114400
rect 225880 114380 226120 114400
rect 226380 114380 226620 114400
rect 226880 114380 227120 114400
rect 227380 114380 227620 114400
rect 227880 114380 228120 114400
rect 228380 114380 228620 114400
rect 228880 114380 229120 114400
rect 229380 114380 229620 114400
rect 229880 114380 230120 114400
rect 230380 114380 230620 114400
rect 230880 114380 231120 114400
rect 231380 114380 231620 114400
rect 231880 114380 232000 114400
rect 214000 114120 214100 114380
rect 214400 114120 214600 114380
rect 214900 114120 215100 114380
rect 215400 114120 215600 114380
rect 215900 114120 216100 114380
rect 216400 114120 216600 114380
rect 216900 114120 217100 114380
rect 217400 114120 217600 114380
rect 217900 114120 218100 114380
rect 218400 114120 218600 114380
rect 218900 114120 219100 114380
rect 219400 114120 219600 114380
rect 219900 114120 220100 114380
rect 220400 114120 220600 114380
rect 220900 114120 221100 114380
rect 221400 114120 221600 114380
rect 221900 114120 222100 114380
rect 222400 114120 222600 114380
rect 222900 114120 223100 114380
rect 223400 114120 223600 114380
rect 223900 114120 224100 114380
rect 224400 114120 224600 114380
rect 224900 114120 225100 114380
rect 225400 114120 225600 114380
rect 225900 114120 226100 114380
rect 226400 114120 226600 114380
rect 226900 114120 227100 114380
rect 227400 114120 227600 114380
rect 227900 114120 228100 114380
rect 228400 114120 228600 114380
rect 228900 114120 229100 114380
rect 229400 114120 229600 114380
rect 229900 114120 230100 114380
rect 230400 114120 230600 114380
rect 230900 114120 231100 114380
rect 231400 114120 231600 114380
rect 231900 114120 232000 114380
rect 214000 114100 214120 114120
rect 214380 114100 214620 114120
rect 214880 114100 215120 114120
rect 215380 114100 215620 114120
rect 215880 114100 216120 114120
rect 216380 114100 216620 114120
rect 216880 114100 217120 114120
rect 217380 114100 217620 114120
rect 217880 114100 218120 114120
rect 218380 114100 218620 114120
rect 218880 114100 219120 114120
rect 219380 114100 219620 114120
rect 219880 114100 220120 114120
rect 220380 114100 220620 114120
rect 220880 114100 221120 114120
rect 221380 114100 221620 114120
rect 221880 114100 222120 114120
rect 222380 114100 222620 114120
rect 222880 114100 223120 114120
rect 223380 114100 223620 114120
rect 223880 114100 224120 114120
rect 224380 114100 224620 114120
rect 224880 114100 225120 114120
rect 225380 114100 225620 114120
rect 225880 114100 226120 114120
rect 226380 114100 226620 114120
rect 226880 114100 227120 114120
rect 227380 114100 227620 114120
rect 227880 114100 228120 114120
rect 228380 114100 228620 114120
rect 228880 114100 229120 114120
rect 229380 114100 229620 114120
rect 229880 114100 230120 114120
rect 230380 114100 230620 114120
rect 230880 114100 231120 114120
rect 231380 114100 231620 114120
rect 231880 114100 232000 114120
rect 214000 114000 232000 114100
rect 178000 113900 232000 114000
rect 178000 113880 178120 113900
rect 178380 113880 178620 113900
rect 178880 113880 179120 113900
rect 179380 113880 179620 113900
rect 179880 113880 180120 113900
rect 180380 113880 180620 113900
rect 180880 113880 181120 113900
rect 181380 113880 181620 113900
rect 181880 113880 182120 113900
rect 182380 113880 182620 113900
rect 182880 113880 183120 113900
rect 183380 113880 183620 113900
rect 183880 113880 184120 113900
rect 184380 113880 184620 113900
rect 184880 113880 185120 113900
rect 185380 113880 185620 113900
rect 185880 113880 186120 113900
rect 186380 113880 186620 113900
rect 186880 113880 187120 113900
rect 187380 113880 187620 113900
rect 187880 113880 188120 113900
rect 188380 113880 188620 113900
rect 188880 113880 189120 113900
rect 189380 113880 189620 113900
rect 189880 113880 190120 113900
rect 190380 113880 190620 113900
rect 190880 113880 191120 113900
rect 191380 113880 191620 113900
rect 191880 113880 192120 113900
rect 192380 113880 192620 113900
rect 192880 113880 193120 113900
rect 193380 113880 193620 113900
rect 193880 113880 194120 113900
rect 194380 113880 194620 113900
rect 194880 113880 195120 113900
rect 195380 113880 195620 113900
rect 195880 113880 196120 113900
rect 196380 113880 196620 113900
rect 196880 113880 197120 113900
rect 197380 113880 197620 113900
rect 197880 113880 198120 113900
rect 198380 113880 198620 113900
rect 198880 113880 199120 113900
rect 199380 113880 199620 113900
rect 199880 113880 200120 113900
rect 200380 113880 200620 113900
rect 200880 113880 201120 113900
rect 201380 113880 201620 113900
rect 201880 113880 202120 113900
rect 202380 113880 202620 113900
rect 202880 113880 203120 113900
rect 203380 113880 203620 113900
rect 203880 113880 204120 113900
rect 204380 113880 204620 113900
rect 204880 113880 205120 113900
rect 205380 113880 205620 113900
rect 205880 113880 206120 113900
rect 206380 113880 206620 113900
rect 206880 113880 207120 113900
rect 207380 113880 207620 113900
rect 207880 113880 208120 113900
rect 208380 113880 208620 113900
rect 208880 113880 209120 113900
rect 209380 113880 209620 113900
rect 209880 113880 210120 113900
rect 210380 113880 210620 113900
rect 210880 113880 211120 113900
rect 211380 113880 211620 113900
rect 211880 113880 212120 113900
rect 212380 113880 212620 113900
rect 212880 113880 213120 113900
rect 213380 113880 213620 113900
rect 213880 113880 214120 113900
rect 214380 113880 214620 113900
rect 214880 113880 215120 113900
rect 215380 113880 215620 113900
rect 215880 113880 216120 113900
rect 216380 113880 216620 113900
rect 216880 113880 217120 113900
rect 217380 113880 217620 113900
rect 217880 113880 218120 113900
rect 218380 113880 218620 113900
rect 218880 113880 219120 113900
rect 219380 113880 219620 113900
rect 219880 113880 220120 113900
rect 220380 113880 220620 113900
rect 220880 113880 221120 113900
rect 221380 113880 221620 113900
rect 221880 113880 222120 113900
rect 222380 113880 222620 113900
rect 222880 113880 223120 113900
rect 223380 113880 223620 113900
rect 223880 113880 224120 113900
rect 224380 113880 224620 113900
rect 224880 113880 225120 113900
rect 225380 113880 225620 113900
rect 225880 113880 226120 113900
rect 226380 113880 226620 113900
rect 226880 113880 227120 113900
rect 227380 113880 227620 113900
rect 227880 113880 228120 113900
rect 228380 113880 228620 113900
rect 228880 113880 229120 113900
rect 229380 113880 229620 113900
rect 229880 113880 230120 113900
rect 230380 113880 230620 113900
rect 230880 113880 231120 113900
rect 231380 113880 231620 113900
rect 231880 113880 232000 113900
rect 178000 113620 178100 113880
rect 178400 113620 178600 113880
rect 178900 113620 179100 113880
rect 179400 113620 179600 113880
rect 179900 113620 180100 113880
rect 180400 113620 180600 113880
rect 180900 113620 181100 113880
rect 181400 113620 181600 113880
rect 181900 113620 182100 113880
rect 182400 113620 182600 113880
rect 182900 113620 183100 113880
rect 183400 113620 183600 113880
rect 183900 113620 184100 113880
rect 184400 113620 184600 113880
rect 184900 113620 185100 113880
rect 185400 113620 185600 113880
rect 185900 113620 186100 113880
rect 186400 113620 186600 113880
rect 186900 113620 187100 113880
rect 187400 113620 187600 113880
rect 187900 113620 188100 113880
rect 188400 113620 188600 113880
rect 188900 113620 189100 113880
rect 189400 113620 189600 113880
rect 189900 113620 190100 113880
rect 190400 113620 190600 113880
rect 190900 113620 191100 113880
rect 191400 113620 191600 113880
rect 191900 113620 192100 113880
rect 192400 113620 192600 113880
rect 192900 113620 193100 113880
rect 193400 113620 193600 113880
rect 193900 113620 194100 113880
rect 194400 113620 194600 113880
rect 194900 113620 195100 113880
rect 195400 113620 195600 113880
rect 195900 113620 196100 113880
rect 196400 113620 196600 113880
rect 196900 113620 197100 113880
rect 197400 113620 197600 113880
rect 197900 113620 198100 113880
rect 198400 113620 198600 113880
rect 198900 113620 199100 113880
rect 199400 113620 199600 113880
rect 199900 113620 200100 113880
rect 200400 113620 200600 113880
rect 200900 113620 201100 113880
rect 201400 113620 201600 113880
rect 201900 113620 202100 113880
rect 202400 113620 202600 113880
rect 202900 113620 203100 113880
rect 203400 113620 203600 113880
rect 203900 113620 204100 113880
rect 204400 113620 204600 113880
rect 204900 113620 205100 113880
rect 205400 113620 205600 113880
rect 205900 113620 206100 113880
rect 206400 113620 206600 113880
rect 206900 113620 207100 113880
rect 207400 113620 207600 113880
rect 207900 113620 208100 113880
rect 208400 113620 208600 113880
rect 208900 113620 209100 113880
rect 209400 113620 209600 113880
rect 209900 113620 210100 113880
rect 210400 113620 210600 113880
rect 210900 113620 211100 113880
rect 211400 113620 211600 113880
rect 211900 113620 212100 113880
rect 212400 113620 212600 113880
rect 212900 113620 213100 113880
rect 213400 113620 213600 113880
rect 213900 113620 214100 113880
rect 214400 113620 214600 113880
rect 214900 113620 215100 113880
rect 215400 113620 215600 113880
rect 215900 113620 216100 113880
rect 216400 113620 216600 113880
rect 216900 113620 217100 113880
rect 217400 113620 217600 113880
rect 217900 113620 218100 113880
rect 218400 113620 218600 113880
rect 218900 113620 219100 113880
rect 219400 113620 219600 113880
rect 219900 113620 220100 113880
rect 220400 113620 220600 113880
rect 220900 113620 221100 113880
rect 221400 113620 221600 113880
rect 221900 113620 222100 113880
rect 222400 113620 222600 113880
rect 222900 113620 223100 113880
rect 223400 113620 223600 113880
rect 223900 113620 224100 113880
rect 224400 113620 224600 113880
rect 224900 113620 225100 113880
rect 225400 113620 225600 113880
rect 225900 113620 226100 113880
rect 226400 113620 226600 113880
rect 226900 113620 227100 113880
rect 227400 113620 227600 113880
rect 227900 113620 228100 113880
rect 228400 113620 228600 113880
rect 228900 113620 229100 113880
rect 229400 113620 229600 113880
rect 229900 113620 230100 113880
rect 230400 113620 230600 113880
rect 230900 113620 231100 113880
rect 231400 113620 231600 113880
rect 231900 113620 232000 113880
rect 178000 113600 178120 113620
rect 178380 113600 178620 113620
rect 178880 113600 179120 113620
rect 179380 113600 179620 113620
rect 179880 113600 180120 113620
rect 180380 113600 180620 113620
rect 180880 113600 181120 113620
rect 181380 113600 181620 113620
rect 181880 113600 182120 113620
rect 182380 113600 182620 113620
rect 182880 113600 183120 113620
rect 183380 113600 183620 113620
rect 183880 113600 184120 113620
rect 184380 113600 184620 113620
rect 184880 113600 185120 113620
rect 185380 113600 185620 113620
rect 185880 113600 186120 113620
rect 186380 113600 186620 113620
rect 186880 113600 187120 113620
rect 187380 113600 187620 113620
rect 187880 113600 188120 113620
rect 188380 113600 188620 113620
rect 188880 113600 189120 113620
rect 189380 113600 189620 113620
rect 189880 113600 190120 113620
rect 190380 113600 190620 113620
rect 190880 113600 191120 113620
rect 191380 113600 191620 113620
rect 191880 113600 192120 113620
rect 192380 113600 192620 113620
rect 192880 113600 193120 113620
rect 193380 113600 193620 113620
rect 193880 113600 194120 113620
rect 194380 113600 194620 113620
rect 194880 113600 195120 113620
rect 195380 113600 195620 113620
rect 195880 113600 196120 113620
rect 196380 113600 196620 113620
rect 196880 113600 197120 113620
rect 197380 113600 197620 113620
rect 197880 113600 198120 113620
rect 198380 113600 198620 113620
rect 198880 113600 199120 113620
rect 199380 113600 199620 113620
rect 199880 113600 200120 113620
rect 200380 113600 200620 113620
rect 200880 113600 201120 113620
rect 201380 113600 201620 113620
rect 201880 113600 202120 113620
rect 202380 113600 202620 113620
rect 202880 113600 203120 113620
rect 203380 113600 203620 113620
rect 203880 113600 204120 113620
rect 204380 113600 204620 113620
rect 204880 113600 205120 113620
rect 205380 113600 205620 113620
rect 205880 113600 206120 113620
rect 206380 113600 206620 113620
rect 206880 113600 207120 113620
rect 207380 113600 207620 113620
rect 207880 113600 208120 113620
rect 208380 113600 208620 113620
rect 208880 113600 209120 113620
rect 209380 113600 209620 113620
rect 209880 113600 210120 113620
rect 210380 113600 210620 113620
rect 210880 113600 211120 113620
rect 211380 113600 211620 113620
rect 211880 113600 212120 113620
rect 212380 113600 212620 113620
rect 212880 113600 213120 113620
rect 213380 113600 213620 113620
rect 213880 113600 214120 113620
rect 214380 113600 214620 113620
rect 214880 113600 215120 113620
rect 215380 113600 215620 113620
rect 215880 113600 216120 113620
rect 216380 113600 216620 113620
rect 216880 113600 217120 113620
rect 217380 113600 217620 113620
rect 217880 113600 218120 113620
rect 218380 113600 218620 113620
rect 218880 113600 219120 113620
rect 219380 113600 219620 113620
rect 219880 113600 220120 113620
rect 220380 113600 220620 113620
rect 220880 113600 221120 113620
rect 221380 113600 221620 113620
rect 221880 113600 222120 113620
rect 222380 113600 222620 113620
rect 222880 113600 223120 113620
rect 223380 113600 223620 113620
rect 223880 113600 224120 113620
rect 224380 113600 224620 113620
rect 224880 113600 225120 113620
rect 225380 113600 225620 113620
rect 225880 113600 226120 113620
rect 226380 113600 226620 113620
rect 226880 113600 227120 113620
rect 227380 113600 227620 113620
rect 227880 113600 228120 113620
rect 228380 113600 228620 113620
rect 228880 113600 229120 113620
rect 229380 113600 229620 113620
rect 229880 113600 230120 113620
rect 230380 113600 230620 113620
rect 230880 113600 231120 113620
rect 231380 113600 231620 113620
rect 231880 113600 232000 113620
rect 178000 113400 232000 113600
rect 178000 113380 178120 113400
rect 178380 113380 178620 113400
rect 178880 113380 179120 113400
rect 179380 113380 179620 113400
rect 179880 113380 180120 113400
rect 180380 113380 180620 113400
rect 180880 113380 181120 113400
rect 181380 113380 181620 113400
rect 181880 113380 182120 113400
rect 182380 113380 182620 113400
rect 182880 113380 183120 113400
rect 183380 113380 183620 113400
rect 183880 113380 184120 113400
rect 184380 113380 184620 113400
rect 184880 113380 185120 113400
rect 185380 113380 185620 113400
rect 185880 113380 186120 113400
rect 186380 113380 186620 113400
rect 186880 113380 187120 113400
rect 187380 113380 187620 113400
rect 187880 113380 188120 113400
rect 188380 113380 188620 113400
rect 188880 113380 189120 113400
rect 189380 113380 189620 113400
rect 189880 113380 190120 113400
rect 190380 113380 190620 113400
rect 190880 113380 191120 113400
rect 191380 113380 191620 113400
rect 191880 113380 192120 113400
rect 192380 113380 192620 113400
rect 192880 113380 193120 113400
rect 193380 113380 193620 113400
rect 193880 113380 194120 113400
rect 194380 113380 194620 113400
rect 194880 113380 195120 113400
rect 195380 113380 195620 113400
rect 195880 113380 196120 113400
rect 196380 113380 196620 113400
rect 196880 113380 197120 113400
rect 197380 113380 197620 113400
rect 197880 113380 198120 113400
rect 198380 113380 198620 113400
rect 198880 113380 199120 113400
rect 199380 113380 199620 113400
rect 199880 113380 200120 113400
rect 200380 113380 200620 113400
rect 200880 113380 201120 113400
rect 201380 113380 201620 113400
rect 201880 113380 202120 113400
rect 202380 113380 202620 113400
rect 202880 113380 203120 113400
rect 203380 113380 203620 113400
rect 203880 113380 204120 113400
rect 204380 113380 204620 113400
rect 204880 113380 205120 113400
rect 205380 113380 205620 113400
rect 205880 113380 206120 113400
rect 206380 113380 206620 113400
rect 206880 113380 207120 113400
rect 207380 113380 207620 113400
rect 207880 113380 208120 113400
rect 208380 113380 208620 113400
rect 208880 113380 209120 113400
rect 209380 113380 209620 113400
rect 209880 113380 210120 113400
rect 210380 113380 210620 113400
rect 210880 113380 211120 113400
rect 211380 113380 211620 113400
rect 211880 113380 212120 113400
rect 212380 113380 212620 113400
rect 212880 113380 213120 113400
rect 213380 113380 213620 113400
rect 213880 113380 214120 113400
rect 214380 113380 214620 113400
rect 214880 113380 215120 113400
rect 215380 113380 215620 113400
rect 215880 113380 216120 113400
rect 216380 113380 216620 113400
rect 216880 113380 217120 113400
rect 217380 113380 217620 113400
rect 217880 113380 218120 113400
rect 218380 113380 218620 113400
rect 218880 113380 219120 113400
rect 219380 113380 219620 113400
rect 219880 113380 220120 113400
rect 220380 113380 220620 113400
rect 220880 113380 221120 113400
rect 221380 113380 221620 113400
rect 221880 113380 222120 113400
rect 222380 113380 222620 113400
rect 222880 113380 223120 113400
rect 223380 113380 223620 113400
rect 223880 113380 224120 113400
rect 224380 113380 224620 113400
rect 224880 113380 225120 113400
rect 225380 113380 225620 113400
rect 225880 113380 226120 113400
rect 226380 113380 226620 113400
rect 226880 113380 227120 113400
rect 227380 113380 227620 113400
rect 227880 113380 228120 113400
rect 228380 113380 228620 113400
rect 228880 113380 229120 113400
rect 229380 113380 229620 113400
rect 229880 113380 230120 113400
rect 230380 113380 230620 113400
rect 230880 113380 231120 113400
rect 231380 113380 231620 113400
rect 231880 113380 232000 113400
rect 178000 113120 178100 113380
rect 178400 113120 178600 113380
rect 178900 113120 179100 113380
rect 179400 113120 179600 113380
rect 179900 113120 180100 113380
rect 180400 113120 180600 113380
rect 180900 113120 181100 113380
rect 181400 113120 181600 113380
rect 181900 113120 182100 113380
rect 182400 113120 182600 113380
rect 182900 113120 183100 113380
rect 183400 113120 183600 113380
rect 183900 113120 184100 113380
rect 184400 113120 184600 113380
rect 184900 113120 185100 113380
rect 185400 113120 185600 113380
rect 185900 113120 186100 113380
rect 186400 113120 186600 113380
rect 186900 113120 187100 113380
rect 187400 113120 187600 113380
rect 187900 113120 188100 113380
rect 188400 113120 188600 113380
rect 188900 113120 189100 113380
rect 189400 113120 189600 113380
rect 189900 113120 190100 113380
rect 190400 113120 190600 113380
rect 190900 113120 191100 113380
rect 191400 113120 191600 113380
rect 191900 113120 192100 113380
rect 192400 113120 192600 113380
rect 192900 113120 193100 113380
rect 193400 113120 193600 113380
rect 193900 113120 194100 113380
rect 194400 113120 194600 113380
rect 194900 113120 195100 113380
rect 195400 113120 195600 113380
rect 195900 113120 196100 113380
rect 196400 113120 196600 113380
rect 196900 113120 197100 113380
rect 197400 113120 197600 113380
rect 197900 113120 198100 113380
rect 198400 113120 198600 113380
rect 198900 113120 199100 113380
rect 199400 113120 199600 113380
rect 199900 113120 200100 113380
rect 200400 113120 200600 113380
rect 200900 113120 201100 113380
rect 201400 113120 201600 113380
rect 201900 113120 202100 113380
rect 202400 113120 202600 113380
rect 202900 113120 203100 113380
rect 203400 113120 203600 113380
rect 203900 113120 204100 113380
rect 204400 113120 204600 113380
rect 204900 113120 205100 113380
rect 205400 113120 205600 113380
rect 205900 113120 206100 113380
rect 206400 113120 206600 113380
rect 206900 113120 207100 113380
rect 207400 113120 207600 113380
rect 207900 113120 208100 113380
rect 208400 113120 208600 113380
rect 208900 113120 209100 113380
rect 209400 113120 209600 113380
rect 209900 113120 210100 113380
rect 210400 113120 210600 113380
rect 210900 113120 211100 113380
rect 211400 113120 211600 113380
rect 211900 113120 212100 113380
rect 212400 113120 212600 113380
rect 212900 113120 213100 113380
rect 213400 113120 213600 113380
rect 213900 113120 214100 113380
rect 214400 113120 214600 113380
rect 214900 113120 215100 113380
rect 215400 113120 215600 113380
rect 215900 113120 216100 113380
rect 216400 113120 216600 113380
rect 216900 113120 217100 113380
rect 217400 113120 217600 113380
rect 217900 113120 218100 113380
rect 218400 113120 218600 113380
rect 218900 113120 219100 113380
rect 219400 113120 219600 113380
rect 219900 113120 220100 113380
rect 220400 113120 220600 113380
rect 220900 113120 221100 113380
rect 221400 113120 221600 113380
rect 221900 113120 222100 113380
rect 222400 113120 222600 113380
rect 222900 113120 223100 113380
rect 223400 113120 223600 113380
rect 223900 113120 224100 113380
rect 224400 113120 224600 113380
rect 224900 113120 225100 113380
rect 225400 113120 225600 113380
rect 225900 113120 226100 113380
rect 226400 113120 226600 113380
rect 226900 113120 227100 113380
rect 227400 113120 227600 113380
rect 227900 113120 228100 113380
rect 228400 113120 228600 113380
rect 228900 113120 229100 113380
rect 229400 113120 229600 113380
rect 229900 113120 230100 113380
rect 230400 113120 230600 113380
rect 230900 113120 231100 113380
rect 231400 113120 231600 113380
rect 231900 113120 232000 113380
rect 178000 113100 178120 113120
rect 178380 113100 178620 113120
rect 178880 113100 179120 113120
rect 179380 113100 179620 113120
rect 179880 113100 180120 113120
rect 180380 113100 180620 113120
rect 180880 113100 181120 113120
rect 181380 113100 181620 113120
rect 181880 113100 182120 113120
rect 182380 113100 182620 113120
rect 182880 113100 183120 113120
rect 183380 113100 183620 113120
rect 183880 113100 184120 113120
rect 184380 113100 184620 113120
rect 184880 113100 185120 113120
rect 185380 113100 185620 113120
rect 185880 113100 186120 113120
rect 186380 113100 186620 113120
rect 186880 113100 187120 113120
rect 187380 113100 187620 113120
rect 187880 113100 188120 113120
rect 188380 113100 188620 113120
rect 188880 113100 189120 113120
rect 189380 113100 189620 113120
rect 189880 113100 190120 113120
rect 190380 113100 190620 113120
rect 190880 113100 191120 113120
rect 191380 113100 191620 113120
rect 191880 113100 192120 113120
rect 192380 113100 192620 113120
rect 192880 113100 193120 113120
rect 193380 113100 193620 113120
rect 193880 113100 194120 113120
rect 194380 113100 194620 113120
rect 194880 113100 195120 113120
rect 195380 113100 195620 113120
rect 195880 113100 196120 113120
rect 196380 113100 196620 113120
rect 196880 113100 197120 113120
rect 197380 113100 197620 113120
rect 197880 113100 198120 113120
rect 198380 113100 198620 113120
rect 198880 113100 199120 113120
rect 199380 113100 199620 113120
rect 199880 113100 200120 113120
rect 200380 113100 200620 113120
rect 200880 113100 201120 113120
rect 201380 113100 201620 113120
rect 201880 113100 202120 113120
rect 202380 113100 202620 113120
rect 202880 113100 203120 113120
rect 203380 113100 203620 113120
rect 203880 113100 204120 113120
rect 204380 113100 204620 113120
rect 204880 113100 205120 113120
rect 205380 113100 205620 113120
rect 205880 113100 206120 113120
rect 206380 113100 206620 113120
rect 206880 113100 207120 113120
rect 207380 113100 207620 113120
rect 207880 113100 208120 113120
rect 208380 113100 208620 113120
rect 208880 113100 209120 113120
rect 209380 113100 209620 113120
rect 209880 113100 210120 113120
rect 210380 113100 210620 113120
rect 210880 113100 211120 113120
rect 211380 113100 211620 113120
rect 211880 113100 212120 113120
rect 212380 113100 212620 113120
rect 212880 113100 213120 113120
rect 213380 113100 213620 113120
rect 213880 113100 214120 113120
rect 214380 113100 214620 113120
rect 214880 113100 215120 113120
rect 215380 113100 215620 113120
rect 215880 113100 216120 113120
rect 216380 113100 216620 113120
rect 216880 113100 217120 113120
rect 217380 113100 217620 113120
rect 217880 113100 218120 113120
rect 218380 113100 218620 113120
rect 218880 113100 219120 113120
rect 219380 113100 219620 113120
rect 219880 113100 220120 113120
rect 220380 113100 220620 113120
rect 220880 113100 221120 113120
rect 221380 113100 221620 113120
rect 221880 113100 222120 113120
rect 222380 113100 222620 113120
rect 222880 113100 223120 113120
rect 223380 113100 223620 113120
rect 223880 113100 224120 113120
rect 224380 113100 224620 113120
rect 224880 113100 225120 113120
rect 225380 113100 225620 113120
rect 225880 113100 226120 113120
rect 226380 113100 226620 113120
rect 226880 113100 227120 113120
rect 227380 113100 227620 113120
rect 227880 113100 228120 113120
rect 228380 113100 228620 113120
rect 228880 113100 229120 113120
rect 229380 113100 229620 113120
rect 229880 113100 230120 113120
rect 230380 113100 230620 113120
rect 230880 113100 231120 113120
rect 231380 113100 231620 113120
rect 231880 113100 232000 113120
rect 178000 112900 232000 113100
rect 178000 112880 178120 112900
rect 178380 112880 178620 112900
rect 178880 112880 179120 112900
rect 179380 112880 179620 112900
rect 179880 112880 180120 112900
rect 180380 112880 180620 112900
rect 180880 112880 181120 112900
rect 181380 112880 181620 112900
rect 181880 112880 182120 112900
rect 182380 112880 182620 112900
rect 182880 112880 183120 112900
rect 183380 112880 183620 112900
rect 183880 112880 184120 112900
rect 184380 112880 184620 112900
rect 184880 112880 185120 112900
rect 185380 112880 185620 112900
rect 185880 112880 186120 112900
rect 186380 112880 186620 112900
rect 186880 112880 187120 112900
rect 187380 112880 187620 112900
rect 187880 112880 188120 112900
rect 188380 112880 188620 112900
rect 188880 112880 189120 112900
rect 189380 112880 189620 112900
rect 189880 112880 190120 112900
rect 190380 112880 190620 112900
rect 190880 112880 191120 112900
rect 191380 112880 191620 112900
rect 191880 112880 192120 112900
rect 192380 112880 192620 112900
rect 192880 112880 193120 112900
rect 193380 112880 193620 112900
rect 193880 112880 194120 112900
rect 194380 112880 194620 112900
rect 194880 112880 195120 112900
rect 195380 112880 195620 112900
rect 195880 112880 196120 112900
rect 196380 112880 196620 112900
rect 196880 112880 197120 112900
rect 197380 112880 197620 112900
rect 197880 112880 198120 112900
rect 198380 112880 198620 112900
rect 198880 112880 199120 112900
rect 199380 112880 199620 112900
rect 199880 112880 200120 112900
rect 200380 112880 200620 112900
rect 200880 112880 201120 112900
rect 201380 112880 201620 112900
rect 201880 112880 202120 112900
rect 202380 112880 202620 112900
rect 202880 112880 203120 112900
rect 203380 112880 203620 112900
rect 203880 112880 204120 112900
rect 204380 112880 204620 112900
rect 204880 112880 205120 112900
rect 205380 112880 205620 112900
rect 205880 112880 206120 112900
rect 206380 112880 206620 112900
rect 206880 112880 207120 112900
rect 207380 112880 207620 112900
rect 207880 112880 208120 112900
rect 208380 112880 208620 112900
rect 208880 112880 209120 112900
rect 209380 112880 209620 112900
rect 209880 112880 210120 112900
rect 210380 112880 210620 112900
rect 210880 112880 211120 112900
rect 211380 112880 211620 112900
rect 211880 112880 212120 112900
rect 212380 112880 212620 112900
rect 212880 112880 213120 112900
rect 213380 112880 213620 112900
rect 213880 112880 214120 112900
rect 214380 112880 214620 112900
rect 214880 112880 215120 112900
rect 215380 112880 215620 112900
rect 215880 112880 216120 112900
rect 216380 112880 216620 112900
rect 216880 112880 217120 112900
rect 217380 112880 217620 112900
rect 217880 112880 218120 112900
rect 218380 112880 218620 112900
rect 218880 112880 219120 112900
rect 219380 112880 219620 112900
rect 219880 112880 220120 112900
rect 220380 112880 220620 112900
rect 220880 112880 221120 112900
rect 221380 112880 221620 112900
rect 221880 112880 222120 112900
rect 222380 112880 222620 112900
rect 222880 112880 223120 112900
rect 223380 112880 223620 112900
rect 223880 112880 224120 112900
rect 224380 112880 224620 112900
rect 224880 112880 225120 112900
rect 225380 112880 225620 112900
rect 225880 112880 226120 112900
rect 226380 112880 226620 112900
rect 226880 112880 227120 112900
rect 227380 112880 227620 112900
rect 227880 112880 228120 112900
rect 228380 112880 228620 112900
rect 228880 112880 229120 112900
rect 229380 112880 229620 112900
rect 229880 112880 230120 112900
rect 230380 112880 230620 112900
rect 230880 112880 231120 112900
rect 231380 112880 231620 112900
rect 231880 112880 232000 112900
rect 178000 112620 178100 112880
rect 178400 112620 178600 112880
rect 178900 112620 179100 112880
rect 179400 112620 179600 112880
rect 179900 112620 180100 112880
rect 180400 112620 180600 112880
rect 180900 112620 181100 112880
rect 181400 112620 181600 112880
rect 181900 112620 182100 112880
rect 182400 112620 182600 112880
rect 182900 112620 183100 112880
rect 183400 112620 183600 112880
rect 183900 112620 184100 112880
rect 184400 112620 184600 112880
rect 184900 112620 185100 112880
rect 185400 112620 185600 112880
rect 185900 112620 186100 112880
rect 186400 112620 186600 112880
rect 186900 112620 187100 112880
rect 187400 112620 187600 112880
rect 187900 112620 188100 112880
rect 188400 112620 188600 112880
rect 188900 112620 189100 112880
rect 189400 112620 189600 112880
rect 189900 112620 190100 112880
rect 190400 112620 190600 112880
rect 190900 112620 191100 112880
rect 191400 112620 191600 112880
rect 191900 112620 192100 112880
rect 192400 112620 192600 112880
rect 192900 112620 193100 112880
rect 193400 112620 193600 112880
rect 193900 112620 194100 112880
rect 194400 112620 194600 112880
rect 194900 112620 195100 112880
rect 195400 112620 195600 112880
rect 195900 112620 196100 112880
rect 196400 112620 196600 112880
rect 196900 112620 197100 112880
rect 197400 112620 197600 112880
rect 197900 112620 198100 112880
rect 198400 112620 198600 112880
rect 198900 112620 199100 112880
rect 199400 112620 199600 112880
rect 199900 112620 200100 112880
rect 200400 112620 200600 112880
rect 200900 112620 201100 112880
rect 201400 112620 201600 112880
rect 201900 112620 202100 112880
rect 202400 112620 202600 112880
rect 202900 112620 203100 112880
rect 203400 112620 203600 112880
rect 203900 112620 204100 112880
rect 204400 112620 204600 112880
rect 204900 112620 205100 112880
rect 205400 112620 205600 112880
rect 205900 112620 206100 112880
rect 206400 112620 206600 112880
rect 206900 112620 207100 112880
rect 207400 112620 207600 112880
rect 207900 112620 208100 112880
rect 208400 112620 208600 112880
rect 208900 112620 209100 112880
rect 209400 112620 209600 112880
rect 209900 112620 210100 112880
rect 210400 112620 210600 112880
rect 210900 112620 211100 112880
rect 211400 112620 211600 112880
rect 211900 112620 212100 112880
rect 212400 112620 212600 112880
rect 212900 112620 213100 112880
rect 213400 112620 213600 112880
rect 213900 112620 214100 112880
rect 214400 112620 214600 112880
rect 214900 112620 215100 112880
rect 215400 112620 215600 112880
rect 215900 112620 216100 112880
rect 216400 112620 216600 112880
rect 216900 112620 217100 112880
rect 217400 112620 217600 112880
rect 217900 112620 218100 112880
rect 218400 112620 218600 112880
rect 218900 112620 219100 112880
rect 219400 112620 219600 112880
rect 219900 112620 220100 112880
rect 220400 112620 220600 112880
rect 220900 112620 221100 112880
rect 221400 112620 221600 112880
rect 221900 112620 222100 112880
rect 222400 112620 222600 112880
rect 222900 112620 223100 112880
rect 223400 112620 223600 112880
rect 223900 112620 224100 112880
rect 224400 112620 224600 112880
rect 224900 112620 225100 112880
rect 225400 112620 225600 112880
rect 225900 112620 226100 112880
rect 226400 112620 226600 112880
rect 226900 112620 227100 112880
rect 227400 112620 227600 112880
rect 227900 112620 228100 112880
rect 228400 112620 228600 112880
rect 228900 112620 229100 112880
rect 229400 112620 229600 112880
rect 229900 112620 230100 112880
rect 230400 112620 230600 112880
rect 230900 112620 231100 112880
rect 231400 112620 231600 112880
rect 231900 112620 232000 112880
rect 178000 112600 178120 112620
rect 178380 112600 178620 112620
rect 178880 112600 179120 112620
rect 179380 112600 179620 112620
rect 179880 112600 180120 112620
rect 180380 112600 180620 112620
rect 180880 112600 181120 112620
rect 181380 112600 181620 112620
rect 181880 112600 182120 112620
rect 182380 112600 182620 112620
rect 182880 112600 183120 112620
rect 183380 112600 183620 112620
rect 183880 112600 184120 112620
rect 184380 112600 184620 112620
rect 184880 112600 185120 112620
rect 185380 112600 185620 112620
rect 185880 112600 186120 112620
rect 186380 112600 186620 112620
rect 186880 112600 187120 112620
rect 187380 112600 187620 112620
rect 187880 112600 188120 112620
rect 188380 112600 188620 112620
rect 188880 112600 189120 112620
rect 189380 112600 189620 112620
rect 189880 112600 190120 112620
rect 190380 112600 190620 112620
rect 190880 112600 191120 112620
rect 191380 112600 191620 112620
rect 191880 112600 192120 112620
rect 192380 112600 192620 112620
rect 192880 112600 193120 112620
rect 193380 112600 193620 112620
rect 193880 112600 194120 112620
rect 194380 112600 194620 112620
rect 194880 112600 195120 112620
rect 195380 112600 195620 112620
rect 195880 112600 196120 112620
rect 196380 112600 196620 112620
rect 196880 112600 197120 112620
rect 197380 112600 197620 112620
rect 197880 112600 198120 112620
rect 198380 112600 198620 112620
rect 198880 112600 199120 112620
rect 199380 112600 199620 112620
rect 199880 112600 200120 112620
rect 200380 112600 200620 112620
rect 200880 112600 201120 112620
rect 201380 112600 201620 112620
rect 201880 112600 202120 112620
rect 202380 112600 202620 112620
rect 202880 112600 203120 112620
rect 203380 112600 203620 112620
rect 203880 112600 204120 112620
rect 204380 112600 204620 112620
rect 204880 112600 205120 112620
rect 205380 112600 205620 112620
rect 205880 112600 206120 112620
rect 206380 112600 206620 112620
rect 206880 112600 207120 112620
rect 207380 112600 207620 112620
rect 207880 112600 208120 112620
rect 208380 112600 208620 112620
rect 208880 112600 209120 112620
rect 209380 112600 209620 112620
rect 209880 112600 210120 112620
rect 210380 112600 210620 112620
rect 210880 112600 211120 112620
rect 211380 112600 211620 112620
rect 211880 112600 212120 112620
rect 212380 112600 212620 112620
rect 212880 112600 213120 112620
rect 213380 112600 213620 112620
rect 213880 112600 214120 112620
rect 214380 112600 214620 112620
rect 214880 112600 215120 112620
rect 215380 112600 215620 112620
rect 215880 112600 216120 112620
rect 216380 112600 216620 112620
rect 216880 112600 217120 112620
rect 217380 112600 217620 112620
rect 217880 112600 218120 112620
rect 218380 112600 218620 112620
rect 218880 112600 219120 112620
rect 219380 112600 219620 112620
rect 219880 112600 220120 112620
rect 220380 112600 220620 112620
rect 220880 112600 221120 112620
rect 221380 112600 221620 112620
rect 221880 112600 222120 112620
rect 222380 112600 222620 112620
rect 222880 112600 223120 112620
rect 223380 112600 223620 112620
rect 223880 112600 224120 112620
rect 224380 112600 224620 112620
rect 224880 112600 225120 112620
rect 225380 112600 225620 112620
rect 225880 112600 226120 112620
rect 226380 112600 226620 112620
rect 226880 112600 227120 112620
rect 227380 112600 227620 112620
rect 227880 112600 228120 112620
rect 228380 112600 228620 112620
rect 228880 112600 229120 112620
rect 229380 112600 229620 112620
rect 229880 112600 230120 112620
rect 230380 112600 230620 112620
rect 230880 112600 231120 112620
rect 231380 112600 231620 112620
rect 231880 112600 232000 112620
rect 178000 112400 232000 112600
rect 178000 112380 178120 112400
rect 178380 112380 178620 112400
rect 178880 112380 179120 112400
rect 179380 112380 179620 112400
rect 179880 112380 180120 112400
rect 180380 112380 180620 112400
rect 180880 112380 181120 112400
rect 181380 112380 181620 112400
rect 181880 112380 182120 112400
rect 182380 112380 182620 112400
rect 182880 112380 183120 112400
rect 183380 112380 183620 112400
rect 183880 112380 184120 112400
rect 184380 112380 184620 112400
rect 184880 112380 185120 112400
rect 185380 112380 185620 112400
rect 185880 112380 186120 112400
rect 186380 112380 186620 112400
rect 186880 112380 187120 112400
rect 187380 112380 187620 112400
rect 187880 112380 188120 112400
rect 188380 112380 188620 112400
rect 188880 112380 189120 112400
rect 189380 112380 189620 112400
rect 189880 112380 190120 112400
rect 190380 112380 190620 112400
rect 190880 112380 191120 112400
rect 191380 112380 191620 112400
rect 191880 112380 192120 112400
rect 192380 112380 192620 112400
rect 192880 112380 193120 112400
rect 193380 112380 193620 112400
rect 193880 112380 194120 112400
rect 194380 112380 194620 112400
rect 194880 112380 195120 112400
rect 195380 112380 195620 112400
rect 195880 112380 196120 112400
rect 196380 112380 196620 112400
rect 196880 112380 197120 112400
rect 197380 112380 197620 112400
rect 197880 112380 198120 112400
rect 198380 112380 198620 112400
rect 198880 112380 199120 112400
rect 199380 112380 199620 112400
rect 199880 112380 200120 112400
rect 200380 112380 200620 112400
rect 200880 112380 201120 112400
rect 201380 112380 201620 112400
rect 201880 112380 202120 112400
rect 202380 112380 202620 112400
rect 202880 112380 203120 112400
rect 203380 112380 203620 112400
rect 203880 112380 204120 112400
rect 204380 112380 204620 112400
rect 204880 112380 205120 112400
rect 205380 112380 205620 112400
rect 205880 112380 206120 112400
rect 206380 112380 206620 112400
rect 206880 112380 207120 112400
rect 207380 112380 207620 112400
rect 207880 112380 208120 112400
rect 208380 112380 208620 112400
rect 208880 112380 209120 112400
rect 209380 112380 209620 112400
rect 209880 112380 210120 112400
rect 210380 112380 210620 112400
rect 210880 112380 211120 112400
rect 211380 112380 211620 112400
rect 211880 112380 212120 112400
rect 212380 112380 212620 112400
rect 212880 112380 213120 112400
rect 213380 112380 213620 112400
rect 213880 112380 214120 112400
rect 214380 112380 214620 112400
rect 214880 112380 215120 112400
rect 215380 112380 215620 112400
rect 215880 112380 216120 112400
rect 216380 112380 216620 112400
rect 216880 112380 217120 112400
rect 217380 112380 217620 112400
rect 217880 112380 218120 112400
rect 218380 112380 218620 112400
rect 218880 112380 219120 112400
rect 219380 112380 219620 112400
rect 219880 112380 220120 112400
rect 220380 112380 220620 112400
rect 220880 112380 221120 112400
rect 221380 112380 221620 112400
rect 221880 112380 222120 112400
rect 222380 112380 222620 112400
rect 222880 112380 223120 112400
rect 223380 112380 223620 112400
rect 223880 112380 224120 112400
rect 224380 112380 224620 112400
rect 224880 112380 225120 112400
rect 225380 112380 225620 112400
rect 225880 112380 226120 112400
rect 226380 112380 226620 112400
rect 226880 112380 227120 112400
rect 227380 112380 227620 112400
rect 227880 112380 228120 112400
rect 228380 112380 228620 112400
rect 228880 112380 229120 112400
rect 229380 112380 229620 112400
rect 229880 112380 230120 112400
rect 230380 112380 230620 112400
rect 230880 112380 231120 112400
rect 231380 112380 231620 112400
rect 231880 112380 232000 112400
rect 178000 112120 178100 112380
rect 178400 112120 178600 112380
rect 178900 112120 179100 112380
rect 179400 112120 179600 112380
rect 179900 112120 180100 112380
rect 180400 112120 180600 112380
rect 180900 112120 181100 112380
rect 181400 112120 181600 112380
rect 181900 112120 182100 112380
rect 182400 112120 182600 112380
rect 182900 112120 183100 112380
rect 183400 112120 183600 112380
rect 183900 112120 184100 112380
rect 184400 112120 184600 112380
rect 184900 112120 185100 112380
rect 185400 112120 185600 112380
rect 185900 112120 186100 112380
rect 186400 112120 186600 112380
rect 186900 112120 187100 112380
rect 187400 112120 187600 112380
rect 187900 112120 188100 112380
rect 188400 112120 188600 112380
rect 188900 112120 189100 112380
rect 189400 112120 189600 112380
rect 189900 112120 190100 112380
rect 190400 112120 190600 112380
rect 190900 112120 191100 112380
rect 191400 112120 191600 112380
rect 191900 112120 192100 112380
rect 192400 112120 192600 112380
rect 192900 112120 193100 112380
rect 193400 112120 193600 112380
rect 193900 112120 194100 112380
rect 194400 112120 194600 112380
rect 194900 112120 195100 112380
rect 195400 112120 195600 112380
rect 195900 112120 196100 112380
rect 196400 112120 196600 112380
rect 196900 112120 197100 112380
rect 197400 112120 197600 112380
rect 197900 112120 198100 112380
rect 198400 112120 198600 112380
rect 198900 112120 199100 112380
rect 199400 112120 199600 112380
rect 199900 112120 200100 112380
rect 200400 112120 200600 112380
rect 200900 112120 201100 112380
rect 201400 112120 201600 112380
rect 201900 112120 202100 112380
rect 202400 112120 202600 112380
rect 202900 112120 203100 112380
rect 203400 112120 203600 112380
rect 203900 112120 204100 112380
rect 204400 112120 204600 112380
rect 204900 112120 205100 112380
rect 205400 112120 205600 112380
rect 205900 112120 206100 112380
rect 206400 112120 206600 112380
rect 206900 112120 207100 112380
rect 207400 112120 207600 112380
rect 207900 112120 208100 112380
rect 208400 112120 208600 112380
rect 208900 112120 209100 112380
rect 209400 112120 209600 112380
rect 209900 112120 210100 112380
rect 210400 112120 210600 112380
rect 210900 112120 211100 112380
rect 211400 112120 211600 112380
rect 211900 112120 212100 112380
rect 212400 112120 212600 112380
rect 212900 112120 213100 112380
rect 213400 112120 213600 112380
rect 213900 112120 214100 112380
rect 214400 112120 214600 112380
rect 214900 112120 215100 112380
rect 215400 112120 215600 112380
rect 215900 112120 216100 112380
rect 216400 112120 216600 112380
rect 216900 112120 217100 112380
rect 217400 112120 217600 112380
rect 217900 112120 218100 112380
rect 218400 112120 218600 112380
rect 218900 112120 219100 112380
rect 219400 112120 219600 112380
rect 219900 112120 220100 112380
rect 220400 112120 220600 112380
rect 220900 112120 221100 112380
rect 221400 112120 221600 112380
rect 221900 112120 222100 112380
rect 222400 112120 222600 112380
rect 222900 112120 223100 112380
rect 223400 112120 223600 112380
rect 223900 112120 224100 112380
rect 224400 112120 224600 112380
rect 224900 112120 225100 112380
rect 225400 112120 225600 112380
rect 225900 112120 226100 112380
rect 226400 112120 226600 112380
rect 226900 112120 227100 112380
rect 227400 112120 227600 112380
rect 227900 112120 228100 112380
rect 228400 112120 228600 112380
rect 228900 112120 229100 112380
rect 229400 112120 229600 112380
rect 229900 112120 230100 112380
rect 230400 112120 230600 112380
rect 230900 112120 231100 112380
rect 231400 112120 231600 112380
rect 231900 112120 232000 112380
rect 178000 112100 178120 112120
rect 178380 112100 178620 112120
rect 178880 112100 179120 112120
rect 179380 112100 179620 112120
rect 179880 112100 180120 112120
rect 180380 112100 180620 112120
rect 180880 112100 181120 112120
rect 181380 112100 181620 112120
rect 181880 112100 182120 112120
rect 182380 112100 182620 112120
rect 182880 112100 183120 112120
rect 183380 112100 183620 112120
rect 183880 112100 184120 112120
rect 184380 112100 184620 112120
rect 184880 112100 185120 112120
rect 185380 112100 185620 112120
rect 185880 112100 186120 112120
rect 186380 112100 186620 112120
rect 186880 112100 187120 112120
rect 187380 112100 187620 112120
rect 187880 112100 188120 112120
rect 188380 112100 188620 112120
rect 188880 112100 189120 112120
rect 189380 112100 189620 112120
rect 189880 112100 190120 112120
rect 190380 112100 190620 112120
rect 190880 112100 191120 112120
rect 191380 112100 191620 112120
rect 191880 112100 192120 112120
rect 192380 112100 192620 112120
rect 192880 112100 193120 112120
rect 193380 112100 193620 112120
rect 193880 112100 194120 112120
rect 194380 112100 194620 112120
rect 194880 112100 195120 112120
rect 195380 112100 195620 112120
rect 195880 112100 196120 112120
rect 196380 112100 196620 112120
rect 196880 112100 197120 112120
rect 197380 112100 197620 112120
rect 197880 112100 198120 112120
rect 198380 112100 198620 112120
rect 198880 112100 199120 112120
rect 199380 112100 199620 112120
rect 199880 112100 200120 112120
rect 200380 112100 200620 112120
rect 200880 112100 201120 112120
rect 201380 112100 201620 112120
rect 201880 112100 202120 112120
rect 202380 112100 202620 112120
rect 202880 112100 203120 112120
rect 203380 112100 203620 112120
rect 203880 112100 204120 112120
rect 204380 112100 204620 112120
rect 204880 112100 205120 112120
rect 205380 112100 205620 112120
rect 205880 112100 206120 112120
rect 206380 112100 206620 112120
rect 206880 112100 207120 112120
rect 207380 112100 207620 112120
rect 207880 112100 208120 112120
rect 208380 112100 208620 112120
rect 208880 112100 209120 112120
rect 209380 112100 209620 112120
rect 209880 112100 210120 112120
rect 210380 112100 210620 112120
rect 210880 112100 211120 112120
rect 211380 112100 211620 112120
rect 211880 112100 212120 112120
rect 212380 112100 212620 112120
rect 212880 112100 213120 112120
rect 213380 112100 213620 112120
rect 213880 112100 214120 112120
rect 214380 112100 214620 112120
rect 214880 112100 215120 112120
rect 215380 112100 215620 112120
rect 215880 112100 216120 112120
rect 216380 112100 216620 112120
rect 216880 112100 217120 112120
rect 217380 112100 217620 112120
rect 217880 112100 218120 112120
rect 218380 112100 218620 112120
rect 218880 112100 219120 112120
rect 219380 112100 219620 112120
rect 219880 112100 220120 112120
rect 220380 112100 220620 112120
rect 220880 112100 221120 112120
rect 221380 112100 221620 112120
rect 221880 112100 222120 112120
rect 222380 112100 222620 112120
rect 222880 112100 223120 112120
rect 223380 112100 223620 112120
rect 223880 112100 224120 112120
rect 224380 112100 224620 112120
rect 224880 112100 225120 112120
rect 225380 112100 225620 112120
rect 225880 112100 226120 112120
rect 226380 112100 226620 112120
rect 226880 112100 227120 112120
rect 227380 112100 227620 112120
rect 227880 112100 228120 112120
rect 228380 112100 228620 112120
rect 228880 112100 229120 112120
rect 229380 112100 229620 112120
rect 229880 112100 230120 112120
rect 230380 112100 230620 112120
rect 230880 112100 231120 112120
rect 231380 112100 231620 112120
rect 231880 112100 232000 112120
rect 178000 111900 232000 112100
rect 178000 111880 178120 111900
rect 178380 111880 178620 111900
rect 178880 111880 179120 111900
rect 179380 111880 179620 111900
rect 179880 111880 180120 111900
rect 180380 111880 180620 111900
rect 180880 111880 181120 111900
rect 181380 111880 181620 111900
rect 181880 111880 182120 111900
rect 182380 111880 182620 111900
rect 182880 111880 183120 111900
rect 183380 111880 183620 111900
rect 183880 111880 184120 111900
rect 184380 111880 184620 111900
rect 184880 111880 185120 111900
rect 185380 111880 185620 111900
rect 185880 111880 186120 111900
rect 186380 111880 186620 111900
rect 186880 111880 187120 111900
rect 187380 111880 187620 111900
rect 187880 111880 188120 111900
rect 188380 111880 188620 111900
rect 188880 111880 189120 111900
rect 189380 111880 189620 111900
rect 189880 111880 190120 111900
rect 190380 111880 190620 111900
rect 190880 111880 191120 111900
rect 191380 111880 191620 111900
rect 191880 111880 192120 111900
rect 192380 111880 192620 111900
rect 192880 111880 193120 111900
rect 193380 111880 193620 111900
rect 193880 111880 194120 111900
rect 194380 111880 194620 111900
rect 194880 111880 195120 111900
rect 195380 111880 195620 111900
rect 195880 111880 196120 111900
rect 196380 111880 196620 111900
rect 196880 111880 197120 111900
rect 197380 111880 197620 111900
rect 197880 111880 198120 111900
rect 198380 111880 198620 111900
rect 198880 111880 199120 111900
rect 199380 111880 199620 111900
rect 199880 111880 200120 111900
rect 200380 111880 200620 111900
rect 200880 111880 201120 111900
rect 201380 111880 201620 111900
rect 201880 111880 202120 111900
rect 202380 111880 202620 111900
rect 202880 111880 203120 111900
rect 203380 111880 203620 111900
rect 203880 111880 204120 111900
rect 204380 111880 204620 111900
rect 204880 111880 205120 111900
rect 205380 111880 205620 111900
rect 205880 111880 206120 111900
rect 206380 111880 206620 111900
rect 206880 111880 207120 111900
rect 207380 111880 207620 111900
rect 207880 111880 208120 111900
rect 208380 111880 208620 111900
rect 208880 111880 209120 111900
rect 209380 111880 209620 111900
rect 209880 111880 210120 111900
rect 210380 111880 210620 111900
rect 210880 111880 211120 111900
rect 211380 111880 211620 111900
rect 211880 111880 212120 111900
rect 212380 111880 212620 111900
rect 212880 111880 213120 111900
rect 213380 111880 213620 111900
rect 213880 111880 214120 111900
rect 214380 111880 214620 111900
rect 214880 111880 215120 111900
rect 215380 111880 215620 111900
rect 215880 111880 216120 111900
rect 216380 111880 216620 111900
rect 216880 111880 217120 111900
rect 217380 111880 217620 111900
rect 217880 111880 218120 111900
rect 218380 111880 218620 111900
rect 218880 111880 219120 111900
rect 219380 111880 219620 111900
rect 219880 111880 220120 111900
rect 220380 111880 220620 111900
rect 220880 111880 221120 111900
rect 221380 111880 221620 111900
rect 221880 111880 222120 111900
rect 222380 111880 222620 111900
rect 222880 111880 223120 111900
rect 223380 111880 223620 111900
rect 223880 111880 224120 111900
rect 224380 111880 224620 111900
rect 224880 111880 225120 111900
rect 225380 111880 225620 111900
rect 225880 111880 226120 111900
rect 226380 111880 226620 111900
rect 226880 111880 227120 111900
rect 227380 111880 227620 111900
rect 227880 111880 228120 111900
rect 228380 111880 228620 111900
rect 228880 111880 229120 111900
rect 229380 111880 229620 111900
rect 229880 111880 230120 111900
rect 230380 111880 230620 111900
rect 230880 111880 231120 111900
rect 231380 111880 231620 111900
rect 231880 111880 232000 111900
rect 178000 111620 178100 111880
rect 178400 111620 178600 111880
rect 178900 111620 179100 111880
rect 179400 111620 179600 111880
rect 179900 111620 180100 111880
rect 180400 111620 180600 111880
rect 180900 111620 181100 111880
rect 181400 111620 181600 111880
rect 181900 111620 182100 111880
rect 182400 111620 182600 111880
rect 182900 111620 183100 111880
rect 183400 111620 183600 111880
rect 183900 111620 184100 111880
rect 184400 111620 184600 111880
rect 184900 111620 185100 111880
rect 185400 111620 185600 111880
rect 185900 111620 186100 111880
rect 186400 111620 186600 111880
rect 186900 111620 187100 111880
rect 187400 111620 187600 111880
rect 187900 111620 188100 111880
rect 188400 111620 188600 111880
rect 188900 111620 189100 111880
rect 189400 111620 189600 111880
rect 189900 111620 190100 111880
rect 190400 111620 190600 111880
rect 190900 111620 191100 111880
rect 191400 111620 191600 111880
rect 191900 111620 192100 111880
rect 192400 111620 192600 111880
rect 192900 111620 193100 111880
rect 193400 111620 193600 111880
rect 193900 111620 194100 111880
rect 194400 111620 194600 111880
rect 194900 111620 195100 111880
rect 195400 111620 195600 111880
rect 195900 111620 196100 111880
rect 196400 111620 196600 111880
rect 196900 111620 197100 111880
rect 197400 111620 197600 111880
rect 197900 111620 198100 111880
rect 198400 111620 198600 111880
rect 198900 111620 199100 111880
rect 199400 111620 199600 111880
rect 199900 111620 200100 111880
rect 200400 111620 200600 111880
rect 200900 111620 201100 111880
rect 201400 111620 201600 111880
rect 201900 111620 202100 111880
rect 202400 111620 202600 111880
rect 202900 111620 203100 111880
rect 203400 111620 203600 111880
rect 203900 111620 204100 111880
rect 204400 111620 204600 111880
rect 204900 111620 205100 111880
rect 205400 111620 205600 111880
rect 205900 111620 206100 111880
rect 206400 111620 206600 111880
rect 206900 111620 207100 111880
rect 207400 111620 207600 111880
rect 207900 111620 208100 111880
rect 208400 111620 208600 111880
rect 208900 111620 209100 111880
rect 209400 111620 209600 111880
rect 209900 111620 210100 111880
rect 210400 111620 210600 111880
rect 210900 111620 211100 111880
rect 211400 111620 211600 111880
rect 211900 111620 212100 111880
rect 212400 111620 212600 111880
rect 212900 111620 213100 111880
rect 213400 111620 213600 111880
rect 213900 111620 214100 111880
rect 214400 111620 214600 111880
rect 214900 111620 215100 111880
rect 215400 111620 215600 111880
rect 215900 111620 216100 111880
rect 216400 111620 216600 111880
rect 216900 111620 217100 111880
rect 217400 111620 217600 111880
rect 217900 111620 218100 111880
rect 218400 111620 218600 111880
rect 218900 111620 219100 111880
rect 219400 111620 219600 111880
rect 219900 111620 220100 111880
rect 220400 111620 220600 111880
rect 220900 111620 221100 111880
rect 221400 111620 221600 111880
rect 221900 111620 222100 111880
rect 222400 111620 222600 111880
rect 222900 111620 223100 111880
rect 223400 111620 223600 111880
rect 223900 111620 224100 111880
rect 224400 111620 224600 111880
rect 224900 111620 225100 111880
rect 225400 111620 225600 111880
rect 225900 111620 226100 111880
rect 226400 111620 226600 111880
rect 226900 111620 227100 111880
rect 227400 111620 227600 111880
rect 227900 111620 228100 111880
rect 228400 111620 228600 111880
rect 228900 111620 229100 111880
rect 229400 111620 229600 111880
rect 229900 111620 230100 111880
rect 230400 111620 230600 111880
rect 230900 111620 231100 111880
rect 231400 111620 231600 111880
rect 231900 111620 232000 111880
rect 178000 111600 178120 111620
rect 178380 111600 178620 111620
rect 178880 111600 179120 111620
rect 179380 111600 179620 111620
rect 179880 111600 180120 111620
rect 180380 111600 180620 111620
rect 180880 111600 181120 111620
rect 181380 111600 181620 111620
rect 181880 111600 182120 111620
rect 182380 111600 182620 111620
rect 182880 111600 183120 111620
rect 183380 111600 183620 111620
rect 183880 111600 184120 111620
rect 184380 111600 184620 111620
rect 184880 111600 185120 111620
rect 185380 111600 185620 111620
rect 185880 111600 186120 111620
rect 186380 111600 186620 111620
rect 186880 111600 187120 111620
rect 187380 111600 187620 111620
rect 187880 111600 188120 111620
rect 188380 111600 188620 111620
rect 188880 111600 189120 111620
rect 189380 111600 189620 111620
rect 189880 111600 190120 111620
rect 190380 111600 190620 111620
rect 190880 111600 191120 111620
rect 191380 111600 191620 111620
rect 191880 111600 192120 111620
rect 192380 111600 192620 111620
rect 192880 111600 193120 111620
rect 193380 111600 193620 111620
rect 193880 111600 194120 111620
rect 194380 111600 194620 111620
rect 194880 111600 195120 111620
rect 195380 111600 195620 111620
rect 195880 111600 196120 111620
rect 196380 111600 196620 111620
rect 196880 111600 197120 111620
rect 197380 111600 197620 111620
rect 197880 111600 198120 111620
rect 198380 111600 198620 111620
rect 198880 111600 199120 111620
rect 199380 111600 199620 111620
rect 199880 111600 200120 111620
rect 200380 111600 200620 111620
rect 200880 111600 201120 111620
rect 201380 111600 201620 111620
rect 201880 111600 202120 111620
rect 202380 111600 202620 111620
rect 202880 111600 203120 111620
rect 203380 111600 203620 111620
rect 203880 111600 204120 111620
rect 204380 111600 204620 111620
rect 204880 111600 205120 111620
rect 205380 111600 205620 111620
rect 205880 111600 206120 111620
rect 206380 111600 206620 111620
rect 206880 111600 207120 111620
rect 207380 111600 207620 111620
rect 207880 111600 208120 111620
rect 208380 111600 208620 111620
rect 208880 111600 209120 111620
rect 209380 111600 209620 111620
rect 209880 111600 210120 111620
rect 210380 111600 210620 111620
rect 210880 111600 211120 111620
rect 211380 111600 211620 111620
rect 211880 111600 212120 111620
rect 212380 111600 212620 111620
rect 212880 111600 213120 111620
rect 213380 111600 213620 111620
rect 213880 111600 214120 111620
rect 214380 111600 214620 111620
rect 214880 111600 215120 111620
rect 215380 111600 215620 111620
rect 215880 111600 216120 111620
rect 216380 111600 216620 111620
rect 216880 111600 217120 111620
rect 217380 111600 217620 111620
rect 217880 111600 218120 111620
rect 218380 111600 218620 111620
rect 218880 111600 219120 111620
rect 219380 111600 219620 111620
rect 219880 111600 220120 111620
rect 220380 111600 220620 111620
rect 220880 111600 221120 111620
rect 221380 111600 221620 111620
rect 221880 111600 222120 111620
rect 222380 111600 222620 111620
rect 222880 111600 223120 111620
rect 223380 111600 223620 111620
rect 223880 111600 224120 111620
rect 224380 111600 224620 111620
rect 224880 111600 225120 111620
rect 225380 111600 225620 111620
rect 225880 111600 226120 111620
rect 226380 111600 226620 111620
rect 226880 111600 227120 111620
rect 227380 111600 227620 111620
rect 227880 111600 228120 111620
rect 228380 111600 228620 111620
rect 228880 111600 229120 111620
rect 229380 111600 229620 111620
rect 229880 111600 230120 111620
rect 230380 111600 230620 111620
rect 230880 111600 231120 111620
rect 231380 111600 231620 111620
rect 231880 111600 232000 111620
rect 178000 111400 232000 111600
rect 178000 111380 178120 111400
rect 178380 111380 178620 111400
rect 178880 111380 179120 111400
rect 179380 111380 179620 111400
rect 179880 111380 180120 111400
rect 180380 111380 180620 111400
rect 180880 111380 181120 111400
rect 181380 111380 181620 111400
rect 181880 111380 182120 111400
rect 182380 111380 182620 111400
rect 182880 111380 183120 111400
rect 183380 111380 183620 111400
rect 183880 111380 184120 111400
rect 184380 111380 184620 111400
rect 184880 111380 185120 111400
rect 185380 111380 185620 111400
rect 185880 111380 186120 111400
rect 186380 111380 186620 111400
rect 186880 111380 187120 111400
rect 187380 111380 187620 111400
rect 187880 111380 188120 111400
rect 188380 111380 188620 111400
rect 188880 111380 189120 111400
rect 189380 111380 189620 111400
rect 189880 111380 190120 111400
rect 190380 111380 190620 111400
rect 190880 111380 191120 111400
rect 191380 111380 191620 111400
rect 191880 111380 192120 111400
rect 192380 111380 192620 111400
rect 192880 111380 193120 111400
rect 193380 111380 193620 111400
rect 193880 111380 194120 111400
rect 194380 111380 194620 111400
rect 194880 111380 195120 111400
rect 195380 111380 195620 111400
rect 195880 111380 196120 111400
rect 196380 111380 196620 111400
rect 196880 111380 197120 111400
rect 197380 111380 197620 111400
rect 197880 111380 198120 111400
rect 198380 111380 198620 111400
rect 198880 111380 199120 111400
rect 199380 111380 199620 111400
rect 199880 111380 200120 111400
rect 200380 111380 200620 111400
rect 200880 111380 201120 111400
rect 201380 111380 201620 111400
rect 201880 111380 202120 111400
rect 202380 111380 202620 111400
rect 202880 111380 203120 111400
rect 203380 111380 203620 111400
rect 203880 111380 204120 111400
rect 204380 111380 204620 111400
rect 204880 111380 205120 111400
rect 205380 111380 205620 111400
rect 205880 111380 206120 111400
rect 206380 111380 206620 111400
rect 206880 111380 207120 111400
rect 207380 111380 207620 111400
rect 207880 111380 208120 111400
rect 208380 111380 208620 111400
rect 208880 111380 209120 111400
rect 209380 111380 209620 111400
rect 209880 111380 210120 111400
rect 210380 111380 210620 111400
rect 210880 111380 211120 111400
rect 211380 111380 211620 111400
rect 211880 111380 212120 111400
rect 212380 111380 212620 111400
rect 212880 111380 213120 111400
rect 213380 111380 213620 111400
rect 213880 111380 214120 111400
rect 214380 111380 214620 111400
rect 214880 111380 215120 111400
rect 215380 111380 215620 111400
rect 215880 111380 216120 111400
rect 216380 111380 216620 111400
rect 216880 111380 217120 111400
rect 217380 111380 217620 111400
rect 217880 111380 218120 111400
rect 218380 111380 218620 111400
rect 218880 111380 219120 111400
rect 219380 111380 219620 111400
rect 219880 111380 220120 111400
rect 220380 111380 220620 111400
rect 220880 111380 221120 111400
rect 221380 111380 221620 111400
rect 221880 111380 222120 111400
rect 222380 111380 222620 111400
rect 222880 111380 223120 111400
rect 223380 111380 223620 111400
rect 223880 111380 224120 111400
rect 224380 111380 224620 111400
rect 224880 111380 225120 111400
rect 225380 111380 225620 111400
rect 225880 111380 226120 111400
rect 226380 111380 226620 111400
rect 226880 111380 227120 111400
rect 227380 111380 227620 111400
rect 227880 111380 228120 111400
rect 228380 111380 228620 111400
rect 228880 111380 229120 111400
rect 229380 111380 229620 111400
rect 229880 111380 230120 111400
rect 230380 111380 230620 111400
rect 230880 111380 231120 111400
rect 231380 111380 231620 111400
rect 231880 111380 232000 111400
rect 178000 111120 178100 111380
rect 178400 111120 178600 111380
rect 178900 111120 179100 111380
rect 179400 111120 179600 111380
rect 179900 111120 180100 111380
rect 180400 111120 180600 111380
rect 180900 111120 181100 111380
rect 181400 111120 181600 111380
rect 181900 111120 182100 111380
rect 182400 111120 182600 111380
rect 182900 111120 183100 111380
rect 183400 111120 183600 111380
rect 183900 111120 184100 111380
rect 184400 111120 184600 111380
rect 184900 111120 185100 111380
rect 185400 111120 185600 111380
rect 185900 111120 186100 111380
rect 186400 111120 186600 111380
rect 186900 111120 187100 111380
rect 187400 111120 187600 111380
rect 187900 111120 188100 111380
rect 188400 111120 188600 111380
rect 188900 111120 189100 111380
rect 189400 111120 189600 111380
rect 189900 111120 190100 111380
rect 190400 111120 190600 111380
rect 190900 111120 191100 111380
rect 191400 111120 191600 111380
rect 191900 111120 192100 111380
rect 192400 111120 192600 111380
rect 192900 111120 193100 111380
rect 193400 111120 193600 111380
rect 193900 111120 194100 111380
rect 194400 111120 194600 111380
rect 194900 111120 195100 111380
rect 195400 111120 195600 111380
rect 195900 111120 196100 111380
rect 196400 111120 196600 111380
rect 196900 111120 197100 111380
rect 197400 111120 197600 111380
rect 197900 111120 198100 111380
rect 198400 111120 198600 111380
rect 198900 111120 199100 111380
rect 199400 111120 199600 111380
rect 199900 111120 200100 111380
rect 200400 111120 200600 111380
rect 200900 111120 201100 111380
rect 201400 111120 201600 111380
rect 201900 111120 202100 111380
rect 202400 111120 202600 111380
rect 202900 111120 203100 111380
rect 203400 111120 203600 111380
rect 203900 111120 204100 111380
rect 204400 111120 204600 111380
rect 204900 111120 205100 111380
rect 205400 111120 205600 111380
rect 205900 111120 206100 111380
rect 206400 111120 206600 111380
rect 206900 111120 207100 111380
rect 207400 111120 207600 111380
rect 207900 111120 208100 111380
rect 208400 111120 208600 111380
rect 208900 111120 209100 111380
rect 209400 111120 209600 111380
rect 209900 111120 210100 111380
rect 210400 111120 210600 111380
rect 210900 111120 211100 111380
rect 211400 111120 211600 111380
rect 211900 111120 212100 111380
rect 212400 111120 212600 111380
rect 212900 111120 213100 111380
rect 213400 111120 213600 111380
rect 213900 111120 214100 111380
rect 214400 111120 214600 111380
rect 214900 111120 215100 111380
rect 215400 111120 215600 111380
rect 215900 111120 216100 111380
rect 216400 111120 216600 111380
rect 216900 111120 217100 111380
rect 217400 111120 217600 111380
rect 217900 111120 218100 111380
rect 218400 111120 218600 111380
rect 218900 111120 219100 111380
rect 219400 111120 219600 111380
rect 219900 111120 220100 111380
rect 220400 111120 220600 111380
rect 220900 111120 221100 111380
rect 221400 111120 221600 111380
rect 221900 111120 222100 111380
rect 222400 111120 222600 111380
rect 222900 111120 223100 111380
rect 223400 111120 223600 111380
rect 223900 111120 224100 111380
rect 224400 111120 224600 111380
rect 224900 111120 225100 111380
rect 225400 111120 225600 111380
rect 225900 111120 226100 111380
rect 226400 111120 226600 111380
rect 226900 111120 227100 111380
rect 227400 111120 227600 111380
rect 227900 111120 228100 111380
rect 228400 111120 228600 111380
rect 228900 111120 229100 111380
rect 229400 111120 229600 111380
rect 229900 111120 230100 111380
rect 230400 111120 230600 111380
rect 230900 111120 231100 111380
rect 231400 111120 231600 111380
rect 231900 111120 232000 111380
rect 178000 111100 178120 111120
rect 178380 111100 178620 111120
rect 178880 111100 179120 111120
rect 179380 111100 179620 111120
rect 179880 111100 180120 111120
rect 180380 111100 180620 111120
rect 180880 111100 181120 111120
rect 181380 111100 181620 111120
rect 181880 111100 182120 111120
rect 182380 111100 182620 111120
rect 182880 111100 183120 111120
rect 183380 111100 183620 111120
rect 183880 111100 184120 111120
rect 184380 111100 184620 111120
rect 184880 111100 185120 111120
rect 185380 111100 185620 111120
rect 185880 111100 186120 111120
rect 186380 111100 186620 111120
rect 186880 111100 187120 111120
rect 187380 111100 187620 111120
rect 187880 111100 188120 111120
rect 188380 111100 188620 111120
rect 188880 111100 189120 111120
rect 189380 111100 189620 111120
rect 189880 111100 190120 111120
rect 190380 111100 190620 111120
rect 190880 111100 191120 111120
rect 191380 111100 191620 111120
rect 191880 111100 192120 111120
rect 192380 111100 192620 111120
rect 192880 111100 193120 111120
rect 193380 111100 193620 111120
rect 193880 111100 194120 111120
rect 194380 111100 194620 111120
rect 194880 111100 195120 111120
rect 195380 111100 195620 111120
rect 195880 111100 196120 111120
rect 196380 111100 196620 111120
rect 196880 111100 197120 111120
rect 197380 111100 197620 111120
rect 197880 111100 198120 111120
rect 198380 111100 198620 111120
rect 198880 111100 199120 111120
rect 199380 111100 199620 111120
rect 199880 111100 200120 111120
rect 200380 111100 200620 111120
rect 200880 111100 201120 111120
rect 201380 111100 201620 111120
rect 201880 111100 202120 111120
rect 202380 111100 202620 111120
rect 202880 111100 203120 111120
rect 203380 111100 203620 111120
rect 203880 111100 204120 111120
rect 204380 111100 204620 111120
rect 204880 111100 205120 111120
rect 205380 111100 205620 111120
rect 205880 111100 206120 111120
rect 206380 111100 206620 111120
rect 206880 111100 207120 111120
rect 207380 111100 207620 111120
rect 207880 111100 208120 111120
rect 208380 111100 208620 111120
rect 208880 111100 209120 111120
rect 209380 111100 209620 111120
rect 209880 111100 210120 111120
rect 210380 111100 210620 111120
rect 210880 111100 211120 111120
rect 211380 111100 211620 111120
rect 211880 111100 212120 111120
rect 212380 111100 212620 111120
rect 212880 111100 213120 111120
rect 213380 111100 213620 111120
rect 213880 111100 214120 111120
rect 214380 111100 214620 111120
rect 214880 111100 215120 111120
rect 215380 111100 215620 111120
rect 215880 111100 216120 111120
rect 216380 111100 216620 111120
rect 216880 111100 217120 111120
rect 217380 111100 217620 111120
rect 217880 111100 218120 111120
rect 218380 111100 218620 111120
rect 218880 111100 219120 111120
rect 219380 111100 219620 111120
rect 219880 111100 220120 111120
rect 220380 111100 220620 111120
rect 220880 111100 221120 111120
rect 221380 111100 221620 111120
rect 221880 111100 222120 111120
rect 222380 111100 222620 111120
rect 222880 111100 223120 111120
rect 223380 111100 223620 111120
rect 223880 111100 224120 111120
rect 224380 111100 224620 111120
rect 224880 111100 225120 111120
rect 225380 111100 225620 111120
rect 225880 111100 226120 111120
rect 226380 111100 226620 111120
rect 226880 111100 227120 111120
rect 227380 111100 227620 111120
rect 227880 111100 228120 111120
rect 228380 111100 228620 111120
rect 228880 111100 229120 111120
rect 229380 111100 229620 111120
rect 229880 111100 230120 111120
rect 230380 111100 230620 111120
rect 230880 111100 231120 111120
rect 231380 111100 231620 111120
rect 231880 111100 232000 111120
rect 178000 110900 232000 111100
rect 178000 110880 178120 110900
rect 178380 110880 178620 110900
rect 178880 110880 179120 110900
rect 179380 110880 179620 110900
rect 179880 110880 180120 110900
rect 180380 110880 180620 110900
rect 180880 110880 181120 110900
rect 181380 110880 181620 110900
rect 181880 110880 182120 110900
rect 182380 110880 182620 110900
rect 182880 110880 183120 110900
rect 183380 110880 183620 110900
rect 183880 110880 184120 110900
rect 184380 110880 184620 110900
rect 184880 110880 185120 110900
rect 185380 110880 185620 110900
rect 185880 110880 186120 110900
rect 186380 110880 186620 110900
rect 186880 110880 187120 110900
rect 187380 110880 187620 110900
rect 187880 110880 188120 110900
rect 188380 110880 188620 110900
rect 188880 110880 189120 110900
rect 189380 110880 189620 110900
rect 189880 110880 190120 110900
rect 190380 110880 190620 110900
rect 190880 110880 191120 110900
rect 191380 110880 191620 110900
rect 191880 110880 192120 110900
rect 192380 110880 192620 110900
rect 192880 110880 193120 110900
rect 193380 110880 193620 110900
rect 193880 110880 194120 110900
rect 194380 110880 194620 110900
rect 194880 110880 195120 110900
rect 195380 110880 195620 110900
rect 195880 110880 196120 110900
rect 196380 110880 196620 110900
rect 196880 110880 197120 110900
rect 197380 110880 197620 110900
rect 197880 110880 198120 110900
rect 198380 110880 198620 110900
rect 198880 110880 199120 110900
rect 199380 110880 199620 110900
rect 199880 110880 200120 110900
rect 200380 110880 200620 110900
rect 200880 110880 201120 110900
rect 201380 110880 201620 110900
rect 201880 110880 202120 110900
rect 202380 110880 202620 110900
rect 202880 110880 203120 110900
rect 203380 110880 203620 110900
rect 203880 110880 204120 110900
rect 204380 110880 204620 110900
rect 204880 110880 205120 110900
rect 205380 110880 205620 110900
rect 205880 110880 206120 110900
rect 206380 110880 206620 110900
rect 206880 110880 207120 110900
rect 207380 110880 207620 110900
rect 207880 110880 208120 110900
rect 208380 110880 208620 110900
rect 208880 110880 209120 110900
rect 209380 110880 209620 110900
rect 209880 110880 210120 110900
rect 210380 110880 210620 110900
rect 210880 110880 211120 110900
rect 211380 110880 211620 110900
rect 211880 110880 212120 110900
rect 212380 110880 212620 110900
rect 212880 110880 213120 110900
rect 213380 110880 213620 110900
rect 213880 110880 214120 110900
rect 214380 110880 214620 110900
rect 214880 110880 215120 110900
rect 215380 110880 215620 110900
rect 215880 110880 216120 110900
rect 216380 110880 216620 110900
rect 216880 110880 217120 110900
rect 217380 110880 217620 110900
rect 217880 110880 218120 110900
rect 218380 110880 218620 110900
rect 218880 110880 219120 110900
rect 219380 110880 219620 110900
rect 219880 110880 220120 110900
rect 220380 110880 220620 110900
rect 220880 110880 221120 110900
rect 221380 110880 221620 110900
rect 221880 110880 222120 110900
rect 222380 110880 222620 110900
rect 222880 110880 223120 110900
rect 223380 110880 223620 110900
rect 223880 110880 224120 110900
rect 224380 110880 224620 110900
rect 224880 110880 225120 110900
rect 225380 110880 225620 110900
rect 225880 110880 226120 110900
rect 226380 110880 226620 110900
rect 226880 110880 227120 110900
rect 227380 110880 227620 110900
rect 227880 110880 228120 110900
rect 228380 110880 228620 110900
rect 228880 110880 229120 110900
rect 229380 110880 229620 110900
rect 229880 110880 230120 110900
rect 230380 110880 230620 110900
rect 230880 110880 231120 110900
rect 231380 110880 231620 110900
rect 231880 110880 232000 110900
rect 178000 110620 178100 110880
rect 178400 110620 178600 110880
rect 178900 110620 179100 110880
rect 179400 110620 179600 110880
rect 179900 110620 180100 110880
rect 180400 110620 180600 110880
rect 180900 110620 181100 110880
rect 181400 110620 181600 110880
rect 181900 110620 182100 110880
rect 182400 110620 182600 110880
rect 182900 110620 183100 110880
rect 183400 110620 183600 110880
rect 183900 110620 184100 110880
rect 184400 110620 184600 110880
rect 184900 110620 185100 110880
rect 185400 110620 185600 110880
rect 185900 110620 186100 110880
rect 186400 110620 186600 110880
rect 186900 110620 187100 110880
rect 187400 110620 187600 110880
rect 187900 110620 188100 110880
rect 188400 110620 188600 110880
rect 188900 110620 189100 110880
rect 189400 110620 189600 110880
rect 189900 110620 190100 110880
rect 190400 110620 190600 110880
rect 190900 110620 191100 110880
rect 191400 110620 191600 110880
rect 191900 110620 192100 110880
rect 192400 110620 192600 110880
rect 192900 110620 193100 110880
rect 193400 110620 193600 110880
rect 193900 110620 194100 110880
rect 194400 110620 194600 110880
rect 194900 110620 195100 110880
rect 195400 110620 195600 110880
rect 195900 110620 196100 110880
rect 196400 110620 196600 110880
rect 196900 110620 197100 110880
rect 197400 110620 197600 110880
rect 197900 110620 198100 110880
rect 198400 110620 198600 110880
rect 198900 110620 199100 110880
rect 199400 110620 199600 110880
rect 199900 110620 200100 110880
rect 200400 110620 200600 110880
rect 200900 110620 201100 110880
rect 201400 110620 201600 110880
rect 201900 110620 202100 110880
rect 202400 110620 202600 110880
rect 202900 110620 203100 110880
rect 203400 110620 203600 110880
rect 203900 110620 204100 110880
rect 204400 110620 204600 110880
rect 204900 110620 205100 110880
rect 205400 110620 205600 110880
rect 205900 110620 206100 110880
rect 206400 110620 206600 110880
rect 206900 110620 207100 110880
rect 207400 110620 207600 110880
rect 207900 110620 208100 110880
rect 208400 110620 208600 110880
rect 208900 110620 209100 110880
rect 209400 110620 209600 110880
rect 209900 110620 210100 110880
rect 210400 110620 210600 110880
rect 210900 110620 211100 110880
rect 211400 110620 211600 110880
rect 211900 110620 212100 110880
rect 212400 110620 212600 110880
rect 212900 110620 213100 110880
rect 213400 110620 213600 110880
rect 213900 110620 214100 110880
rect 214400 110620 214600 110880
rect 214900 110620 215100 110880
rect 215400 110620 215600 110880
rect 215900 110620 216100 110880
rect 216400 110620 216600 110880
rect 216900 110620 217100 110880
rect 217400 110620 217600 110880
rect 217900 110620 218100 110880
rect 218400 110620 218600 110880
rect 218900 110620 219100 110880
rect 219400 110620 219600 110880
rect 219900 110620 220100 110880
rect 220400 110620 220600 110880
rect 220900 110620 221100 110880
rect 221400 110620 221600 110880
rect 221900 110620 222100 110880
rect 222400 110620 222600 110880
rect 222900 110620 223100 110880
rect 223400 110620 223600 110880
rect 223900 110620 224100 110880
rect 224400 110620 224600 110880
rect 224900 110620 225100 110880
rect 225400 110620 225600 110880
rect 225900 110620 226100 110880
rect 226400 110620 226600 110880
rect 226900 110620 227100 110880
rect 227400 110620 227600 110880
rect 227900 110620 228100 110880
rect 228400 110620 228600 110880
rect 228900 110620 229100 110880
rect 229400 110620 229600 110880
rect 229900 110620 230100 110880
rect 230400 110620 230600 110880
rect 230900 110620 231100 110880
rect 231400 110620 231600 110880
rect 231900 110620 232000 110880
rect 178000 110600 178120 110620
rect 178380 110600 178620 110620
rect 178880 110600 179120 110620
rect 179380 110600 179620 110620
rect 179880 110600 180120 110620
rect 180380 110600 180620 110620
rect 180880 110600 181120 110620
rect 181380 110600 181620 110620
rect 181880 110600 182120 110620
rect 182380 110600 182620 110620
rect 182880 110600 183120 110620
rect 183380 110600 183620 110620
rect 183880 110600 184120 110620
rect 184380 110600 184620 110620
rect 184880 110600 185120 110620
rect 185380 110600 185620 110620
rect 185880 110600 186120 110620
rect 186380 110600 186620 110620
rect 186880 110600 187120 110620
rect 187380 110600 187620 110620
rect 187880 110600 188120 110620
rect 188380 110600 188620 110620
rect 188880 110600 189120 110620
rect 189380 110600 189620 110620
rect 189880 110600 190120 110620
rect 190380 110600 190620 110620
rect 190880 110600 191120 110620
rect 191380 110600 191620 110620
rect 191880 110600 192120 110620
rect 192380 110600 192620 110620
rect 192880 110600 193120 110620
rect 193380 110600 193620 110620
rect 193880 110600 194120 110620
rect 194380 110600 194620 110620
rect 194880 110600 195120 110620
rect 195380 110600 195620 110620
rect 195880 110600 196120 110620
rect 196380 110600 196620 110620
rect 196880 110600 197120 110620
rect 197380 110600 197620 110620
rect 197880 110600 198120 110620
rect 198380 110600 198620 110620
rect 198880 110600 199120 110620
rect 199380 110600 199620 110620
rect 199880 110600 200120 110620
rect 200380 110600 200620 110620
rect 200880 110600 201120 110620
rect 201380 110600 201620 110620
rect 201880 110600 202120 110620
rect 202380 110600 202620 110620
rect 202880 110600 203120 110620
rect 203380 110600 203620 110620
rect 203880 110600 204120 110620
rect 204380 110600 204620 110620
rect 204880 110600 205120 110620
rect 205380 110600 205620 110620
rect 205880 110600 206120 110620
rect 206380 110600 206620 110620
rect 206880 110600 207120 110620
rect 207380 110600 207620 110620
rect 207880 110600 208120 110620
rect 208380 110600 208620 110620
rect 208880 110600 209120 110620
rect 209380 110600 209620 110620
rect 209880 110600 210120 110620
rect 210380 110600 210620 110620
rect 210880 110600 211120 110620
rect 211380 110600 211620 110620
rect 211880 110600 212120 110620
rect 212380 110600 212620 110620
rect 212880 110600 213120 110620
rect 213380 110600 213620 110620
rect 213880 110600 214120 110620
rect 214380 110600 214620 110620
rect 214880 110600 215120 110620
rect 215380 110600 215620 110620
rect 215880 110600 216120 110620
rect 216380 110600 216620 110620
rect 216880 110600 217120 110620
rect 217380 110600 217620 110620
rect 217880 110600 218120 110620
rect 218380 110600 218620 110620
rect 218880 110600 219120 110620
rect 219380 110600 219620 110620
rect 219880 110600 220120 110620
rect 220380 110600 220620 110620
rect 220880 110600 221120 110620
rect 221380 110600 221620 110620
rect 221880 110600 222120 110620
rect 222380 110600 222620 110620
rect 222880 110600 223120 110620
rect 223380 110600 223620 110620
rect 223880 110600 224120 110620
rect 224380 110600 224620 110620
rect 224880 110600 225120 110620
rect 225380 110600 225620 110620
rect 225880 110600 226120 110620
rect 226380 110600 226620 110620
rect 226880 110600 227120 110620
rect 227380 110600 227620 110620
rect 227880 110600 228120 110620
rect 228380 110600 228620 110620
rect 228880 110600 229120 110620
rect 229380 110600 229620 110620
rect 229880 110600 230120 110620
rect 230380 110600 230620 110620
rect 230880 110600 231120 110620
rect 231380 110600 231620 110620
rect 231880 110600 232000 110620
rect 178000 110400 232000 110600
rect 178000 110380 178120 110400
rect 178380 110380 178620 110400
rect 178880 110380 179120 110400
rect 179380 110380 179620 110400
rect 179880 110380 180120 110400
rect 180380 110380 180620 110400
rect 180880 110380 181120 110400
rect 181380 110380 181620 110400
rect 181880 110380 182120 110400
rect 182380 110380 182620 110400
rect 182880 110380 183120 110400
rect 183380 110380 183620 110400
rect 183880 110380 184120 110400
rect 184380 110380 184620 110400
rect 184880 110380 185120 110400
rect 185380 110380 185620 110400
rect 185880 110380 186120 110400
rect 186380 110380 186620 110400
rect 186880 110380 187120 110400
rect 187380 110380 187620 110400
rect 187880 110380 188120 110400
rect 188380 110380 188620 110400
rect 188880 110380 189120 110400
rect 189380 110380 189620 110400
rect 189880 110380 190120 110400
rect 190380 110380 190620 110400
rect 190880 110380 191120 110400
rect 191380 110380 191620 110400
rect 191880 110380 192120 110400
rect 192380 110380 192620 110400
rect 192880 110380 193120 110400
rect 193380 110380 193620 110400
rect 193880 110380 194120 110400
rect 194380 110380 194620 110400
rect 194880 110380 195120 110400
rect 195380 110380 195620 110400
rect 195880 110380 196120 110400
rect 196380 110380 196620 110400
rect 196880 110380 197120 110400
rect 197380 110380 197620 110400
rect 197880 110380 198120 110400
rect 198380 110380 198620 110400
rect 198880 110380 199120 110400
rect 199380 110380 199620 110400
rect 199880 110380 200120 110400
rect 200380 110380 200620 110400
rect 200880 110380 201120 110400
rect 201380 110380 201620 110400
rect 201880 110380 202120 110400
rect 202380 110380 202620 110400
rect 202880 110380 203120 110400
rect 203380 110380 203620 110400
rect 203880 110380 204120 110400
rect 204380 110380 204620 110400
rect 204880 110380 205120 110400
rect 205380 110380 205620 110400
rect 205880 110380 206120 110400
rect 206380 110380 206620 110400
rect 206880 110380 207120 110400
rect 207380 110380 207620 110400
rect 207880 110380 208120 110400
rect 208380 110380 208620 110400
rect 208880 110380 209120 110400
rect 209380 110380 209620 110400
rect 209880 110380 210120 110400
rect 210380 110380 210620 110400
rect 210880 110380 211120 110400
rect 211380 110380 211620 110400
rect 211880 110380 212120 110400
rect 212380 110380 212620 110400
rect 212880 110380 213120 110400
rect 213380 110380 213620 110400
rect 213880 110380 214120 110400
rect 214380 110380 214620 110400
rect 214880 110380 215120 110400
rect 215380 110380 215620 110400
rect 215880 110380 216120 110400
rect 216380 110380 216620 110400
rect 216880 110380 217120 110400
rect 217380 110380 217620 110400
rect 217880 110380 218120 110400
rect 218380 110380 218620 110400
rect 218880 110380 219120 110400
rect 219380 110380 219620 110400
rect 219880 110380 220120 110400
rect 220380 110380 220620 110400
rect 220880 110380 221120 110400
rect 221380 110380 221620 110400
rect 221880 110380 222120 110400
rect 222380 110380 222620 110400
rect 222880 110380 223120 110400
rect 223380 110380 223620 110400
rect 223880 110380 224120 110400
rect 224380 110380 224620 110400
rect 224880 110380 225120 110400
rect 225380 110380 225620 110400
rect 225880 110380 226120 110400
rect 226380 110380 226620 110400
rect 226880 110380 227120 110400
rect 227380 110380 227620 110400
rect 227880 110380 228120 110400
rect 228380 110380 228620 110400
rect 228880 110380 229120 110400
rect 229380 110380 229620 110400
rect 229880 110380 230120 110400
rect 230380 110380 230620 110400
rect 230880 110380 231120 110400
rect 231380 110380 231620 110400
rect 231880 110380 232000 110400
rect 178000 110120 178100 110380
rect 178400 110120 178600 110380
rect 178900 110120 179100 110380
rect 179400 110120 179600 110380
rect 179900 110120 180100 110380
rect 180400 110120 180600 110380
rect 180900 110120 181100 110380
rect 181400 110120 181600 110380
rect 181900 110120 182100 110380
rect 182400 110120 182600 110380
rect 182900 110120 183100 110380
rect 183400 110120 183600 110380
rect 183900 110120 184100 110380
rect 184400 110120 184600 110380
rect 184900 110120 185100 110380
rect 185400 110120 185600 110380
rect 185900 110120 186100 110380
rect 186400 110120 186600 110380
rect 186900 110120 187100 110380
rect 187400 110120 187600 110380
rect 187900 110120 188100 110380
rect 188400 110120 188600 110380
rect 188900 110120 189100 110380
rect 189400 110120 189600 110380
rect 189900 110120 190100 110380
rect 190400 110120 190600 110380
rect 190900 110120 191100 110380
rect 191400 110120 191600 110380
rect 191900 110120 192100 110380
rect 192400 110120 192600 110380
rect 192900 110120 193100 110380
rect 193400 110120 193600 110380
rect 193900 110120 194100 110380
rect 194400 110120 194600 110380
rect 194900 110120 195100 110380
rect 195400 110120 195600 110380
rect 195900 110120 196100 110380
rect 196400 110120 196600 110380
rect 196900 110120 197100 110380
rect 197400 110120 197600 110380
rect 197900 110120 198100 110380
rect 198400 110120 198600 110380
rect 198900 110120 199100 110380
rect 199400 110120 199600 110380
rect 199900 110120 200100 110380
rect 200400 110120 200600 110380
rect 200900 110120 201100 110380
rect 201400 110120 201600 110380
rect 201900 110120 202100 110380
rect 202400 110120 202600 110380
rect 202900 110120 203100 110380
rect 203400 110120 203600 110380
rect 203900 110120 204100 110380
rect 204400 110120 204600 110380
rect 204900 110120 205100 110380
rect 205400 110120 205600 110380
rect 205900 110120 206100 110380
rect 206400 110120 206600 110380
rect 206900 110120 207100 110380
rect 207400 110120 207600 110380
rect 207900 110120 208100 110380
rect 208400 110120 208600 110380
rect 208900 110120 209100 110380
rect 209400 110120 209600 110380
rect 209900 110120 210100 110380
rect 210400 110120 210600 110380
rect 210900 110120 211100 110380
rect 211400 110120 211600 110380
rect 211900 110120 212100 110380
rect 212400 110120 212600 110380
rect 212900 110120 213100 110380
rect 213400 110120 213600 110380
rect 213900 110120 214100 110380
rect 214400 110120 214600 110380
rect 214900 110120 215100 110380
rect 215400 110120 215600 110380
rect 215900 110120 216100 110380
rect 216400 110120 216600 110380
rect 216900 110120 217100 110380
rect 217400 110120 217600 110380
rect 217900 110120 218100 110380
rect 218400 110120 218600 110380
rect 218900 110120 219100 110380
rect 219400 110120 219600 110380
rect 219900 110120 220100 110380
rect 220400 110120 220600 110380
rect 220900 110120 221100 110380
rect 221400 110120 221600 110380
rect 221900 110120 222100 110380
rect 222400 110120 222600 110380
rect 222900 110120 223100 110380
rect 223400 110120 223600 110380
rect 223900 110120 224100 110380
rect 224400 110120 224600 110380
rect 224900 110120 225100 110380
rect 225400 110120 225600 110380
rect 225900 110120 226100 110380
rect 226400 110120 226600 110380
rect 226900 110120 227100 110380
rect 227400 110120 227600 110380
rect 227900 110120 228100 110380
rect 228400 110120 228600 110380
rect 228900 110120 229100 110380
rect 229400 110120 229600 110380
rect 229900 110120 230100 110380
rect 230400 110120 230600 110380
rect 230900 110120 231100 110380
rect 231400 110120 231600 110380
rect 231900 110120 232000 110380
rect 178000 110100 178120 110120
rect 178380 110100 178620 110120
rect 178880 110100 179120 110120
rect 179380 110100 179620 110120
rect 179880 110100 180120 110120
rect 180380 110100 180620 110120
rect 180880 110100 181120 110120
rect 181380 110100 181620 110120
rect 181880 110100 182120 110120
rect 182380 110100 182620 110120
rect 182880 110100 183120 110120
rect 183380 110100 183620 110120
rect 183880 110100 184120 110120
rect 184380 110100 184620 110120
rect 184880 110100 185120 110120
rect 185380 110100 185620 110120
rect 185880 110100 186120 110120
rect 186380 110100 186620 110120
rect 186880 110100 187120 110120
rect 187380 110100 187620 110120
rect 187880 110100 188120 110120
rect 188380 110100 188620 110120
rect 188880 110100 189120 110120
rect 189380 110100 189620 110120
rect 189880 110100 190120 110120
rect 190380 110100 190620 110120
rect 190880 110100 191120 110120
rect 191380 110100 191620 110120
rect 191880 110100 192120 110120
rect 192380 110100 192620 110120
rect 192880 110100 193120 110120
rect 193380 110100 193620 110120
rect 193880 110100 194120 110120
rect 194380 110100 194620 110120
rect 194880 110100 195120 110120
rect 195380 110100 195620 110120
rect 195880 110100 196120 110120
rect 196380 110100 196620 110120
rect 196880 110100 197120 110120
rect 197380 110100 197620 110120
rect 197880 110100 198120 110120
rect 198380 110100 198620 110120
rect 198880 110100 199120 110120
rect 199380 110100 199620 110120
rect 199880 110100 200120 110120
rect 200380 110100 200620 110120
rect 200880 110100 201120 110120
rect 201380 110100 201620 110120
rect 201880 110100 202120 110120
rect 202380 110100 202620 110120
rect 202880 110100 203120 110120
rect 203380 110100 203620 110120
rect 203880 110100 204120 110120
rect 204380 110100 204620 110120
rect 204880 110100 205120 110120
rect 205380 110100 205620 110120
rect 205880 110100 206120 110120
rect 206380 110100 206620 110120
rect 206880 110100 207120 110120
rect 207380 110100 207620 110120
rect 207880 110100 208120 110120
rect 208380 110100 208620 110120
rect 208880 110100 209120 110120
rect 209380 110100 209620 110120
rect 209880 110100 210120 110120
rect 210380 110100 210620 110120
rect 210880 110100 211120 110120
rect 211380 110100 211620 110120
rect 211880 110100 212120 110120
rect 212380 110100 212620 110120
rect 212880 110100 213120 110120
rect 213380 110100 213620 110120
rect 213880 110100 214120 110120
rect 214380 110100 214620 110120
rect 214880 110100 215120 110120
rect 215380 110100 215620 110120
rect 215880 110100 216120 110120
rect 216380 110100 216620 110120
rect 216880 110100 217120 110120
rect 217380 110100 217620 110120
rect 217880 110100 218120 110120
rect 218380 110100 218620 110120
rect 218880 110100 219120 110120
rect 219380 110100 219620 110120
rect 219880 110100 220120 110120
rect 220380 110100 220620 110120
rect 220880 110100 221120 110120
rect 221380 110100 221620 110120
rect 221880 110100 222120 110120
rect 222380 110100 222620 110120
rect 222880 110100 223120 110120
rect 223380 110100 223620 110120
rect 223880 110100 224120 110120
rect 224380 110100 224620 110120
rect 224880 110100 225120 110120
rect 225380 110100 225620 110120
rect 225880 110100 226120 110120
rect 226380 110100 226620 110120
rect 226880 110100 227120 110120
rect 227380 110100 227620 110120
rect 227880 110100 228120 110120
rect 228380 110100 228620 110120
rect 228880 110100 229120 110120
rect 229380 110100 229620 110120
rect 229880 110100 230120 110120
rect 230380 110100 230620 110120
rect 230880 110100 231120 110120
rect 231380 110100 231620 110120
rect 231880 110100 232000 110120
rect 178000 109900 232000 110100
rect 178000 109880 178120 109900
rect 178380 109880 178620 109900
rect 178880 109880 179120 109900
rect 179380 109880 179620 109900
rect 179880 109880 180120 109900
rect 180380 109880 180620 109900
rect 180880 109880 181120 109900
rect 181380 109880 181620 109900
rect 181880 109880 182120 109900
rect 182380 109880 182620 109900
rect 182880 109880 183120 109900
rect 183380 109880 183620 109900
rect 183880 109880 184120 109900
rect 184380 109880 184620 109900
rect 184880 109880 185120 109900
rect 185380 109880 185620 109900
rect 185880 109880 186120 109900
rect 186380 109880 186620 109900
rect 186880 109880 187120 109900
rect 187380 109880 187620 109900
rect 187880 109880 188120 109900
rect 188380 109880 188620 109900
rect 188880 109880 189120 109900
rect 189380 109880 189620 109900
rect 189880 109880 190120 109900
rect 190380 109880 190620 109900
rect 190880 109880 191120 109900
rect 191380 109880 191620 109900
rect 191880 109880 192120 109900
rect 192380 109880 192620 109900
rect 192880 109880 193120 109900
rect 193380 109880 193620 109900
rect 193880 109880 194120 109900
rect 194380 109880 194620 109900
rect 194880 109880 195120 109900
rect 195380 109880 195620 109900
rect 195880 109880 196120 109900
rect 196380 109880 196620 109900
rect 196880 109880 197120 109900
rect 197380 109880 197620 109900
rect 197880 109880 198120 109900
rect 198380 109880 198620 109900
rect 198880 109880 199120 109900
rect 199380 109880 199620 109900
rect 199880 109880 200120 109900
rect 200380 109880 200620 109900
rect 200880 109880 201120 109900
rect 201380 109880 201620 109900
rect 201880 109880 202120 109900
rect 202380 109880 202620 109900
rect 202880 109880 203120 109900
rect 203380 109880 203620 109900
rect 203880 109880 204120 109900
rect 204380 109880 204620 109900
rect 204880 109880 205120 109900
rect 205380 109880 205620 109900
rect 205880 109880 206120 109900
rect 206380 109880 206620 109900
rect 206880 109880 207120 109900
rect 207380 109880 207620 109900
rect 207880 109880 208120 109900
rect 208380 109880 208620 109900
rect 208880 109880 209120 109900
rect 209380 109880 209620 109900
rect 209880 109880 210120 109900
rect 210380 109880 210620 109900
rect 210880 109880 211120 109900
rect 211380 109880 211620 109900
rect 211880 109880 212120 109900
rect 212380 109880 212620 109900
rect 212880 109880 213120 109900
rect 213380 109880 213620 109900
rect 213880 109880 214120 109900
rect 214380 109880 214620 109900
rect 214880 109880 215120 109900
rect 215380 109880 215620 109900
rect 215880 109880 216120 109900
rect 216380 109880 216620 109900
rect 216880 109880 217120 109900
rect 217380 109880 217620 109900
rect 217880 109880 218120 109900
rect 218380 109880 218620 109900
rect 218880 109880 219120 109900
rect 219380 109880 219620 109900
rect 219880 109880 220120 109900
rect 220380 109880 220620 109900
rect 220880 109880 221120 109900
rect 221380 109880 221620 109900
rect 221880 109880 222120 109900
rect 222380 109880 222620 109900
rect 222880 109880 223120 109900
rect 223380 109880 223620 109900
rect 223880 109880 224120 109900
rect 224380 109880 224620 109900
rect 224880 109880 225120 109900
rect 225380 109880 225620 109900
rect 225880 109880 226120 109900
rect 226380 109880 226620 109900
rect 226880 109880 227120 109900
rect 227380 109880 227620 109900
rect 227880 109880 228120 109900
rect 228380 109880 228620 109900
rect 228880 109880 229120 109900
rect 229380 109880 229620 109900
rect 229880 109880 230120 109900
rect 230380 109880 230620 109900
rect 230880 109880 231120 109900
rect 231380 109880 231620 109900
rect 231880 109880 232000 109900
rect 178000 109620 178100 109880
rect 178400 109620 178600 109880
rect 178900 109620 179100 109880
rect 179400 109620 179600 109880
rect 179900 109620 180100 109880
rect 180400 109620 180600 109880
rect 180900 109620 181100 109880
rect 181400 109620 181600 109880
rect 181900 109620 182100 109880
rect 182400 109620 182600 109880
rect 182900 109620 183100 109880
rect 183400 109620 183600 109880
rect 183900 109620 184100 109880
rect 184400 109620 184600 109880
rect 184900 109620 185100 109880
rect 185400 109620 185600 109880
rect 185900 109620 186100 109880
rect 186400 109620 186600 109880
rect 186900 109620 187100 109880
rect 187400 109620 187600 109880
rect 187900 109620 188100 109880
rect 188400 109620 188600 109880
rect 188900 109620 189100 109880
rect 189400 109620 189600 109880
rect 189900 109620 190100 109880
rect 190400 109620 190600 109880
rect 190900 109620 191100 109880
rect 191400 109620 191600 109880
rect 191900 109620 192100 109880
rect 192400 109620 192600 109880
rect 192900 109620 193100 109880
rect 193400 109620 193600 109880
rect 193900 109620 194100 109880
rect 194400 109620 194600 109880
rect 194900 109620 195100 109880
rect 195400 109620 195600 109880
rect 195900 109620 196100 109880
rect 196400 109620 196600 109880
rect 196900 109620 197100 109880
rect 197400 109620 197600 109880
rect 197900 109620 198100 109880
rect 198400 109620 198600 109880
rect 198900 109620 199100 109880
rect 199400 109620 199600 109880
rect 199900 109620 200100 109880
rect 200400 109620 200600 109880
rect 200900 109620 201100 109880
rect 201400 109620 201600 109880
rect 201900 109620 202100 109880
rect 202400 109620 202600 109880
rect 202900 109620 203100 109880
rect 203400 109620 203600 109880
rect 203900 109620 204100 109880
rect 204400 109620 204600 109880
rect 204900 109620 205100 109880
rect 205400 109620 205600 109880
rect 205900 109620 206100 109880
rect 206400 109620 206600 109880
rect 206900 109620 207100 109880
rect 207400 109620 207600 109880
rect 207900 109620 208100 109880
rect 208400 109620 208600 109880
rect 208900 109620 209100 109880
rect 209400 109620 209600 109880
rect 209900 109620 210100 109880
rect 210400 109620 210600 109880
rect 210900 109620 211100 109880
rect 211400 109620 211600 109880
rect 211900 109620 212100 109880
rect 212400 109620 212600 109880
rect 212900 109620 213100 109880
rect 213400 109620 213600 109880
rect 213900 109620 214100 109880
rect 214400 109620 214600 109880
rect 214900 109620 215100 109880
rect 215400 109620 215600 109880
rect 215900 109620 216100 109880
rect 216400 109620 216600 109880
rect 216900 109620 217100 109880
rect 217400 109620 217600 109880
rect 217900 109620 218100 109880
rect 218400 109620 218600 109880
rect 218900 109620 219100 109880
rect 219400 109620 219600 109880
rect 219900 109620 220100 109880
rect 220400 109620 220600 109880
rect 220900 109620 221100 109880
rect 221400 109620 221600 109880
rect 221900 109620 222100 109880
rect 222400 109620 222600 109880
rect 222900 109620 223100 109880
rect 223400 109620 223600 109880
rect 223900 109620 224100 109880
rect 224400 109620 224600 109880
rect 224900 109620 225100 109880
rect 225400 109620 225600 109880
rect 225900 109620 226100 109880
rect 226400 109620 226600 109880
rect 226900 109620 227100 109880
rect 227400 109620 227600 109880
rect 227900 109620 228100 109880
rect 228400 109620 228600 109880
rect 228900 109620 229100 109880
rect 229400 109620 229600 109880
rect 229900 109620 230100 109880
rect 230400 109620 230600 109880
rect 230900 109620 231100 109880
rect 231400 109620 231600 109880
rect 231900 109620 232000 109880
rect 178000 109600 178120 109620
rect 178380 109600 178620 109620
rect 178880 109600 179120 109620
rect 179380 109600 179620 109620
rect 179880 109600 180120 109620
rect 180380 109600 180620 109620
rect 180880 109600 181120 109620
rect 181380 109600 181620 109620
rect 181880 109600 182120 109620
rect 182380 109600 182620 109620
rect 182880 109600 183120 109620
rect 183380 109600 183620 109620
rect 183880 109600 184120 109620
rect 184380 109600 184620 109620
rect 184880 109600 185120 109620
rect 185380 109600 185620 109620
rect 185880 109600 186120 109620
rect 186380 109600 186620 109620
rect 186880 109600 187120 109620
rect 187380 109600 187620 109620
rect 187880 109600 188120 109620
rect 188380 109600 188620 109620
rect 188880 109600 189120 109620
rect 189380 109600 189620 109620
rect 189880 109600 190120 109620
rect 190380 109600 190620 109620
rect 190880 109600 191120 109620
rect 191380 109600 191620 109620
rect 191880 109600 192120 109620
rect 192380 109600 192620 109620
rect 192880 109600 193120 109620
rect 193380 109600 193620 109620
rect 193880 109600 194120 109620
rect 194380 109600 194620 109620
rect 194880 109600 195120 109620
rect 195380 109600 195620 109620
rect 195880 109600 196120 109620
rect 196380 109600 196620 109620
rect 196880 109600 197120 109620
rect 197380 109600 197620 109620
rect 197880 109600 198120 109620
rect 198380 109600 198620 109620
rect 198880 109600 199120 109620
rect 199380 109600 199620 109620
rect 199880 109600 200120 109620
rect 200380 109600 200620 109620
rect 200880 109600 201120 109620
rect 201380 109600 201620 109620
rect 201880 109600 202120 109620
rect 202380 109600 202620 109620
rect 202880 109600 203120 109620
rect 203380 109600 203620 109620
rect 203880 109600 204120 109620
rect 204380 109600 204620 109620
rect 204880 109600 205120 109620
rect 205380 109600 205620 109620
rect 205880 109600 206120 109620
rect 206380 109600 206620 109620
rect 206880 109600 207120 109620
rect 207380 109600 207620 109620
rect 207880 109600 208120 109620
rect 208380 109600 208620 109620
rect 208880 109600 209120 109620
rect 209380 109600 209620 109620
rect 209880 109600 210120 109620
rect 210380 109600 210620 109620
rect 210880 109600 211120 109620
rect 211380 109600 211620 109620
rect 211880 109600 212120 109620
rect 212380 109600 212620 109620
rect 212880 109600 213120 109620
rect 213380 109600 213620 109620
rect 213880 109600 214120 109620
rect 214380 109600 214620 109620
rect 214880 109600 215120 109620
rect 215380 109600 215620 109620
rect 215880 109600 216120 109620
rect 216380 109600 216620 109620
rect 216880 109600 217120 109620
rect 217380 109600 217620 109620
rect 217880 109600 218120 109620
rect 218380 109600 218620 109620
rect 218880 109600 219120 109620
rect 219380 109600 219620 109620
rect 219880 109600 220120 109620
rect 220380 109600 220620 109620
rect 220880 109600 221120 109620
rect 221380 109600 221620 109620
rect 221880 109600 222120 109620
rect 222380 109600 222620 109620
rect 222880 109600 223120 109620
rect 223380 109600 223620 109620
rect 223880 109600 224120 109620
rect 224380 109600 224620 109620
rect 224880 109600 225120 109620
rect 225380 109600 225620 109620
rect 225880 109600 226120 109620
rect 226380 109600 226620 109620
rect 226880 109600 227120 109620
rect 227380 109600 227620 109620
rect 227880 109600 228120 109620
rect 228380 109600 228620 109620
rect 228880 109600 229120 109620
rect 229380 109600 229620 109620
rect 229880 109600 230120 109620
rect 230380 109600 230620 109620
rect 230880 109600 231120 109620
rect 231380 109600 231620 109620
rect 231880 109600 232000 109620
rect 178000 109400 232000 109600
rect 178000 109380 178120 109400
rect 178380 109380 178620 109400
rect 178880 109380 179120 109400
rect 179380 109380 179620 109400
rect 179880 109380 180120 109400
rect 180380 109380 180620 109400
rect 180880 109380 181120 109400
rect 181380 109380 181620 109400
rect 181880 109380 182120 109400
rect 182380 109380 182620 109400
rect 182880 109380 183120 109400
rect 183380 109380 183620 109400
rect 183880 109380 184120 109400
rect 184380 109380 184620 109400
rect 184880 109380 185120 109400
rect 185380 109380 185620 109400
rect 185880 109380 186120 109400
rect 186380 109380 186620 109400
rect 186880 109380 187120 109400
rect 187380 109380 187620 109400
rect 187880 109380 188120 109400
rect 188380 109380 188620 109400
rect 188880 109380 189120 109400
rect 189380 109380 189620 109400
rect 189880 109380 190120 109400
rect 190380 109380 190620 109400
rect 190880 109380 191120 109400
rect 191380 109380 191620 109400
rect 191880 109380 192120 109400
rect 192380 109380 192620 109400
rect 192880 109380 193120 109400
rect 193380 109380 193620 109400
rect 193880 109380 194120 109400
rect 194380 109380 194620 109400
rect 194880 109380 195120 109400
rect 195380 109380 195620 109400
rect 195880 109380 196120 109400
rect 196380 109380 196620 109400
rect 196880 109380 197120 109400
rect 197380 109380 197620 109400
rect 197880 109380 198120 109400
rect 198380 109380 198620 109400
rect 198880 109380 199120 109400
rect 199380 109380 199620 109400
rect 199880 109380 200120 109400
rect 200380 109380 200620 109400
rect 200880 109380 201120 109400
rect 201380 109380 201620 109400
rect 201880 109380 202120 109400
rect 202380 109380 202620 109400
rect 202880 109380 203120 109400
rect 203380 109380 203620 109400
rect 203880 109380 204120 109400
rect 204380 109380 204620 109400
rect 204880 109380 205120 109400
rect 205380 109380 205620 109400
rect 205880 109380 206120 109400
rect 206380 109380 206620 109400
rect 206880 109380 207120 109400
rect 207380 109380 207620 109400
rect 207880 109380 208120 109400
rect 208380 109380 208620 109400
rect 208880 109380 209120 109400
rect 209380 109380 209620 109400
rect 209880 109380 210120 109400
rect 210380 109380 210620 109400
rect 210880 109380 211120 109400
rect 211380 109380 211620 109400
rect 211880 109380 212120 109400
rect 212380 109380 212620 109400
rect 212880 109380 213120 109400
rect 213380 109380 213620 109400
rect 213880 109380 214120 109400
rect 214380 109380 214620 109400
rect 214880 109380 215120 109400
rect 215380 109380 215620 109400
rect 215880 109380 216120 109400
rect 216380 109380 216620 109400
rect 216880 109380 217120 109400
rect 217380 109380 217620 109400
rect 217880 109380 218120 109400
rect 218380 109380 218620 109400
rect 218880 109380 219120 109400
rect 219380 109380 219620 109400
rect 219880 109380 220120 109400
rect 220380 109380 220620 109400
rect 220880 109380 221120 109400
rect 221380 109380 221620 109400
rect 221880 109380 222120 109400
rect 222380 109380 222620 109400
rect 222880 109380 223120 109400
rect 223380 109380 223620 109400
rect 223880 109380 224120 109400
rect 224380 109380 224620 109400
rect 224880 109380 225120 109400
rect 225380 109380 225620 109400
rect 225880 109380 226120 109400
rect 226380 109380 226620 109400
rect 226880 109380 227120 109400
rect 227380 109380 227620 109400
rect 227880 109380 228120 109400
rect 228380 109380 228620 109400
rect 228880 109380 229120 109400
rect 229380 109380 229620 109400
rect 229880 109380 230120 109400
rect 230380 109380 230620 109400
rect 230880 109380 231120 109400
rect 231380 109380 231620 109400
rect 231880 109380 232000 109400
rect 178000 109120 178100 109380
rect 178400 109120 178600 109380
rect 178900 109120 179100 109380
rect 179400 109120 179600 109380
rect 179900 109120 180100 109380
rect 180400 109120 180600 109380
rect 180900 109120 181100 109380
rect 181400 109120 181600 109380
rect 181900 109120 182100 109380
rect 182400 109120 182600 109380
rect 182900 109120 183100 109380
rect 183400 109120 183600 109380
rect 183900 109120 184100 109380
rect 184400 109120 184600 109380
rect 184900 109120 185100 109380
rect 185400 109120 185600 109380
rect 185900 109120 186100 109380
rect 186400 109120 186600 109380
rect 186900 109120 187100 109380
rect 187400 109120 187600 109380
rect 187900 109120 188100 109380
rect 188400 109120 188600 109380
rect 188900 109120 189100 109380
rect 189400 109120 189600 109380
rect 189900 109120 190100 109380
rect 190400 109120 190600 109380
rect 190900 109120 191100 109380
rect 191400 109120 191600 109380
rect 191900 109120 192100 109380
rect 192400 109120 192600 109380
rect 192900 109120 193100 109380
rect 193400 109120 193600 109380
rect 193900 109120 194100 109380
rect 194400 109120 194600 109380
rect 194900 109120 195100 109380
rect 195400 109120 195600 109380
rect 195900 109120 196100 109380
rect 196400 109120 196600 109380
rect 196900 109120 197100 109380
rect 197400 109120 197600 109380
rect 197900 109120 198100 109380
rect 198400 109120 198600 109380
rect 198900 109120 199100 109380
rect 199400 109120 199600 109380
rect 199900 109120 200100 109380
rect 200400 109120 200600 109380
rect 200900 109120 201100 109380
rect 201400 109120 201600 109380
rect 201900 109120 202100 109380
rect 202400 109120 202600 109380
rect 202900 109120 203100 109380
rect 203400 109120 203600 109380
rect 203900 109120 204100 109380
rect 204400 109120 204600 109380
rect 204900 109120 205100 109380
rect 205400 109120 205600 109380
rect 205900 109120 206100 109380
rect 206400 109120 206600 109380
rect 206900 109120 207100 109380
rect 207400 109120 207600 109380
rect 207900 109120 208100 109380
rect 208400 109120 208600 109380
rect 208900 109120 209100 109380
rect 209400 109120 209600 109380
rect 209900 109120 210100 109380
rect 210400 109120 210600 109380
rect 210900 109120 211100 109380
rect 211400 109120 211600 109380
rect 211900 109120 212100 109380
rect 212400 109120 212600 109380
rect 212900 109120 213100 109380
rect 213400 109120 213600 109380
rect 213900 109120 214100 109380
rect 214400 109120 214600 109380
rect 214900 109120 215100 109380
rect 215400 109120 215600 109380
rect 215900 109120 216100 109380
rect 216400 109120 216600 109380
rect 216900 109120 217100 109380
rect 217400 109120 217600 109380
rect 217900 109120 218100 109380
rect 218400 109120 218600 109380
rect 218900 109120 219100 109380
rect 219400 109120 219600 109380
rect 219900 109120 220100 109380
rect 220400 109120 220600 109380
rect 220900 109120 221100 109380
rect 221400 109120 221600 109380
rect 221900 109120 222100 109380
rect 222400 109120 222600 109380
rect 222900 109120 223100 109380
rect 223400 109120 223600 109380
rect 223900 109120 224100 109380
rect 224400 109120 224600 109380
rect 224900 109120 225100 109380
rect 225400 109120 225600 109380
rect 225900 109120 226100 109380
rect 226400 109120 226600 109380
rect 226900 109120 227100 109380
rect 227400 109120 227600 109380
rect 227900 109120 228100 109380
rect 228400 109120 228600 109380
rect 228900 109120 229100 109380
rect 229400 109120 229600 109380
rect 229900 109120 230100 109380
rect 230400 109120 230600 109380
rect 230900 109120 231100 109380
rect 231400 109120 231600 109380
rect 231900 109120 232000 109380
rect 178000 109100 178120 109120
rect 178380 109100 178620 109120
rect 178880 109100 179120 109120
rect 179380 109100 179620 109120
rect 179880 109100 180120 109120
rect 180380 109100 180620 109120
rect 180880 109100 181120 109120
rect 181380 109100 181620 109120
rect 181880 109100 182120 109120
rect 182380 109100 182620 109120
rect 182880 109100 183120 109120
rect 183380 109100 183620 109120
rect 183880 109100 184120 109120
rect 184380 109100 184620 109120
rect 184880 109100 185120 109120
rect 185380 109100 185620 109120
rect 185880 109100 186120 109120
rect 186380 109100 186620 109120
rect 186880 109100 187120 109120
rect 187380 109100 187620 109120
rect 187880 109100 188120 109120
rect 188380 109100 188620 109120
rect 188880 109100 189120 109120
rect 189380 109100 189620 109120
rect 189880 109100 190120 109120
rect 190380 109100 190620 109120
rect 190880 109100 191120 109120
rect 191380 109100 191620 109120
rect 191880 109100 192120 109120
rect 192380 109100 192620 109120
rect 192880 109100 193120 109120
rect 193380 109100 193620 109120
rect 193880 109100 194120 109120
rect 194380 109100 194620 109120
rect 194880 109100 195120 109120
rect 195380 109100 195620 109120
rect 195880 109100 196120 109120
rect 196380 109100 196620 109120
rect 196880 109100 197120 109120
rect 197380 109100 197620 109120
rect 197880 109100 198120 109120
rect 198380 109100 198620 109120
rect 198880 109100 199120 109120
rect 199380 109100 199620 109120
rect 199880 109100 200120 109120
rect 200380 109100 200620 109120
rect 200880 109100 201120 109120
rect 201380 109100 201620 109120
rect 201880 109100 202120 109120
rect 202380 109100 202620 109120
rect 202880 109100 203120 109120
rect 203380 109100 203620 109120
rect 203880 109100 204120 109120
rect 204380 109100 204620 109120
rect 204880 109100 205120 109120
rect 205380 109100 205620 109120
rect 205880 109100 206120 109120
rect 206380 109100 206620 109120
rect 206880 109100 207120 109120
rect 207380 109100 207620 109120
rect 207880 109100 208120 109120
rect 208380 109100 208620 109120
rect 208880 109100 209120 109120
rect 209380 109100 209620 109120
rect 209880 109100 210120 109120
rect 210380 109100 210620 109120
rect 210880 109100 211120 109120
rect 211380 109100 211620 109120
rect 211880 109100 212120 109120
rect 212380 109100 212620 109120
rect 212880 109100 213120 109120
rect 213380 109100 213620 109120
rect 213880 109100 214120 109120
rect 214380 109100 214620 109120
rect 214880 109100 215120 109120
rect 215380 109100 215620 109120
rect 215880 109100 216120 109120
rect 216380 109100 216620 109120
rect 216880 109100 217120 109120
rect 217380 109100 217620 109120
rect 217880 109100 218120 109120
rect 218380 109100 218620 109120
rect 218880 109100 219120 109120
rect 219380 109100 219620 109120
rect 219880 109100 220120 109120
rect 220380 109100 220620 109120
rect 220880 109100 221120 109120
rect 221380 109100 221620 109120
rect 221880 109100 222120 109120
rect 222380 109100 222620 109120
rect 222880 109100 223120 109120
rect 223380 109100 223620 109120
rect 223880 109100 224120 109120
rect 224380 109100 224620 109120
rect 224880 109100 225120 109120
rect 225380 109100 225620 109120
rect 225880 109100 226120 109120
rect 226380 109100 226620 109120
rect 226880 109100 227120 109120
rect 227380 109100 227620 109120
rect 227880 109100 228120 109120
rect 228380 109100 228620 109120
rect 228880 109100 229120 109120
rect 229380 109100 229620 109120
rect 229880 109100 230120 109120
rect 230380 109100 230620 109120
rect 230880 109100 231120 109120
rect 231380 109100 231620 109120
rect 231880 109100 232000 109120
rect 178000 108900 232000 109100
rect 178000 108880 178120 108900
rect 178380 108880 178620 108900
rect 178880 108880 179120 108900
rect 179380 108880 179620 108900
rect 179880 108880 180120 108900
rect 180380 108880 180620 108900
rect 180880 108880 181120 108900
rect 181380 108880 181620 108900
rect 181880 108880 182120 108900
rect 182380 108880 182620 108900
rect 182880 108880 183120 108900
rect 183380 108880 183620 108900
rect 183880 108880 184120 108900
rect 184380 108880 184620 108900
rect 184880 108880 185120 108900
rect 185380 108880 185620 108900
rect 185880 108880 186120 108900
rect 186380 108880 186620 108900
rect 186880 108880 187120 108900
rect 187380 108880 187620 108900
rect 187880 108880 188120 108900
rect 188380 108880 188620 108900
rect 188880 108880 189120 108900
rect 189380 108880 189620 108900
rect 189880 108880 190120 108900
rect 190380 108880 190620 108900
rect 190880 108880 191120 108900
rect 191380 108880 191620 108900
rect 191880 108880 192120 108900
rect 192380 108880 192620 108900
rect 192880 108880 193120 108900
rect 193380 108880 193620 108900
rect 193880 108880 194120 108900
rect 194380 108880 194620 108900
rect 194880 108880 195120 108900
rect 195380 108880 195620 108900
rect 195880 108880 196120 108900
rect 196380 108880 196620 108900
rect 196880 108880 197120 108900
rect 197380 108880 197620 108900
rect 197880 108880 198120 108900
rect 198380 108880 198620 108900
rect 198880 108880 199120 108900
rect 199380 108880 199620 108900
rect 199880 108880 200120 108900
rect 200380 108880 200620 108900
rect 200880 108880 201120 108900
rect 201380 108880 201620 108900
rect 201880 108880 202120 108900
rect 202380 108880 202620 108900
rect 202880 108880 203120 108900
rect 203380 108880 203620 108900
rect 203880 108880 204120 108900
rect 204380 108880 204620 108900
rect 204880 108880 205120 108900
rect 205380 108880 205620 108900
rect 205880 108880 206120 108900
rect 206380 108880 206620 108900
rect 206880 108880 207120 108900
rect 207380 108880 207620 108900
rect 207880 108880 208120 108900
rect 208380 108880 208620 108900
rect 208880 108880 209120 108900
rect 209380 108880 209620 108900
rect 209880 108880 210120 108900
rect 210380 108880 210620 108900
rect 210880 108880 211120 108900
rect 211380 108880 211620 108900
rect 211880 108880 212120 108900
rect 212380 108880 212620 108900
rect 212880 108880 213120 108900
rect 213380 108880 213620 108900
rect 213880 108880 214120 108900
rect 214380 108880 214620 108900
rect 214880 108880 215120 108900
rect 215380 108880 215620 108900
rect 215880 108880 216120 108900
rect 216380 108880 216620 108900
rect 216880 108880 217120 108900
rect 217380 108880 217620 108900
rect 217880 108880 218120 108900
rect 218380 108880 218620 108900
rect 218880 108880 219120 108900
rect 219380 108880 219620 108900
rect 219880 108880 220120 108900
rect 220380 108880 220620 108900
rect 220880 108880 221120 108900
rect 221380 108880 221620 108900
rect 221880 108880 222120 108900
rect 222380 108880 222620 108900
rect 222880 108880 223120 108900
rect 223380 108880 223620 108900
rect 223880 108880 224120 108900
rect 224380 108880 224620 108900
rect 224880 108880 225120 108900
rect 225380 108880 225620 108900
rect 225880 108880 226120 108900
rect 226380 108880 226620 108900
rect 226880 108880 227120 108900
rect 227380 108880 227620 108900
rect 227880 108880 228120 108900
rect 228380 108880 228620 108900
rect 228880 108880 229120 108900
rect 229380 108880 229620 108900
rect 229880 108880 230120 108900
rect 230380 108880 230620 108900
rect 230880 108880 231120 108900
rect 231380 108880 231620 108900
rect 231880 108880 232000 108900
rect 178000 108620 178100 108880
rect 178400 108620 178600 108880
rect 178900 108620 179100 108880
rect 179400 108620 179600 108880
rect 179900 108620 180100 108880
rect 180400 108620 180600 108880
rect 180900 108620 181100 108880
rect 181400 108620 181600 108880
rect 181900 108620 182100 108880
rect 182400 108620 182600 108880
rect 182900 108620 183100 108880
rect 183400 108620 183600 108880
rect 183900 108620 184100 108880
rect 184400 108620 184600 108880
rect 184900 108620 185100 108880
rect 185400 108620 185600 108880
rect 185900 108620 186100 108880
rect 186400 108620 186600 108880
rect 186900 108620 187100 108880
rect 187400 108620 187600 108880
rect 187900 108620 188100 108880
rect 188400 108620 188600 108880
rect 188900 108620 189100 108880
rect 189400 108620 189600 108880
rect 189900 108620 190100 108880
rect 190400 108620 190600 108880
rect 190900 108620 191100 108880
rect 191400 108620 191600 108880
rect 191900 108620 192100 108880
rect 192400 108620 192600 108880
rect 192900 108620 193100 108880
rect 193400 108620 193600 108880
rect 193900 108620 194100 108880
rect 194400 108620 194600 108880
rect 194900 108620 195100 108880
rect 195400 108620 195600 108880
rect 195900 108620 196100 108880
rect 196400 108620 196600 108880
rect 196900 108620 197100 108880
rect 197400 108620 197600 108880
rect 197900 108620 198100 108880
rect 198400 108620 198600 108880
rect 198900 108620 199100 108880
rect 199400 108620 199600 108880
rect 199900 108620 200100 108880
rect 200400 108620 200600 108880
rect 200900 108620 201100 108880
rect 201400 108620 201600 108880
rect 201900 108620 202100 108880
rect 202400 108620 202600 108880
rect 202900 108620 203100 108880
rect 203400 108620 203600 108880
rect 203900 108620 204100 108880
rect 204400 108620 204600 108880
rect 204900 108620 205100 108880
rect 205400 108620 205600 108880
rect 205900 108620 206100 108880
rect 206400 108620 206600 108880
rect 206900 108620 207100 108880
rect 207400 108620 207600 108880
rect 207900 108620 208100 108880
rect 208400 108620 208600 108880
rect 208900 108620 209100 108880
rect 209400 108620 209600 108880
rect 209900 108620 210100 108880
rect 210400 108620 210600 108880
rect 210900 108620 211100 108880
rect 211400 108620 211600 108880
rect 211900 108620 212100 108880
rect 212400 108620 212600 108880
rect 212900 108620 213100 108880
rect 213400 108620 213600 108880
rect 213900 108620 214100 108880
rect 214400 108620 214600 108880
rect 214900 108620 215100 108880
rect 215400 108620 215600 108880
rect 215900 108620 216100 108880
rect 216400 108620 216600 108880
rect 216900 108620 217100 108880
rect 217400 108620 217600 108880
rect 217900 108620 218100 108880
rect 218400 108620 218600 108880
rect 218900 108620 219100 108880
rect 219400 108620 219600 108880
rect 219900 108620 220100 108880
rect 220400 108620 220600 108880
rect 220900 108620 221100 108880
rect 221400 108620 221600 108880
rect 221900 108620 222100 108880
rect 222400 108620 222600 108880
rect 222900 108620 223100 108880
rect 223400 108620 223600 108880
rect 223900 108620 224100 108880
rect 224400 108620 224600 108880
rect 224900 108620 225100 108880
rect 225400 108620 225600 108880
rect 225900 108620 226100 108880
rect 226400 108620 226600 108880
rect 226900 108620 227100 108880
rect 227400 108620 227600 108880
rect 227900 108620 228100 108880
rect 228400 108620 228600 108880
rect 228900 108620 229100 108880
rect 229400 108620 229600 108880
rect 229900 108620 230100 108880
rect 230400 108620 230600 108880
rect 230900 108620 231100 108880
rect 231400 108620 231600 108880
rect 231900 108620 232000 108880
rect 178000 108600 178120 108620
rect 178380 108600 178620 108620
rect 178880 108600 179120 108620
rect 179380 108600 179620 108620
rect 179880 108600 180120 108620
rect 180380 108600 180620 108620
rect 180880 108600 181120 108620
rect 181380 108600 181620 108620
rect 181880 108600 182120 108620
rect 182380 108600 182620 108620
rect 182880 108600 183120 108620
rect 183380 108600 183620 108620
rect 183880 108600 184120 108620
rect 184380 108600 184620 108620
rect 184880 108600 185120 108620
rect 185380 108600 185620 108620
rect 185880 108600 186120 108620
rect 186380 108600 186620 108620
rect 186880 108600 187120 108620
rect 187380 108600 187620 108620
rect 187880 108600 188120 108620
rect 188380 108600 188620 108620
rect 188880 108600 189120 108620
rect 189380 108600 189620 108620
rect 189880 108600 190120 108620
rect 190380 108600 190620 108620
rect 190880 108600 191120 108620
rect 191380 108600 191620 108620
rect 191880 108600 192120 108620
rect 192380 108600 192620 108620
rect 192880 108600 193120 108620
rect 193380 108600 193620 108620
rect 193880 108600 194120 108620
rect 194380 108600 194620 108620
rect 194880 108600 195120 108620
rect 195380 108600 195620 108620
rect 195880 108600 196120 108620
rect 196380 108600 196620 108620
rect 196880 108600 197120 108620
rect 197380 108600 197620 108620
rect 197880 108600 198120 108620
rect 198380 108600 198620 108620
rect 198880 108600 199120 108620
rect 199380 108600 199620 108620
rect 199880 108600 200120 108620
rect 200380 108600 200620 108620
rect 200880 108600 201120 108620
rect 201380 108600 201620 108620
rect 201880 108600 202120 108620
rect 202380 108600 202620 108620
rect 202880 108600 203120 108620
rect 203380 108600 203620 108620
rect 203880 108600 204120 108620
rect 204380 108600 204620 108620
rect 204880 108600 205120 108620
rect 205380 108600 205620 108620
rect 205880 108600 206120 108620
rect 206380 108600 206620 108620
rect 206880 108600 207120 108620
rect 207380 108600 207620 108620
rect 207880 108600 208120 108620
rect 208380 108600 208620 108620
rect 208880 108600 209120 108620
rect 209380 108600 209620 108620
rect 209880 108600 210120 108620
rect 210380 108600 210620 108620
rect 210880 108600 211120 108620
rect 211380 108600 211620 108620
rect 211880 108600 212120 108620
rect 212380 108600 212620 108620
rect 212880 108600 213120 108620
rect 213380 108600 213620 108620
rect 213880 108600 214120 108620
rect 214380 108600 214620 108620
rect 214880 108600 215120 108620
rect 215380 108600 215620 108620
rect 215880 108600 216120 108620
rect 216380 108600 216620 108620
rect 216880 108600 217120 108620
rect 217380 108600 217620 108620
rect 217880 108600 218120 108620
rect 218380 108600 218620 108620
rect 218880 108600 219120 108620
rect 219380 108600 219620 108620
rect 219880 108600 220120 108620
rect 220380 108600 220620 108620
rect 220880 108600 221120 108620
rect 221380 108600 221620 108620
rect 221880 108600 222120 108620
rect 222380 108600 222620 108620
rect 222880 108600 223120 108620
rect 223380 108600 223620 108620
rect 223880 108600 224120 108620
rect 224380 108600 224620 108620
rect 224880 108600 225120 108620
rect 225380 108600 225620 108620
rect 225880 108600 226120 108620
rect 226380 108600 226620 108620
rect 226880 108600 227120 108620
rect 227380 108600 227620 108620
rect 227880 108600 228120 108620
rect 228380 108600 228620 108620
rect 228880 108600 229120 108620
rect 229380 108600 229620 108620
rect 229880 108600 230120 108620
rect 230380 108600 230620 108620
rect 230880 108600 231120 108620
rect 231380 108600 231620 108620
rect 231880 108600 232000 108620
rect 178000 108400 232000 108600
rect 178000 108380 178120 108400
rect 178380 108380 178620 108400
rect 178880 108380 179120 108400
rect 179380 108380 179620 108400
rect 179880 108380 180120 108400
rect 180380 108380 180620 108400
rect 180880 108380 181120 108400
rect 181380 108380 181620 108400
rect 181880 108380 182120 108400
rect 182380 108380 182620 108400
rect 182880 108380 183120 108400
rect 183380 108380 183620 108400
rect 183880 108380 184120 108400
rect 184380 108380 184620 108400
rect 184880 108380 185120 108400
rect 185380 108380 185620 108400
rect 185880 108380 186120 108400
rect 186380 108380 186620 108400
rect 186880 108380 187120 108400
rect 187380 108380 187620 108400
rect 187880 108380 188120 108400
rect 188380 108380 188620 108400
rect 188880 108380 189120 108400
rect 189380 108380 189620 108400
rect 189880 108380 190120 108400
rect 190380 108380 190620 108400
rect 190880 108380 191120 108400
rect 191380 108380 191620 108400
rect 191880 108380 192120 108400
rect 192380 108380 192620 108400
rect 192880 108380 193120 108400
rect 193380 108380 193620 108400
rect 193880 108380 194120 108400
rect 194380 108380 194620 108400
rect 194880 108380 195120 108400
rect 195380 108380 195620 108400
rect 195880 108380 196120 108400
rect 196380 108380 196620 108400
rect 196880 108380 197120 108400
rect 197380 108380 197620 108400
rect 197880 108380 198120 108400
rect 198380 108380 198620 108400
rect 198880 108380 199120 108400
rect 199380 108380 199620 108400
rect 199880 108380 200120 108400
rect 200380 108380 200620 108400
rect 200880 108380 201120 108400
rect 201380 108380 201620 108400
rect 201880 108380 202120 108400
rect 202380 108380 202620 108400
rect 202880 108380 203120 108400
rect 203380 108380 203620 108400
rect 203880 108380 204120 108400
rect 204380 108380 204620 108400
rect 204880 108380 205120 108400
rect 205380 108380 205620 108400
rect 205880 108380 206120 108400
rect 206380 108380 206620 108400
rect 206880 108380 207120 108400
rect 207380 108380 207620 108400
rect 207880 108380 208120 108400
rect 208380 108380 208620 108400
rect 208880 108380 209120 108400
rect 209380 108380 209620 108400
rect 209880 108380 210120 108400
rect 210380 108380 210620 108400
rect 210880 108380 211120 108400
rect 211380 108380 211620 108400
rect 211880 108380 212120 108400
rect 212380 108380 212620 108400
rect 212880 108380 213120 108400
rect 213380 108380 213620 108400
rect 213880 108380 214120 108400
rect 214380 108380 214620 108400
rect 214880 108380 215120 108400
rect 215380 108380 215620 108400
rect 215880 108380 216120 108400
rect 216380 108380 216620 108400
rect 216880 108380 217120 108400
rect 217380 108380 217620 108400
rect 217880 108380 218120 108400
rect 218380 108380 218620 108400
rect 218880 108380 219120 108400
rect 219380 108380 219620 108400
rect 219880 108380 220120 108400
rect 220380 108380 220620 108400
rect 220880 108380 221120 108400
rect 221380 108380 221620 108400
rect 221880 108380 222120 108400
rect 222380 108380 222620 108400
rect 222880 108380 223120 108400
rect 223380 108380 223620 108400
rect 223880 108380 224120 108400
rect 224380 108380 224620 108400
rect 224880 108380 225120 108400
rect 225380 108380 225620 108400
rect 225880 108380 226120 108400
rect 226380 108380 226620 108400
rect 226880 108380 227120 108400
rect 227380 108380 227620 108400
rect 227880 108380 228120 108400
rect 228380 108380 228620 108400
rect 228880 108380 229120 108400
rect 229380 108380 229620 108400
rect 229880 108380 230120 108400
rect 230380 108380 230620 108400
rect 230880 108380 231120 108400
rect 231380 108380 231620 108400
rect 231880 108380 232000 108400
rect 178000 108120 178100 108380
rect 178400 108120 178600 108380
rect 178900 108120 179100 108380
rect 179400 108120 179600 108380
rect 179900 108120 180100 108380
rect 180400 108120 180600 108380
rect 180900 108120 181100 108380
rect 181400 108120 181600 108380
rect 181900 108120 182100 108380
rect 182400 108120 182600 108380
rect 182900 108120 183100 108380
rect 183400 108120 183600 108380
rect 183900 108120 184100 108380
rect 184400 108120 184600 108380
rect 184900 108120 185100 108380
rect 185400 108120 185600 108380
rect 185900 108120 186100 108380
rect 186400 108120 186600 108380
rect 186900 108120 187100 108380
rect 187400 108120 187600 108380
rect 187900 108120 188100 108380
rect 188400 108120 188600 108380
rect 188900 108120 189100 108380
rect 189400 108120 189600 108380
rect 189900 108120 190100 108380
rect 190400 108120 190600 108380
rect 190900 108120 191100 108380
rect 191400 108120 191600 108380
rect 191900 108120 192100 108380
rect 192400 108120 192600 108380
rect 192900 108120 193100 108380
rect 193400 108120 193600 108380
rect 193900 108120 194100 108380
rect 194400 108120 194600 108380
rect 194900 108120 195100 108380
rect 195400 108120 195600 108380
rect 195900 108120 196100 108380
rect 196400 108120 196600 108380
rect 196900 108120 197100 108380
rect 197400 108120 197600 108380
rect 197900 108120 198100 108380
rect 198400 108120 198600 108380
rect 198900 108120 199100 108380
rect 199400 108120 199600 108380
rect 199900 108120 200100 108380
rect 200400 108120 200600 108380
rect 200900 108120 201100 108380
rect 201400 108120 201600 108380
rect 201900 108120 202100 108380
rect 202400 108120 202600 108380
rect 202900 108120 203100 108380
rect 203400 108120 203600 108380
rect 203900 108120 204100 108380
rect 204400 108120 204600 108380
rect 204900 108120 205100 108380
rect 205400 108120 205600 108380
rect 205900 108120 206100 108380
rect 206400 108120 206600 108380
rect 206900 108120 207100 108380
rect 207400 108120 207600 108380
rect 207900 108120 208100 108380
rect 208400 108120 208600 108380
rect 208900 108120 209100 108380
rect 209400 108120 209600 108380
rect 209900 108120 210100 108380
rect 210400 108120 210600 108380
rect 210900 108120 211100 108380
rect 211400 108120 211600 108380
rect 211900 108120 212100 108380
rect 212400 108120 212600 108380
rect 212900 108120 213100 108380
rect 213400 108120 213600 108380
rect 213900 108120 214100 108380
rect 214400 108120 214600 108380
rect 214900 108120 215100 108380
rect 215400 108120 215600 108380
rect 215900 108120 216100 108380
rect 216400 108120 216600 108380
rect 216900 108120 217100 108380
rect 217400 108120 217600 108380
rect 217900 108120 218100 108380
rect 218400 108120 218600 108380
rect 218900 108120 219100 108380
rect 219400 108120 219600 108380
rect 219900 108120 220100 108380
rect 220400 108120 220600 108380
rect 220900 108120 221100 108380
rect 221400 108120 221600 108380
rect 221900 108120 222100 108380
rect 222400 108120 222600 108380
rect 222900 108120 223100 108380
rect 223400 108120 223600 108380
rect 223900 108120 224100 108380
rect 224400 108120 224600 108380
rect 224900 108120 225100 108380
rect 225400 108120 225600 108380
rect 225900 108120 226100 108380
rect 226400 108120 226600 108380
rect 226900 108120 227100 108380
rect 227400 108120 227600 108380
rect 227900 108120 228100 108380
rect 228400 108120 228600 108380
rect 228900 108120 229100 108380
rect 229400 108120 229600 108380
rect 229900 108120 230100 108380
rect 230400 108120 230600 108380
rect 230900 108120 231100 108380
rect 231400 108120 231600 108380
rect 231900 108120 232000 108380
rect 178000 108100 178120 108120
rect 178380 108100 178620 108120
rect 178880 108100 179120 108120
rect 179380 108100 179620 108120
rect 179880 108100 180120 108120
rect 180380 108100 180620 108120
rect 180880 108100 181120 108120
rect 181380 108100 181620 108120
rect 181880 108100 182120 108120
rect 182380 108100 182620 108120
rect 182880 108100 183120 108120
rect 183380 108100 183620 108120
rect 183880 108100 184120 108120
rect 184380 108100 184620 108120
rect 184880 108100 185120 108120
rect 185380 108100 185620 108120
rect 185880 108100 186120 108120
rect 186380 108100 186620 108120
rect 186880 108100 187120 108120
rect 187380 108100 187620 108120
rect 187880 108100 188120 108120
rect 188380 108100 188620 108120
rect 188880 108100 189120 108120
rect 189380 108100 189620 108120
rect 189880 108100 190120 108120
rect 190380 108100 190620 108120
rect 190880 108100 191120 108120
rect 191380 108100 191620 108120
rect 191880 108100 192120 108120
rect 192380 108100 192620 108120
rect 192880 108100 193120 108120
rect 193380 108100 193620 108120
rect 193880 108100 194120 108120
rect 194380 108100 194620 108120
rect 194880 108100 195120 108120
rect 195380 108100 195620 108120
rect 195880 108100 196120 108120
rect 196380 108100 196620 108120
rect 196880 108100 197120 108120
rect 197380 108100 197620 108120
rect 197880 108100 198120 108120
rect 198380 108100 198620 108120
rect 198880 108100 199120 108120
rect 199380 108100 199620 108120
rect 199880 108100 200120 108120
rect 200380 108100 200620 108120
rect 200880 108100 201120 108120
rect 201380 108100 201620 108120
rect 201880 108100 202120 108120
rect 202380 108100 202620 108120
rect 202880 108100 203120 108120
rect 203380 108100 203620 108120
rect 203880 108100 204120 108120
rect 204380 108100 204620 108120
rect 204880 108100 205120 108120
rect 205380 108100 205620 108120
rect 205880 108100 206120 108120
rect 206380 108100 206620 108120
rect 206880 108100 207120 108120
rect 207380 108100 207620 108120
rect 207880 108100 208120 108120
rect 208380 108100 208620 108120
rect 208880 108100 209120 108120
rect 209380 108100 209620 108120
rect 209880 108100 210120 108120
rect 210380 108100 210620 108120
rect 210880 108100 211120 108120
rect 211380 108100 211620 108120
rect 211880 108100 212120 108120
rect 212380 108100 212620 108120
rect 212880 108100 213120 108120
rect 213380 108100 213620 108120
rect 213880 108100 214120 108120
rect 214380 108100 214620 108120
rect 214880 108100 215120 108120
rect 215380 108100 215620 108120
rect 215880 108100 216120 108120
rect 216380 108100 216620 108120
rect 216880 108100 217120 108120
rect 217380 108100 217620 108120
rect 217880 108100 218120 108120
rect 218380 108100 218620 108120
rect 218880 108100 219120 108120
rect 219380 108100 219620 108120
rect 219880 108100 220120 108120
rect 220380 108100 220620 108120
rect 220880 108100 221120 108120
rect 221380 108100 221620 108120
rect 221880 108100 222120 108120
rect 222380 108100 222620 108120
rect 222880 108100 223120 108120
rect 223380 108100 223620 108120
rect 223880 108100 224120 108120
rect 224380 108100 224620 108120
rect 224880 108100 225120 108120
rect 225380 108100 225620 108120
rect 225880 108100 226120 108120
rect 226380 108100 226620 108120
rect 226880 108100 227120 108120
rect 227380 108100 227620 108120
rect 227880 108100 228120 108120
rect 228380 108100 228620 108120
rect 228880 108100 229120 108120
rect 229380 108100 229620 108120
rect 229880 108100 230120 108120
rect 230380 108100 230620 108120
rect 230880 108100 231120 108120
rect 231380 108100 231620 108120
rect 231880 108100 232000 108120
rect 178000 107900 232000 108100
rect 178000 107880 178120 107900
rect 178380 107880 178620 107900
rect 178880 107880 179120 107900
rect 179380 107880 179620 107900
rect 179880 107880 180120 107900
rect 180380 107880 180620 107900
rect 180880 107880 181120 107900
rect 181380 107880 181620 107900
rect 181880 107880 182120 107900
rect 182380 107880 182620 107900
rect 182880 107880 183120 107900
rect 183380 107880 183620 107900
rect 183880 107880 184120 107900
rect 184380 107880 184620 107900
rect 184880 107880 185120 107900
rect 185380 107880 185620 107900
rect 185880 107880 186120 107900
rect 186380 107880 186620 107900
rect 186880 107880 187120 107900
rect 187380 107880 187620 107900
rect 187880 107880 188120 107900
rect 188380 107880 188620 107900
rect 188880 107880 189120 107900
rect 189380 107880 189620 107900
rect 189880 107880 190120 107900
rect 190380 107880 190620 107900
rect 190880 107880 191120 107900
rect 191380 107880 191620 107900
rect 191880 107880 192120 107900
rect 192380 107880 192620 107900
rect 192880 107880 193120 107900
rect 193380 107880 193620 107900
rect 193880 107880 194120 107900
rect 194380 107880 194620 107900
rect 194880 107880 195120 107900
rect 195380 107880 195620 107900
rect 195880 107880 196120 107900
rect 196380 107880 196620 107900
rect 196880 107880 197120 107900
rect 197380 107880 197620 107900
rect 197880 107880 198120 107900
rect 198380 107880 198620 107900
rect 198880 107880 199120 107900
rect 199380 107880 199620 107900
rect 199880 107880 200120 107900
rect 200380 107880 200620 107900
rect 200880 107880 201120 107900
rect 201380 107880 201620 107900
rect 201880 107880 202120 107900
rect 202380 107880 202620 107900
rect 202880 107880 203120 107900
rect 203380 107880 203620 107900
rect 203880 107880 204120 107900
rect 204380 107880 204620 107900
rect 204880 107880 205120 107900
rect 205380 107880 205620 107900
rect 205880 107880 206120 107900
rect 206380 107880 206620 107900
rect 206880 107880 207120 107900
rect 207380 107880 207620 107900
rect 207880 107880 208120 107900
rect 208380 107880 208620 107900
rect 208880 107880 209120 107900
rect 209380 107880 209620 107900
rect 209880 107880 210120 107900
rect 210380 107880 210620 107900
rect 210880 107880 211120 107900
rect 211380 107880 211620 107900
rect 211880 107880 212120 107900
rect 212380 107880 212620 107900
rect 212880 107880 213120 107900
rect 213380 107880 213620 107900
rect 213880 107880 214120 107900
rect 214380 107880 214620 107900
rect 214880 107880 215120 107900
rect 215380 107880 215620 107900
rect 215880 107880 216120 107900
rect 216380 107880 216620 107900
rect 216880 107880 217120 107900
rect 217380 107880 217620 107900
rect 217880 107880 218120 107900
rect 218380 107880 218620 107900
rect 218880 107880 219120 107900
rect 219380 107880 219620 107900
rect 219880 107880 220120 107900
rect 220380 107880 220620 107900
rect 220880 107880 221120 107900
rect 221380 107880 221620 107900
rect 221880 107880 222120 107900
rect 222380 107880 222620 107900
rect 222880 107880 223120 107900
rect 223380 107880 223620 107900
rect 223880 107880 224120 107900
rect 224380 107880 224620 107900
rect 224880 107880 225120 107900
rect 225380 107880 225620 107900
rect 225880 107880 226120 107900
rect 226380 107880 226620 107900
rect 226880 107880 227120 107900
rect 227380 107880 227620 107900
rect 227880 107880 228120 107900
rect 228380 107880 228620 107900
rect 228880 107880 229120 107900
rect 229380 107880 229620 107900
rect 229880 107880 230120 107900
rect 230380 107880 230620 107900
rect 230880 107880 231120 107900
rect 231380 107880 231620 107900
rect 231880 107880 232000 107900
rect 178000 107620 178100 107880
rect 178400 107620 178600 107880
rect 178900 107620 179100 107880
rect 179400 107620 179600 107880
rect 179900 107620 180100 107880
rect 180400 107620 180600 107880
rect 180900 107620 181100 107880
rect 181400 107620 181600 107880
rect 181900 107620 182100 107880
rect 182400 107620 182600 107880
rect 182900 107620 183100 107880
rect 183400 107620 183600 107880
rect 183900 107620 184100 107880
rect 184400 107620 184600 107880
rect 184900 107620 185100 107880
rect 185400 107620 185600 107880
rect 185900 107620 186100 107880
rect 186400 107620 186600 107880
rect 186900 107620 187100 107880
rect 187400 107620 187600 107880
rect 187900 107620 188100 107880
rect 188400 107620 188600 107880
rect 188900 107620 189100 107880
rect 189400 107620 189600 107880
rect 189900 107620 190100 107880
rect 190400 107620 190600 107880
rect 190900 107620 191100 107880
rect 191400 107620 191600 107880
rect 191900 107620 192100 107880
rect 192400 107620 192600 107880
rect 192900 107620 193100 107880
rect 193400 107620 193600 107880
rect 193900 107620 194100 107880
rect 194400 107620 194600 107880
rect 194900 107620 195100 107880
rect 195400 107620 195600 107880
rect 195900 107620 196100 107880
rect 196400 107620 196600 107880
rect 196900 107620 197100 107880
rect 197400 107620 197600 107880
rect 197900 107620 198100 107880
rect 198400 107620 198600 107880
rect 198900 107620 199100 107880
rect 199400 107620 199600 107880
rect 199900 107620 200100 107880
rect 200400 107620 200600 107880
rect 200900 107620 201100 107880
rect 201400 107620 201600 107880
rect 201900 107620 202100 107880
rect 202400 107620 202600 107880
rect 202900 107620 203100 107880
rect 203400 107620 203600 107880
rect 203900 107620 204100 107880
rect 204400 107620 204600 107880
rect 204900 107620 205100 107880
rect 205400 107620 205600 107880
rect 205900 107620 206100 107880
rect 206400 107620 206600 107880
rect 206900 107620 207100 107880
rect 207400 107620 207600 107880
rect 207900 107620 208100 107880
rect 208400 107620 208600 107880
rect 208900 107620 209100 107880
rect 209400 107620 209600 107880
rect 209900 107620 210100 107880
rect 210400 107620 210600 107880
rect 210900 107620 211100 107880
rect 211400 107620 211600 107880
rect 211900 107620 212100 107880
rect 212400 107620 212600 107880
rect 212900 107620 213100 107880
rect 213400 107620 213600 107880
rect 213900 107620 214100 107880
rect 214400 107620 214600 107880
rect 214900 107620 215100 107880
rect 215400 107620 215600 107880
rect 215900 107620 216100 107880
rect 216400 107620 216600 107880
rect 216900 107620 217100 107880
rect 217400 107620 217600 107880
rect 217900 107620 218100 107880
rect 218400 107620 218600 107880
rect 218900 107620 219100 107880
rect 219400 107620 219600 107880
rect 219900 107620 220100 107880
rect 220400 107620 220600 107880
rect 220900 107620 221100 107880
rect 221400 107620 221600 107880
rect 221900 107620 222100 107880
rect 222400 107620 222600 107880
rect 222900 107620 223100 107880
rect 223400 107620 223600 107880
rect 223900 107620 224100 107880
rect 224400 107620 224600 107880
rect 224900 107620 225100 107880
rect 225400 107620 225600 107880
rect 225900 107620 226100 107880
rect 226400 107620 226600 107880
rect 226900 107620 227100 107880
rect 227400 107620 227600 107880
rect 227900 107620 228100 107880
rect 228400 107620 228600 107880
rect 228900 107620 229100 107880
rect 229400 107620 229600 107880
rect 229900 107620 230100 107880
rect 230400 107620 230600 107880
rect 230900 107620 231100 107880
rect 231400 107620 231600 107880
rect 231900 107620 232000 107880
rect 178000 107600 178120 107620
rect 178380 107600 178620 107620
rect 178880 107600 179120 107620
rect 179380 107600 179620 107620
rect 179880 107600 180120 107620
rect 180380 107600 180620 107620
rect 180880 107600 181120 107620
rect 181380 107600 181620 107620
rect 181880 107600 182120 107620
rect 182380 107600 182620 107620
rect 182880 107600 183120 107620
rect 183380 107600 183620 107620
rect 183880 107600 184120 107620
rect 184380 107600 184620 107620
rect 184880 107600 185120 107620
rect 185380 107600 185620 107620
rect 185880 107600 186120 107620
rect 186380 107600 186620 107620
rect 186880 107600 187120 107620
rect 187380 107600 187620 107620
rect 187880 107600 188120 107620
rect 188380 107600 188620 107620
rect 188880 107600 189120 107620
rect 189380 107600 189620 107620
rect 189880 107600 190120 107620
rect 190380 107600 190620 107620
rect 190880 107600 191120 107620
rect 191380 107600 191620 107620
rect 191880 107600 192120 107620
rect 192380 107600 192620 107620
rect 192880 107600 193120 107620
rect 193380 107600 193620 107620
rect 193880 107600 194120 107620
rect 194380 107600 194620 107620
rect 194880 107600 195120 107620
rect 195380 107600 195620 107620
rect 195880 107600 196120 107620
rect 196380 107600 196620 107620
rect 196880 107600 197120 107620
rect 197380 107600 197620 107620
rect 197880 107600 198120 107620
rect 198380 107600 198620 107620
rect 198880 107600 199120 107620
rect 199380 107600 199620 107620
rect 199880 107600 200120 107620
rect 200380 107600 200620 107620
rect 200880 107600 201120 107620
rect 201380 107600 201620 107620
rect 201880 107600 202120 107620
rect 202380 107600 202620 107620
rect 202880 107600 203120 107620
rect 203380 107600 203620 107620
rect 203880 107600 204120 107620
rect 204380 107600 204620 107620
rect 204880 107600 205120 107620
rect 205380 107600 205620 107620
rect 205880 107600 206120 107620
rect 206380 107600 206620 107620
rect 206880 107600 207120 107620
rect 207380 107600 207620 107620
rect 207880 107600 208120 107620
rect 208380 107600 208620 107620
rect 208880 107600 209120 107620
rect 209380 107600 209620 107620
rect 209880 107600 210120 107620
rect 210380 107600 210620 107620
rect 210880 107600 211120 107620
rect 211380 107600 211620 107620
rect 211880 107600 212120 107620
rect 212380 107600 212620 107620
rect 212880 107600 213120 107620
rect 213380 107600 213620 107620
rect 213880 107600 214120 107620
rect 214380 107600 214620 107620
rect 214880 107600 215120 107620
rect 215380 107600 215620 107620
rect 215880 107600 216120 107620
rect 216380 107600 216620 107620
rect 216880 107600 217120 107620
rect 217380 107600 217620 107620
rect 217880 107600 218120 107620
rect 218380 107600 218620 107620
rect 218880 107600 219120 107620
rect 219380 107600 219620 107620
rect 219880 107600 220120 107620
rect 220380 107600 220620 107620
rect 220880 107600 221120 107620
rect 221380 107600 221620 107620
rect 221880 107600 222120 107620
rect 222380 107600 222620 107620
rect 222880 107600 223120 107620
rect 223380 107600 223620 107620
rect 223880 107600 224120 107620
rect 224380 107600 224620 107620
rect 224880 107600 225120 107620
rect 225380 107600 225620 107620
rect 225880 107600 226120 107620
rect 226380 107600 226620 107620
rect 226880 107600 227120 107620
rect 227380 107600 227620 107620
rect 227880 107600 228120 107620
rect 228380 107600 228620 107620
rect 228880 107600 229120 107620
rect 229380 107600 229620 107620
rect 229880 107600 230120 107620
rect 230380 107600 230620 107620
rect 230880 107600 231120 107620
rect 231380 107600 231620 107620
rect 231880 107600 232000 107620
rect 178000 107400 232000 107600
rect 178000 107380 178120 107400
rect 178380 107380 178620 107400
rect 178880 107380 179120 107400
rect 179380 107380 179620 107400
rect 179880 107380 180120 107400
rect 180380 107380 180620 107400
rect 180880 107380 181120 107400
rect 181380 107380 181620 107400
rect 181880 107380 182120 107400
rect 182380 107380 182620 107400
rect 182880 107380 183120 107400
rect 183380 107380 183620 107400
rect 183880 107380 184120 107400
rect 184380 107380 184620 107400
rect 184880 107380 185120 107400
rect 185380 107380 185620 107400
rect 185880 107380 186120 107400
rect 186380 107380 186620 107400
rect 186880 107380 187120 107400
rect 187380 107380 187620 107400
rect 187880 107380 188120 107400
rect 188380 107380 188620 107400
rect 188880 107380 189120 107400
rect 189380 107380 189620 107400
rect 189880 107380 190120 107400
rect 190380 107380 190620 107400
rect 190880 107380 191120 107400
rect 191380 107380 191620 107400
rect 191880 107380 192120 107400
rect 192380 107380 192620 107400
rect 192880 107380 193120 107400
rect 193380 107380 193620 107400
rect 193880 107380 194120 107400
rect 194380 107380 194620 107400
rect 194880 107380 195120 107400
rect 195380 107380 195620 107400
rect 195880 107380 196120 107400
rect 196380 107380 196620 107400
rect 196880 107380 197120 107400
rect 197380 107380 197620 107400
rect 197880 107380 198120 107400
rect 198380 107380 198620 107400
rect 198880 107380 199120 107400
rect 199380 107380 199620 107400
rect 199880 107380 200120 107400
rect 200380 107380 200620 107400
rect 200880 107380 201120 107400
rect 201380 107380 201620 107400
rect 201880 107380 202120 107400
rect 202380 107380 202620 107400
rect 202880 107380 203120 107400
rect 203380 107380 203620 107400
rect 203880 107380 204120 107400
rect 204380 107380 204620 107400
rect 204880 107380 205120 107400
rect 205380 107380 205620 107400
rect 205880 107380 206120 107400
rect 206380 107380 206620 107400
rect 206880 107380 207120 107400
rect 207380 107380 207620 107400
rect 207880 107380 208120 107400
rect 208380 107380 208620 107400
rect 208880 107380 209120 107400
rect 209380 107380 209620 107400
rect 209880 107380 210120 107400
rect 210380 107380 210620 107400
rect 210880 107380 211120 107400
rect 211380 107380 211620 107400
rect 211880 107380 212120 107400
rect 212380 107380 212620 107400
rect 212880 107380 213120 107400
rect 213380 107380 213620 107400
rect 213880 107380 214120 107400
rect 214380 107380 214620 107400
rect 214880 107380 215120 107400
rect 215380 107380 215620 107400
rect 215880 107380 216120 107400
rect 216380 107380 216620 107400
rect 216880 107380 217120 107400
rect 217380 107380 217620 107400
rect 217880 107380 218120 107400
rect 218380 107380 218620 107400
rect 218880 107380 219120 107400
rect 219380 107380 219620 107400
rect 219880 107380 220120 107400
rect 220380 107380 220620 107400
rect 220880 107380 221120 107400
rect 221380 107380 221620 107400
rect 221880 107380 222120 107400
rect 222380 107380 222620 107400
rect 222880 107380 223120 107400
rect 223380 107380 223620 107400
rect 223880 107380 224120 107400
rect 224380 107380 224620 107400
rect 224880 107380 225120 107400
rect 225380 107380 225620 107400
rect 225880 107380 226120 107400
rect 226380 107380 226620 107400
rect 226880 107380 227120 107400
rect 227380 107380 227620 107400
rect 227880 107380 228120 107400
rect 228380 107380 228620 107400
rect 228880 107380 229120 107400
rect 229380 107380 229620 107400
rect 229880 107380 230120 107400
rect 230380 107380 230620 107400
rect 230880 107380 231120 107400
rect 231380 107380 231620 107400
rect 231880 107380 232000 107400
rect 178000 107120 178100 107380
rect 178400 107120 178600 107380
rect 178900 107120 179100 107380
rect 179400 107120 179600 107380
rect 179900 107120 180100 107380
rect 180400 107120 180600 107380
rect 180900 107120 181100 107380
rect 181400 107120 181600 107380
rect 181900 107120 182100 107380
rect 182400 107120 182600 107380
rect 182900 107120 183100 107380
rect 183400 107120 183600 107380
rect 183900 107120 184100 107380
rect 184400 107120 184600 107380
rect 184900 107120 185100 107380
rect 185400 107120 185600 107380
rect 185900 107120 186100 107380
rect 186400 107120 186600 107380
rect 186900 107120 187100 107380
rect 187400 107120 187600 107380
rect 187900 107120 188100 107380
rect 188400 107120 188600 107380
rect 188900 107120 189100 107380
rect 189400 107120 189600 107380
rect 189900 107120 190100 107380
rect 190400 107120 190600 107380
rect 190900 107120 191100 107380
rect 191400 107120 191600 107380
rect 191900 107120 192100 107380
rect 192400 107120 192600 107380
rect 192900 107120 193100 107380
rect 193400 107120 193600 107380
rect 193900 107120 194100 107380
rect 194400 107120 194600 107380
rect 194900 107120 195100 107380
rect 195400 107120 195600 107380
rect 195900 107120 196100 107380
rect 196400 107120 196600 107380
rect 196900 107120 197100 107380
rect 197400 107120 197600 107380
rect 197900 107120 198100 107380
rect 198400 107120 198600 107380
rect 198900 107120 199100 107380
rect 199400 107120 199600 107380
rect 199900 107120 200100 107380
rect 200400 107120 200600 107380
rect 200900 107120 201100 107380
rect 201400 107120 201600 107380
rect 201900 107120 202100 107380
rect 202400 107120 202600 107380
rect 202900 107120 203100 107380
rect 203400 107120 203600 107380
rect 203900 107120 204100 107380
rect 204400 107120 204600 107380
rect 204900 107120 205100 107380
rect 205400 107120 205600 107380
rect 205900 107120 206100 107380
rect 206400 107120 206600 107380
rect 206900 107120 207100 107380
rect 207400 107120 207600 107380
rect 207900 107120 208100 107380
rect 208400 107120 208600 107380
rect 208900 107120 209100 107380
rect 209400 107120 209600 107380
rect 209900 107120 210100 107380
rect 210400 107120 210600 107380
rect 210900 107120 211100 107380
rect 211400 107120 211600 107380
rect 211900 107120 212100 107380
rect 212400 107120 212600 107380
rect 212900 107120 213100 107380
rect 213400 107120 213600 107380
rect 213900 107120 214100 107380
rect 214400 107120 214600 107380
rect 214900 107120 215100 107380
rect 215400 107120 215600 107380
rect 215900 107120 216100 107380
rect 216400 107120 216600 107380
rect 216900 107120 217100 107380
rect 217400 107120 217600 107380
rect 217900 107120 218100 107380
rect 218400 107120 218600 107380
rect 218900 107120 219100 107380
rect 219400 107120 219600 107380
rect 219900 107120 220100 107380
rect 220400 107120 220600 107380
rect 220900 107120 221100 107380
rect 221400 107120 221600 107380
rect 221900 107120 222100 107380
rect 222400 107120 222600 107380
rect 222900 107120 223100 107380
rect 223400 107120 223600 107380
rect 223900 107120 224100 107380
rect 224400 107120 224600 107380
rect 224900 107120 225100 107380
rect 225400 107120 225600 107380
rect 225900 107120 226100 107380
rect 226400 107120 226600 107380
rect 226900 107120 227100 107380
rect 227400 107120 227600 107380
rect 227900 107120 228100 107380
rect 228400 107120 228600 107380
rect 228900 107120 229100 107380
rect 229400 107120 229600 107380
rect 229900 107120 230100 107380
rect 230400 107120 230600 107380
rect 230900 107120 231100 107380
rect 231400 107120 231600 107380
rect 231900 107120 232000 107380
rect 178000 107100 178120 107120
rect 178380 107100 178620 107120
rect 178880 107100 179120 107120
rect 179380 107100 179620 107120
rect 179880 107100 180120 107120
rect 180380 107100 180620 107120
rect 180880 107100 181120 107120
rect 181380 107100 181620 107120
rect 181880 107100 182120 107120
rect 182380 107100 182620 107120
rect 182880 107100 183120 107120
rect 183380 107100 183620 107120
rect 183880 107100 184120 107120
rect 184380 107100 184620 107120
rect 184880 107100 185120 107120
rect 185380 107100 185620 107120
rect 185880 107100 186120 107120
rect 186380 107100 186620 107120
rect 186880 107100 187120 107120
rect 187380 107100 187620 107120
rect 187880 107100 188120 107120
rect 188380 107100 188620 107120
rect 188880 107100 189120 107120
rect 189380 107100 189620 107120
rect 189880 107100 190120 107120
rect 190380 107100 190620 107120
rect 190880 107100 191120 107120
rect 191380 107100 191620 107120
rect 191880 107100 192120 107120
rect 192380 107100 192620 107120
rect 192880 107100 193120 107120
rect 193380 107100 193620 107120
rect 193880 107100 194120 107120
rect 194380 107100 194620 107120
rect 194880 107100 195120 107120
rect 195380 107100 195620 107120
rect 195880 107100 196120 107120
rect 196380 107100 196620 107120
rect 196880 107100 197120 107120
rect 197380 107100 197620 107120
rect 197880 107100 198120 107120
rect 198380 107100 198620 107120
rect 198880 107100 199120 107120
rect 199380 107100 199620 107120
rect 199880 107100 200120 107120
rect 200380 107100 200620 107120
rect 200880 107100 201120 107120
rect 201380 107100 201620 107120
rect 201880 107100 202120 107120
rect 202380 107100 202620 107120
rect 202880 107100 203120 107120
rect 203380 107100 203620 107120
rect 203880 107100 204120 107120
rect 204380 107100 204620 107120
rect 204880 107100 205120 107120
rect 205380 107100 205620 107120
rect 205880 107100 206120 107120
rect 206380 107100 206620 107120
rect 206880 107100 207120 107120
rect 207380 107100 207620 107120
rect 207880 107100 208120 107120
rect 208380 107100 208620 107120
rect 208880 107100 209120 107120
rect 209380 107100 209620 107120
rect 209880 107100 210120 107120
rect 210380 107100 210620 107120
rect 210880 107100 211120 107120
rect 211380 107100 211620 107120
rect 211880 107100 212120 107120
rect 212380 107100 212620 107120
rect 212880 107100 213120 107120
rect 213380 107100 213620 107120
rect 213880 107100 214120 107120
rect 214380 107100 214620 107120
rect 214880 107100 215120 107120
rect 215380 107100 215620 107120
rect 215880 107100 216120 107120
rect 216380 107100 216620 107120
rect 216880 107100 217120 107120
rect 217380 107100 217620 107120
rect 217880 107100 218120 107120
rect 218380 107100 218620 107120
rect 218880 107100 219120 107120
rect 219380 107100 219620 107120
rect 219880 107100 220120 107120
rect 220380 107100 220620 107120
rect 220880 107100 221120 107120
rect 221380 107100 221620 107120
rect 221880 107100 222120 107120
rect 222380 107100 222620 107120
rect 222880 107100 223120 107120
rect 223380 107100 223620 107120
rect 223880 107100 224120 107120
rect 224380 107100 224620 107120
rect 224880 107100 225120 107120
rect 225380 107100 225620 107120
rect 225880 107100 226120 107120
rect 226380 107100 226620 107120
rect 226880 107100 227120 107120
rect 227380 107100 227620 107120
rect 227880 107100 228120 107120
rect 228380 107100 228620 107120
rect 228880 107100 229120 107120
rect 229380 107100 229620 107120
rect 229880 107100 230120 107120
rect 230380 107100 230620 107120
rect 230880 107100 231120 107120
rect 231380 107100 231620 107120
rect 231880 107100 232000 107120
rect 178000 106900 232000 107100
rect 178000 106880 178120 106900
rect 178380 106880 178620 106900
rect 178880 106880 179120 106900
rect 179380 106880 179620 106900
rect 179880 106880 180120 106900
rect 180380 106880 180620 106900
rect 180880 106880 181120 106900
rect 181380 106880 181620 106900
rect 181880 106880 182120 106900
rect 182380 106880 182620 106900
rect 182880 106880 183120 106900
rect 183380 106880 183620 106900
rect 183880 106880 184120 106900
rect 184380 106880 184620 106900
rect 184880 106880 185120 106900
rect 185380 106880 185620 106900
rect 185880 106880 186120 106900
rect 186380 106880 186620 106900
rect 186880 106880 187120 106900
rect 187380 106880 187620 106900
rect 187880 106880 188120 106900
rect 188380 106880 188620 106900
rect 188880 106880 189120 106900
rect 189380 106880 189620 106900
rect 189880 106880 190120 106900
rect 190380 106880 190620 106900
rect 190880 106880 191120 106900
rect 191380 106880 191620 106900
rect 191880 106880 192120 106900
rect 192380 106880 192620 106900
rect 192880 106880 193120 106900
rect 193380 106880 193620 106900
rect 193880 106880 194120 106900
rect 194380 106880 194620 106900
rect 194880 106880 195120 106900
rect 195380 106880 195620 106900
rect 195880 106880 196120 106900
rect 196380 106880 196620 106900
rect 196880 106880 197120 106900
rect 197380 106880 197620 106900
rect 197880 106880 198120 106900
rect 198380 106880 198620 106900
rect 198880 106880 199120 106900
rect 199380 106880 199620 106900
rect 199880 106880 200120 106900
rect 200380 106880 200620 106900
rect 200880 106880 201120 106900
rect 201380 106880 201620 106900
rect 201880 106880 202120 106900
rect 202380 106880 202620 106900
rect 202880 106880 203120 106900
rect 203380 106880 203620 106900
rect 203880 106880 204120 106900
rect 204380 106880 204620 106900
rect 204880 106880 205120 106900
rect 205380 106880 205620 106900
rect 205880 106880 206120 106900
rect 206380 106880 206620 106900
rect 206880 106880 207120 106900
rect 207380 106880 207620 106900
rect 207880 106880 208120 106900
rect 208380 106880 208620 106900
rect 208880 106880 209120 106900
rect 209380 106880 209620 106900
rect 209880 106880 210120 106900
rect 210380 106880 210620 106900
rect 210880 106880 211120 106900
rect 211380 106880 211620 106900
rect 211880 106880 212120 106900
rect 212380 106880 212620 106900
rect 212880 106880 213120 106900
rect 213380 106880 213620 106900
rect 213880 106880 214120 106900
rect 214380 106880 214620 106900
rect 214880 106880 215120 106900
rect 215380 106880 215620 106900
rect 215880 106880 216120 106900
rect 216380 106880 216620 106900
rect 216880 106880 217120 106900
rect 217380 106880 217620 106900
rect 217880 106880 218120 106900
rect 218380 106880 218620 106900
rect 218880 106880 219120 106900
rect 219380 106880 219620 106900
rect 219880 106880 220120 106900
rect 220380 106880 220620 106900
rect 220880 106880 221120 106900
rect 221380 106880 221620 106900
rect 221880 106880 222120 106900
rect 222380 106880 222620 106900
rect 222880 106880 223120 106900
rect 223380 106880 223620 106900
rect 223880 106880 224120 106900
rect 224380 106880 224620 106900
rect 224880 106880 225120 106900
rect 225380 106880 225620 106900
rect 225880 106880 226120 106900
rect 226380 106880 226620 106900
rect 226880 106880 227120 106900
rect 227380 106880 227620 106900
rect 227880 106880 228120 106900
rect 228380 106880 228620 106900
rect 228880 106880 229120 106900
rect 229380 106880 229620 106900
rect 229880 106880 230120 106900
rect 230380 106880 230620 106900
rect 230880 106880 231120 106900
rect 231380 106880 231620 106900
rect 231880 106880 232000 106900
rect 178000 106620 178100 106880
rect 178400 106620 178600 106880
rect 178900 106620 179100 106880
rect 179400 106620 179600 106880
rect 179900 106620 180100 106880
rect 180400 106620 180600 106880
rect 180900 106620 181100 106880
rect 181400 106620 181600 106880
rect 181900 106620 182100 106880
rect 182400 106620 182600 106880
rect 182900 106620 183100 106880
rect 183400 106620 183600 106880
rect 183900 106620 184100 106880
rect 184400 106620 184600 106880
rect 184900 106620 185100 106880
rect 185400 106620 185600 106880
rect 185900 106620 186100 106880
rect 186400 106620 186600 106880
rect 186900 106620 187100 106880
rect 187400 106620 187600 106880
rect 187900 106620 188100 106880
rect 188400 106620 188600 106880
rect 188900 106620 189100 106880
rect 189400 106620 189600 106880
rect 189900 106620 190100 106880
rect 190400 106620 190600 106880
rect 190900 106620 191100 106880
rect 191400 106620 191600 106880
rect 191900 106620 192100 106880
rect 192400 106620 192600 106880
rect 192900 106620 193100 106880
rect 193400 106620 193600 106880
rect 193900 106620 194100 106880
rect 194400 106620 194600 106880
rect 194900 106620 195100 106880
rect 195400 106620 195600 106880
rect 195900 106620 196100 106880
rect 196400 106620 196600 106880
rect 196900 106620 197100 106880
rect 197400 106620 197600 106880
rect 197900 106620 198100 106880
rect 198400 106620 198600 106880
rect 198900 106620 199100 106880
rect 199400 106620 199600 106880
rect 199900 106620 200100 106880
rect 200400 106620 200600 106880
rect 200900 106620 201100 106880
rect 201400 106620 201600 106880
rect 201900 106620 202100 106880
rect 202400 106620 202600 106880
rect 202900 106620 203100 106880
rect 203400 106620 203600 106880
rect 203900 106620 204100 106880
rect 204400 106620 204600 106880
rect 204900 106620 205100 106880
rect 205400 106620 205600 106880
rect 205900 106620 206100 106880
rect 206400 106620 206600 106880
rect 206900 106620 207100 106880
rect 207400 106620 207600 106880
rect 207900 106620 208100 106880
rect 208400 106620 208600 106880
rect 208900 106620 209100 106880
rect 209400 106620 209600 106880
rect 209900 106620 210100 106880
rect 210400 106620 210600 106880
rect 210900 106620 211100 106880
rect 211400 106620 211600 106880
rect 211900 106620 212100 106880
rect 212400 106620 212600 106880
rect 212900 106620 213100 106880
rect 213400 106620 213600 106880
rect 213900 106620 214100 106880
rect 214400 106620 214600 106880
rect 214900 106620 215100 106880
rect 215400 106620 215600 106880
rect 215900 106620 216100 106880
rect 216400 106620 216600 106880
rect 216900 106620 217100 106880
rect 217400 106620 217600 106880
rect 217900 106620 218100 106880
rect 218400 106620 218600 106880
rect 218900 106620 219100 106880
rect 219400 106620 219600 106880
rect 219900 106620 220100 106880
rect 220400 106620 220600 106880
rect 220900 106620 221100 106880
rect 221400 106620 221600 106880
rect 221900 106620 222100 106880
rect 222400 106620 222600 106880
rect 222900 106620 223100 106880
rect 223400 106620 223600 106880
rect 223900 106620 224100 106880
rect 224400 106620 224600 106880
rect 224900 106620 225100 106880
rect 225400 106620 225600 106880
rect 225900 106620 226100 106880
rect 226400 106620 226600 106880
rect 226900 106620 227100 106880
rect 227400 106620 227600 106880
rect 227900 106620 228100 106880
rect 228400 106620 228600 106880
rect 228900 106620 229100 106880
rect 229400 106620 229600 106880
rect 229900 106620 230100 106880
rect 230400 106620 230600 106880
rect 230900 106620 231100 106880
rect 231400 106620 231600 106880
rect 231900 106620 232000 106880
rect 178000 106600 178120 106620
rect 178380 106600 178620 106620
rect 178880 106600 179120 106620
rect 179380 106600 179620 106620
rect 179880 106600 180120 106620
rect 180380 106600 180620 106620
rect 180880 106600 181120 106620
rect 181380 106600 181620 106620
rect 181880 106600 182120 106620
rect 182380 106600 182620 106620
rect 182880 106600 183120 106620
rect 183380 106600 183620 106620
rect 183880 106600 184120 106620
rect 184380 106600 184620 106620
rect 184880 106600 185120 106620
rect 185380 106600 185620 106620
rect 185880 106600 186120 106620
rect 186380 106600 186620 106620
rect 186880 106600 187120 106620
rect 187380 106600 187620 106620
rect 187880 106600 188120 106620
rect 188380 106600 188620 106620
rect 188880 106600 189120 106620
rect 189380 106600 189620 106620
rect 189880 106600 190120 106620
rect 190380 106600 190620 106620
rect 190880 106600 191120 106620
rect 191380 106600 191620 106620
rect 191880 106600 192120 106620
rect 192380 106600 192620 106620
rect 192880 106600 193120 106620
rect 193380 106600 193620 106620
rect 193880 106600 194120 106620
rect 194380 106600 194620 106620
rect 194880 106600 195120 106620
rect 195380 106600 195620 106620
rect 195880 106600 196120 106620
rect 196380 106600 196620 106620
rect 196880 106600 197120 106620
rect 197380 106600 197620 106620
rect 197880 106600 198120 106620
rect 198380 106600 198620 106620
rect 198880 106600 199120 106620
rect 199380 106600 199620 106620
rect 199880 106600 200120 106620
rect 200380 106600 200620 106620
rect 200880 106600 201120 106620
rect 201380 106600 201620 106620
rect 201880 106600 202120 106620
rect 202380 106600 202620 106620
rect 202880 106600 203120 106620
rect 203380 106600 203620 106620
rect 203880 106600 204120 106620
rect 204380 106600 204620 106620
rect 204880 106600 205120 106620
rect 205380 106600 205620 106620
rect 205880 106600 206120 106620
rect 206380 106600 206620 106620
rect 206880 106600 207120 106620
rect 207380 106600 207620 106620
rect 207880 106600 208120 106620
rect 208380 106600 208620 106620
rect 208880 106600 209120 106620
rect 209380 106600 209620 106620
rect 209880 106600 210120 106620
rect 210380 106600 210620 106620
rect 210880 106600 211120 106620
rect 211380 106600 211620 106620
rect 211880 106600 212120 106620
rect 212380 106600 212620 106620
rect 212880 106600 213120 106620
rect 213380 106600 213620 106620
rect 213880 106600 214120 106620
rect 214380 106600 214620 106620
rect 214880 106600 215120 106620
rect 215380 106600 215620 106620
rect 215880 106600 216120 106620
rect 216380 106600 216620 106620
rect 216880 106600 217120 106620
rect 217380 106600 217620 106620
rect 217880 106600 218120 106620
rect 218380 106600 218620 106620
rect 218880 106600 219120 106620
rect 219380 106600 219620 106620
rect 219880 106600 220120 106620
rect 220380 106600 220620 106620
rect 220880 106600 221120 106620
rect 221380 106600 221620 106620
rect 221880 106600 222120 106620
rect 222380 106600 222620 106620
rect 222880 106600 223120 106620
rect 223380 106600 223620 106620
rect 223880 106600 224120 106620
rect 224380 106600 224620 106620
rect 224880 106600 225120 106620
rect 225380 106600 225620 106620
rect 225880 106600 226120 106620
rect 226380 106600 226620 106620
rect 226880 106600 227120 106620
rect 227380 106600 227620 106620
rect 227880 106600 228120 106620
rect 228380 106600 228620 106620
rect 228880 106600 229120 106620
rect 229380 106600 229620 106620
rect 229880 106600 230120 106620
rect 230380 106600 230620 106620
rect 230880 106600 231120 106620
rect 231380 106600 231620 106620
rect 231880 106600 232000 106620
rect 178000 106400 232000 106600
rect 178000 106380 178120 106400
rect 178380 106380 178620 106400
rect 178880 106380 179120 106400
rect 179380 106380 179620 106400
rect 179880 106380 180120 106400
rect 180380 106380 180620 106400
rect 180880 106380 181120 106400
rect 181380 106380 181620 106400
rect 181880 106380 182120 106400
rect 182380 106380 182620 106400
rect 182880 106380 183120 106400
rect 183380 106380 183620 106400
rect 183880 106380 184120 106400
rect 184380 106380 184620 106400
rect 184880 106380 185120 106400
rect 185380 106380 185620 106400
rect 185880 106380 186120 106400
rect 186380 106380 186620 106400
rect 186880 106380 187120 106400
rect 187380 106380 187620 106400
rect 187880 106380 188120 106400
rect 188380 106380 188620 106400
rect 188880 106380 189120 106400
rect 189380 106380 189620 106400
rect 189880 106380 190120 106400
rect 190380 106380 190620 106400
rect 190880 106380 191120 106400
rect 191380 106380 191620 106400
rect 191880 106380 192120 106400
rect 192380 106380 192620 106400
rect 192880 106380 193120 106400
rect 193380 106380 193620 106400
rect 193880 106380 194120 106400
rect 194380 106380 194620 106400
rect 194880 106380 195120 106400
rect 195380 106380 195620 106400
rect 195880 106380 196120 106400
rect 196380 106380 196620 106400
rect 196880 106380 197120 106400
rect 197380 106380 197620 106400
rect 197880 106380 198120 106400
rect 198380 106380 198620 106400
rect 198880 106380 199120 106400
rect 199380 106380 199620 106400
rect 199880 106380 200120 106400
rect 200380 106380 200620 106400
rect 200880 106380 201120 106400
rect 201380 106380 201620 106400
rect 201880 106380 202120 106400
rect 202380 106380 202620 106400
rect 202880 106380 203120 106400
rect 203380 106380 203620 106400
rect 203880 106380 204120 106400
rect 204380 106380 204620 106400
rect 204880 106380 205120 106400
rect 205380 106380 205620 106400
rect 205880 106380 206120 106400
rect 206380 106380 206620 106400
rect 206880 106380 207120 106400
rect 207380 106380 207620 106400
rect 207880 106380 208120 106400
rect 208380 106380 208620 106400
rect 208880 106380 209120 106400
rect 209380 106380 209620 106400
rect 209880 106380 210120 106400
rect 210380 106380 210620 106400
rect 210880 106380 211120 106400
rect 211380 106380 211620 106400
rect 211880 106380 212120 106400
rect 212380 106380 212620 106400
rect 212880 106380 213120 106400
rect 213380 106380 213620 106400
rect 213880 106380 214120 106400
rect 214380 106380 214620 106400
rect 214880 106380 215120 106400
rect 215380 106380 215620 106400
rect 215880 106380 216120 106400
rect 216380 106380 216620 106400
rect 216880 106380 217120 106400
rect 217380 106380 217620 106400
rect 217880 106380 218120 106400
rect 218380 106380 218620 106400
rect 218880 106380 219120 106400
rect 219380 106380 219620 106400
rect 219880 106380 220120 106400
rect 220380 106380 220620 106400
rect 220880 106380 221120 106400
rect 221380 106380 221620 106400
rect 221880 106380 222120 106400
rect 222380 106380 222620 106400
rect 222880 106380 223120 106400
rect 223380 106380 223620 106400
rect 223880 106380 224120 106400
rect 224380 106380 224620 106400
rect 224880 106380 225120 106400
rect 225380 106380 225620 106400
rect 225880 106380 226120 106400
rect 226380 106380 226620 106400
rect 226880 106380 227120 106400
rect 227380 106380 227620 106400
rect 227880 106380 228120 106400
rect 228380 106380 228620 106400
rect 228880 106380 229120 106400
rect 229380 106380 229620 106400
rect 229880 106380 230120 106400
rect 230380 106380 230620 106400
rect 230880 106380 231120 106400
rect 231380 106380 231620 106400
rect 231880 106380 232000 106400
rect 178000 106120 178100 106380
rect 178400 106120 178600 106380
rect 178900 106120 179100 106380
rect 179400 106120 179600 106380
rect 179900 106120 180100 106380
rect 180400 106120 180600 106380
rect 180900 106120 181100 106380
rect 181400 106120 181600 106380
rect 181900 106120 182100 106380
rect 182400 106120 182600 106380
rect 182900 106120 183100 106380
rect 183400 106120 183600 106380
rect 183900 106120 184100 106380
rect 184400 106120 184600 106380
rect 184900 106120 185100 106380
rect 185400 106120 185600 106380
rect 185900 106120 186100 106380
rect 186400 106120 186600 106380
rect 186900 106120 187100 106380
rect 187400 106120 187600 106380
rect 187900 106120 188100 106380
rect 188400 106120 188600 106380
rect 188900 106120 189100 106380
rect 189400 106120 189600 106380
rect 189900 106120 190100 106380
rect 190400 106120 190600 106380
rect 190900 106120 191100 106380
rect 191400 106120 191600 106380
rect 191900 106120 192100 106380
rect 192400 106120 192600 106380
rect 192900 106120 193100 106380
rect 193400 106120 193600 106380
rect 193900 106120 194100 106380
rect 194400 106120 194600 106380
rect 194900 106120 195100 106380
rect 195400 106120 195600 106380
rect 195900 106120 196100 106380
rect 196400 106120 196600 106380
rect 196900 106120 197100 106380
rect 197400 106120 197600 106380
rect 197900 106120 198100 106380
rect 198400 106120 198600 106380
rect 198900 106120 199100 106380
rect 199400 106120 199600 106380
rect 199900 106120 200100 106380
rect 200400 106120 200600 106380
rect 200900 106120 201100 106380
rect 201400 106120 201600 106380
rect 201900 106120 202100 106380
rect 202400 106120 202600 106380
rect 202900 106120 203100 106380
rect 203400 106120 203600 106380
rect 203900 106120 204100 106380
rect 204400 106120 204600 106380
rect 204900 106120 205100 106380
rect 205400 106120 205600 106380
rect 205900 106120 206100 106380
rect 206400 106120 206600 106380
rect 206900 106120 207100 106380
rect 207400 106120 207600 106380
rect 207900 106120 208100 106380
rect 208400 106120 208600 106380
rect 208900 106120 209100 106380
rect 209400 106120 209600 106380
rect 209900 106120 210100 106380
rect 210400 106120 210600 106380
rect 210900 106120 211100 106380
rect 211400 106120 211600 106380
rect 211900 106120 212100 106380
rect 212400 106120 212600 106380
rect 212900 106120 213100 106380
rect 213400 106120 213600 106380
rect 213900 106120 214100 106380
rect 214400 106120 214600 106380
rect 214900 106120 215100 106380
rect 215400 106120 215600 106380
rect 215900 106120 216100 106380
rect 216400 106120 216600 106380
rect 216900 106120 217100 106380
rect 217400 106120 217600 106380
rect 217900 106120 218100 106380
rect 218400 106120 218600 106380
rect 218900 106120 219100 106380
rect 219400 106120 219600 106380
rect 219900 106120 220100 106380
rect 220400 106120 220600 106380
rect 220900 106120 221100 106380
rect 221400 106120 221600 106380
rect 221900 106120 222100 106380
rect 222400 106120 222600 106380
rect 222900 106120 223100 106380
rect 223400 106120 223600 106380
rect 223900 106120 224100 106380
rect 224400 106120 224600 106380
rect 224900 106120 225100 106380
rect 225400 106120 225600 106380
rect 225900 106120 226100 106380
rect 226400 106120 226600 106380
rect 226900 106120 227100 106380
rect 227400 106120 227600 106380
rect 227900 106120 228100 106380
rect 228400 106120 228600 106380
rect 228900 106120 229100 106380
rect 229400 106120 229600 106380
rect 229900 106120 230100 106380
rect 230400 106120 230600 106380
rect 230900 106120 231100 106380
rect 231400 106120 231600 106380
rect 231900 106120 232000 106380
rect 178000 106100 178120 106120
rect 178380 106100 178620 106120
rect 178880 106100 179120 106120
rect 179380 106100 179620 106120
rect 179880 106100 180120 106120
rect 180380 106100 180620 106120
rect 180880 106100 181120 106120
rect 181380 106100 181620 106120
rect 181880 106100 182120 106120
rect 182380 106100 182620 106120
rect 182880 106100 183120 106120
rect 183380 106100 183620 106120
rect 183880 106100 184120 106120
rect 184380 106100 184620 106120
rect 184880 106100 185120 106120
rect 185380 106100 185620 106120
rect 185880 106100 186120 106120
rect 186380 106100 186620 106120
rect 186880 106100 187120 106120
rect 187380 106100 187620 106120
rect 187880 106100 188120 106120
rect 188380 106100 188620 106120
rect 188880 106100 189120 106120
rect 189380 106100 189620 106120
rect 189880 106100 190120 106120
rect 190380 106100 190620 106120
rect 190880 106100 191120 106120
rect 191380 106100 191620 106120
rect 191880 106100 192120 106120
rect 192380 106100 192620 106120
rect 192880 106100 193120 106120
rect 193380 106100 193620 106120
rect 193880 106100 194120 106120
rect 194380 106100 194620 106120
rect 194880 106100 195120 106120
rect 195380 106100 195620 106120
rect 195880 106100 196120 106120
rect 196380 106100 196620 106120
rect 196880 106100 197120 106120
rect 197380 106100 197620 106120
rect 197880 106100 198120 106120
rect 198380 106100 198620 106120
rect 198880 106100 199120 106120
rect 199380 106100 199620 106120
rect 199880 106100 200120 106120
rect 200380 106100 200620 106120
rect 200880 106100 201120 106120
rect 201380 106100 201620 106120
rect 201880 106100 202120 106120
rect 202380 106100 202620 106120
rect 202880 106100 203120 106120
rect 203380 106100 203620 106120
rect 203880 106100 204120 106120
rect 204380 106100 204620 106120
rect 204880 106100 205120 106120
rect 205380 106100 205620 106120
rect 205880 106100 206120 106120
rect 206380 106100 206620 106120
rect 206880 106100 207120 106120
rect 207380 106100 207620 106120
rect 207880 106100 208120 106120
rect 208380 106100 208620 106120
rect 208880 106100 209120 106120
rect 209380 106100 209620 106120
rect 209880 106100 210120 106120
rect 210380 106100 210620 106120
rect 210880 106100 211120 106120
rect 211380 106100 211620 106120
rect 211880 106100 212120 106120
rect 212380 106100 212620 106120
rect 212880 106100 213120 106120
rect 213380 106100 213620 106120
rect 213880 106100 214120 106120
rect 214380 106100 214620 106120
rect 214880 106100 215120 106120
rect 215380 106100 215620 106120
rect 215880 106100 216120 106120
rect 216380 106100 216620 106120
rect 216880 106100 217120 106120
rect 217380 106100 217620 106120
rect 217880 106100 218120 106120
rect 218380 106100 218620 106120
rect 218880 106100 219120 106120
rect 219380 106100 219620 106120
rect 219880 106100 220120 106120
rect 220380 106100 220620 106120
rect 220880 106100 221120 106120
rect 221380 106100 221620 106120
rect 221880 106100 222120 106120
rect 222380 106100 222620 106120
rect 222880 106100 223120 106120
rect 223380 106100 223620 106120
rect 223880 106100 224120 106120
rect 224380 106100 224620 106120
rect 224880 106100 225120 106120
rect 225380 106100 225620 106120
rect 225880 106100 226120 106120
rect 226380 106100 226620 106120
rect 226880 106100 227120 106120
rect 227380 106100 227620 106120
rect 227880 106100 228120 106120
rect 228380 106100 228620 106120
rect 228880 106100 229120 106120
rect 229380 106100 229620 106120
rect 229880 106100 230120 106120
rect 230380 106100 230620 106120
rect 230880 106100 231120 106120
rect 231380 106100 231620 106120
rect 231880 106100 232000 106120
rect 178000 105900 232000 106100
rect 178000 105880 178120 105900
rect 178380 105880 178620 105900
rect 178880 105880 179120 105900
rect 179380 105880 179620 105900
rect 179880 105880 180120 105900
rect 180380 105880 180620 105900
rect 180880 105880 181120 105900
rect 181380 105880 181620 105900
rect 181880 105880 182120 105900
rect 182380 105880 182620 105900
rect 182880 105880 183120 105900
rect 183380 105880 183620 105900
rect 183880 105880 184120 105900
rect 184380 105880 184620 105900
rect 184880 105880 185120 105900
rect 185380 105880 185620 105900
rect 185880 105880 186120 105900
rect 186380 105880 186620 105900
rect 186880 105880 187120 105900
rect 187380 105880 187620 105900
rect 187880 105880 188120 105900
rect 188380 105880 188620 105900
rect 188880 105880 189120 105900
rect 189380 105880 189620 105900
rect 189880 105880 190120 105900
rect 190380 105880 190620 105900
rect 190880 105880 191120 105900
rect 191380 105880 191620 105900
rect 191880 105880 192120 105900
rect 192380 105880 192620 105900
rect 192880 105880 193120 105900
rect 193380 105880 193620 105900
rect 193880 105880 194120 105900
rect 194380 105880 194620 105900
rect 194880 105880 195120 105900
rect 195380 105880 195620 105900
rect 195880 105880 196120 105900
rect 196380 105880 196620 105900
rect 196880 105880 197120 105900
rect 197380 105880 197620 105900
rect 197880 105880 198120 105900
rect 198380 105880 198620 105900
rect 198880 105880 199120 105900
rect 199380 105880 199620 105900
rect 199880 105880 200120 105900
rect 200380 105880 200620 105900
rect 200880 105880 201120 105900
rect 201380 105880 201620 105900
rect 201880 105880 202120 105900
rect 202380 105880 202620 105900
rect 202880 105880 203120 105900
rect 203380 105880 203620 105900
rect 203880 105880 204120 105900
rect 204380 105880 204620 105900
rect 204880 105880 205120 105900
rect 205380 105880 205620 105900
rect 205880 105880 206120 105900
rect 206380 105880 206620 105900
rect 206880 105880 207120 105900
rect 207380 105880 207620 105900
rect 207880 105880 208120 105900
rect 208380 105880 208620 105900
rect 208880 105880 209120 105900
rect 209380 105880 209620 105900
rect 209880 105880 210120 105900
rect 210380 105880 210620 105900
rect 210880 105880 211120 105900
rect 211380 105880 211620 105900
rect 211880 105880 212120 105900
rect 212380 105880 212620 105900
rect 212880 105880 213120 105900
rect 213380 105880 213620 105900
rect 213880 105880 214120 105900
rect 214380 105880 214620 105900
rect 214880 105880 215120 105900
rect 215380 105880 215620 105900
rect 215880 105880 216120 105900
rect 216380 105880 216620 105900
rect 216880 105880 217120 105900
rect 217380 105880 217620 105900
rect 217880 105880 218120 105900
rect 218380 105880 218620 105900
rect 218880 105880 219120 105900
rect 219380 105880 219620 105900
rect 219880 105880 220120 105900
rect 220380 105880 220620 105900
rect 220880 105880 221120 105900
rect 221380 105880 221620 105900
rect 221880 105880 222120 105900
rect 222380 105880 222620 105900
rect 222880 105880 223120 105900
rect 223380 105880 223620 105900
rect 223880 105880 224120 105900
rect 224380 105880 224620 105900
rect 224880 105880 225120 105900
rect 225380 105880 225620 105900
rect 225880 105880 226120 105900
rect 226380 105880 226620 105900
rect 226880 105880 227120 105900
rect 227380 105880 227620 105900
rect 227880 105880 228120 105900
rect 228380 105880 228620 105900
rect 228880 105880 229120 105900
rect 229380 105880 229620 105900
rect 229880 105880 230120 105900
rect 230380 105880 230620 105900
rect 230880 105880 231120 105900
rect 231380 105880 231620 105900
rect 231880 105880 232000 105900
rect 178000 105620 178100 105880
rect 178400 105620 178600 105880
rect 178900 105620 179100 105880
rect 179400 105620 179600 105880
rect 179900 105620 180100 105880
rect 180400 105620 180600 105880
rect 180900 105620 181100 105880
rect 181400 105620 181600 105880
rect 181900 105620 182100 105880
rect 182400 105620 182600 105880
rect 182900 105620 183100 105880
rect 183400 105620 183600 105880
rect 183900 105620 184100 105880
rect 184400 105620 184600 105880
rect 184900 105620 185100 105880
rect 185400 105620 185600 105880
rect 185900 105620 186100 105880
rect 186400 105620 186600 105880
rect 186900 105620 187100 105880
rect 187400 105620 187600 105880
rect 187900 105620 188100 105880
rect 188400 105620 188600 105880
rect 188900 105620 189100 105880
rect 189400 105620 189600 105880
rect 189900 105620 190100 105880
rect 190400 105620 190600 105880
rect 190900 105620 191100 105880
rect 191400 105620 191600 105880
rect 191900 105620 192100 105880
rect 192400 105620 192600 105880
rect 192900 105620 193100 105880
rect 193400 105620 193600 105880
rect 193900 105620 194100 105880
rect 194400 105620 194600 105880
rect 194900 105620 195100 105880
rect 195400 105620 195600 105880
rect 195900 105620 196100 105880
rect 196400 105620 196600 105880
rect 196900 105620 197100 105880
rect 197400 105620 197600 105880
rect 197900 105620 198100 105880
rect 198400 105620 198600 105880
rect 198900 105620 199100 105880
rect 199400 105620 199600 105880
rect 199900 105620 200100 105880
rect 200400 105620 200600 105880
rect 200900 105620 201100 105880
rect 201400 105620 201600 105880
rect 201900 105620 202100 105880
rect 202400 105620 202600 105880
rect 202900 105620 203100 105880
rect 203400 105620 203600 105880
rect 203900 105620 204100 105880
rect 204400 105620 204600 105880
rect 204900 105620 205100 105880
rect 205400 105620 205600 105880
rect 205900 105620 206100 105880
rect 206400 105620 206600 105880
rect 206900 105620 207100 105880
rect 207400 105620 207600 105880
rect 207900 105620 208100 105880
rect 208400 105620 208600 105880
rect 208900 105620 209100 105880
rect 209400 105620 209600 105880
rect 209900 105620 210100 105880
rect 210400 105620 210600 105880
rect 210900 105620 211100 105880
rect 211400 105620 211600 105880
rect 211900 105620 212100 105880
rect 212400 105620 212600 105880
rect 212900 105620 213100 105880
rect 213400 105620 213600 105880
rect 213900 105620 214100 105880
rect 214400 105620 214600 105880
rect 214900 105620 215100 105880
rect 215400 105620 215600 105880
rect 215900 105620 216100 105880
rect 216400 105620 216600 105880
rect 216900 105620 217100 105880
rect 217400 105620 217600 105880
rect 217900 105620 218100 105880
rect 218400 105620 218600 105880
rect 218900 105620 219100 105880
rect 219400 105620 219600 105880
rect 219900 105620 220100 105880
rect 220400 105620 220600 105880
rect 220900 105620 221100 105880
rect 221400 105620 221600 105880
rect 221900 105620 222100 105880
rect 222400 105620 222600 105880
rect 222900 105620 223100 105880
rect 223400 105620 223600 105880
rect 223900 105620 224100 105880
rect 224400 105620 224600 105880
rect 224900 105620 225100 105880
rect 225400 105620 225600 105880
rect 225900 105620 226100 105880
rect 226400 105620 226600 105880
rect 226900 105620 227100 105880
rect 227400 105620 227600 105880
rect 227900 105620 228100 105880
rect 228400 105620 228600 105880
rect 228900 105620 229100 105880
rect 229400 105620 229600 105880
rect 229900 105620 230100 105880
rect 230400 105620 230600 105880
rect 230900 105620 231100 105880
rect 231400 105620 231600 105880
rect 231900 105620 232000 105880
rect 178000 105600 178120 105620
rect 178380 105600 178620 105620
rect 178880 105600 179120 105620
rect 179380 105600 179620 105620
rect 179880 105600 180120 105620
rect 180380 105600 180620 105620
rect 180880 105600 181120 105620
rect 181380 105600 181620 105620
rect 181880 105600 182120 105620
rect 182380 105600 182620 105620
rect 182880 105600 183120 105620
rect 183380 105600 183620 105620
rect 183880 105600 184120 105620
rect 184380 105600 184620 105620
rect 184880 105600 185120 105620
rect 185380 105600 185620 105620
rect 185880 105600 186120 105620
rect 186380 105600 186620 105620
rect 186880 105600 187120 105620
rect 187380 105600 187620 105620
rect 187880 105600 188120 105620
rect 188380 105600 188620 105620
rect 188880 105600 189120 105620
rect 189380 105600 189620 105620
rect 189880 105600 190120 105620
rect 190380 105600 190620 105620
rect 190880 105600 191120 105620
rect 191380 105600 191620 105620
rect 191880 105600 192120 105620
rect 192380 105600 192620 105620
rect 192880 105600 193120 105620
rect 193380 105600 193620 105620
rect 193880 105600 194120 105620
rect 194380 105600 194620 105620
rect 194880 105600 195120 105620
rect 195380 105600 195620 105620
rect 195880 105600 196120 105620
rect 196380 105600 196620 105620
rect 196880 105600 197120 105620
rect 197380 105600 197620 105620
rect 197880 105600 198120 105620
rect 198380 105600 198620 105620
rect 198880 105600 199120 105620
rect 199380 105600 199620 105620
rect 199880 105600 200120 105620
rect 200380 105600 200620 105620
rect 200880 105600 201120 105620
rect 201380 105600 201620 105620
rect 201880 105600 202120 105620
rect 202380 105600 202620 105620
rect 202880 105600 203120 105620
rect 203380 105600 203620 105620
rect 203880 105600 204120 105620
rect 204380 105600 204620 105620
rect 204880 105600 205120 105620
rect 205380 105600 205620 105620
rect 205880 105600 206120 105620
rect 206380 105600 206620 105620
rect 206880 105600 207120 105620
rect 207380 105600 207620 105620
rect 207880 105600 208120 105620
rect 208380 105600 208620 105620
rect 208880 105600 209120 105620
rect 209380 105600 209620 105620
rect 209880 105600 210120 105620
rect 210380 105600 210620 105620
rect 210880 105600 211120 105620
rect 211380 105600 211620 105620
rect 211880 105600 212120 105620
rect 212380 105600 212620 105620
rect 212880 105600 213120 105620
rect 213380 105600 213620 105620
rect 213880 105600 214120 105620
rect 214380 105600 214620 105620
rect 214880 105600 215120 105620
rect 215380 105600 215620 105620
rect 215880 105600 216120 105620
rect 216380 105600 216620 105620
rect 216880 105600 217120 105620
rect 217380 105600 217620 105620
rect 217880 105600 218120 105620
rect 218380 105600 218620 105620
rect 218880 105600 219120 105620
rect 219380 105600 219620 105620
rect 219880 105600 220120 105620
rect 220380 105600 220620 105620
rect 220880 105600 221120 105620
rect 221380 105600 221620 105620
rect 221880 105600 222120 105620
rect 222380 105600 222620 105620
rect 222880 105600 223120 105620
rect 223380 105600 223620 105620
rect 223880 105600 224120 105620
rect 224380 105600 224620 105620
rect 224880 105600 225120 105620
rect 225380 105600 225620 105620
rect 225880 105600 226120 105620
rect 226380 105600 226620 105620
rect 226880 105600 227120 105620
rect 227380 105600 227620 105620
rect 227880 105600 228120 105620
rect 228380 105600 228620 105620
rect 228880 105600 229120 105620
rect 229380 105600 229620 105620
rect 229880 105600 230120 105620
rect 230380 105600 230620 105620
rect 230880 105600 231120 105620
rect 231380 105600 231620 105620
rect 231880 105600 232000 105620
rect 178000 105400 232000 105600
rect 178000 105380 178120 105400
rect 178380 105380 178620 105400
rect 178880 105380 179120 105400
rect 179380 105380 179620 105400
rect 179880 105380 180120 105400
rect 180380 105380 180620 105400
rect 180880 105380 181120 105400
rect 181380 105380 181620 105400
rect 181880 105380 182120 105400
rect 182380 105380 182620 105400
rect 182880 105380 183120 105400
rect 183380 105380 183620 105400
rect 183880 105380 184120 105400
rect 184380 105380 184620 105400
rect 184880 105380 185120 105400
rect 185380 105380 185620 105400
rect 185880 105380 186120 105400
rect 186380 105380 186620 105400
rect 186880 105380 187120 105400
rect 187380 105380 187620 105400
rect 187880 105380 188120 105400
rect 188380 105380 188620 105400
rect 188880 105380 189120 105400
rect 189380 105380 189620 105400
rect 189880 105380 190120 105400
rect 190380 105380 190620 105400
rect 190880 105380 191120 105400
rect 191380 105380 191620 105400
rect 191880 105380 192120 105400
rect 192380 105380 192620 105400
rect 192880 105380 193120 105400
rect 193380 105380 193620 105400
rect 193880 105380 194120 105400
rect 194380 105380 194620 105400
rect 194880 105380 195120 105400
rect 195380 105380 195620 105400
rect 195880 105380 196120 105400
rect 196380 105380 196620 105400
rect 196880 105380 197120 105400
rect 197380 105380 197620 105400
rect 197880 105380 198120 105400
rect 198380 105380 198620 105400
rect 198880 105380 199120 105400
rect 199380 105380 199620 105400
rect 199880 105380 200120 105400
rect 200380 105380 200620 105400
rect 200880 105380 201120 105400
rect 201380 105380 201620 105400
rect 201880 105380 202120 105400
rect 202380 105380 202620 105400
rect 202880 105380 203120 105400
rect 203380 105380 203620 105400
rect 203880 105380 204120 105400
rect 204380 105380 204620 105400
rect 204880 105380 205120 105400
rect 205380 105380 205620 105400
rect 205880 105380 206120 105400
rect 206380 105380 206620 105400
rect 206880 105380 207120 105400
rect 207380 105380 207620 105400
rect 207880 105380 208120 105400
rect 208380 105380 208620 105400
rect 208880 105380 209120 105400
rect 209380 105380 209620 105400
rect 209880 105380 210120 105400
rect 210380 105380 210620 105400
rect 210880 105380 211120 105400
rect 211380 105380 211620 105400
rect 211880 105380 212120 105400
rect 212380 105380 212620 105400
rect 212880 105380 213120 105400
rect 213380 105380 213620 105400
rect 213880 105380 214120 105400
rect 214380 105380 214620 105400
rect 214880 105380 215120 105400
rect 215380 105380 215620 105400
rect 215880 105380 216120 105400
rect 216380 105380 216620 105400
rect 216880 105380 217120 105400
rect 217380 105380 217620 105400
rect 217880 105380 218120 105400
rect 218380 105380 218620 105400
rect 218880 105380 219120 105400
rect 219380 105380 219620 105400
rect 219880 105380 220120 105400
rect 220380 105380 220620 105400
rect 220880 105380 221120 105400
rect 221380 105380 221620 105400
rect 221880 105380 222120 105400
rect 222380 105380 222620 105400
rect 222880 105380 223120 105400
rect 223380 105380 223620 105400
rect 223880 105380 224120 105400
rect 224380 105380 224620 105400
rect 224880 105380 225120 105400
rect 225380 105380 225620 105400
rect 225880 105380 226120 105400
rect 226380 105380 226620 105400
rect 226880 105380 227120 105400
rect 227380 105380 227620 105400
rect 227880 105380 228120 105400
rect 228380 105380 228620 105400
rect 228880 105380 229120 105400
rect 229380 105380 229620 105400
rect 229880 105380 230120 105400
rect 230380 105380 230620 105400
rect 230880 105380 231120 105400
rect 231380 105380 231620 105400
rect 231880 105380 232000 105400
rect 178000 105120 178100 105380
rect 178400 105120 178600 105380
rect 178900 105120 179100 105380
rect 179400 105120 179600 105380
rect 179900 105120 180100 105380
rect 180400 105120 180600 105380
rect 180900 105120 181100 105380
rect 181400 105120 181600 105380
rect 181900 105120 182100 105380
rect 182400 105120 182600 105380
rect 182900 105120 183100 105380
rect 183400 105120 183600 105380
rect 183900 105120 184100 105380
rect 184400 105120 184600 105380
rect 184900 105120 185100 105380
rect 185400 105120 185600 105380
rect 185900 105120 186100 105380
rect 186400 105120 186600 105380
rect 186900 105120 187100 105380
rect 187400 105120 187600 105380
rect 187900 105120 188100 105380
rect 188400 105120 188600 105380
rect 188900 105120 189100 105380
rect 189400 105120 189600 105380
rect 189900 105120 190100 105380
rect 190400 105120 190600 105380
rect 190900 105120 191100 105380
rect 191400 105120 191600 105380
rect 191900 105120 192100 105380
rect 192400 105120 192600 105380
rect 192900 105120 193100 105380
rect 193400 105120 193600 105380
rect 193900 105120 194100 105380
rect 194400 105120 194600 105380
rect 194900 105120 195100 105380
rect 195400 105120 195600 105380
rect 195900 105120 196100 105380
rect 196400 105120 196600 105380
rect 196900 105120 197100 105380
rect 197400 105120 197600 105380
rect 197900 105120 198100 105380
rect 198400 105120 198600 105380
rect 198900 105120 199100 105380
rect 199400 105120 199600 105380
rect 199900 105120 200100 105380
rect 200400 105120 200600 105380
rect 200900 105120 201100 105380
rect 201400 105120 201600 105380
rect 201900 105120 202100 105380
rect 202400 105120 202600 105380
rect 202900 105120 203100 105380
rect 203400 105120 203600 105380
rect 203900 105120 204100 105380
rect 204400 105120 204600 105380
rect 204900 105120 205100 105380
rect 205400 105120 205600 105380
rect 205900 105120 206100 105380
rect 206400 105120 206600 105380
rect 206900 105120 207100 105380
rect 207400 105120 207600 105380
rect 207900 105120 208100 105380
rect 208400 105120 208600 105380
rect 208900 105120 209100 105380
rect 209400 105120 209600 105380
rect 209900 105120 210100 105380
rect 210400 105120 210600 105380
rect 210900 105120 211100 105380
rect 211400 105120 211600 105380
rect 211900 105120 212100 105380
rect 212400 105120 212600 105380
rect 212900 105120 213100 105380
rect 213400 105120 213600 105380
rect 213900 105120 214100 105380
rect 214400 105120 214600 105380
rect 214900 105120 215100 105380
rect 215400 105120 215600 105380
rect 215900 105120 216100 105380
rect 216400 105120 216600 105380
rect 216900 105120 217100 105380
rect 217400 105120 217600 105380
rect 217900 105120 218100 105380
rect 218400 105120 218600 105380
rect 218900 105120 219100 105380
rect 219400 105120 219600 105380
rect 219900 105120 220100 105380
rect 220400 105120 220600 105380
rect 220900 105120 221100 105380
rect 221400 105120 221600 105380
rect 221900 105120 222100 105380
rect 222400 105120 222600 105380
rect 222900 105120 223100 105380
rect 223400 105120 223600 105380
rect 223900 105120 224100 105380
rect 224400 105120 224600 105380
rect 224900 105120 225100 105380
rect 225400 105120 225600 105380
rect 225900 105120 226100 105380
rect 226400 105120 226600 105380
rect 226900 105120 227100 105380
rect 227400 105120 227600 105380
rect 227900 105120 228100 105380
rect 228400 105120 228600 105380
rect 228900 105120 229100 105380
rect 229400 105120 229600 105380
rect 229900 105120 230100 105380
rect 230400 105120 230600 105380
rect 230900 105120 231100 105380
rect 231400 105120 231600 105380
rect 231900 105120 232000 105380
rect 178000 105100 178120 105120
rect 178380 105100 178620 105120
rect 178880 105100 179120 105120
rect 179380 105100 179620 105120
rect 179880 105100 180120 105120
rect 180380 105100 180620 105120
rect 180880 105100 181120 105120
rect 181380 105100 181620 105120
rect 181880 105100 182120 105120
rect 182380 105100 182620 105120
rect 182880 105100 183120 105120
rect 183380 105100 183620 105120
rect 183880 105100 184120 105120
rect 184380 105100 184620 105120
rect 184880 105100 185120 105120
rect 185380 105100 185620 105120
rect 185880 105100 186120 105120
rect 186380 105100 186620 105120
rect 186880 105100 187120 105120
rect 187380 105100 187620 105120
rect 187880 105100 188120 105120
rect 188380 105100 188620 105120
rect 188880 105100 189120 105120
rect 189380 105100 189620 105120
rect 189880 105100 190120 105120
rect 190380 105100 190620 105120
rect 190880 105100 191120 105120
rect 191380 105100 191620 105120
rect 191880 105100 192120 105120
rect 192380 105100 192620 105120
rect 192880 105100 193120 105120
rect 193380 105100 193620 105120
rect 193880 105100 194120 105120
rect 194380 105100 194620 105120
rect 194880 105100 195120 105120
rect 195380 105100 195620 105120
rect 195880 105100 196120 105120
rect 196380 105100 196620 105120
rect 196880 105100 197120 105120
rect 197380 105100 197620 105120
rect 197880 105100 198120 105120
rect 198380 105100 198620 105120
rect 198880 105100 199120 105120
rect 199380 105100 199620 105120
rect 199880 105100 200120 105120
rect 200380 105100 200620 105120
rect 200880 105100 201120 105120
rect 201380 105100 201620 105120
rect 201880 105100 202120 105120
rect 202380 105100 202620 105120
rect 202880 105100 203120 105120
rect 203380 105100 203620 105120
rect 203880 105100 204120 105120
rect 204380 105100 204620 105120
rect 204880 105100 205120 105120
rect 205380 105100 205620 105120
rect 205880 105100 206120 105120
rect 206380 105100 206620 105120
rect 206880 105100 207120 105120
rect 207380 105100 207620 105120
rect 207880 105100 208120 105120
rect 208380 105100 208620 105120
rect 208880 105100 209120 105120
rect 209380 105100 209620 105120
rect 209880 105100 210120 105120
rect 210380 105100 210620 105120
rect 210880 105100 211120 105120
rect 211380 105100 211620 105120
rect 211880 105100 212120 105120
rect 212380 105100 212620 105120
rect 212880 105100 213120 105120
rect 213380 105100 213620 105120
rect 213880 105100 214120 105120
rect 214380 105100 214620 105120
rect 214880 105100 215120 105120
rect 215380 105100 215620 105120
rect 215880 105100 216120 105120
rect 216380 105100 216620 105120
rect 216880 105100 217120 105120
rect 217380 105100 217620 105120
rect 217880 105100 218120 105120
rect 218380 105100 218620 105120
rect 218880 105100 219120 105120
rect 219380 105100 219620 105120
rect 219880 105100 220120 105120
rect 220380 105100 220620 105120
rect 220880 105100 221120 105120
rect 221380 105100 221620 105120
rect 221880 105100 222120 105120
rect 222380 105100 222620 105120
rect 222880 105100 223120 105120
rect 223380 105100 223620 105120
rect 223880 105100 224120 105120
rect 224380 105100 224620 105120
rect 224880 105100 225120 105120
rect 225380 105100 225620 105120
rect 225880 105100 226120 105120
rect 226380 105100 226620 105120
rect 226880 105100 227120 105120
rect 227380 105100 227620 105120
rect 227880 105100 228120 105120
rect 228380 105100 228620 105120
rect 228880 105100 229120 105120
rect 229380 105100 229620 105120
rect 229880 105100 230120 105120
rect 230380 105100 230620 105120
rect 230880 105100 231120 105120
rect 231380 105100 231620 105120
rect 231880 105100 232000 105120
rect 178000 104900 232000 105100
rect 178000 104880 178120 104900
rect 178380 104880 178620 104900
rect 178880 104880 179120 104900
rect 179380 104880 179620 104900
rect 179880 104880 180120 104900
rect 180380 104880 180620 104900
rect 180880 104880 181120 104900
rect 181380 104880 181620 104900
rect 181880 104880 182120 104900
rect 182380 104880 182620 104900
rect 182880 104880 183120 104900
rect 183380 104880 183620 104900
rect 183880 104880 184120 104900
rect 184380 104880 184620 104900
rect 184880 104880 185120 104900
rect 185380 104880 185620 104900
rect 185880 104880 186120 104900
rect 186380 104880 186620 104900
rect 186880 104880 187120 104900
rect 187380 104880 187620 104900
rect 187880 104880 188120 104900
rect 188380 104880 188620 104900
rect 188880 104880 189120 104900
rect 189380 104880 189620 104900
rect 189880 104880 190120 104900
rect 190380 104880 190620 104900
rect 190880 104880 191120 104900
rect 191380 104880 191620 104900
rect 191880 104880 192120 104900
rect 192380 104880 192620 104900
rect 192880 104880 193120 104900
rect 193380 104880 193620 104900
rect 193880 104880 194120 104900
rect 194380 104880 194620 104900
rect 194880 104880 195120 104900
rect 195380 104880 195620 104900
rect 195880 104880 196120 104900
rect 196380 104880 196620 104900
rect 196880 104880 197120 104900
rect 197380 104880 197620 104900
rect 197880 104880 198120 104900
rect 198380 104880 198620 104900
rect 198880 104880 199120 104900
rect 199380 104880 199620 104900
rect 199880 104880 200120 104900
rect 200380 104880 200620 104900
rect 200880 104880 201120 104900
rect 201380 104880 201620 104900
rect 201880 104880 202120 104900
rect 202380 104880 202620 104900
rect 202880 104880 203120 104900
rect 203380 104880 203620 104900
rect 203880 104880 204120 104900
rect 204380 104880 204620 104900
rect 204880 104880 205120 104900
rect 205380 104880 205620 104900
rect 205880 104880 206120 104900
rect 206380 104880 206620 104900
rect 206880 104880 207120 104900
rect 207380 104880 207620 104900
rect 207880 104880 208120 104900
rect 208380 104880 208620 104900
rect 208880 104880 209120 104900
rect 209380 104880 209620 104900
rect 209880 104880 210120 104900
rect 210380 104880 210620 104900
rect 210880 104880 211120 104900
rect 211380 104880 211620 104900
rect 211880 104880 212120 104900
rect 212380 104880 212620 104900
rect 212880 104880 213120 104900
rect 213380 104880 213620 104900
rect 213880 104880 214120 104900
rect 214380 104880 214620 104900
rect 214880 104880 215120 104900
rect 215380 104880 215620 104900
rect 215880 104880 216120 104900
rect 216380 104880 216620 104900
rect 216880 104880 217120 104900
rect 217380 104880 217620 104900
rect 217880 104880 218120 104900
rect 218380 104880 218620 104900
rect 218880 104880 219120 104900
rect 219380 104880 219620 104900
rect 219880 104880 220120 104900
rect 220380 104880 220620 104900
rect 220880 104880 221120 104900
rect 221380 104880 221620 104900
rect 221880 104880 222120 104900
rect 222380 104880 222620 104900
rect 222880 104880 223120 104900
rect 223380 104880 223620 104900
rect 223880 104880 224120 104900
rect 224380 104880 224620 104900
rect 224880 104880 225120 104900
rect 225380 104880 225620 104900
rect 225880 104880 226120 104900
rect 226380 104880 226620 104900
rect 226880 104880 227120 104900
rect 227380 104880 227620 104900
rect 227880 104880 228120 104900
rect 228380 104880 228620 104900
rect 228880 104880 229120 104900
rect 229380 104880 229620 104900
rect 229880 104880 230120 104900
rect 230380 104880 230620 104900
rect 230880 104880 231120 104900
rect 231380 104880 231620 104900
rect 231880 104880 232000 104900
rect 178000 104620 178100 104880
rect 178400 104620 178600 104880
rect 178900 104620 179100 104880
rect 179400 104620 179600 104880
rect 179900 104620 180100 104880
rect 180400 104620 180600 104880
rect 180900 104620 181100 104880
rect 181400 104620 181600 104880
rect 181900 104620 182100 104880
rect 182400 104620 182600 104880
rect 182900 104620 183100 104880
rect 183400 104620 183600 104880
rect 183900 104620 184100 104880
rect 184400 104620 184600 104880
rect 184900 104620 185100 104880
rect 185400 104620 185600 104880
rect 185900 104620 186100 104880
rect 186400 104620 186600 104880
rect 186900 104620 187100 104880
rect 187400 104620 187600 104880
rect 187900 104620 188100 104880
rect 188400 104620 188600 104880
rect 188900 104620 189100 104880
rect 189400 104620 189600 104880
rect 189900 104620 190100 104880
rect 190400 104620 190600 104880
rect 190900 104620 191100 104880
rect 191400 104620 191600 104880
rect 191900 104620 192100 104880
rect 192400 104620 192600 104880
rect 192900 104620 193100 104880
rect 193400 104620 193600 104880
rect 193900 104620 194100 104880
rect 194400 104620 194600 104880
rect 194900 104620 195100 104880
rect 195400 104620 195600 104880
rect 195900 104620 196100 104880
rect 196400 104620 196600 104880
rect 196900 104620 197100 104880
rect 197400 104620 197600 104880
rect 197900 104620 198100 104880
rect 198400 104620 198600 104880
rect 198900 104620 199100 104880
rect 199400 104620 199600 104880
rect 199900 104620 200100 104880
rect 200400 104620 200600 104880
rect 200900 104620 201100 104880
rect 201400 104620 201600 104880
rect 201900 104620 202100 104880
rect 202400 104620 202600 104880
rect 202900 104620 203100 104880
rect 203400 104620 203600 104880
rect 203900 104620 204100 104880
rect 204400 104620 204600 104880
rect 204900 104620 205100 104880
rect 205400 104620 205600 104880
rect 205900 104620 206100 104880
rect 206400 104620 206600 104880
rect 206900 104620 207100 104880
rect 207400 104620 207600 104880
rect 207900 104620 208100 104880
rect 208400 104620 208600 104880
rect 208900 104620 209100 104880
rect 209400 104620 209600 104880
rect 209900 104620 210100 104880
rect 210400 104620 210600 104880
rect 210900 104620 211100 104880
rect 211400 104620 211600 104880
rect 211900 104620 212100 104880
rect 212400 104620 212600 104880
rect 212900 104620 213100 104880
rect 213400 104620 213600 104880
rect 213900 104620 214100 104880
rect 214400 104620 214600 104880
rect 214900 104620 215100 104880
rect 215400 104620 215600 104880
rect 215900 104620 216100 104880
rect 216400 104620 216600 104880
rect 216900 104620 217100 104880
rect 217400 104620 217600 104880
rect 217900 104620 218100 104880
rect 218400 104620 218600 104880
rect 218900 104620 219100 104880
rect 219400 104620 219600 104880
rect 219900 104620 220100 104880
rect 220400 104620 220600 104880
rect 220900 104620 221100 104880
rect 221400 104620 221600 104880
rect 221900 104620 222100 104880
rect 222400 104620 222600 104880
rect 222900 104620 223100 104880
rect 223400 104620 223600 104880
rect 223900 104620 224100 104880
rect 224400 104620 224600 104880
rect 224900 104620 225100 104880
rect 225400 104620 225600 104880
rect 225900 104620 226100 104880
rect 226400 104620 226600 104880
rect 226900 104620 227100 104880
rect 227400 104620 227600 104880
rect 227900 104620 228100 104880
rect 228400 104620 228600 104880
rect 228900 104620 229100 104880
rect 229400 104620 229600 104880
rect 229900 104620 230100 104880
rect 230400 104620 230600 104880
rect 230900 104620 231100 104880
rect 231400 104620 231600 104880
rect 231900 104620 232000 104880
rect 178000 104600 178120 104620
rect 178380 104600 178620 104620
rect 178880 104600 179120 104620
rect 179380 104600 179620 104620
rect 179880 104600 180120 104620
rect 180380 104600 180620 104620
rect 180880 104600 181120 104620
rect 181380 104600 181620 104620
rect 181880 104600 182120 104620
rect 182380 104600 182620 104620
rect 182880 104600 183120 104620
rect 183380 104600 183620 104620
rect 183880 104600 184120 104620
rect 184380 104600 184620 104620
rect 184880 104600 185120 104620
rect 185380 104600 185620 104620
rect 185880 104600 186120 104620
rect 186380 104600 186620 104620
rect 186880 104600 187120 104620
rect 187380 104600 187620 104620
rect 187880 104600 188120 104620
rect 188380 104600 188620 104620
rect 188880 104600 189120 104620
rect 189380 104600 189620 104620
rect 189880 104600 190120 104620
rect 190380 104600 190620 104620
rect 190880 104600 191120 104620
rect 191380 104600 191620 104620
rect 191880 104600 192120 104620
rect 192380 104600 192620 104620
rect 192880 104600 193120 104620
rect 193380 104600 193620 104620
rect 193880 104600 194120 104620
rect 194380 104600 194620 104620
rect 194880 104600 195120 104620
rect 195380 104600 195620 104620
rect 195880 104600 196120 104620
rect 196380 104600 196620 104620
rect 196880 104600 197120 104620
rect 197380 104600 197620 104620
rect 197880 104600 198120 104620
rect 198380 104600 198620 104620
rect 198880 104600 199120 104620
rect 199380 104600 199620 104620
rect 199880 104600 200120 104620
rect 200380 104600 200620 104620
rect 200880 104600 201120 104620
rect 201380 104600 201620 104620
rect 201880 104600 202120 104620
rect 202380 104600 202620 104620
rect 202880 104600 203120 104620
rect 203380 104600 203620 104620
rect 203880 104600 204120 104620
rect 204380 104600 204620 104620
rect 204880 104600 205120 104620
rect 205380 104600 205620 104620
rect 205880 104600 206120 104620
rect 206380 104600 206620 104620
rect 206880 104600 207120 104620
rect 207380 104600 207620 104620
rect 207880 104600 208120 104620
rect 208380 104600 208620 104620
rect 208880 104600 209120 104620
rect 209380 104600 209620 104620
rect 209880 104600 210120 104620
rect 210380 104600 210620 104620
rect 210880 104600 211120 104620
rect 211380 104600 211620 104620
rect 211880 104600 212120 104620
rect 212380 104600 212620 104620
rect 212880 104600 213120 104620
rect 213380 104600 213620 104620
rect 213880 104600 214120 104620
rect 214380 104600 214620 104620
rect 214880 104600 215120 104620
rect 215380 104600 215620 104620
rect 215880 104600 216120 104620
rect 216380 104600 216620 104620
rect 216880 104600 217120 104620
rect 217380 104600 217620 104620
rect 217880 104600 218120 104620
rect 218380 104600 218620 104620
rect 218880 104600 219120 104620
rect 219380 104600 219620 104620
rect 219880 104600 220120 104620
rect 220380 104600 220620 104620
rect 220880 104600 221120 104620
rect 221380 104600 221620 104620
rect 221880 104600 222120 104620
rect 222380 104600 222620 104620
rect 222880 104600 223120 104620
rect 223380 104600 223620 104620
rect 223880 104600 224120 104620
rect 224380 104600 224620 104620
rect 224880 104600 225120 104620
rect 225380 104600 225620 104620
rect 225880 104600 226120 104620
rect 226380 104600 226620 104620
rect 226880 104600 227120 104620
rect 227380 104600 227620 104620
rect 227880 104600 228120 104620
rect 228380 104600 228620 104620
rect 228880 104600 229120 104620
rect 229380 104600 229620 104620
rect 229880 104600 230120 104620
rect 230380 104600 230620 104620
rect 230880 104600 231120 104620
rect 231380 104600 231620 104620
rect 231880 104600 232000 104620
rect 178000 104400 232000 104600
rect 178000 104380 178120 104400
rect 178380 104380 178620 104400
rect 178880 104380 179120 104400
rect 179380 104380 179620 104400
rect 179880 104380 180120 104400
rect 180380 104380 180620 104400
rect 180880 104380 181120 104400
rect 181380 104380 181620 104400
rect 181880 104380 182120 104400
rect 182380 104380 182620 104400
rect 182880 104380 183120 104400
rect 183380 104380 183620 104400
rect 183880 104380 184120 104400
rect 184380 104380 184620 104400
rect 184880 104380 185120 104400
rect 185380 104380 185620 104400
rect 185880 104380 186120 104400
rect 186380 104380 186620 104400
rect 186880 104380 187120 104400
rect 187380 104380 187620 104400
rect 187880 104380 188120 104400
rect 188380 104380 188620 104400
rect 188880 104380 189120 104400
rect 189380 104380 189620 104400
rect 189880 104380 190120 104400
rect 190380 104380 190620 104400
rect 190880 104380 191120 104400
rect 191380 104380 191620 104400
rect 191880 104380 192120 104400
rect 192380 104380 192620 104400
rect 192880 104380 193120 104400
rect 193380 104380 193620 104400
rect 193880 104380 194120 104400
rect 194380 104380 194620 104400
rect 194880 104380 195120 104400
rect 195380 104380 195620 104400
rect 195880 104380 196120 104400
rect 196380 104380 196620 104400
rect 196880 104380 197120 104400
rect 197380 104380 197620 104400
rect 197880 104380 198120 104400
rect 198380 104380 198620 104400
rect 198880 104380 199120 104400
rect 199380 104380 199620 104400
rect 199880 104380 200120 104400
rect 200380 104380 200620 104400
rect 200880 104380 201120 104400
rect 201380 104380 201620 104400
rect 201880 104380 202120 104400
rect 202380 104380 202620 104400
rect 202880 104380 203120 104400
rect 203380 104380 203620 104400
rect 203880 104380 204120 104400
rect 204380 104380 204620 104400
rect 204880 104380 205120 104400
rect 205380 104380 205620 104400
rect 205880 104380 206120 104400
rect 206380 104380 206620 104400
rect 206880 104380 207120 104400
rect 207380 104380 207620 104400
rect 207880 104380 208120 104400
rect 208380 104380 208620 104400
rect 208880 104380 209120 104400
rect 209380 104380 209620 104400
rect 209880 104380 210120 104400
rect 210380 104380 210620 104400
rect 210880 104380 211120 104400
rect 211380 104380 211620 104400
rect 211880 104380 212120 104400
rect 212380 104380 212620 104400
rect 212880 104380 213120 104400
rect 213380 104380 213620 104400
rect 213880 104380 214120 104400
rect 214380 104380 214620 104400
rect 214880 104380 215120 104400
rect 215380 104380 215620 104400
rect 215880 104380 216120 104400
rect 216380 104380 216620 104400
rect 216880 104380 217120 104400
rect 217380 104380 217620 104400
rect 217880 104380 218120 104400
rect 218380 104380 218620 104400
rect 218880 104380 219120 104400
rect 219380 104380 219620 104400
rect 219880 104380 220120 104400
rect 220380 104380 220620 104400
rect 220880 104380 221120 104400
rect 221380 104380 221620 104400
rect 221880 104380 222120 104400
rect 222380 104380 222620 104400
rect 222880 104380 223120 104400
rect 223380 104380 223620 104400
rect 223880 104380 224120 104400
rect 224380 104380 224620 104400
rect 224880 104380 225120 104400
rect 225380 104380 225620 104400
rect 225880 104380 226120 104400
rect 226380 104380 226620 104400
rect 226880 104380 227120 104400
rect 227380 104380 227620 104400
rect 227880 104380 228120 104400
rect 228380 104380 228620 104400
rect 228880 104380 229120 104400
rect 229380 104380 229620 104400
rect 229880 104380 230120 104400
rect 230380 104380 230620 104400
rect 230880 104380 231120 104400
rect 231380 104380 231620 104400
rect 231880 104380 232000 104400
rect 178000 104120 178100 104380
rect 178400 104120 178600 104380
rect 178900 104120 179100 104380
rect 179400 104120 179600 104380
rect 179900 104120 180100 104380
rect 180400 104120 180600 104380
rect 180900 104120 181100 104380
rect 181400 104120 181600 104380
rect 181900 104120 182100 104380
rect 182400 104120 182600 104380
rect 182900 104120 183100 104380
rect 183400 104120 183600 104380
rect 183900 104120 184100 104380
rect 184400 104120 184600 104380
rect 184900 104120 185100 104380
rect 185400 104120 185600 104380
rect 185900 104120 186100 104380
rect 186400 104120 186600 104380
rect 186900 104120 187100 104380
rect 187400 104120 187600 104380
rect 187900 104120 188100 104380
rect 188400 104120 188600 104380
rect 188900 104120 189100 104380
rect 189400 104120 189600 104380
rect 189900 104120 190100 104380
rect 190400 104120 190600 104380
rect 190900 104120 191100 104380
rect 191400 104120 191600 104380
rect 191900 104120 192100 104380
rect 192400 104120 192600 104380
rect 192900 104120 193100 104380
rect 193400 104120 193600 104380
rect 193900 104120 194100 104380
rect 194400 104120 194600 104380
rect 194900 104120 195100 104380
rect 195400 104120 195600 104380
rect 195900 104120 196100 104380
rect 196400 104120 196600 104380
rect 196900 104120 197100 104380
rect 197400 104120 197600 104380
rect 197900 104120 198100 104380
rect 198400 104120 198600 104380
rect 198900 104120 199100 104380
rect 199400 104120 199600 104380
rect 199900 104120 200100 104380
rect 200400 104120 200600 104380
rect 200900 104120 201100 104380
rect 201400 104120 201600 104380
rect 201900 104120 202100 104380
rect 202400 104120 202600 104380
rect 202900 104120 203100 104380
rect 203400 104120 203600 104380
rect 203900 104120 204100 104380
rect 204400 104120 204600 104380
rect 204900 104120 205100 104380
rect 205400 104120 205600 104380
rect 205900 104120 206100 104380
rect 206400 104120 206600 104380
rect 206900 104120 207100 104380
rect 207400 104120 207600 104380
rect 207900 104120 208100 104380
rect 208400 104120 208600 104380
rect 208900 104120 209100 104380
rect 209400 104120 209600 104380
rect 209900 104120 210100 104380
rect 210400 104120 210600 104380
rect 210900 104120 211100 104380
rect 211400 104120 211600 104380
rect 211900 104120 212100 104380
rect 212400 104120 212600 104380
rect 212900 104120 213100 104380
rect 213400 104120 213600 104380
rect 213900 104120 214100 104380
rect 214400 104120 214600 104380
rect 214900 104120 215100 104380
rect 215400 104120 215600 104380
rect 215900 104120 216100 104380
rect 216400 104120 216600 104380
rect 216900 104120 217100 104380
rect 217400 104120 217600 104380
rect 217900 104120 218100 104380
rect 218400 104120 218600 104380
rect 218900 104120 219100 104380
rect 219400 104120 219600 104380
rect 219900 104120 220100 104380
rect 220400 104120 220600 104380
rect 220900 104120 221100 104380
rect 221400 104120 221600 104380
rect 221900 104120 222100 104380
rect 222400 104120 222600 104380
rect 222900 104120 223100 104380
rect 223400 104120 223600 104380
rect 223900 104120 224100 104380
rect 224400 104120 224600 104380
rect 224900 104120 225100 104380
rect 225400 104120 225600 104380
rect 225900 104120 226100 104380
rect 226400 104120 226600 104380
rect 226900 104120 227100 104380
rect 227400 104120 227600 104380
rect 227900 104120 228100 104380
rect 228400 104120 228600 104380
rect 228900 104120 229100 104380
rect 229400 104120 229600 104380
rect 229900 104120 230100 104380
rect 230400 104120 230600 104380
rect 230900 104120 231100 104380
rect 231400 104120 231600 104380
rect 231900 104120 232000 104380
rect 178000 104100 178120 104120
rect 178380 104100 178620 104120
rect 178880 104100 179120 104120
rect 179380 104100 179620 104120
rect 179880 104100 180120 104120
rect 180380 104100 180620 104120
rect 180880 104100 181120 104120
rect 181380 104100 181620 104120
rect 181880 104100 182120 104120
rect 182380 104100 182620 104120
rect 182880 104100 183120 104120
rect 183380 104100 183620 104120
rect 183880 104100 184120 104120
rect 184380 104100 184620 104120
rect 184880 104100 185120 104120
rect 185380 104100 185620 104120
rect 185880 104100 186120 104120
rect 186380 104100 186620 104120
rect 186880 104100 187120 104120
rect 187380 104100 187620 104120
rect 187880 104100 188120 104120
rect 188380 104100 188620 104120
rect 188880 104100 189120 104120
rect 189380 104100 189620 104120
rect 189880 104100 190120 104120
rect 190380 104100 190620 104120
rect 190880 104100 191120 104120
rect 191380 104100 191620 104120
rect 191880 104100 192120 104120
rect 192380 104100 192620 104120
rect 192880 104100 193120 104120
rect 193380 104100 193620 104120
rect 193880 104100 194120 104120
rect 194380 104100 194620 104120
rect 194880 104100 195120 104120
rect 195380 104100 195620 104120
rect 195880 104100 196120 104120
rect 196380 104100 196620 104120
rect 196880 104100 197120 104120
rect 197380 104100 197620 104120
rect 197880 104100 198120 104120
rect 198380 104100 198620 104120
rect 198880 104100 199120 104120
rect 199380 104100 199620 104120
rect 199880 104100 200120 104120
rect 200380 104100 200620 104120
rect 200880 104100 201120 104120
rect 201380 104100 201620 104120
rect 201880 104100 202120 104120
rect 202380 104100 202620 104120
rect 202880 104100 203120 104120
rect 203380 104100 203620 104120
rect 203880 104100 204120 104120
rect 204380 104100 204620 104120
rect 204880 104100 205120 104120
rect 205380 104100 205620 104120
rect 205880 104100 206120 104120
rect 206380 104100 206620 104120
rect 206880 104100 207120 104120
rect 207380 104100 207620 104120
rect 207880 104100 208120 104120
rect 208380 104100 208620 104120
rect 208880 104100 209120 104120
rect 209380 104100 209620 104120
rect 209880 104100 210120 104120
rect 210380 104100 210620 104120
rect 210880 104100 211120 104120
rect 211380 104100 211620 104120
rect 211880 104100 212120 104120
rect 212380 104100 212620 104120
rect 212880 104100 213120 104120
rect 213380 104100 213620 104120
rect 213880 104100 214120 104120
rect 214380 104100 214620 104120
rect 214880 104100 215120 104120
rect 215380 104100 215620 104120
rect 215880 104100 216120 104120
rect 216380 104100 216620 104120
rect 216880 104100 217120 104120
rect 217380 104100 217620 104120
rect 217880 104100 218120 104120
rect 218380 104100 218620 104120
rect 218880 104100 219120 104120
rect 219380 104100 219620 104120
rect 219880 104100 220120 104120
rect 220380 104100 220620 104120
rect 220880 104100 221120 104120
rect 221380 104100 221620 104120
rect 221880 104100 222120 104120
rect 222380 104100 222620 104120
rect 222880 104100 223120 104120
rect 223380 104100 223620 104120
rect 223880 104100 224120 104120
rect 224380 104100 224620 104120
rect 224880 104100 225120 104120
rect 225380 104100 225620 104120
rect 225880 104100 226120 104120
rect 226380 104100 226620 104120
rect 226880 104100 227120 104120
rect 227380 104100 227620 104120
rect 227880 104100 228120 104120
rect 228380 104100 228620 104120
rect 228880 104100 229120 104120
rect 229380 104100 229620 104120
rect 229880 104100 230120 104120
rect 230380 104100 230620 104120
rect 230880 104100 231120 104120
rect 231380 104100 231620 104120
rect 231880 104100 232000 104120
rect 178000 103900 232000 104100
rect 178000 103880 178120 103900
rect 178380 103880 178620 103900
rect 178880 103880 179120 103900
rect 179380 103880 179620 103900
rect 179880 103880 180120 103900
rect 180380 103880 180620 103900
rect 180880 103880 181120 103900
rect 181380 103880 181620 103900
rect 181880 103880 182120 103900
rect 182380 103880 182620 103900
rect 182880 103880 183120 103900
rect 183380 103880 183620 103900
rect 183880 103880 184120 103900
rect 184380 103880 184620 103900
rect 184880 103880 185120 103900
rect 185380 103880 185620 103900
rect 185880 103880 186120 103900
rect 186380 103880 186620 103900
rect 186880 103880 187120 103900
rect 187380 103880 187620 103900
rect 187880 103880 188120 103900
rect 188380 103880 188620 103900
rect 188880 103880 189120 103900
rect 189380 103880 189620 103900
rect 189880 103880 190120 103900
rect 190380 103880 190620 103900
rect 190880 103880 191120 103900
rect 191380 103880 191620 103900
rect 191880 103880 192120 103900
rect 192380 103880 192620 103900
rect 192880 103880 193120 103900
rect 193380 103880 193620 103900
rect 193880 103880 194120 103900
rect 194380 103880 194620 103900
rect 194880 103880 195120 103900
rect 195380 103880 195620 103900
rect 195880 103880 196120 103900
rect 196380 103880 196620 103900
rect 196880 103880 197120 103900
rect 197380 103880 197620 103900
rect 197880 103880 198120 103900
rect 198380 103880 198620 103900
rect 198880 103880 199120 103900
rect 199380 103880 199620 103900
rect 199880 103880 200120 103900
rect 200380 103880 200620 103900
rect 200880 103880 201120 103900
rect 201380 103880 201620 103900
rect 201880 103880 202120 103900
rect 202380 103880 202620 103900
rect 202880 103880 203120 103900
rect 203380 103880 203620 103900
rect 203880 103880 204120 103900
rect 204380 103880 204620 103900
rect 204880 103880 205120 103900
rect 205380 103880 205620 103900
rect 205880 103880 206120 103900
rect 206380 103880 206620 103900
rect 206880 103880 207120 103900
rect 207380 103880 207620 103900
rect 207880 103880 208120 103900
rect 208380 103880 208620 103900
rect 208880 103880 209120 103900
rect 209380 103880 209620 103900
rect 209880 103880 210120 103900
rect 210380 103880 210620 103900
rect 210880 103880 211120 103900
rect 211380 103880 211620 103900
rect 211880 103880 212120 103900
rect 212380 103880 212620 103900
rect 212880 103880 213120 103900
rect 213380 103880 213620 103900
rect 213880 103880 214120 103900
rect 214380 103880 214620 103900
rect 214880 103880 215120 103900
rect 215380 103880 215620 103900
rect 215880 103880 216120 103900
rect 216380 103880 216620 103900
rect 216880 103880 217120 103900
rect 217380 103880 217620 103900
rect 217880 103880 218120 103900
rect 218380 103880 218620 103900
rect 218880 103880 219120 103900
rect 219380 103880 219620 103900
rect 219880 103880 220120 103900
rect 220380 103880 220620 103900
rect 220880 103880 221120 103900
rect 221380 103880 221620 103900
rect 221880 103880 222120 103900
rect 222380 103880 222620 103900
rect 222880 103880 223120 103900
rect 223380 103880 223620 103900
rect 223880 103880 224120 103900
rect 224380 103880 224620 103900
rect 224880 103880 225120 103900
rect 225380 103880 225620 103900
rect 225880 103880 226120 103900
rect 226380 103880 226620 103900
rect 226880 103880 227120 103900
rect 227380 103880 227620 103900
rect 227880 103880 228120 103900
rect 228380 103880 228620 103900
rect 228880 103880 229120 103900
rect 229380 103880 229620 103900
rect 229880 103880 230120 103900
rect 230380 103880 230620 103900
rect 230880 103880 231120 103900
rect 231380 103880 231620 103900
rect 231880 103880 232000 103900
rect 9740 103750 9900 103760
rect 9740 103650 9750 103750
rect 9570 103600 9750 103650
rect 9740 103030 9750 103600
rect 9570 102980 9750 103030
rect 9500 102910 9660 102920
rect 9500 102260 9510 102910
rect 9570 102870 9660 102910
rect 9570 102840 9590 102870
rect 9740 102840 9750 102980
rect 9570 102340 9580 102840
rect 9640 102340 9750 102840
rect 9570 102300 9590 102340
rect 9570 102260 9660 102300
rect 9500 102250 9660 102260
rect 9740 102190 9750 102340
rect 9560 102150 9750 102190
rect 9740 101580 9750 102150
rect 9570 101530 9750 101580
rect 9740 101410 9750 101530
rect 9890 101410 9900 103750
rect 178000 103620 178100 103880
rect 178400 103620 178600 103880
rect 178900 103620 179100 103880
rect 179400 103620 179600 103880
rect 179900 103620 180100 103880
rect 180400 103620 180600 103880
rect 180900 103620 181100 103880
rect 181400 103620 181600 103880
rect 181900 103620 182100 103880
rect 182400 103620 182600 103880
rect 182900 103620 183100 103880
rect 183400 103620 183600 103880
rect 183900 103620 184100 103880
rect 184400 103620 184600 103880
rect 184900 103620 185100 103880
rect 185400 103620 185600 103880
rect 185900 103620 186100 103880
rect 186400 103620 186600 103880
rect 186900 103620 187100 103880
rect 187400 103620 187600 103880
rect 187900 103620 188100 103880
rect 188400 103620 188600 103880
rect 188900 103620 189100 103880
rect 189400 103620 189600 103880
rect 189900 103620 190100 103880
rect 190400 103620 190600 103880
rect 190900 103620 191100 103880
rect 191400 103620 191600 103880
rect 191900 103620 192100 103880
rect 192400 103620 192600 103880
rect 192900 103620 193100 103880
rect 193400 103620 193600 103880
rect 193900 103620 194100 103880
rect 194400 103620 194600 103880
rect 194900 103620 195100 103880
rect 195400 103620 195600 103880
rect 195900 103620 196100 103880
rect 196400 103620 196600 103880
rect 196900 103620 197100 103880
rect 197400 103620 197600 103880
rect 197900 103620 198100 103880
rect 198400 103620 198600 103880
rect 198900 103620 199100 103880
rect 199400 103620 199600 103880
rect 199900 103620 200100 103880
rect 200400 103620 200600 103880
rect 200900 103620 201100 103880
rect 201400 103620 201600 103880
rect 201900 103620 202100 103880
rect 202400 103620 202600 103880
rect 202900 103620 203100 103880
rect 203400 103620 203600 103880
rect 203900 103620 204100 103880
rect 204400 103620 204600 103880
rect 204900 103620 205100 103880
rect 205400 103620 205600 103880
rect 205900 103620 206100 103880
rect 206400 103620 206600 103880
rect 206900 103620 207100 103880
rect 207400 103620 207600 103880
rect 207900 103620 208100 103880
rect 208400 103620 208600 103880
rect 208900 103620 209100 103880
rect 209400 103620 209600 103880
rect 209900 103620 210100 103880
rect 210400 103620 210600 103880
rect 210900 103620 211100 103880
rect 211400 103620 211600 103880
rect 211900 103620 212100 103880
rect 212400 103620 212600 103880
rect 212900 103620 213100 103880
rect 213400 103620 213600 103880
rect 213900 103620 214100 103880
rect 214400 103620 214600 103880
rect 214900 103620 215100 103880
rect 215400 103620 215600 103880
rect 215900 103620 216100 103880
rect 216400 103620 216600 103880
rect 216900 103620 217100 103880
rect 217400 103620 217600 103880
rect 217900 103620 218100 103880
rect 218400 103620 218600 103880
rect 218900 103620 219100 103880
rect 219400 103620 219600 103880
rect 219900 103620 220100 103880
rect 220400 103620 220600 103880
rect 220900 103620 221100 103880
rect 221400 103620 221600 103880
rect 221900 103620 222100 103880
rect 222400 103620 222600 103880
rect 222900 103620 223100 103880
rect 223400 103620 223600 103880
rect 223900 103620 224100 103880
rect 224400 103620 224600 103880
rect 224900 103620 225100 103880
rect 225400 103620 225600 103880
rect 225900 103620 226100 103880
rect 226400 103620 226600 103880
rect 226900 103620 227100 103880
rect 227400 103620 227600 103880
rect 227900 103620 228100 103880
rect 228400 103620 228600 103880
rect 228900 103620 229100 103880
rect 229400 103620 229600 103880
rect 229900 103620 230100 103880
rect 230400 103620 230600 103880
rect 230900 103620 231100 103880
rect 231400 103620 231600 103880
rect 231900 103620 232000 103880
rect 178000 103600 178120 103620
rect 178380 103600 178620 103620
rect 178880 103600 179120 103620
rect 179380 103600 179620 103620
rect 179880 103600 180120 103620
rect 180380 103600 180620 103620
rect 180880 103600 181120 103620
rect 181380 103600 181620 103620
rect 181880 103600 182120 103620
rect 182380 103600 182620 103620
rect 182880 103600 183120 103620
rect 183380 103600 183620 103620
rect 183880 103600 184120 103620
rect 184380 103600 184620 103620
rect 184880 103600 185120 103620
rect 185380 103600 185620 103620
rect 185880 103600 186120 103620
rect 186380 103600 186620 103620
rect 186880 103600 187120 103620
rect 187380 103600 187620 103620
rect 187880 103600 188120 103620
rect 188380 103600 188620 103620
rect 188880 103600 189120 103620
rect 189380 103600 189620 103620
rect 189880 103600 190120 103620
rect 190380 103600 190620 103620
rect 190880 103600 191120 103620
rect 191380 103600 191620 103620
rect 191880 103600 192120 103620
rect 192380 103600 192620 103620
rect 192880 103600 193120 103620
rect 193380 103600 193620 103620
rect 193880 103600 194120 103620
rect 194380 103600 194620 103620
rect 194880 103600 195120 103620
rect 195380 103600 195620 103620
rect 195880 103600 196120 103620
rect 196380 103600 196620 103620
rect 196880 103600 197120 103620
rect 197380 103600 197620 103620
rect 197880 103600 198120 103620
rect 198380 103600 198620 103620
rect 198880 103600 199120 103620
rect 199380 103600 199620 103620
rect 199880 103600 200120 103620
rect 200380 103600 200620 103620
rect 200880 103600 201120 103620
rect 201380 103600 201620 103620
rect 201880 103600 202120 103620
rect 202380 103600 202620 103620
rect 202880 103600 203120 103620
rect 203380 103600 203620 103620
rect 203880 103600 204120 103620
rect 204380 103600 204620 103620
rect 204880 103600 205120 103620
rect 205380 103600 205620 103620
rect 205880 103600 206120 103620
rect 206380 103600 206620 103620
rect 206880 103600 207120 103620
rect 207380 103600 207620 103620
rect 207880 103600 208120 103620
rect 208380 103600 208620 103620
rect 208880 103600 209120 103620
rect 209380 103600 209620 103620
rect 209880 103600 210120 103620
rect 210380 103600 210620 103620
rect 210880 103600 211120 103620
rect 211380 103600 211620 103620
rect 211880 103600 212120 103620
rect 212380 103600 212620 103620
rect 212880 103600 213120 103620
rect 213380 103600 213620 103620
rect 213880 103600 214120 103620
rect 214380 103600 214620 103620
rect 214880 103600 215120 103620
rect 215380 103600 215620 103620
rect 215880 103600 216120 103620
rect 216380 103600 216620 103620
rect 216880 103600 217120 103620
rect 217380 103600 217620 103620
rect 217880 103600 218120 103620
rect 218380 103600 218620 103620
rect 218880 103600 219120 103620
rect 219380 103600 219620 103620
rect 219880 103600 220120 103620
rect 220380 103600 220620 103620
rect 220880 103600 221120 103620
rect 221380 103600 221620 103620
rect 221880 103600 222120 103620
rect 222380 103600 222620 103620
rect 222880 103600 223120 103620
rect 223380 103600 223620 103620
rect 223880 103600 224120 103620
rect 224380 103600 224620 103620
rect 224880 103600 225120 103620
rect 225380 103600 225620 103620
rect 225880 103600 226120 103620
rect 226380 103600 226620 103620
rect 226880 103600 227120 103620
rect 227380 103600 227620 103620
rect 227880 103600 228120 103620
rect 228380 103600 228620 103620
rect 228880 103600 229120 103620
rect 229380 103600 229620 103620
rect 229880 103600 230120 103620
rect 230380 103600 230620 103620
rect 230880 103600 231120 103620
rect 231380 103600 231620 103620
rect 231880 103600 232000 103620
rect 178000 103400 232000 103600
rect 178000 103380 178120 103400
rect 178380 103380 178620 103400
rect 178880 103380 179120 103400
rect 179380 103380 179620 103400
rect 179880 103380 180120 103400
rect 180380 103380 180620 103400
rect 180880 103380 181120 103400
rect 181380 103380 181620 103400
rect 181880 103380 182120 103400
rect 182380 103380 182620 103400
rect 182880 103380 183120 103400
rect 183380 103380 183620 103400
rect 183880 103380 184120 103400
rect 184380 103380 184620 103400
rect 184880 103380 185120 103400
rect 185380 103380 185620 103400
rect 185880 103380 186120 103400
rect 186380 103380 186620 103400
rect 186880 103380 187120 103400
rect 187380 103380 187620 103400
rect 187880 103380 188120 103400
rect 188380 103380 188620 103400
rect 188880 103380 189120 103400
rect 189380 103380 189620 103400
rect 189880 103380 190120 103400
rect 190380 103380 190620 103400
rect 190880 103380 191120 103400
rect 191380 103380 191620 103400
rect 191880 103380 192120 103400
rect 192380 103380 192620 103400
rect 192880 103380 193120 103400
rect 193380 103380 193620 103400
rect 193880 103380 194120 103400
rect 194380 103380 194620 103400
rect 194880 103380 195120 103400
rect 195380 103380 195620 103400
rect 195880 103380 196120 103400
rect 196380 103380 196620 103400
rect 196880 103380 197120 103400
rect 197380 103380 197620 103400
rect 197880 103380 198120 103400
rect 198380 103380 198620 103400
rect 198880 103380 199120 103400
rect 199380 103380 199620 103400
rect 199880 103380 200120 103400
rect 200380 103380 200620 103400
rect 200880 103380 201120 103400
rect 201380 103380 201620 103400
rect 201880 103380 202120 103400
rect 202380 103380 202620 103400
rect 202880 103380 203120 103400
rect 203380 103380 203620 103400
rect 203880 103380 204120 103400
rect 204380 103380 204620 103400
rect 204880 103380 205120 103400
rect 205380 103380 205620 103400
rect 205880 103380 206120 103400
rect 206380 103380 206620 103400
rect 206880 103380 207120 103400
rect 207380 103380 207620 103400
rect 207880 103380 208120 103400
rect 208380 103380 208620 103400
rect 208880 103380 209120 103400
rect 209380 103380 209620 103400
rect 209880 103380 210120 103400
rect 210380 103380 210620 103400
rect 210880 103380 211120 103400
rect 211380 103380 211620 103400
rect 211880 103380 212120 103400
rect 212380 103380 212620 103400
rect 212880 103380 213120 103400
rect 213380 103380 213620 103400
rect 213880 103380 214120 103400
rect 214380 103380 214620 103400
rect 214880 103380 215120 103400
rect 215380 103380 215620 103400
rect 215880 103380 216120 103400
rect 216380 103380 216620 103400
rect 216880 103380 217120 103400
rect 217380 103380 217620 103400
rect 217880 103380 218120 103400
rect 218380 103380 218620 103400
rect 218880 103380 219120 103400
rect 219380 103380 219620 103400
rect 219880 103380 220120 103400
rect 220380 103380 220620 103400
rect 220880 103380 221120 103400
rect 221380 103380 221620 103400
rect 221880 103380 222120 103400
rect 222380 103380 222620 103400
rect 222880 103380 223120 103400
rect 223380 103380 223620 103400
rect 223880 103380 224120 103400
rect 224380 103380 224620 103400
rect 224880 103380 225120 103400
rect 225380 103380 225620 103400
rect 225880 103380 226120 103400
rect 226380 103380 226620 103400
rect 226880 103380 227120 103400
rect 227380 103380 227620 103400
rect 227880 103380 228120 103400
rect 228380 103380 228620 103400
rect 228880 103380 229120 103400
rect 229380 103380 229620 103400
rect 229880 103380 230120 103400
rect 230380 103380 230620 103400
rect 230880 103380 231120 103400
rect 231380 103380 231620 103400
rect 231880 103380 232000 103400
rect 178000 103120 178100 103380
rect 178400 103120 178600 103380
rect 178900 103120 179100 103380
rect 179400 103120 179600 103380
rect 179900 103120 180100 103380
rect 180400 103120 180600 103380
rect 180900 103120 181100 103380
rect 181400 103120 181600 103380
rect 181900 103120 182100 103380
rect 182400 103120 182600 103380
rect 182900 103120 183100 103380
rect 183400 103120 183600 103380
rect 183900 103120 184100 103380
rect 184400 103120 184600 103380
rect 184900 103120 185100 103380
rect 185400 103120 185600 103380
rect 185900 103120 186100 103380
rect 186400 103120 186600 103380
rect 186900 103120 187100 103380
rect 187400 103120 187600 103380
rect 187900 103120 188100 103380
rect 188400 103120 188600 103380
rect 188900 103120 189100 103380
rect 189400 103120 189600 103380
rect 189900 103120 190100 103380
rect 190400 103120 190600 103380
rect 190900 103120 191100 103380
rect 191400 103120 191600 103380
rect 191900 103120 192100 103380
rect 192400 103120 192600 103380
rect 192900 103120 193100 103380
rect 193400 103120 193600 103380
rect 193900 103120 194100 103380
rect 194400 103120 194600 103380
rect 194900 103120 195100 103380
rect 195400 103120 195600 103380
rect 195900 103120 196100 103380
rect 196400 103120 196600 103380
rect 196900 103120 197100 103380
rect 197400 103120 197600 103380
rect 197900 103120 198100 103380
rect 198400 103120 198600 103380
rect 198900 103120 199100 103380
rect 199400 103120 199600 103380
rect 199900 103120 200100 103380
rect 200400 103120 200600 103380
rect 200900 103120 201100 103380
rect 201400 103120 201600 103380
rect 201900 103120 202100 103380
rect 202400 103120 202600 103380
rect 202900 103120 203100 103380
rect 203400 103120 203600 103380
rect 203900 103120 204100 103380
rect 204400 103120 204600 103380
rect 204900 103120 205100 103380
rect 205400 103120 205600 103380
rect 205900 103120 206100 103380
rect 206400 103120 206600 103380
rect 206900 103120 207100 103380
rect 207400 103120 207600 103380
rect 207900 103120 208100 103380
rect 208400 103120 208600 103380
rect 208900 103120 209100 103380
rect 209400 103120 209600 103380
rect 209900 103120 210100 103380
rect 210400 103120 210600 103380
rect 210900 103120 211100 103380
rect 211400 103120 211600 103380
rect 211900 103120 212100 103380
rect 212400 103120 212600 103380
rect 212900 103120 213100 103380
rect 213400 103120 213600 103380
rect 213900 103120 214100 103380
rect 214400 103120 214600 103380
rect 214900 103120 215100 103380
rect 215400 103120 215600 103380
rect 215900 103120 216100 103380
rect 216400 103120 216600 103380
rect 216900 103120 217100 103380
rect 217400 103120 217600 103380
rect 217900 103120 218100 103380
rect 218400 103120 218600 103380
rect 218900 103120 219100 103380
rect 219400 103120 219600 103380
rect 219900 103120 220100 103380
rect 220400 103120 220600 103380
rect 220900 103120 221100 103380
rect 221400 103120 221600 103380
rect 221900 103120 222100 103380
rect 222400 103120 222600 103380
rect 222900 103120 223100 103380
rect 223400 103120 223600 103380
rect 223900 103120 224100 103380
rect 224400 103120 224600 103380
rect 224900 103120 225100 103380
rect 225400 103120 225600 103380
rect 225900 103120 226100 103380
rect 226400 103120 226600 103380
rect 226900 103120 227100 103380
rect 227400 103120 227600 103380
rect 227900 103120 228100 103380
rect 228400 103120 228600 103380
rect 228900 103120 229100 103380
rect 229400 103120 229600 103380
rect 229900 103120 230100 103380
rect 230400 103120 230600 103380
rect 230900 103120 231100 103380
rect 231400 103120 231600 103380
rect 231900 103120 232000 103380
rect 178000 103100 178120 103120
rect 178380 103100 178620 103120
rect 178880 103100 179120 103120
rect 179380 103100 179620 103120
rect 179880 103100 180120 103120
rect 180380 103100 180620 103120
rect 180880 103100 181120 103120
rect 181380 103100 181620 103120
rect 181880 103100 182120 103120
rect 182380 103100 182620 103120
rect 182880 103100 183120 103120
rect 183380 103100 183620 103120
rect 183880 103100 184120 103120
rect 184380 103100 184620 103120
rect 184880 103100 185120 103120
rect 185380 103100 185620 103120
rect 185880 103100 186120 103120
rect 186380 103100 186620 103120
rect 186880 103100 187120 103120
rect 187380 103100 187620 103120
rect 187880 103100 188120 103120
rect 188380 103100 188620 103120
rect 188880 103100 189120 103120
rect 189380 103100 189620 103120
rect 189880 103100 190120 103120
rect 190380 103100 190620 103120
rect 190880 103100 191120 103120
rect 191380 103100 191620 103120
rect 191880 103100 192120 103120
rect 192380 103100 192620 103120
rect 192880 103100 193120 103120
rect 193380 103100 193620 103120
rect 193880 103100 194120 103120
rect 194380 103100 194620 103120
rect 194880 103100 195120 103120
rect 195380 103100 195620 103120
rect 195880 103100 196120 103120
rect 196380 103100 196620 103120
rect 196880 103100 197120 103120
rect 197380 103100 197620 103120
rect 197880 103100 198120 103120
rect 198380 103100 198620 103120
rect 198880 103100 199120 103120
rect 199380 103100 199620 103120
rect 199880 103100 200120 103120
rect 200380 103100 200620 103120
rect 200880 103100 201120 103120
rect 201380 103100 201620 103120
rect 201880 103100 202120 103120
rect 202380 103100 202620 103120
rect 202880 103100 203120 103120
rect 203380 103100 203620 103120
rect 203880 103100 204120 103120
rect 204380 103100 204620 103120
rect 204880 103100 205120 103120
rect 205380 103100 205620 103120
rect 205880 103100 206120 103120
rect 206380 103100 206620 103120
rect 206880 103100 207120 103120
rect 207380 103100 207620 103120
rect 207880 103100 208120 103120
rect 208380 103100 208620 103120
rect 208880 103100 209120 103120
rect 209380 103100 209620 103120
rect 209880 103100 210120 103120
rect 210380 103100 210620 103120
rect 210880 103100 211120 103120
rect 211380 103100 211620 103120
rect 211880 103100 212120 103120
rect 212380 103100 212620 103120
rect 212880 103100 213120 103120
rect 213380 103100 213620 103120
rect 213880 103100 214120 103120
rect 214380 103100 214620 103120
rect 214880 103100 215120 103120
rect 215380 103100 215620 103120
rect 215880 103100 216120 103120
rect 216380 103100 216620 103120
rect 216880 103100 217120 103120
rect 217380 103100 217620 103120
rect 217880 103100 218120 103120
rect 218380 103100 218620 103120
rect 218880 103100 219120 103120
rect 219380 103100 219620 103120
rect 219880 103100 220120 103120
rect 220380 103100 220620 103120
rect 220880 103100 221120 103120
rect 221380 103100 221620 103120
rect 221880 103100 222120 103120
rect 222380 103100 222620 103120
rect 222880 103100 223120 103120
rect 223380 103100 223620 103120
rect 223880 103100 224120 103120
rect 224380 103100 224620 103120
rect 224880 103100 225120 103120
rect 225380 103100 225620 103120
rect 225880 103100 226120 103120
rect 226380 103100 226620 103120
rect 226880 103100 227120 103120
rect 227380 103100 227620 103120
rect 227880 103100 228120 103120
rect 228380 103100 228620 103120
rect 228880 103100 229120 103120
rect 229380 103100 229620 103120
rect 229880 103100 230120 103120
rect 230380 103100 230620 103120
rect 230880 103100 231120 103120
rect 231380 103100 231620 103120
rect 231880 103100 232000 103120
rect 178000 102900 232000 103100
rect 178000 102880 178120 102900
rect 178380 102880 178620 102900
rect 178880 102880 179120 102900
rect 179380 102880 179620 102900
rect 179880 102880 180120 102900
rect 180380 102880 180620 102900
rect 180880 102880 181120 102900
rect 181380 102880 181620 102900
rect 181880 102880 182120 102900
rect 182380 102880 182620 102900
rect 182880 102880 183120 102900
rect 183380 102880 183620 102900
rect 183880 102880 184120 102900
rect 184380 102880 184620 102900
rect 184880 102880 185120 102900
rect 185380 102880 185620 102900
rect 185880 102880 186120 102900
rect 186380 102880 186620 102900
rect 186880 102880 187120 102900
rect 187380 102880 187620 102900
rect 187880 102880 188120 102900
rect 188380 102880 188620 102900
rect 188880 102880 189120 102900
rect 189380 102880 189620 102900
rect 189880 102880 190120 102900
rect 190380 102880 190620 102900
rect 190880 102880 191120 102900
rect 191380 102880 191620 102900
rect 191880 102880 192120 102900
rect 192380 102880 192620 102900
rect 192880 102880 193120 102900
rect 193380 102880 193620 102900
rect 193880 102880 194120 102900
rect 194380 102880 194620 102900
rect 194880 102880 195120 102900
rect 195380 102880 195620 102900
rect 195880 102880 196120 102900
rect 196380 102880 196620 102900
rect 196880 102880 197120 102900
rect 197380 102880 197620 102900
rect 197880 102880 198120 102900
rect 198380 102880 198620 102900
rect 198880 102880 199120 102900
rect 199380 102880 199620 102900
rect 199880 102880 200120 102900
rect 200380 102880 200620 102900
rect 200880 102880 201120 102900
rect 201380 102880 201620 102900
rect 201880 102880 202120 102900
rect 202380 102880 202620 102900
rect 202880 102880 203120 102900
rect 203380 102880 203620 102900
rect 203880 102880 204120 102900
rect 204380 102880 204620 102900
rect 204880 102880 205120 102900
rect 205380 102880 205620 102900
rect 205880 102880 206120 102900
rect 206380 102880 206620 102900
rect 206880 102880 207120 102900
rect 207380 102880 207620 102900
rect 207880 102880 208120 102900
rect 208380 102880 208620 102900
rect 208880 102880 209120 102900
rect 209380 102880 209620 102900
rect 209880 102880 210120 102900
rect 210380 102880 210620 102900
rect 210880 102880 211120 102900
rect 211380 102880 211620 102900
rect 211880 102880 212120 102900
rect 212380 102880 212620 102900
rect 212880 102880 213120 102900
rect 213380 102880 213620 102900
rect 213880 102880 214120 102900
rect 214380 102880 214620 102900
rect 214880 102880 215120 102900
rect 215380 102880 215620 102900
rect 215880 102880 216120 102900
rect 216380 102880 216620 102900
rect 216880 102880 217120 102900
rect 217380 102880 217620 102900
rect 217880 102880 218120 102900
rect 218380 102880 218620 102900
rect 218880 102880 219120 102900
rect 219380 102880 219620 102900
rect 219880 102880 220120 102900
rect 220380 102880 220620 102900
rect 220880 102880 221120 102900
rect 221380 102880 221620 102900
rect 221880 102880 222120 102900
rect 222380 102880 222620 102900
rect 222880 102880 223120 102900
rect 223380 102880 223620 102900
rect 223880 102880 224120 102900
rect 224380 102880 224620 102900
rect 224880 102880 225120 102900
rect 225380 102880 225620 102900
rect 225880 102880 226120 102900
rect 226380 102880 226620 102900
rect 226880 102880 227120 102900
rect 227380 102880 227620 102900
rect 227880 102880 228120 102900
rect 228380 102880 228620 102900
rect 228880 102880 229120 102900
rect 229380 102880 229620 102900
rect 229880 102880 230120 102900
rect 230380 102880 230620 102900
rect 230880 102880 231120 102900
rect 231380 102880 231620 102900
rect 231880 102880 232000 102900
rect 178000 102620 178100 102880
rect 178400 102620 178600 102880
rect 178900 102620 179100 102880
rect 179400 102620 179600 102880
rect 179900 102620 180100 102880
rect 180400 102620 180600 102880
rect 180900 102620 181100 102880
rect 181400 102620 181600 102880
rect 181900 102620 182100 102880
rect 182400 102620 182600 102880
rect 182900 102620 183100 102880
rect 183400 102620 183600 102880
rect 183900 102620 184100 102880
rect 184400 102620 184600 102880
rect 184900 102620 185100 102880
rect 185400 102620 185600 102880
rect 185900 102620 186100 102880
rect 186400 102620 186600 102880
rect 186900 102620 187100 102880
rect 187400 102620 187600 102880
rect 187900 102620 188100 102880
rect 188400 102620 188600 102880
rect 188900 102620 189100 102880
rect 189400 102620 189600 102880
rect 189900 102620 190100 102880
rect 190400 102620 190600 102880
rect 190900 102620 191100 102880
rect 191400 102620 191600 102880
rect 191900 102620 192100 102880
rect 192400 102620 192600 102880
rect 192900 102620 193100 102880
rect 193400 102620 193600 102880
rect 193900 102620 194100 102880
rect 194400 102620 194600 102880
rect 194900 102620 195100 102880
rect 195400 102620 195600 102880
rect 195900 102620 196100 102880
rect 196400 102620 196600 102880
rect 196900 102620 197100 102880
rect 197400 102620 197600 102880
rect 197900 102620 198100 102880
rect 198400 102620 198600 102880
rect 198900 102620 199100 102880
rect 199400 102620 199600 102880
rect 199900 102620 200100 102880
rect 200400 102620 200600 102880
rect 200900 102620 201100 102880
rect 201400 102620 201600 102880
rect 201900 102620 202100 102880
rect 202400 102620 202600 102880
rect 202900 102620 203100 102880
rect 203400 102620 203600 102880
rect 203900 102620 204100 102880
rect 204400 102620 204600 102880
rect 204900 102620 205100 102880
rect 205400 102620 205600 102880
rect 205900 102620 206100 102880
rect 206400 102620 206600 102880
rect 206900 102620 207100 102880
rect 207400 102620 207600 102880
rect 207900 102620 208100 102880
rect 208400 102620 208600 102880
rect 208900 102620 209100 102880
rect 209400 102620 209600 102880
rect 209900 102620 210100 102880
rect 210400 102620 210600 102880
rect 210900 102620 211100 102880
rect 211400 102620 211600 102880
rect 211900 102620 212100 102880
rect 212400 102620 212600 102880
rect 212900 102620 213100 102880
rect 213400 102620 213600 102880
rect 213900 102620 214100 102880
rect 214400 102620 214600 102880
rect 214900 102620 215100 102880
rect 215400 102620 215600 102880
rect 215900 102620 216100 102880
rect 216400 102620 216600 102880
rect 216900 102620 217100 102880
rect 217400 102620 217600 102880
rect 217900 102620 218100 102880
rect 218400 102620 218600 102880
rect 218900 102620 219100 102880
rect 219400 102620 219600 102880
rect 219900 102620 220100 102880
rect 220400 102620 220600 102880
rect 220900 102620 221100 102880
rect 221400 102620 221600 102880
rect 221900 102620 222100 102880
rect 222400 102620 222600 102880
rect 222900 102620 223100 102880
rect 223400 102620 223600 102880
rect 223900 102620 224100 102880
rect 224400 102620 224600 102880
rect 224900 102620 225100 102880
rect 225400 102620 225600 102880
rect 225900 102620 226100 102880
rect 226400 102620 226600 102880
rect 226900 102620 227100 102880
rect 227400 102620 227600 102880
rect 227900 102620 228100 102880
rect 228400 102620 228600 102880
rect 228900 102620 229100 102880
rect 229400 102620 229600 102880
rect 229900 102620 230100 102880
rect 230400 102620 230600 102880
rect 230900 102620 231100 102880
rect 231400 102620 231600 102880
rect 231900 102620 232000 102880
rect 178000 102600 178120 102620
rect 178380 102600 178620 102620
rect 178880 102600 179120 102620
rect 179380 102600 179620 102620
rect 179880 102600 180120 102620
rect 180380 102600 180620 102620
rect 180880 102600 181120 102620
rect 181380 102600 181620 102620
rect 181880 102600 182120 102620
rect 182380 102600 182620 102620
rect 182880 102600 183120 102620
rect 183380 102600 183620 102620
rect 183880 102600 184120 102620
rect 184380 102600 184620 102620
rect 184880 102600 185120 102620
rect 185380 102600 185620 102620
rect 185880 102600 186120 102620
rect 186380 102600 186620 102620
rect 186880 102600 187120 102620
rect 187380 102600 187620 102620
rect 187880 102600 188120 102620
rect 188380 102600 188620 102620
rect 188880 102600 189120 102620
rect 189380 102600 189620 102620
rect 189880 102600 190120 102620
rect 190380 102600 190620 102620
rect 190880 102600 191120 102620
rect 191380 102600 191620 102620
rect 191880 102600 192120 102620
rect 192380 102600 192620 102620
rect 192880 102600 193120 102620
rect 193380 102600 193620 102620
rect 193880 102600 194120 102620
rect 194380 102600 194620 102620
rect 194880 102600 195120 102620
rect 195380 102600 195620 102620
rect 195880 102600 196120 102620
rect 196380 102600 196620 102620
rect 196880 102600 197120 102620
rect 197380 102600 197620 102620
rect 197880 102600 198120 102620
rect 198380 102600 198620 102620
rect 198880 102600 199120 102620
rect 199380 102600 199620 102620
rect 199880 102600 200120 102620
rect 200380 102600 200620 102620
rect 200880 102600 201120 102620
rect 201380 102600 201620 102620
rect 201880 102600 202120 102620
rect 202380 102600 202620 102620
rect 202880 102600 203120 102620
rect 203380 102600 203620 102620
rect 203880 102600 204120 102620
rect 204380 102600 204620 102620
rect 204880 102600 205120 102620
rect 205380 102600 205620 102620
rect 205880 102600 206120 102620
rect 206380 102600 206620 102620
rect 206880 102600 207120 102620
rect 207380 102600 207620 102620
rect 207880 102600 208120 102620
rect 208380 102600 208620 102620
rect 208880 102600 209120 102620
rect 209380 102600 209620 102620
rect 209880 102600 210120 102620
rect 210380 102600 210620 102620
rect 210880 102600 211120 102620
rect 211380 102600 211620 102620
rect 211880 102600 212120 102620
rect 212380 102600 212620 102620
rect 212880 102600 213120 102620
rect 213380 102600 213620 102620
rect 213880 102600 214120 102620
rect 214380 102600 214620 102620
rect 214880 102600 215120 102620
rect 215380 102600 215620 102620
rect 215880 102600 216120 102620
rect 216380 102600 216620 102620
rect 216880 102600 217120 102620
rect 217380 102600 217620 102620
rect 217880 102600 218120 102620
rect 218380 102600 218620 102620
rect 218880 102600 219120 102620
rect 219380 102600 219620 102620
rect 219880 102600 220120 102620
rect 220380 102600 220620 102620
rect 220880 102600 221120 102620
rect 221380 102600 221620 102620
rect 221880 102600 222120 102620
rect 222380 102600 222620 102620
rect 222880 102600 223120 102620
rect 223380 102600 223620 102620
rect 223880 102600 224120 102620
rect 224380 102600 224620 102620
rect 224880 102600 225120 102620
rect 225380 102600 225620 102620
rect 225880 102600 226120 102620
rect 226380 102600 226620 102620
rect 226880 102600 227120 102620
rect 227380 102600 227620 102620
rect 227880 102600 228120 102620
rect 228380 102600 228620 102620
rect 228880 102600 229120 102620
rect 229380 102600 229620 102620
rect 229880 102600 230120 102620
rect 230380 102600 230620 102620
rect 230880 102600 231120 102620
rect 231380 102600 231620 102620
rect 231880 102600 232000 102620
rect 178000 102400 232000 102600
rect 178000 102380 178120 102400
rect 178380 102380 178620 102400
rect 178880 102380 179120 102400
rect 179380 102380 179620 102400
rect 179880 102380 180120 102400
rect 180380 102380 180620 102400
rect 180880 102380 181120 102400
rect 181380 102380 181620 102400
rect 181880 102380 182120 102400
rect 182380 102380 182620 102400
rect 182880 102380 183120 102400
rect 183380 102380 183620 102400
rect 183880 102380 184120 102400
rect 184380 102380 184620 102400
rect 184880 102380 185120 102400
rect 185380 102380 185620 102400
rect 185880 102380 186120 102400
rect 186380 102380 186620 102400
rect 186880 102380 187120 102400
rect 187380 102380 187620 102400
rect 187880 102380 188120 102400
rect 188380 102380 188620 102400
rect 188880 102380 189120 102400
rect 189380 102380 189620 102400
rect 189880 102380 190120 102400
rect 190380 102380 190620 102400
rect 190880 102380 191120 102400
rect 191380 102380 191620 102400
rect 191880 102380 192120 102400
rect 192380 102380 192620 102400
rect 192880 102380 193120 102400
rect 193380 102380 193620 102400
rect 193880 102380 194120 102400
rect 194380 102380 194620 102400
rect 194880 102380 195120 102400
rect 195380 102380 195620 102400
rect 195880 102380 196120 102400
rect 196380 102380 196620 102400
rect 196880 102380 197120 102400
rect 197380 102380 197620 102400
rect 197880 102380 198120 102400
rect 198380 102380 198620 102400
rect 198880 102380 199120 102400
rect 199380 102380 199620 102400
rect 199880 102380 200120 102400
rect 200380 102380 200620 102400
rect 200880 102380 201120 102400
rect 201380 102380 201620 102400
rect 201880 102380 202120 102400
rect 202380 102380 202620 102400
rect 202880 102380 203120 102400
rect 203380 102380 203620 102400
rect 203880 102380 204120 102400
rect 204380 102380 204620 102400
rect 204880 102380 205120 102400
rect 205380 102380 205620 102400
rect 205880 102380 206120 102400
rect 206380 102380 206620 102400
rect 206880 102380 207120 102400
rect 207380 102380 207620 102400
rect 207880 102380 208120 102400
rect 208380 102380 208620 102400
rect 208880 102380 209120 102400
rect 209380 102380 209620 102400
rect 209880 102380 210120 102400
rect 210380 102380 210620 102400
rect 210880 102380 211120 102400
rect 211380 102380 211620 102400
rect 211880 102380 212120 102400
rect 212380 102380 212620 102400
rect 212880 102380 213120 102400
rect 213380 102380 213620 102400
rect 213880 102380 214120 102400
rect 214380 102380 214620 102400
rect 214880 102380 215120 102400
rect 215380 102380 215620 102400
rect 215880 102380 216120 102400
rect 216380 102380 216620 102400
rect 216880 102380 217120 102400
rect 217380 102380 217620 102400
rect 217880 102380 218120 102400
rect 218380 102380 218620 102400
rect 218880 102380 219120 102400
rect 219380 102380 219620 102400
rect 219880 102380 220120 102400
rect 220380 102380 220620 102400
rect 220880 102380 221120 102400
rect 221380 102380 221620 102400
rect 221880 102380 222120 102400
rect 222380 102380 222620 102400
rect 222880 102380 223120 102400
rect 223380 102380 223620 102400
rect 223880 102380 224120 102400
rect 224380 102380 224620 102400
rect 224880 102380 225120 102400
rect 225380 102380 225620 102400
rect 225880 102380 226120 102400
rect 226380 102380 226620 102400
rect 226880 102380 227120 102400
rect 227380 102380 227620 102400
rect 227880 102380 228120 102400
rect 228380 102380 228620 102400
rect 228880 102380 229120 102400
rect 229380 102380 229620 102400
rect 229880 102380 230120 102400
rect 230380 102380 230620 102400
rect 230880 102380 231120 102400
rect 231380 102380 231620 102400
rect 231880 102380 232000 102400
rect 178000 102120 178100 102380
rect 178400 102120 178600 102380
rect 178900 102120 179100 102380
rect 179400 102120 179600 102380
rect 179900 102120 180100 102380
rect 180400 102120 180600 102380
rect 180900 102120 181100 102380
rect 181400 102120 181600 102380
rect 181900 102120 182100 102380
rect 182400 102120 182600 102380
rect 182900 102120 183100 102380
rect 183400 102120 183600 102380
rect 183900 102120 184100 102380
rect 184400 102120 184600 102380
rect 184900 102120 185100 102380
rect 185400 102120 185600 102380
rect 185900 102120 186100 102380
rect 186400 102120 186600 102380
rect 186900 102120 187100 102380
rect 187400 102120 187600 102380
rect 187900 102120 188100 102380
rect 188400 102120 188600 102380
rect 188900 102120 189100 102380
rect 189400 102120 189600 102380
rect 189900 102120 190100 102380
rect 190400 102120 190600 102380
rect 190900 102120 191100 102380
rect 191400 102120 191600 102380
rect 191900 102120 192100 102380
rect 192400 102120 192600 102380
rect 192900 102120 193100 102380
rect 193400 102120 193600 102380
rect 193900 102120 194100 102380
rect 194400 102120 194600 102380
rect 194900 102120 195100 102380
rect 195400 102120 195600 102380
rect 195900 102120 196100 102380
rect 196400 102120 196600 102380
rect 196900 102120 197100 102380
rect 197400 102120 197600 102380
rect 197900 102120 198100 102380
rect 198400 102120 198600 102380
rect 198900 102120 199100 102380
rect 199400 102120 199600 102380
rect 199900 102120 200100 102380
rect 200400 102120 200600 102380
rect 200900 102120 201100 102380
rect 201400 102120 201600 102380
rect 201900 102120 202100 102380
rect 202400 102120 202600 102380
rect 202900 102120 203100 102380
rect 203400 102120 203600 102380
rect 203900 102120 204100 102380
rect 204400 102120 204600 102380
rect 204900 102120 205100 102380
rect 205400 102120 205600 102380
rect 205900 102120 206100 102380
rect 206400 102120 206600 102380
rect 206900 102120 207100 102380
rect 207400 102120 207600 102380
rect 207900 102120 208100 102380
rect 208400 102120 208600 102380
rect 208900 102120 209100 102380
rect 209400 102120 209600 102380
rect 209900 102120 210100 102380
rect 210400 102120 210600 102380
rect 210900 102120 211100 102380
rect 211400 102120 211600 102380
rect 211900 102120 212100 102380
rect 212400 102120 212600 102380
rect 212900 102120 213100 102380
rect 213400 102120 213600 102380
rect 213900 102120 214100 102380
rect 214400 102120 214600 102380
rect 214900 102120 215100 102380
rect 215400 102120 215600 102380
rect 215900 102120 216100 102380
rect 216400 102120 216600 102380
rect 216900 102120 217100 102380
rect 217400 102120 217600 102380
rect 217900 102120 218100 102380
rect 218400 102120 218600 102380
rect 218900 102120 219100 102380
rect 219400 102120 219600 102380
rect 219900 102120 220100 102380
rect 220400 102120 220600 102380
rect 220900 102120 221100 102380
rect 221400 102120 221600 102380
rect 221900 102120 222100 102380
rect 222400 102120 222600 102380
rect 222900 102120 223100 102380
rect 223400 102120 223600 102380
rect 223900 102120 224100 102380
rect 224400 102120 224600 102380
rect 224900 102120 225100 102380
rect 225400 102120 225600 102380
rect 225900 102120 226100 102380
rect 226400 102120 226600 102380
rect 226900 102120 227100 102380
rect 227400 102120 227600 102380
rect 227900 102120 228100 102380
rect 228400 102120 228600 102380
rect 228900 102120 229100 102380
rect 229400 102120 229600 102380
rect 229900 102120 230100 102380
rect 230400 102120 230600 102380
rect 230900 102120 231100 102380
rect 231400 102120 231600 102380
rect 231900 102120 232000 102380
rect 178000 102100 178120 102120
rect 178380 102100 178620 102120
rect 178880 102100 179120 102120
rect 179380 102100 179620 102120
rect 179880 102100 180120 102120
rect 180380 102100 180620 102120
rect 180880 102100 181120 102120
rect 181380 102100 181620 102120
rect 181880 102100 182120 102120
rect 182380 102100 182620 102120
rect 182880 102100 183120 102120
rect 183380 102100 183620 102120
rect 183880 102100 184120 102120
rect 184380 102100 184620 102120
rect 184880 102100 185120 102120
rect 185380 102100 185620 102120
rect 185880 102100 186120 102120
rect 186380 102100 186620 102120
rect 186880 102100 187120 102120
rect 187380 102100 187620 102120
rect 187880 102100 188120 102120
rect 188380 102100 188620 102120
rect 188880 102100 189120 102120
rect 189380 102100 189620 102120
rect 189880 102100 190120 102120
rect 190380 102100 190620 102120
rect 190880 102100 191120 102120
rect 191380 102100 191620 102120
rect 191880 102100 192120 102120
rect 192380 102100 192620 102120
rect 192880 102100 193120 102120
rect 193380 102100 193620 102120
rect 193880 102100 194120 102120
rect 194380 102100 194620 102120
rect 194880 102100 195120 102120
rect 195380 102100 195620 102120
rect 195880 102100 196120 102120
rect 196380 102100 196620 102120
rect 196880 102100 197120 102120
rect 197380 102100 197620 102120
rect 197880 102100 198120 102120
rect 198380 102100 198620 102120
rect 198880 102100 199120 102120
rect 199380 102100 199620 102120
rect 199880 102100 200120 102120
rect 200380 102100 200620 102120
rect 200880 102100 201120 102120
rect 201380 102100 201620 102120
rect 201880 102100 202120 102120
rect 202380 102100 202620 102120
rect 202880 102100 203120 102120
rect 203380 102100 203620 102120
rect 203880 102100 204120 102120
rect 204380 102100 204620 102120
rect 204880 102100 205120 102120
rect 205380 102100 205620 102120
rect 205880 102100 206120 102120
rect 206380 102100 206620 102120
rect 206880 102100 207120 102120
rect 207380 102100 207620 102120
rect 207880 102100 208120 102120
rect 208380 102100 208620 102120
rect 208880 102100 209120 102120
rect 209380 102100 209620 102120
rect 209880 102100 210120 102120
rect 210380 102100 210620 102120
rect 210880 102100 211120 102120
rect 211380 102100 211620 102120
rect 211880 102100 212120 102120
rect 212380 102100 212620 102120
rect 212880 102100 213120 102120
rect 213380 102100 213620 102120
rect 213880 102100 214120 102120
rect 214380 102100 214620 102120
rect 214880 102100 215120 102120
rect 215380 102100 215620 102120
rect 215880 102100 216120 102120
rect 216380 102100 216620 102120
rect 216880 102100 217120 102120
rect 217380 102100 217620 102120
rect 217880 102100 218120 102120
rect 218380 102100 218620 102120
rect 218880 102100 219120 102120
rect 219380 102100 219620 102120
rect 219880 102100 220120 102120
rect 220380 102100 220620 102120
rect 220880 102100 221120 102120
rect 221380 102100 221620 102120
rect 221880 102100 222120 102120
rect 222380 102100 222620 102120
rect 222880 102100 223120 102120
rect 223380 102100 223620 102120
rect 223880 102100 224120 102120
rect 224380 102100 224620 102120
rect 224880 102100 225120 102120
rect 225380 102100 225620 102120
rect 225880 102100 226120 102120
rect 226380 102100 226620 102120
rect 226880 102100 227120 102120
rect 227380 102100 227620 102120
rect 227880 102100 228120 102120
rect 228380 102100 228620 102120
rect 228880 102100 229120 102120
rect 229380 102100 229620 102120
rect 229880 102100 230120 102120
rect 230380 102100 230620 102120
rect 230880 102100 231120 102120
rect 231380 102100 231620 102120
rect 231880 102100 232000 102120
rect 178000 102000 232000 102100
rect 9740 101400 9900 101410
<< via1 >>
rect 9750 103740 9890 103750
rect 9510 102260 9570 102910
rect 9750 101420 9760 103740
rect 9760 101420 9840 103740
rect 9840 101420 9890 103740
rect 9750 101410 9890 101420
<< metal2 >>
rect 9800 103760 10000 103800
rect 9740 103750 10000 103760
rect 9500 102910 9580 102920
rect 9500 102260 9510 102910
rect 9570 102260 9580 102910
rect 9500 102250 9580 102260
rect 9740 101410 9750 103750
rect 9890 101410 10000 103750
rect 9740 101400 10000 101410
<< via2 >>
rect 9510 102260 9570 102910
<< metal3 >>
rect 16000 121800 22000 124000
rect 68194 123800 73194 124000
rect 68194 122300 73200 123800
rect 68200 122000 73200 122300
rect 16000 116200 16200 121800
rect 21800 116200 22000 121800
rect 16000 116000 22000 116200
rect 120000 121800 126000 124000
rect 165594 122300 170594 124000
rect 170894 122300 173094 124000
rect 173394 122300 175594 124000
rect 175894 122300 180894 124000
rect 217294 122300 222294 124000
rect 222594 122300 224794 124000
rect 225094 122300 227294 124000
rect 227594 122300 232594 124000
rect 318994 122300 323994 124000
rect 324294 122300 326494 124000
rect 326794 122300 328994 124000
rect 329294 122300 334294 124000
rect 413394 122300 418394 124000
rect 465394 123600 470400 124000
rect 465394 122300 465600 123600
rect 120000 116200 120200 121800
rect 125800 116200 126000 121800
rect 120000 116000 126000 116200
rect 166000 121800 170000 122300
rect 166000 115200 166200 121800
rect 169800 115200 170000 121800
rect 166000 115000 170000 115200
rect 218000 121800 222000 122300
rect 218000 115200 218200 121800
rect 221800 115200 222000 121800
rect 465400 121400 465600 122300
rect 469800 121400 470400 123600
rect 510594 123200 515394 124000
rect 510594 122340 515400 123200
rect 520594 122340 525394 124000
rect 465400 121200 470400 121400
rect 510600 122200 515400 122340
rect 566594 122300 571594 124000
rect 510600 116200 510800 122200
rect 515200 116200 515400 122200
rect 510600 115800 515400 116200
rect 218000 115000 222000 115200
rect 0 103000 1700 105242
rect 0 102920 9500 103000
rect 0 102910 9580 102920
rect 0 102260 9510 102910
rect 9570 102260 9580 102910
rect 0 102250 9580 102260
rect 0 102200 9500 102250
rect 0 100242 1700 102200
rect 3000 99000 8000 102200
rect 1000 72000 9000 99000
rect 582300 97984 584000 102984
rect 3000 69800 8000 72000
rect 0 63842 1660 68642
rect 3000 67200 3200 69800
rect 7800 67600 8000 69800
rect 7800 67200 9800 67600
rect 3000 67000 9800 67200
rect 582340 59784 584000 64584
rect 0 53842 1660 58642
rect 582340 49784 584000 54584
rect 583520 9472 584800 9584
rect 583520 8290 584800 8402
rect 583520 7108 584800 7220
rect 583520 5926 584800 6038
rect 583520 4744 584800 4856
rect 583520 3562 584800 3674
rect 20000 0 20112 400
rect 25400 0 25512 400
rect 30800 0 30912 400
rect 36200 0 36312 400
rect 41600 0 41712 400
rect 47000 0 47112 400
rect 52400 0 52512 400
rect 57800 0 57912 400
rect 63200 0 63312 400
rect 68600 0 68712 400
rect 74000 0 74112 400
rect 79400 0 79512 400
rect 84800 0 84912 400
rect 90200 0 90312 400
rect 95600 0 95712 400
rect 101000 0 101112 400
rect 106400 0 106512 400
rect 111800 0 111912 400
rect 117200 0 117312 400
rect 122600 0 122712 400
rect 128000 0 128112 400
rect 133400 0 133512 400
rect 138800 0 138912 400
rect 144200 0 144312 400
rect 149600 0 149712 400
rect 155000 0 155112 400
rect 160400 0 160512 400
rect 165800 0 165912 400
rect 171200 0 171312 400
rect 176600 0 176712 400
rect 182000 0 182112 400
rect 187400 0 187512 400
rect 192800 0 192912 400
rect 198200 0 198312 400
rect 203600 0 203712 400
rect 209000 0 209112 400
rect 214400 0 214512 400
rect 219800 0 219912 400
rect 225200 0 225312 400
rect 230600 0 230712 400
rect 236000 0 236112 400
rect 241400 0 241512 400
rect 246800 0 246912 400
rect 252200 0 252312 400
rect 257600 0 257712 400
rect 263000 0 263112 400
rect 268400 0 268512 400
rect 273800 0 273912 400
rect 279200 0 279312 400
rect 284600 0 284712 400
rect 290000 0 290112 400
rect 295400 0 295512 400
rect 300800 0 300912 400
rect 306200 0 306312 400
rect 311600 0 311712 400
rect 317000 0 317112 400
rect 322400 0 322512 400
rect 327800 0 327912 400
rect 333200 0 333312 400
rect 338600 0 338712 400
rect 344000 0 344112 400
rect 349400 0 349512 400
rect 354800 0 354912 400
rect 360200 0 360312 400
rect 365600 0 365712 400
rect 371000 0 371112 400
rect 376400 0 376512 400
rect 381800 0 381912 400
rect 387200 0 387312 400
rect 392600 0 392712 400
rect 398000 0 398112 400
rect 403400 0 403512 400
rect 408800 0 408912 400
rect 414200 0 414312 400
rect 419600 0 419712 400
rect 425000 0 425112 400
rect 430400 0 430512 400
rect 435800 0 435912 400
rect 441200 0 441312 400
rect 446600 0 446712 400
rect 452000 0 452112 400
rect 457400 0 457512 400
rect 462800 0 462912 400
rect 468200 0 468312 400
rect 473600 0 473712 400
rect 479000 0 479112 400
rect 484400 0 484512 400
rect 489800 0 489912 400
rect 495200 0 495312 400
rect 500600 0 500712 400
rect 506000 0 506112 400
rect 511400 0 511512 400
<< via3 >>
rect 16200 116200 21800 121800
rect 120200 116200 125800 121800
rect 166200 115200 169800 121800
rect 218200 115200 221800 121800
rect 465600 121400 469800 123600
rect 510800 116200 515200 122200
rect 3200 67200 7800 69800
<< mimcap >>
rect 1200 98600 8800 98800
rect 1200 72400 1400 98600
rect 8600 72400 8800 98600
rect 1200 72200 8800 72400
<< mimcapcontact >>
rect 1400 72400 8600 98600
<< metal4 >>
rect 465400 123600 470000 123800
rect 16000 121800 22000 122000
rect 16000 116200 16200 121800
rect 21800 116200 22000 121800
rect 16000 116000 22000 116200
rect 120000 121800 126000 122000
rect 120000 116200 120200 121800
rect 125800 116200 126000 121800
rect 120000 116000 126000 116200
rect 166000 121800 170000 122000
rect 166000 115200 166200 121800
rect 169800 115200 170000 121800
rect 166000 110000 170000 115200
rect 218000 121800 222000 122000
rect 218000 115200 218200 121800
rect 221800 115200 222000 121800
rect 465400 121400 465600 123600
rect 469800 121400 470000 123600
rect 465400 121200 470000 121400
rect 510600 122200 515400 122400
rect 510600 116200 510800 122200
rect 515200 116200 515400 122200
rect 510600 115800 515400 116200
rect 218000 108000 222000 115200
rect 170000 105000 222000 108000
rect 1000 98600 9000 99000
rect 1000 72400 1400 98600
rect 8600 72400 9000 98600
rect 1000 72000 9000 72400
rect 3000 69800 8000 70000
rect 3000 67200 3200 69800
rect 7800 67200 8000 69800
rect 3000 67000 8000 67200
rect 6098 0 13798 800
rect 14458 0 22158 800
rect 24098 0 31798 800
rect 564098 0 571798 800
rect 572458 0 580158 800
<< via4 >>
rect 16200 116200 21800 121800
rect 120200 116200 125800 121800
rect 465600 121400 469800 123600
rect 3200 67200 7800 69800
<< mimcap2 >>
rect 1200 98600 8800 98800
rect 1200 72400 1400 98600
rect 8600 72400 8800 98600
rect 1200 72200 8800 72400
<< mimcap2contact >>
rect 1400 72400 8600 98600
<< metal5 >>
rect 465400 123600 470000 123800
rect 16000 121800 22000 122000
rect 16000 116200 16200 121800
rect 21800 120000 22000 121800
rect 120000 121800 126000 122000
rect 21800 116200 56000 120000
rect 16000 116000 56000 116200
rect 120000 116200 120200 121800
rect 125800 120000 126000 121800
rect 465400 121400 465600 123600
rect 469800 121400 470000 123600
rect 465400 121200 470000 121400
rect 125800 116200 138000 120000
rect 466000 119800 469400 121200
rect 120000 116000 138000 116200
rect 52000 110000 56000 116000
rect 134000 110000 138000 116000
rect 1000 98600 9000 99000
rect 1000 72400 1400 98600
rect 8600 72400 9000 98600
rect 1000 72000 9000 72400
rect 3000 69800 8000 72000
rect 3000 67200 3200 69800
rect 7800 67200 8000 69800
rect 3000 67000 8000 67200
use RX_top  RX_top_0
timestamp 1662175719
transform 1 0 38000 0 -1 100000
box -37000 -23800 168000 99600
use TX_top  TX_top_0
timestamp 1662096097
transform 1 0 439300 0 -1 83800
box -83500 -36200 96500 55900
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501637
transform 1 0 10000 0 -1 122000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_38
timestamp 1659501637
transform 1 0 10000 0 -1 118000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660792292
transform 1 0 66000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_1
timestamp 1660792292
transform 1 0 74000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_2
timestamp 1660792292
transform 1 0 82000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_3
timestamp 1660792292
transform 1 0 90000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_4
timestamp 1660792292
transform 1 0 98000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_5
timestamp 1660792292
transform 1 0 106000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_6
timestamp 1660792292
transform 1 0 110000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_7
timestamp 1660792292
transform 1 0 142000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_8
timestamp 1660792292
transform 1 0 150000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_9
timestamp 1660792292
transform 1 0 154000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_10
timestamp 1660792292
transform 1 0 194000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_11
timestamp 1660792292
transform 1 0 186000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_12
timestamp 1660792292
transform 1 0 182000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_13
timestamp 1660792292
transform 1 0 202000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_14
timestamp 1660792292
transform 1 0 206000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_15
timestamp 1660792292
transform 1 0 214000 0 -1 22000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_16
timestamp 1660792292
transform 1 0 222000 0 -1 22000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_17
timestamp 1660792292
transform 1 0 230000 0 -1 22000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_70
timestamp 1660792292
transform 1 0 58000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_80
timestamp 1660792292
transform 1 0 206000 0 -1 22000
box 0 0 8000 8000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1662168084
transform 1 0 206000 0 1 86000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_1
timestamp 1662168084
transform 1 0 222000 0 1 86000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_2
timestamp 1662168084
transform 1 0 222000 0 1 70000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_3
timestamp 1662168084
transform 1 0 206000 0 1 70000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_4
timestamp 1662168084
transform 1 0 222000 0 1 54000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_5
timestamp 1662168084
transform 1 0 206000 0 1 54000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_6
timestamp 1662168084
transform 1 0 222000 0 1 38000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_7
timestamp 1662168084
transform 1 0 206000 0 1 38000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_8
timestamp 1662168084
transform 1 0 222000 0 1 22000
box 0 0 16000 16000
use hash_m1m2m3m4_W160L160_flat  hash_m1m2m3m4_W160L160_flat_9
timestamp 1662168084
transform 1 0 206000 0 1 22000
box 0 0 16000 16000
use sky130_fd_pr__nfet_01v8_NLRNVT  sky130_fd_pr__nfet_01v8_NLRNVT_0
timestamp 1662175719
transform 1 0 9611 0 1 102587
box -211 -1187 211 1187
<< labels >>
rlabel metal3 s 583520 3562 584800 3674 4 gpio_analog[6]
port 1 nsew
rlabel metal3 s 583520 4744 584800 4856 4 gpio_noesd[6]
port 2 nsew
rlabel metal3 s 582300 97984 584000 102984 4 io_analog[0]
port 3 nsew
rlabel metal3 s 566594 122300 571594 124000 4 io_analog[1]
port 4 nsew
rlabel metal3 s 465394 122300 470394 124000 4 io_analog[2]
port 5 nsew
rlabel metal3 s 413394 122300 418394 124000 4 io_analog[3]
port 6 nsew
rlabel metal3 s 318994 122300 323994 124000 4 io_analog[4]
port 7 nsew
rlabel metal3 s 326794 122300 328994 124000 4 io_clamp_high[0]
port 8 nsew
rlabel metal3 s 324294 122300 326494 124000 4 io_clamp_low[0]
port 9 nsew
rlabel metal3 s 583520 7108 584800 7220 4 io_in[13]
port 10 nsew
rlabel metal3 s 583520 5926 584800 6038 4 io_in_3v3[13]
port 11 nsew
rlabel metal3 s 583520 9472 584800 9584 4 io_oeb[13]
port 12 nsew
rlabel metal3 s 583520 8290 584800 8402 4 io_out[13]
port 13 nsew
rlabel metal3 s 582340 49784 584000 54584 4 vccd1
port 14 nsew
rlabel metal3 s 510594 122340 515394 124000 4 vssa1
port 15 nsew
rlabel metal3 s 173394 122300 175594 124000 4 io_clamp_high[2]
port 16 nsew
rlabel metal3 s 217294 122300 222294 124000 4 io_analog[5]
port 17 nsew
rlabel metal3 s 222594 122300 224794 124000 4 io_clamp_low[1]
port 18 nsew
rlabel metal3 s 170894 122300 173094 124000 4 io_clamp_low[2]
port 19 nsew
rlabel metal3 s 165594 122300 170594 124000 4 io_analog[6]
port 20 nsew
rlabel metal3 s 120194 122300 125194 124000 4 io_analog[7]
port 21 nsew
rlabel metal3 s 68194 122300 73194 124000 4 io_analog[8]
port 22 nsew
rlabel metal3 s 16194 122300 21194 124000 4 io_analog[9]
port 23 nsew
rlabel metal3 s 0 100242 1700 105242 4 io_analog[10]
port 24 nsew
rlabel metal3 s 0 53842 1660 58642 4 vccd2
port 25 nsew
rlabel metal3 s 225094 122300 227294 124000 4 io_clamp_high[1]
port 26 nsew
rlabel metal3 s 160400 0 160512 400 4 analog_la_out[26]
port 27 nsew
rlabel metal3 s 165800 0 165912 400 4 analog_la_out[27]
port 28 nsew
rlabel metal3 s 171200 0 171312 400 4 analog_la_out[28]
port 29 nsew
rlabel metal3 s 176600 0 176712 400 4 analog_la_out[29]
port 30 nsew
rlabel metal3 s 182000 0 182112 400 4 analog_la_in[0]
port 31 nsew
rlabel metal3 s 187400 0 187512 400 4 analog_la_in[1]
port 32 nsew
rlabel metal3 s 192800 0 192912 400 4 analog_la_in[2]
port 33 nsew
rlabel metal3 s 198200 0 198312 400 4 analog_la_in[3]
port 34 nsew
rlabel metal3 s 203600 0 203712 400 4 analog_la_in[4]
port 35 nsew
rlabel metal3 s 209000 0 209112 400 4 analog_la_in[5]
port 36 nsew
rlabel metal3 s 214400 0 214512 400 4 analog_la_in[6]
port 37 nsew
rlabel metal3 s 219800 0 219912 400 4 analog_la_in[7]
port 38 nsew
rlabel metal3 s 225200 0 225312 400 4 analog_la_in[8]
port 39 nsew
rlabel metal3 s 230600 0 230712 400 4 analog_la_in[9]
port 40 nsew
rlabel metal3 s 236000 0 236112 400 4 analog_la_in[10]
port 41 nsew
rlabel metal3 s 241400 0 241512 400 4 analog_la_in[11]
port 42 nsew
rlabel metal3 s 246800 0 246912 400 4 analog_la_in[12]
port 43 nsew
rlabel metal3 s 252200 0 252312 400 4 analog_la_in[13]
port 44 nsew
rlabel metal3 s 257600 0 257712 400 4 analog_la_in[14]
port 45 nsew
rlabel metal3 s 263000 0 263112 400 4 analog_la_in[15]
port 46 nsew
rlabel metal3 s 268400 0 268512 400 4 analog_la_in[16]
port 47 nsew
rlabel metal3 s 273800 0 273912 400 4 analog_la_in[17]
port 48 nsew
rlabel metal3 s 279200 0 279312 400 4 analog_la_in[18]
port 49 nsew
rlabel metal3 s 284600 0 284712 400 4 analog_la_in[19]
port 50 nsew
rlabel metal3 s 290000 0 290112 400 4 analog_la_in[20]
port 51 nsew
rlabel metal3 s 20000 0 20112 400 4 analog_la_out[0]
port 52 nsew
rlabel metal3 s 25400 0 25512 400 4 analog_la_out[1]
port 53 nsew
rlabel metal3 s 30800 0 30912 400 4 analog_la_out[2]
port 54 nsew
rlabel metal3 s 36200 0 36312 400 4 analog_la_out[3]
port 55 nsew
rlabel metal3 s 41600 0 41712 400 4 analog_la_out[4]
port 56 nsew
rlabel metal3 s 47000 0 47112 400 4 analog_la_out[5]
port 57 nsew
rlabel metal3 s 52400 0 52512 400 4 analog_la_out[6]
port 58 nsew
rlabel metal3 s 57800 0 57912 400 4 analog_la_out[7]
port 59 nsew
rlabel metal3 s 63200 0 63312 400 4 analog_la_out[8]
port 60 nsew
rlabel metal3 s 68600 0 68712 400 4 analog_la_out[9]
port 61 nsew
rlabel metal3 s 74000 0 74112 400 4 analog_la_out[10]
port 62 nsew
rlabel metal3 s 79400 0 79512 400 4 analog_la_out[11]
port 63 nsew
rlabel metal3 s 84800 0 84912 400 4 analog_la_out[12]
port 64 nsew
rlabel metal3 s 90200 0 90312 400 4 analog_la_out[13]
port 65 nsew
rlabel metal3 s 95600 0 95712 400 4 analog_la_out[14]
port 66 nsew
rlabel metal3 s 101000 0 101112 400 4 analog_la_out[15]
port 67 nsew
rlabel metal3 s 106400 0 106512 400 4 analog_la_out[16]
port 68 nsew
rlabel metal3 s 111800 0 111912 400 4 analog_la_out[17]
port 69 nsew
rlabel metal3 s 117200 0 117312 400 4 analog_la_out[18]
port 70 nsew
rlabel metal3 s 122600 0 122712 400 4 analog_la_out[19]
port 71 nsew
rlabel metal3 s 128000 0 128112 400 4 analog_la_out[20]
port 72 nsew
rlabel metal3 s 133400 0 133512 400 4 analog_la_out[21]
port 73 nsew
rlabel metal3 s 138800 0 138912 400 4 analog_la_out[22]
port 74 nsew
rlabel metal3 s 144200 0 144312 400 4 analog_la_out[23]
port 75 nsew
rlabel metal3 s 149600 0 149712 400 4 analog_la_out[24]
port 76 nsew
rlabel metal3 s 155000 0 155112 400 4 analog_la_out[25]
port 77 nsew
rlabel metal3 s 446600 0 446712 400 4 ctln[7]
port 78 nsew
rlabel metal3 s 452000 0 452112 400 4 ctln[8]
port 79 nsew
rlabel metal3 s 457400 0 457512 400 4 ctln[9]
port 80 nsew
rlabel metal3 s 462800 0 462912 400 4 trim[0]
port 81 nsew
rlabel metal3 s 468200 0 468312 400 4 trim[1]
port 82 nsew
rlabel metal3 s 473600 0 473712 400 4 trim[2]
port 83 nsew
rlabel metal3 s 479000 0 479112 400 4 trim[3]
port 84 nsew
rlabel metal3 s 484400 0 484512 400 4 trim[4]
port 85 nsew
rlabel metal3 s 489800 0 489912 400 4 trimb[0]
port 86 nsew
rlabel metal3 s 495200 0 495312 400 4 trimb[1]
port 87 nsew
rlabel metal3 s 500600 0 500712 400 4 trimb[2]
port 88 nsew
rlabel metal3 s 506000 0 506112 400 4 trimb[3]
port 89 nsew
rlabel metal3 s 511400 0 511512 400 4 trimb[4]
port 90 nsew
rlabel metal3 s 295400 0 295512 400 4 analog_la_in[21]
port 91 nsew
rlabel metal3 s 300800 0 300912 400 4 analog_la_in[22]
port 92 nsew
rlabel metal3 s 306200 0 306312 400 4 analog_la_in[23]
port 93 nsew
rlabel metal3 s 311600 0 311712 400 4 analog_la_in[24]
port 94 nsew
rlabel metal3 s 317000 0 317112 400 4 analog_la_in[25]
port 95 nsew
rlabel metal3 s 322400 0 322512 400 4 analog_la_in[26]
port 96 nsew
rlabel metal3 s 327800 0 327912 400 4 analog_la_in[27]
port 97 nsew
rlabel metal3 s 333200 0 333312 400 4 analog_la_in[28]
port 98 nsew
rlabel metal3 s 349400 0 349512 400 4 analog_la_in[29]
port 99 nsew
rlabel metal3 s 354800 0 354912 400 4 ctlp[0]
port 100 nsew
rlabel metal3 s 360200 0 360312 400 4 ctlp[1]
port 101 nsew
rlabel metal3 s 365600 0 365712 400 4 ctlp[2]
port 102 nsew
rlabel metal3 s 371000 0 371112 400 4 ctlp[3]
port 103 nsew
rlabel metal3 s 376400 0 376512 400 4 ctlp[4]
port 104 nsew
rlabel metal3 s 381800 0 381912 400 4 ctlp[5]
port 105 nsew
rlabel metal3 s 387200 0 387312 400 4 ctlp[6]
port 106 nsew
rlabel metal3 s 392600 0 392712 400 4 ctlp[7]
port 107 nsew
rlabel metal3 s 398000 0 398112 400 4 ctlp[8]
port 108 nsew
rlabel metal3 s 403400 0 403512 400 4 ctlp[9]
port 109 nsew
rlabel metal3 s 408800 0 408912 400 4 ctln[0]
port 110 nsew
rlabel metal3 s 414200 0 414312 400 4 ctln[1]
port 111 nsew
rlabel metal3 s 419600 0 419712 400 4 ctln[2]
port 112 nsew
rlabel metal3 s 425000 0 425112 400 4 ctln[3]
port 113 nsew
rlabel metal3 s 430400 0 430512 400 4 ctln[4]
port 114 nsew
rlabel metal3 s 435800 0 435912 400 4 ctln[5]
port 115 nsew
rlabel metal3 s 441200 0 441312 400 4 ctln[6]
port 116 nsew
rlabel metal4 s 572458 0 580158 800 4 vssa1
port 15 nsew
rlabel metal4 s 6098 0 13798 800 4 vdda2
port 117 nsew
rlabel metal4 s 14458 0 22158 800 4 vssd2
port 118 nsew
rlabel metal4 s 24098 0 31798 800 4 vssa2
port 119 nsew
rlabel metal4 s 564098 0 571798 800 4 vdda1
port 120 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 164000
string path 1929.280 0.000 1929.280 2.000 
<< end >>
