magic
tech sky130B
timestamp 1662654558
<< metal1 >>
rect -695 1555 -675 1560
rect -695 1000 -690 1555
rect -695 995 -675 1000
rect -605 875 -600 915
rect -105 875 -100 905
rect -605 870 -100 875
rect 155 750 1330 755
rect -605 705 -80 710
rect -605 675 -600 705
rect -85 675 -80 705
rect 155 695 160 750
rect 1320 695 1330 750
rect 155 690 1330 695
rect -605 670 -80 675
rect -695 580 -675 585
rect -695 25 -690 580
rect -695 20 -675 25
<< via1 >>
rect -690 1000 -640 1555
rect 1360 1000 1420 1465
rect -600 875 -105 905
rect 170 855 1330 910
rect -600 675 -85 705
rect 160 695 1320 750
rect -690 25 -620 580
rect 1360 130 1420 595
<< metal2 >>
rect -720 1555 -635 1560
rect -720 1000 -690 1555
rect -640 1000 -635 1555
rect 1355 1465 1425 1470
rect -720 990 -635 1000
rect -85 995 0 1005
rect -720 590 -645 990
rect -85 935 -80 995
rect -5 935 0 995
rect -85 930 0 935
rect 1355 1000 1360 1465
rect 1420 1000 1425 1465
rect -605 910 1335 915
rect -605 905 50 910
rect -605 875 -600 905
rect -105 875 50 905
rect -605 860 50 875
rect 125 860 170 910
rect -605 855 170 860
rect 1330 855 1335 910
rect -605 845 1335 855
rect 155 750 1330 755
rect 155 745 160 750
rect -5 740 160 745
rect -605 735 160 740
rect -605 705 -80 735
rect -605 675 -600 705
rect -85 685 -80 705
rect -5 695 160 735
rect 1320 695 1330 750
rect -5 690 1330 695
rect -5 685 0 690
rect -85 680 0 685
rect -85 675 -65 680
rect -605 670 -65 675
rect 30 665 130 670
rect 30 655 50 665
rect -75 615 50 655
rect 125 615 130 665
rect -75 610 130 615
rect 1355 595 1425 1000
rect -720 580 -615 590
rect -720 25 -690 580
rect -620 25 -615 580
rect 1355 130 1360 595
rect 1420 130 1425 595
rect 1355 125 1425 130
rect -720 20 -615 25
<< via2 >>
rect -80 935 -5 995
rect 50 860 125 910
rect -80 685 -5 735
rect 50 615 125 665
<< metal3 >>
rect -85 995 55 1015
rect -85 935 -80 995
rect -5 955 55 995
rect -5 935 0 955
rect -85 735 0 935
rect -85 685 -80 735
rect -5 685 0 735
rect -85 680 0 685
rect 45 910 130 915
rect 45 860 50 910
rect 125 860 130 910
rect 45 665 130 860
rect 45 625 50 665
rect 35 615 50 625
rect 125 615 130 665
rect 35 580 130 615
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659929390
transform 1 0 -435 0 1 -1100
box -253 1105 435 1790
use RF_nfet_8xW5p0L0p15  RF_nfet_8xW5p0L0p15_1
timestamp 1659929390
transform 1 0 -435 0 -1 2680
box -253 1105 435 1790
use RF_pfet_28xW5p0L0p15  RF_pfet_28xW5p0L0p15_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1662654558
transform 1 0 -490 0 1 50
box 490 -50 1940 693
use RF_pfet_28xW5p0L0p15  RF_pfet_28xW5p0L0p15_1
timestamp 1662654558
transform 1 0 -481 0 -1 1545
box 490 -50 1940 693
<< labels >>
rlabel metal3 -85 780 0 830 1 G1
rlabel metal3 45 780 130 830 1 G2
rlabel metal2 1355 755 1425 840 1 VH
rlabel metal2 -720 725 -645 835 1 VL
<< end >>
