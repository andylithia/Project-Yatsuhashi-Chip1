* NGSPICE file created from q1.ext - technology: sky130A

.subckt NMOS_30_0p5_30_1 SD2 G SD1 SUB
X0 SD2.t29 G SD1.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X1 SD1.t0 G SD2.t28 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X2 SD1.t6 G SD2.t27 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X3 SD2.t26 G SD1.t22 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X4 SD2.t25 G SD1.t1 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X5 SD1.t14 G SD2.t24 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X6 SD1.t7 G SD2.t23 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X7 SD1.t2 G SD2.t22 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X8 SD1.t15 G SD2.t21 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X9 SD2.t20 G SD1.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X10 SD2.t19 G SD1.t17 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X11 SD2.t18 G SD1.t8 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X12 SD1.t3 G SD2.t17 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X13 SD1.t16 G SD2.t16 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X14 SD1.t26 G SD2.t15 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X15 SD2.t14 G SD1.t18 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X16 SD2.t13 G SD1.t10 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X17 SD1.t19 G SD2.t12 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X18 SD1.t9 G SD2.t11 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X19 SD2.t10 G SD1.t4 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X20 SD1.t5 G SD2.t9 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X21 SD1.t20 G SD2.t8 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X22 SD2.t7 G SD1.t24 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X23 SD2.t6 G SD1.t25 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X24 SD2.t5 G SD1.t29 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X25 SD1.t28 G SD2.t4 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X26 SD2.t3 G SD1.t11 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X27 SD1.t13 G SD2.t2 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X28 SD2.t1 G SD1.t21 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
X29 SD2.t0 G SD1.t23 SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+07u l=500000u
C0 G SD2 19.79fF
C1 SD1 SD2 198.43fF
C2 G SD1 20.02fF
R0 SD1.n2 SD1.n16 1.435
R1 SD1 SD1.n4 1.428
R2 SD1 SD1.n5 1.428
R3 SD1 SD1.n6 1.428
R4 SD1.n0 SD1.n7 1.428
R5 SD1.n0 SD1.n8 1.428
R6 SD1.n0 SD1.n9 1.428
R7 SD1.n1 SD1.n10 1.428
R8 SD1.n1 SD1.n11 1.428
R9 SD1.n1 SD1.n12 1.428
R10 SD1.n1 SD1.n13 1.428
R11 SD1.n2 SD1.n14 1.428
R12 SD1.n2 SD1.n15 1.428
R13 SD1 SD1.n3 1.427
R14 SD1.n0 SD1.n17 1.427
R15 SD1.n3 SD1.t18 0.551
R16 SD1.n3 SD1.t28 0.551
R17 SD1.n4 SD1.t24 0.551
R18 SD1.n4 SD1.t5 0.551
R19 SD1.n5 SD1.t25 0.551
R20 SD1.n5 SD1.t3 0.551
R21 SD1.n6 SD1.t10 0.551
R22 SD1.n6 SD1.t16 0.551
R23 SD1.n7 SD1.t17 0.551
R24 SD1.n7 SD1.t15 0.551
R25 SD1.n8 SD1.t12 0.551
R26 SD1.n8 SD1.t19 0.551
R27 SD1.n9 SD1.t21 0.551
R28 SD1.n9 SD1.t14 0.551
R29 SD1.n10 SD1.t27 0.551
R30 SD1.n10 SD1.t13 0.551
R31 SD1.n11 SD1.t29 0.551
R32 SD1.n11 SD1.t9 0.551
R33 SD1.n12 SD1.t4 0.551
R34 SD1.n12 SD1.t26 0.551
R35 SD1.n13 SD1.t8 0.551
R36 SD1.n13 SD1.t20 0.551
R37 SD1.n14 SD1.t22 0.551
R38 SD1.n14 SD1.t2 0.551
R39 SD1.n15 SD1.t23 0.551
R40 SD1.n15 SD1.t7 0.551
R41 SD1.n16 SD1.t1 0.551
R42 SD1.n16 SD1.t6 0.551
R43 SD1.n17 SD1.t11 0.551
R44 SD1.n17 SD1.t0 0.551
R45 SD1 SD1.n0 0.042
R46 SD1.n0 SD1.n1 0.028
R47 SD1.n1 SD1.n2 0.021
R48 SD2.n13 SD2.t25 1.972
R49 SD2 SD2.t4 1.965
R50 SD2.n27 SD2.n0 1.414
R51 SD2.n26 SD2.n1 1.414
R52 SD2.n25 SD2.n2 1.414
R53 SD2.n24 SD2.n3 1.414
R54 SD2.n23 SD2.n4 1.414
R55 SD2.n22 SD2.n5 1.414
R56 SD2.n19 SD2.n6 1.414
R57 SD2.n18 SD2.n7 1.414
R58 SD2.n17 SD2.n8 1.414
R59 SD2.n16 SD2.n9 1.414
R60 SD2.n15 SD2.n10 1.414
R61 SD2.n14 SD2.n11 1.414
R62 SD2.n13 SD2.n12 1.414
R63 SD2.n21 SD2.n20 1.413
R64 SD2.n0 SD2.t9 0.551
R65 SD2.n0 SD2.t14 0.551
R66 SD2.n1 SD2.t17 0.551
R67 SD2.n1 SD2.t7 0.551
R68 SD2.n2 SD2.t16 0.551
R69 SD2.n2 SD2.t6 0.551
R70 SD2.n3 SD2.t21 0.551
R71 SD2.n3 SD2.t13 0.551
R72 SD2.n4 SD2.t12 0.551
R73 SD2.n4 SD2.t19 0.551
R74 SD2.n5 SD2.t24 0.551
R75 SD2.n5 SD2.t20 0.551
R76 SD2.n6 SD2.t2 0.551
R77 SD2.n6 SD2.t3 0.551
R78 SD2.n7 SD2.t11 0.551
R79 SD2.n7 SD2.t29 0.551
R80 SD2.n8 SD2.t15 0.551
R81 SD2.n8 SD2.t5 0.551
R82 SD2.n9 SD2.t8 0.551
R83 SD2.n9 SD2.t10 0.551
R84 SD2.n10 SD2.t22 0.551
R85 SD2.n10 SD2.t18 0.551
R86 SD2.n11 SD2.t23 0.551
R87 SD2.n11 SD2.t26 0.551
R88 SD2.n12 SD2.t27 0.551
R89 SD2.n12 SD2.t0 0.551
R90 SD2.n20 SD2.t28 0.551
R91 SD2.n20 SD2.t1 0.551
R92 SD2.n14 SD2.n13 0.007
R93 SD2.n15 SD2.n14 0.007
R94 SD2.n16 SD2.n15 0.007
R95 SD2.n17 SD2.n16 0.007
R96 SD2.n18 SD2.n17 0.007
R97 SD2.n19 SD2.n18 0.007
R98 SD2.n21 SD2.n19 0.007
R99 SD2.n22 SD2.n21 0.007
R100 SD2.n23 SD2.n22 0.007
R101 SD2.n24 SD2.n23 0.007
R102 SD2.n25 SD2.n24 0.007
R103 SD2.n26 SD2.n25 0.007
R104 SD2.n27 SD2.n26 0.007
R105 SD2 SD2.n27 0.007
C3 SD1 SUB 32.55fF
C4 SD2 SUB 24.38fF
C5 G SUB 24.46fF $ **FLOATING
C6 SD2.t4 SUB 5.46fF $ **FLOATING
C7 SD2.n0 SUB 6.06fF
C8 SD2.n1 SUB 6.06fF
C9 SD2.n2 SUB 6.06fF
C10 SD2.n3 SUB 6.06fF
C11 SD2.n4 SUB 6.06fF
C12 SD2.n5 SUB 6.06fF
C13 SD2.n6 SUB 6.06fF
C14 SD2.n7 SUB 6.06fF
C15 SD2.n8 SUB 6.06fF
C16 SD2.n9 SUB 6.06fF
C17 SD2.n10 SUB 6.06fF
C18 SD2.n11 SUB 6.06fF
C19 SD2.n12 SUB 6.06fF
C20 SD2.t25 SUB 5.49fF $ **FLOATING
C21 SD2.n13 SUB 16.50fF
C22 SD2.n14 SUB 7.22fF
C23 SD2.n15 SUB 7.22fF
C24 SD2.n16 SUB 7.22fF
C25 SD2.n17 SUB 7.22fF
C26 SD2.n18 SUB 7.22fF
C27 SD2.n19 SUB 7.22fF
C28 SD2.n20 SUB 6.06fF
C29 SD2.n21 SUB 7.22fF
C30 SD2.n22 SUB 7.22fF
C31 SD2.n23 SUB 7.22fF
C32 SD2.n24 SUB 7.22fF
C33 SD2.n25 SUB 7.22fF
C34 SD2.n26 SUB 7.22fF
C35 SD2.n27 SUB 7.22fF
C36 SD1.n0 SUB 28.23fF
C37 SD1.n1 SUB 28.23fF
C38 SD1.n2 SUB 23.60fF
C39 SD1.n3 SUB 5.93fF
C40 SD1.n4 SUB 5.93fF
C41 SD1.n5 SUB 5.93fF
C42 SD1.n6 SUB 5.93fF
C43 SD1.n7 SUB 5.93fF
C44 SD1.n8 SUB 5.93fF
C45 SD1.n9 SUB 5.93fF
C46 SD1.n10 SUB 5.93fF
C47 SD1.n11 SUB 5.93fF
C48 SD1.n12 SUB 5.93fF
C49 SD1.n13 SUB 5.93fF
C50 SD1.n14 SUB 5.93fF
C51 SD1.n15 SUB 5.93fF
C52 SD1.n16 SUB 5.97fF
C53 SD1.n17 SUB 5.93fF
.ends
