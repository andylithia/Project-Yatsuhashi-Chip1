magic
tech sky130B
magscale 1 2
timestamp 1661296025
<< pwell >>
rect -26 -26 176 174
<< scnmos >>
rect 60 0 90 148
<< ndiff >>
rect 0 0 60 148
rect 90 0 150 148
<< poly >>
rect 60 148 90 174
rect 60 -26 90 0
<< locali >>
rect 108 41 142 107
use sky130_sram_1r1w_24x128_8_contact_10  sky130_sram_1r1w_24x128_8_contact_10_0
timestamp 1661296025
transform 1 0 100 0 1 41
box -26 -22 76 88
<< labels >>
rlabel poly s 75 74 75 74 4 G
port 1 nsew
rlabel mvpsubdiff s 25 74 25 74 4 S
rlabel locali s 125 74 125 74 4 D
port 2 nsew
<< properties >>
string FIXED_BBOX -25 -26 175 174
<< end >>
